magic
tech ihp-sg13g2
magscale 1 2
timestamp 1753877633
<< metal1 >>
rect 1152 41600 20452 41624
rect 1152 41560 4928 41600
rect 4968 41560 5010 41600
rect 5050 41560 5092 41600
rect 5132 41560 5174 41600
rect 5214 41560 5256 41600
rect 5296 41560 20048 41600
rect 20088 41560 20130 41600
rect 20170 41560 20212 41600
rect 20252 41560 20294 41600
rect 20334 41560 20376 41600
rect 20416 41560 20452 41600
rect 1152 41536 20452 41560
rect 1515 41432 1557 41441
rect 1515 41392 1516 41432
rect 1556 41392 1557 41432
rect 1515 41383 1557 41392
rect 19563 41432 19605 41441
rect 19563 41392 19564 41432
rect 19604 41392 19605 41432
rect 19563 41383 19605 41392
rect 19947 41432 19989 41441
rect 19947 41392 19948 41432
rect 19988 41392 19989 41432
rect 19947 41383 19989 41392
rect 1699 41264 1757 41265
rect 1699 41224 1708 41264
rect 1748 41224 1757 41264
rect 1699 41223 1757 41224
rect 2947 41264 3005 41265
rect 2947 41224 2956 41264
rect 2996 41224 3005 41264
rect 2947 41223 3005 41224
rect 3331 41264 3389 41265
rect 3331 41224 3340 41264
rect 3380 41224 3389 41264
rect 3331 41223 3389 41224
rect 4579 41264 4637 41265
rect 4579 41224 4588 41264
rect 4628 41224 4637 41264
rect 4579 41223 4637 41224
rect 4963 41264 5021 41265
rect 4963 41224 4972 41264
rect 5012 41224 5021 41264
rect 4963 41223 5021 41224
rect 6211 41264 6269 41265
rect 6211 41224 6220 41264
rect 6260 41224 6269 41264
rect 6211 41223 6269 41224
rect 6595 41264 6653 41265
rect 6595 41224 6604 41264
rect 6644 41224 6653 41264
rect 6595 41223 6653 41224
rect 7843 41264 7901 41265
rect 7843 41224 7852 41264
rect 7892 41224 7901 41264
rect 7843 41223 7901 41224
rect 8227 41264 8285 41265
rect 8227 41224 8236 41264
rect 8276 41224 8285 41264
rect 8227 41223 8285 41224
rect 9475 41264 9533 41265
rect 9475 41224 9484 41264
rect 9524 41224 9533 41264
rect 9475 41223 9533 41224
rect 10243 41264 10301 41265
rect 10243 41224 10252 41264
rect 10292 41224 10301 41264
rect 10243 41223 10301 41224
rect 10627 41264 10685 41265
rect 10627 41224 10636 41264
rect 10676 41224 10685 41264
rect 10627 41223 10685 41224
rect 11875 41264 11933 41265
rect 11875 41224 11884 41264
rect 11924 41224 11933 41264
rect 11875 41223 11933 41224
rect 12451 41264 12509 41265
rect 12451 41224 12460 41264
rect 12500 41224 12509 41264
rect 12451 41223 12509 41224
rect 13699 41264 13757 41265
rect 13699 41224 13708 41264
rect 13748 41224 13757 41264
rect 13699 41223 13757 41224
rect 14083 41264 14141 41265
rect 14083 41224 14092 41264
rect 14132 41224 14141 41264
rect 14083 41223 14141 41224
rect 15331 41264 15389 41265
rect 15331 41224 15340 41264
rect 15380 41224 15389 41264
rect 15331 41223 15389 41224
rect 15715 41264 15773 41265
rect 15715 41224 15724 41264
rect 15764 41224 15773 41264
rect 15715 41223 15773 41224
rect 16963 41264 17021 41265
rect 16963 41224 16972 41264
rect 17012 41224 17021 41264
rect 16963 41223 17021 41224
rect 1315 41180 1373 41181
rect 1315 41140 1324 41180
rect 1364 41140 1373 41180
rect 1315 41139 1373 41140
rect 17347 41180 17405 41181
rect 17347 41140 17356 41180
rect 17396 41140 17405 41180
rect 17347 41139 17405 41140
rect 17731 41180 17789 41181
rect 17731 41140 17740 41180
rect 17780 41140 17789 41180
rect 17731 41139 17789 41140
rect 18115 41180 18173 41181
rect 18115 41140 18124 41180
rect 18164 41140 18173 41180
rect 18115 41139 18173 41140
rect 18499 41180 18557 41181
rect 18499 41140 18508 41180
rect 18548 41140 18557 41180
rect 18499 41139 18557 41140
rect 18883 41180 18941 41181
rect 18883 41140 18892 41180
rect 18932 41140 18941 41180
rect 18883 41139 18941 41140
rect 19363 41180 19421 41181
rect 19363 41140 19372 41180
rect 19412 41140 19421 41180
rect 19363 41139 19421 41140
rect 19747 41180 19805 41181
rect 19747 41140 19756 41180
rect 19796 41140 19805 41180
rect 19747 41139 19805 41140
rect 20120 41177 20162 41186
rect 20120 41137 20121 41177
rect 20161 41137 20162 41177
rect 20120 41128 20162 41137
rect 9867 41096 9909 41105
rect 9867 41056 9868 41096
rect 9908 41056 9909 41096
rect 9867 41047 9909 41056
rect 19179 41096 19221 41105
rect 19179 41056 19180 41096
rect 19220 41056 19221 41096
rect 19179 41047 19221 41056
rect 3147 41012 3189 41021
rect 3147 40972 3148 41012
rect 3188 40972 3189 41012
rect 3147 40963 3189 40972
rect 4779 41012 4821 41021
rect 4779 40972 4780 41012
rect 4820 40972 4821 41012
rect 4779 40963 4821 40972
rect 6411 41012 6453 41021
rect 6411 40972 6412 41012
rect 6452 40972 6453 41012
rect 6411 40963 6453 40972
rect 8043 41012 8085 41021
rect 8043 40972 8044 41012
rect 8084 40972 8085 41012
rect 8043 40963 8085 40972
rect 9675 41012 9717 41021
rect 9675 40972 9676 41012
rect 9716 40972 9717 41012
rect 9675 40963 9717 40972
rect 10155 41012 10197 41021
rect 10155 40972 10156 41012
rect 10196 40972 10197 41012
rect 10155 40963 10197 40972
rect 12075 41012 12117 41021
rect 12075 40972 12076 41012
rect 12116 40972 12117 41012
rect 12075 40963 12117 40972
rect 12267 41012 12309 41021
rect 12267 40972 12268 41012
rect 12308 40972 12309 41012
rect 12267 40963 12309 40972
rect 13899 41012 13941 41021
rect 13899 40972 13900 41012
rect 13940 40972 13941 41012
rect 13899 40963 13941 40972
rect 15531 41012 15573 41021
rect 15531 40972 15532 41012
rect 15572 40972 15573 41012
rect 15531 40963 15573 40972
rect 17163 41012 17205 41021
rect 17163 40972 17164 41012
rect 17204 40972 17205 41012
rect 17163 40963 17205 40972
rect 17547 41012 17589 41021
rect 17547 40972 17548 41012
rect 17588 40972 17589 41012
rect 17547 40963 17589 40972
rect 17931 41012 17973 41021
rect 17931 40972 17932 41012
rect 17972 40972 17973 41012
rect 17931 40963 17973 40972
rect 18315 41012 18357 41021
rect 18315 40972 18316 41012
rect 18356 40972 18357 41012
rect 18315 40963 18357 40972
rect 18699 41012 18741 41021
rect 18699 40972 18700 41012
rect 18740 40972 18741 41012
rect 18699 40963 18741 40972
rect 1152 40844 20352 40868
rect 1152 40804 3688 40844
rect 3728 40804 3770 40844
rect 3810 40804 3852 40844
rect 3892 40804 3934 40844
rect 3974 40804 4016 40844
rect 4056 40804 18808 40844
rect 18848 40804 18890 40844
rect 18930 40804 18972 40844
rect 19012 40804 19054 40844
rect 19094 40804 19136 40844
rect 19176 40804 20352 40844
rect 1152 40780 20352 40804
rect 1611 40676 1653 40685
rect 1611 40636 1612 40676
rect 1652 40636 1653 40676
rect 1611 40627 1653 40636
rect 5835 40676 5877 40685
rect 5835 40636 5836 40676
rect 5876 40636 5877 40676
rect 5835 40627 5877 40636
rect 7659 40676 7701 40685
rect 7659 40636 7660 40676
rect 7700 40636 7701 40676
rect 7659 40627 7701 40636
rect 14283 40676 14325 40685
rect 14283 40636 14284 40676
rect 14324 40636 14325 40676
rect 14283 40627 14325 40636
rect 18411 40676 18453 40685
rect 18411 40636 18412 40676
rect 18452 40636 18453 40676
rect 18411 40627 18453 40636
rect 18795 40676 18837 40685
rect 18795 40636 18796 40676
rect 18836 40636 18837 40676
rect 18795 40627 18837 40636
rect 19947 40676 19989 40685
rect 19947 40636 19948 40676
rect 19988 40636 19989 40676
rect 19947 40627 19989 40636
rect 2091 40592 2133 40601
rect 2091 40552 2092 40592
rect 2132 40552 2133 40592
rect 2091 40543 2133 40552
rect 14571 40592 14613 40601
rect 14571 40552 14572 40592
rect 14612 40552 14613 40592
rect 14571 40543 14613 40552
rect 17163 40592 17205 40601
rect 17163 40552 17164 40592
rect 17204 40552 17205 40592
rect 17163 40543 17205 40552
rect 17547 40592 17589 40601
rect 17547 40552 17548 40592
rect 17588 40552 17589 40592
rect 17547 40543 17589 40552
rect 17931 40592 17973 40601
rect 17931 40552 17932 40592
rect 17972 40552 17973 40592
rect 17931 40543 17973 40552
rect 19371 40592 19413 40601
rect 19371 40552 19372 40592
rect 19412 40552 19413 40592
rect 19371 40543 19413 40552
rect 1411 40508 1469 40509
rect 1411 40468 1420 40508
rect 1460 40468 1469 40508
rect 1411 40467 1469 40468
rect 1891 40508 1949 40509
rect 1891 40468 1900 40508
rect 1940 40468 1949 40508
rect 1891 40467 1949 40468
rect 5635 40508 5693 40509
rect 5635 40468 5644 40508
rect 5684 40468 5693 40508
rect 5635 40467 5693 40468
rect 7843 40508 7901 40509
rect 7843 40468 7852 40508
rect 7892 40468 7901 40508
rect 7843 40467 7901 40468
rect 10443 40508 10485 40517
rect 10443 40468 10444 40508
rect 10484 40468 10485 40508
rect 10443 40459 10485 40468
rect 10539 40508 10581 40517
rect 10539 40468 10540 40508
rect 10580 40468 10581 40508
rect 10539 40459 10581 40468
rect 16579 40508 16637 40509
rect 16579 40468 16588 40508
rect 16628 40468 16637 40508
rect 16579 40467 16637 40468
rect 16963 40508 17021 40509
rect 16963 40468 16972 40508
rect 17012 40468 17021 40508
rect 16963 40467 17021 40468
rect 17347 40508 17405 40509
rect 17347 40468 17356 40508
rect 17396 40468 17405 40508
rect 17347 40467 17405 40468
rect 17731 40508 17789 40509
rect 17731 40468 17740 40508
rect 17780 40468 17789 40508
rect 17731 40467 17789 40468
rect 18115 40508 18173 40509
rect 18115 40468 18124 40508
rect 18164 40468 18173 40508
rect 18115 40467 18173 40468
rect 18595 40508 18653 40509
rect 18595 40468 18604 40508
rect 18644 40468 18653 40508
rect 18595 40467 18653 40468
rect 18979 40508 19037 40509
rect 18979 40468 18988 40508
rect 19028 40468 19037 40508
rect 18979 40467 19037 40468
rect 19171 40508 19229 40509
rect 19171 40468 19180 40508
rect 19220 40468 19229 40508
rect 19171 40467 19229 40468
rect 20120 40508 20162 40517
rect 20120 40468 20121 40508
rect 20161 40468 20162 40508
rect 20120 40459 20162 40468
rect 11499 40438 11541 40447
rect 2275 40424 2333 40425
rect 2275 40384 2284 40424
rect 2324 40384 2333 40424
rect 2275 40383 2333 40384
rect 3523 40424 3581 40425
rect 3523 40384 3532 40424
rect 3572 40384 3581 40424
rect 3523 40383 3581 40384
rect 3907 40424 3965 40425
rect 3907 40384 3916 40424
rect 3956 40384 3965 40424
rect 3907 40383 3965 40384
rect 5155 40424 5213 40425
rect 5155 40384 5164 40424
rect 5204 40384 5213 40424
rect 5155 40383 5213 40384
rect 6019 40424 6077 40425
rect 6019 40384 6028 40424
rect 6068 40384 6077 40424
rect 6019 40383 6077 40384
rect 7267 40424 7325 40425
rect 7267 40384 7276 40424
rect 7316 40384 7325 40424
rect 7267 40383 7325 40384
rect 8035 40424 8093 40425
rect 8035 40384 8044 40424
rect 8084 40384 8093 40424
rect 8035 40383 8093 40384
rect 9283 40424 9341 40425
rect 9283 40384 9292 40424
rect 9332 40384 9341 40424
rect 9283 40383 9341 40384
rect 9963 40424 10005 40433
rect 9963 40384 9964 40424
rect 10004 40384 10005 40424
rect 9963 40375 10005 40384
rect 10059 40424 10101 40433
rect 10059 40384 10060 40424
rect 10100 40384 10101 40424
rect 10059 40375 10101 40384
rect 11011 40424 11069 40425
rect 11011 40384 11020 40424
rect 11060 40384 11069 40424
rect 11499 40398 11500 40438
rect 11540 40398 11541 40438
rect 13315 40445 13373 40446
rect 11499 40389 11541 40398
rect 12067 40424 12125 40425
rect 11011 40383 11069 40384
rect 12067 40384 12076 40424
rect 12116 40384 12125 40424
rect 13315 40405 13324 40445
rect 13364 40405 13373 40445
rect 13315 40404 13373 40405
rect 13741 40431 13783 40440
rect 12067 40383 12125 40384
rect 13741 40391 13742 40431
rect 13782 40391 13783 40431
rect 13741 40382 13783 40391
rect 13899 40424 13941 40433
rect 13899 40384 13900 40424
rect 13940 40384 13941 40424
rect 13899 40375 13941 40384
rect 13995 40424 14037 40433
rect 13995 40384 13996 40424
rect 14036 40384 14037 40424
rect 13995 40375 14037 40384
rect 14179 40424 14237 40425
rect 14179 40384 14188 40424
rect 14228 40384 14237 40424
rect 14179 40383 14237 40384
rect 14275 40424 14333 40425
rect 14275 40384 14284 40424
rect 14324 40384 14333 40424
rect 14275 40383 14333 40384
rect 14467 40424 14525 40425
rect 14467 40384 14476 40424
rect 14516 40384 14525 40424
rect 14467 40383 14525 40384
rect 14755 40424 14813 40425
rect 14755 40384 14764 40424
rect 14804 40384 14813 40424
rect 14755 40383 14813 40384
rect 16003 40424 16061 40425
rect 16003 40384 16012 40424
rect 16052 40384 16061 40424
rect 16003 40383 16061 40384
rect 19563 40424 19605 40433
rect 19563 40384 19564 40424
rect 19604 40384 19605 40424
rect 19563 40375 19605 40384
rect 19755 40424 19797 40433
rect 19755 40384 19756 40424
rect 19796 40384 19797 40424
rect 19755 40375 19797 40384
rect 5355 40340 5397 40349
rect 5355 40300 5356 40340
rect 5396 40300 5397 40340
rect 5355 40291 5397 40300
rect 9483 40340 9525 40349
rect 9483 40300 9484 40340
rect 9524 40300 9525 40340
rect 9483 40291 9525 40300
rect 13515 40340 13557 40349
rect 13515 40300 13516 40340
rect 13556 40300 13557 40340
rect 13515 40291 13557 40300
rect 3723 40256 3765 40265
rect 3723 40216 3724 40256
rect 3764 40216 3765 40256
rect 3723 40207 3765 40216
rect 7467 40256 7509 40265
rect 7467 40216 7468 40256
rect 7508 40216 7509 40256
rect 7467 40207 7509 40216
rect 11691 40256 11733 40265
rect 11691 40216 11692 40256
rect 11732 40216 11733 40256
rect 11691 40207 11733 40216
rect 16203 40256 16245 40265
rect 16203 40216 16204 40256
rect 16244 40216 16245 40256
rect 16203 40207 16245 40216
rect 16395 40256 16437 40265
rect 16395 40216 16396 40256
rect 16436 40216 16437 40256
rect 16395 40207 16437 40216
rect 16779 40256 16821 40265
rect 16779 40216 16780 40256
rect 16820 40216 16821 40256
rect 16779 40207 16821 40216
rect 19659 40256 19701 40265
rect 19659 40216 19660 40256
rect 19700 40216 19701 40256
rect 19659 40207 19701 40216
rect 1152 40088 20452 40112
rect 1152 40048 4928 40088
rect 4968 40048 5010 40088
rect 5050 40048 5092 40088
rect 5132 40048 5174 40088
rect 5214 40048 5256 40088
rect 5296 40048 20048 40088
rect 20088 40048 20130 40088
rect 20170 40048 20212 40088
rect 20252 40048 20294 40088
rect 20334 40048 20376 40088
rect 20416 40048 20452 40088
rect 1152 40024 20452 40048
rect 3915 39920 3957 39929
rect 3915 39880 3916 39920
rect 3956 39880 3957 39920
rect 3915 39871 3957 39880
rect 4299 39920 4341 39929
rect 4299 39880 4300 39920
rect 4340 39880 4341 39920
rect 4299 39871 4341 39880
rect 4683 39920 4725 39929
rect 4683 39880 4684 39920
rect 4724 39880 4725 39920
rect 4683 39871 4725 39880
rect 5067 39920 5109 39929
rect 5067 39880 5068 39920
rect 5108 39880 5109 39920
rect 5067 39871 5109 39880
rect 7843 39920 7901 39921
rect 7843 39880 7852 39920
rect 7892 39880 7901 39920
rect 7843 39879 7901 39880
rect 10531 39920 10589 39921
rect 10531 39880 10540 39920
rect 10580 39880 10589 39920
rect 10531 39879 10589 39880
rect 10819 39920 10877 39921
rect 10819 39880 10828 39920
rect 10868 39880 10877 39920
rect 10819 39879 10877 39880
rect 14667 39920 14709 39929
rect 14667 39880 14668 39920
rect 14708 39880 14709 39920
rect 14667 39871 14709 39880
rect 15331 39920 15389 39921
rect 15331 39880 15340 39920
rect 15380 39880 15389 39920
rect 15331 39879 15389 39880
rect 17835 39920 17877 39929
rect 17835 39880 17836 39920
rect 17876 39880 17877 39920
rect 17835 39871 17877 39880
rect 18027 39920 18069 39929
rect 18027 39880 18028 39920
rect 18068 39880 18069 39920
rect 18027 39871 18069 39880
rect 1419 39836 1461 39845
rect 1419 39796 1420 39836
rect 1460 39796 1461 39836
rect 1419 39787 1461 39796
rect 3531 39836 3573 39845
rect 3531 39796 3532 39836
rect 3572 39796 3573 39836
rect 3531 39787 3573 39796
rect 7371 39836 7413 39845
rect 7371 39796 7372 39836
rect 7412 39796 7413 39836
rect 7371 39787 7413 39796
rect 14379 39836 14421 39845
rect 14379 39796 14380 39836
rect 14420 39796 14421 39836
rect 14379 39787 14421 39796
rect 2083 39752 2141 39753
rect 1611 39738 1653 39747
rect 1611 39698 1612 39738
rect 1652 39698 1653 39738
rect 2083 39712 2092 39752
rect 2132 39712 2141 39752
rect 2083 39711 2141 39712
rect 2667 39752 2709 39761
rect 2667 39712 2668 39752
rect 2708 39712 2709 39752
rect 2667 39703 2709 39712
rect 3051 39752 3093 39761
rect 3051 39712 3052 39752
rect 3092 39712 3093 39752
rect 3051 39703 3093 39712
rect 3147 39752 3189 39761
rect 3147 39712 3148 39752
rect 3188 39712 3189 39752
rect 3147 39703 3189 39712
rect 5347 39752 5405 39753
rect 5347 39712 5356 39752
rect 5396 39712 5405 39752
rect 5347 39711 5405 39712
rect 5643 39752 5685 39761
rect 5643 39712 5644 39752
rect 5684 39712 5685 39752
rect 5643 39703 5685 39712
rect 5739 39752 5781 39761
rect 5739 39712 5740 39752
rect 5780 39712 5781 39752
rect 5739 39703 5781 39712
rect 6691 39752 6749 39753
rect 6691 39712 6700 39752
rect 6740 39712 6749 39752
rect 6691 39711 6749 39712
rect 7179 39747 7221 39756
rect 7179 39707 7180 39747
rect 7220 39707 7221 39747
rect 7179 39698 7221 39707
rect 7563 39752 7605 39761
rect 7563 39712 7564 39752
rect 7604 39712 7605 39752
rect 7563 39703 7605 39712
rect 7659 39752 7701 39761
rect 7659 39712 7660 39752
rect 7700 39712 7701 39752
rect 7659 39703 7701 39712
rect 8227 39752 8285 39753
rect 8227 39712 8236 39752
rect 8276 39712 8285 39752
rect 8227 39711 8285 39712
rect 9475 39752 9533 39753
rect 9475 39712 9484 39752
rect 9524 39712 9533 39752
rect 9475 39711 9533 39712
rect 11299 39752 11357 39753
rect 11299 39712 11308 39752
rect 11348 39712 11357 39752
rect 11299 39711 11357 39712
rect 12547 39752 12605 39753
rect 12547 39712 12556 39752
rect 12596 39712 12605 39752
rect 12547 39711 12605 39712
rect 12931 39752 12989 39753
rect 12931 39712 12940 39752
rect 12980 39712 12989 39752
rect 12931 39711 12989 39712
rect 14179 39752 14237 39753
rect 14179 39712 14188 39752
rect 14228 39712 14237 39752
rect 14179 39711 14237 39712
rect 14571 39752 14613 39761
rect 14571 39712 14572 39752
rect 14612 39712 14613 39752
rect 14571 39703 14613 39712
rect 14763 39752 14805 39761
rect 14763 39712 14764 39752
rect 14804 39712 14805 39752
rect 14763 39703 14805 39712
rect 14859 39752 14901 39761
rect 14859 39712 14860 39752
rect 14900 39712 14901 39752
rect 14859 39703 14901 39712
rect 15051 39752 15093 39761
rect 15051 39712 15052 39752
rect 15092 39712 15093 39752
rect 15051 39703 15093 39712
rect 15147 39752 15189 39761
rect 15147 39712 15148 39752
rect 15188 39712 15189 39752
rect 15147 39703 15189 39712
rect 16107 39752 16149 39761
rect 16107 39712 16108 39752
rect 16148 39712 16149 39752
rect 16107 39703 16149 39712
rect 16203 39752 16245 39761
rect 16203 39712 16204 39752
rect 16244 39712 16245 39752
rect 16203 39703 16245 39712
rect 17155 39752 17213 39753
rect 17155 39712 17164 39752
rect 17204 39712 17213 39752
rect 19947 39752 19989 39761
rect 17155 39711 17213 39712
rect 17691 39710 17733 39719
rect 1611 39689 1653 39698
rect 2571 39668 2613 39677
rect 2571 39628 2572 39668
rect 2612 39628 2613 39668
rect 2571 39619 2613 39628
rect 3715 39668 3773 39669
rect 3715 39628 3724 39668
rect 3764 39628 3773 39668
rect 3715 39627 3773 39628
rect 4099 39668 4157 39669
rect 4099 39628 4108 39668
rect 4148 39628 4157 39668
rect 4099 39627 4157 39628
rect 4483 39668 4541 39669
rect 4483 39628 4492 39668
rect 4532 39628 4541 39668
rect 4483 39627 4541 39628
rect 4867 39668 4925 39669
rect 4867 39628 4876 39668
rect 4916 39628 4925 39668
rect 4867 39627 4925 39628
rect 6123 39668 6165 39677
rect 6123 39628 6124 39668
rect 6164 39628 6165 39668
rect 6123 39619 6165 39628
rect 6219 39668 6261 39677
rect 6219 39628 6220 39668
rect 6260 39628 6261 39668
rect 15715 39668 15773 39669
rect 6219 39619 6261 39628
rect 10147 39665 10205 39666
rect 10147 39625 10156 39665
rect 10196 39625 10205 39665
rect 15715 39628 15724 39668
rect 15764 39628 15773 39668
rect 15715 39627 15773 39628
rect 16587 39668 16629 39677
rect 16587 39628 16588 39668
rect 16628 39628 16629 39668
rect 10147 39624 10205 39625
rect 16587 39619 16629 39628
rect 16683 39668 16725 39677
rect 16683 39628 16684 39668
rect 16724 39628 16725 39668
rect 17691 39670 17692 39710
rect 17732 39670 17733 39710
rect 19947 39712 19948 39752
rect 19988 39712 19989 39752
rect 19947 39703 19989 39712
rect 20139 39739 20181 39748
rect 20139 39699 20140 39739
rect 20180 39699 20181 39739
rect 20139 39690 20181 39699
rect 17691 39661 17733 39670
rect 18211 39668 18269 39669
rect 16683 39619 16725 39628
rect 18211 39628 18220 39668
rect 18260 39628 18269 39668
rect 18211 39627 18269 39628
rect 18595 39668 18653 39669
rect 18595 39628 18604 39668
rect 18644 39628 18653 39668
rect 18595 39627 18653 39628
rect 18787 39668 18845 39669
rect 18787 39628 18796 39668
rect 18836 39628 18845 39668
rect 18787 39627 18845 39628
rect 19171 39668 19229 39669
rect 19171 39628 19180 39668
rect 19220 39628 19229 39668
rect 19171 39627 19229 39628
rect 19555 39668 19613 39669
rect 19555 39628 19564 39668
rect 19604 39628 19613 39668
rect 19555 39627 19613 39628
rect 20043 39668 20085 39677
rect 20043 39628 20044 39668
rect 20084 39628 20085 39668
rect 20043 39619 20085 39628
rect 9867 39584 9909 39593
rect 9867 39544 9868 39584
rect 9908 39544 9909 39584
rect 9867 39535 9909 39544
rect 10923 39584 10965 39593
rect 10923 39544 10924 39584
rect 10964 39544 10965 39584
rect 10923 39535 10965 39544
rect 5259 39500 5301 39509
rect 5259 39460 5260 39500
rect 5300 39460 5301 39500
rect 5259 39451 5301 39460
rect 9675 39500 9717 39509
rect 9675 39460 9676 39500
rect 9716 39460 9717 39500
rect 9675 39451 9717 39460
rect 10347 39500 10389 39509
rect 10347 39460 10348 39500
rect 10388 39460 10389 39500
rect 10347 39451 10389 39460
rect 12747 39500 12789 39509
rect 12747 39460 12748 39500
rect 12788 39460 12789 39500
rect 12747 39451 12789 39460
rect 15531 39500 15573 39509
rect 15531 39460 15532 39500
rect 15572 39460 15573 39500
rect 15531 39451 15573 39460
rect 18411 39500 18453 39509
rect 18411 39460 18412 39500
rect 18452 39460 18453 39500
rect 18411 39451 18453 39460
rect 18987 39500 19029 39509
rect 18987 39460 18988 39500
rect 19028 39460 19029 39500
rect 18987 39451 19029 39460
rect 19371 39500 19413 39509
rect 19371 39460 19372 39500
rect 19412 39460 19413 39500
rect 19371 39451 19413 39460
rect 19755 39500 19797 39509
rect 19755 39460 19756 39500
rect 19796 39460 19797 39500
rect 19755 39451 19797 39460
rect 1152 39332 20352 39356
rect 1152 39292 3688 39332
rect 3728 39292 3770 39332
rect 3810 39292 3852 39332
rect 3892 39292 3934 39332
rect 3974 39292 4016 39332
rect 4056 39292 18808 39332
rect 18848 39292 18890 39332
rect 18930 39292 18972 39332
rect 19012 39292 19054 39332
rect 19094 39292 19136 39332
rect 19176 39292 20352 39332
rect 1152 39268 20352 39292
rect 17739 39164 17781 39173
rect 17739 39124 17740 39164
rect 17780 39124 17781 39164
rect 17739 39115 17781 39124
rect 1419 39080 1461 39089
rect 1419 39040 1420 39080
rect 1460 39040 1461 39080
rect 1419 39031 1461 39040
rect 2187 39080 2229 39089
rect 2187 39040 2188 39080
rect 2228 39040 2229 39080
rect 2187 39031 2229 39040
rect 1219 38996 1277 38997
rect 1219 38956 1228 38996
rect 1268 38956 1277 38996
rect 1219 38955 1277 38956
rect 1603 38996 1661 38997
rect 1603 38956 1612 38996
rect 1652 38956 1661 38996
rect 1603 38955 1661 38956
rect 1987 38996 2045 38997
rect 1987 38956 1996 38996
rect 2036 38956 2045 38996
rect 1987 38955 2045 38956
rect 2371 38996 2429 38997
rect 2371 38956 2380 38996
rect 2420 38956 2429 38996
rect 2371 38955 2429 38956
rect 2755 38996 2813 38997
rect 2755 38956 2764 38996
rect 2804 38956 2813 38996
rect 2755 38955 2813 38956
rect 3139 38996 3197 38997
rect 3139 38956 3148 38996
rect 3188 38956 3197 38996
rect 3139 38955 3197 38956
rect 3523 38996 3581 38997
rect 3523 38956 3532 38996
rect 3572 38956 3581 38996
rect 3523 38955 3581 38956
rect 4587 38996 4629 39005
rect 4587 38956 4588 38996
rect 4628 38956 4629 38996
rect 4587 38947 4629 38956
rect 7747 38996 7805 38997
rect 7747 38956 7756 38996
rect 7796 38956 7805 38996
rect 7747 38955 7805 38956
rect 8715 38996 8757 39005
rect 8715 38956 8716 38996
rect 8756 38956 8757 38996
rect 8715 38947 8757 38956
rect 10531 38996 10589 38997
rect 10531 38956 10540 38996
rect 10580 38956 10589 38996
rect 10531 38955 10589 38956
rect 11403 38996 11445 39005
rect 11403 38956 11404 38996
rect 11444 38956 11445 38996
rect 11403 38947 11445 38956
rect 18403 38996 18461 38997
rect 18403 38956 18412 38996
rect 18452 38956 18461 38996
rect 18403 38955 18461 38956
rect 19363 38996 19421 38997
rect 19363 38956 19372 38996
rect 19412 38956 19421 38996
rect 19363 38955 19421 38956
rect 19843 38996 19901 38997
rect 19843 38956 19852 38996
rect 19892 38956 19901 38996
rect 19843 38955 19901 38956
rect 4011 38931 4053 38940
rect 4011 38891 4012 38931
rect 4052 38891 4053 38931
rect 5547 38926 5589 38935
rect 4011 38882 4053 38891
rect 4107 38912 4149 38921
rect 4107 38872 4108 38912
rect 4148 38872 4149 38912
rect 4107 38863 4149 38872
rect 4491 38912 4533 38921
rect 4491 38872 4492 38912
rect 4532 38872 4533 38912
rect 4491 38863 4533 38872
rect 5059 38912 5117 38913
rect 5059 38872 5068 38912
rect 5108 38872 5117 38912
rect 5547 38886 5548 38926
rect 5588 38886 5589 38926
rect 9675 38926 9717 38935
rect 5547 38877 5589 38886
rect 5923 38912 5981 38913
rect 5059 38871 5117 38872
rect 5923 38872 5932 38912
rect 5972 38872 5981 38912
rect 5923 38871 5981 38872
rect 7171 38912 7229 38913
rect 7171 38872 7180 38912
rect 7220 38872 7229 38912
rect 7171 38871 7229 38872
rect 8139 38912 8181 38921
rect 8139 38872 8140 38912
rect 8180 38872 8181 38912
rect 8139 38863 8181 38872
rect 8235 38912 8277 38921
rect 8235 38872 8236 38912
rect 8276 38872 8277 38912
rect 8235 38863 8277 38872
rect 8619 38912 8661 38921
rect 8619 38872 8620 38912
rect 8660 38872 8661 38912
rect 8619 38863 8661 38872
rect 9187 38912 9245 38913
rect 9187 38872 9196 38912
rect 9236 38872 9245 38912
rect 9675 38886 9676 38926
rect 9716 38886 9717 38926
rect 12363 38926 12405 38935
rect 9675 38877 9717 38886
rect 10827 38912 10869 38921
rect 9187 38871 9245 38872
rect 10827 38872 10828 38912
rect 10868 38872 10869 38912
rect 10827 38863 10869 38872
rect 10923 38912 10965 38921
rect 10923 38872 10924 38912
rect 10964 38872 10965 38912
rect 10923 38863 10965 38872
rect 11307 38912 11349 38921
rect 11307 38872 11308 38912
rect 11348 38872 11349 38912
rect 11307 38863 11349 38872
rect 11875 38912 11933 38913
rect 11875 38872 11884 38912
rect 11924 38872 11933 38912
rect 12363 38886 12364 38926
rect 12404 38886 12405 38926
rect 12363 38877 12405 38886
rect 12931 38912 12989 38913
rect 11875 38871 11933 38872
rect 12931 38872 12940 38912
rect 12980 38872 12989 38912
rect 12931 38871 12989 38872
rect 14179 38912 14237 38913
rect 14179 38872 14188 38912
rect 14228 38872 14237 38912
rect 14179 38871 14237 38872
rect 14371 38912 14429 38913
rect 14371 38872 14380 38912
rect 14420 38872 14429 38912
rect 14371 38871 14429 38872
rect 15619 38912 15677 38913
rect 15619 38872 15628 38912
rect 15668 38872 15677 38912
rect 15619 38871 15677 38872
rect 16291 38912 16349 38913
rect 16291 38872 16300 38912
rect 16340 38872 16349 38912
rect 16291 38871 16349 38872
rect 17539 38912 17597 38913
rect 17539 38872 17548 38912
rect 17588 38872 17597 38912
rect 17539 38871 17597 38872
rect 17923 38912 17981 38913
rect 17923 38872 17932 38912
rect 17972 38872 17981 38912
rect 17923 38871 17981 38872
rect 18027 38912 18069 38921
rect 18027 38872 18028 38912
rect 18068 38872 18069 38912
rect 18027 38863 18069 38872
rect 18219 38912 18261 38921
rect 18219 38872 18220 38912
rect 18260 38872 18261 38912
rect 18219 38863 18261 38872
rect 18795 38912 18837 38921
rect 18795 38872 18796 38912
rect 18836 38872 18837 38912
rect 18795 38863 18837 38872
rect 18987 38912 19029 38921
rect 18987 38872 18988 38912
rect 19028 38872 19029 38912
rect 18987 38863 19029 38872
rect 9867 38828 9909 38837
rect 9867 38788 9868 38828
rect 9908 38788 9909 38828
rect 9867 38779 9909 38788
rect 1803 38744 1845 38753
rect 1803 38704 1804 38744
rect 1844 38704 1845 38744
rect 1803 38695 1845 38704
rect 2571 38744 2613 38753
rect 2571 38704 2572 38744
rect 2612 38704 2613 38744
rect 2571 38695 2613 38704
rect 2955 38744 2997 38753
rect 2955 38704 2956 38744
rect 2996 38704 2997 38744
rect 2955 38695 2997 38704
rect 3339 38744 3381 38753
rect 3339 38704 3340 38744
rect 3380 38704 3381 38744
rect 3339 38695 3381 38704
rect 3723 38744 3765 38753
rect 3723 38704 3724 38744
rect 3764 38704 3765 38744
rect 3723 38695 3765 38704
rect 5739 38744 5781 38753
rect 5739 38704 5740 38744
rect 5780 38704 5781 38744
rect 5739 38695 5781 38704
rect 7371 38744 7413 38753
rect 7371 38704 7372 38744
rect 7412 38704 7413 38744
rect 7371 38695 7413 38704
rect 7563 38744 7605 38753
rect 7563 38704 7564 38744
rect 7604 38704 7605 38744
rect 7563 38695 7605 38704
rect 10051 38744 10109 38745
rect 10051 38704 10060 38744
rect 10100 38704 10109 38744
rect 10051 38703 10109 38704
rect 10347 38744 10389 38753
rect 10347 38704 10348 38744
rect 10388 38704 10389 38744
rect 10347 38695 10389 38704
rect 12555 38744 12597 38753
rect 12555 38704 12556 38744
rect 12596 38704 12597 38744
rect 12555 38695 12597 38704
rect 12747 38744 12789 38753
rect 12747 38704 12748 38744
rect 12788 38704 12789 38744
rect 12747 38695 12789 38704
rect 15819 38744 15861 38753
rect 15819 38704 15820 38744
rect 15860 38704 15861 38744
rect 15819 38695 15861 38704
rect 16003 38744 16061 38745
rect 16003 38704 16012 38744
rect 16052 38704 16061 38744
rect 16003 38703 16061 38704
rect 18115 38744 18173 38745
rect 18115 38704 18124 38744
rect 18164 38704 18173 38744
rect 18115 38703 18173 38704
rect 18603 38744 18645 38753
rect 18603 38704 18604 38744
rect 18644 38704 18645 38744
rect 18603 38695 18645 38704
rect 18891 38744 18933 38753
rect 18891 38704 18892 38744
rect 18932 38704 18933 38744
rect 18891 38695 18933 38704
rect 19563 38744 19605 38753
rect 19563 38704 19564 38744
rect 19604 38704 19605 38744
rect 19563 38695 19605 38704
rect 20043 38744 20085 38753
rect 20043 38704 20044 38744
rect 20084 38704 20085 38744
rect 20043 38695 20085 38704
rect 1152 38576 20452 38600
rect 1152 38536 4928 38576
rect 4968 38536 5010 38576
rect 5050 38536 5092 38576
rect 5132 38536 5174 38576
rect 5214 38536 5256 38576
rect 5296 38536 20048 38576
rect 20088 38536 20130 38576
rect 20170 38536 20212 38576
rect 20252 38536 20294 38576
rect 20334 38536 20376 38576
rect 20416 38536 20452 38576
rect 1152 38512 20452 38536
rect 1707 38408 1749 38417
rect 1707 38368 1708 38408
rect 1748 38368 1749 38408
rect 1707 38359 1749 38368
rect 2955 38408 2997 38417
rect 2955 38368 2956 38408
rect 2996 38368 2997 38408
rect 2955 38359 2997 38368
rect 7083 38408 7125 38417
rect 7083 38368 7084 38408
rect 7124 38368 7125 38408
rect 7083 38359 7125 38368
rect 7843 38408 7901 38409
rect 7843 38368 7852 38408
rect 7892 38368 7901 38408
rect 7843 38367 7901 38368
rect 10827 38408 10869 38417
rect 10827 38368 10828 38408
rect 10868 38368 10869 38408
rect 10827 38359 10869 38368
rect 13227 38408 13269 38417
rect 13227 38368 13228 38408
rect 13268 38368 13269 38408
rect 13227 38359 13269 38368
rect 13611 38408 13653 38417
rect 13611 38368 13612 38408
rect 13652 38368 13653 38408
rect 13611 38359 13653 38368
rect 20227 38408 20285 38409
rect 20227 38368 20236 38408
rect 20276 38368 20285 38408
rect 20227 38367 20285 38368
rect 8043 38324 8085 38333
rect 8043 38284 8044 38324
rect 8084 38284 8085 38324
rect 8043 38275 8085 38284
rect 12843 38324 12885 38333
rect 12843 38284 12844 38324
rect 12884 38284 12885 38324
rect 12843 38275 12885 38284
rect 19083 38324 19125 38333
rect 19083 38284 19084 38324
rect 19124 38284 19125 38324
rect 19083 38275 19125 38284
rect 20139 38261 20181 38270
rect 3139 38240 3197 38241
rect 3139 38200 3148 38240
rect 3188 38200 3197 38240
rect 3139 38199 3197 38200
rect 4387 38240 4445 38241
rect 4387 38200 4396 38240
rect 4436 38200 4445 38240
rect 4387 38199 4445 38200
rect 5059 38240 5117 38241
rect 5059 38200 5068 38240
rect 5108 38200 5117 38240
rect 5059 38199 5117 38200
rect 6307 38240 6365 38241
rect 6307 38200 6316 38240
rect 6356 38200 6365 38240
rect 6307 38199 6365 38200
rect 8323 38240 8381 38241
rect 8323 38200 8332 38240
rect 8372 38200 8381 38240
rect 8323 38199 8381 38200
rect 9571 38240 9629 38241
rect 9571 38200 9580 38240
rect 9620 38200 9629 38240
rect 9571 38199 9629 38200
rect 10051 38240 10109 38241
rect 10051 38200 10060 38240
rect 10100 38200 10109 38240
rect 10051 38199 10109 38200
rect 10251 38240 10293 38249
rect 10251 38200 10252 38240
rect 10292 38200 10293 38240
rect 10251 38191 10293 38200
rect 10443 38240 10485 38249
rect 10443 38200 10444 38240
rect 10484 38200 10485 38240
rect 10443 38191 10485 38200
rect 11115 38240 11157 38249
rect 11115 38200 11116 38240
rect 11156 38200 11157 38240
rect 11115 38191 11157 38200
rect 11211 38240 11253 38249
rect 11211 38200 11212 38240
rect 11252 38200 11253 38240
rect 11211 38191 11253 38200
rect 11691 38240 11733 38249
rect 11691 38200 11692 38240
rect 11732 38200 11733 38240
rect 11691 38191 11733 38200
rect 12163 38240 12221 38241
rect 12163 38200 12172 38240
rect 12212 38200 12221 38240
rect 12163 38199 12221 38200
rect 12651 38235 12693 38244
rect 12651 38195 12652 38235
rect 12692 38195 12693 38235
rect 13795 38240 13853 38241
rect 13795 38200 13804 38240
rect 13844 38200 13853 38240
rect 13795 38199 13853 38200
rect 15043 38240 15101 38241
rect 15043 38200 15052 38240
rect 15092 38200 15101 38240
rect 15043 38199 15101 38200
rect 15531 38240 15573 38249
rect 15531 38200 15532 38240
rect 15572 38200 15573 38240
rect 12651 38186 12693 38195
rect 15531 38191 15573 38200
rect 15915 38240 15957 38249
rect 15915 38200 15916 38240
rect 15956 38200 15957 38240
rect 15915 38191 15957 38200
rect 16011 38240 16053 38249
rect 16011 38200 16012 38240
rect 16052 38200 16053 38240
rect 16011 38191 16053 38200
rect 16107 38240 16149 38249
rect 16107 38200 16108 38240
rect 16148 38200 16149 38240
rect 16107 38191 16149 38200
rect 16203 38240 16245 38249
rect 16203 38200 16204 38240
rect 16244 38200 16245 38240
rect 16203 38191 16245 38200
rect 16395 38240 16437 38249
rect 16395 38200 16396 38240
rect 16436 38200 16437 38240
rect 16675 38240 16733 38241
rect 16395 38191 16437 38200
rect 16579 38226 16637 38227
rect 16579 38186 16588 38226
rect 16628 38186 16637 38226
rect 16675 38200 16684 38240
rect 16724 38200 16733 38240
rect 16675 38199 16733 38200
rect 17067 38240 17109 38249
rect 17067 38200 17068 38240
rect 17108 38200 17109 38240
rect 17067 38191 17109 38200
rect 17259 38240 17301 38249
rect 17259 38200 17260 38240
rect 17300 38200 17301 38240
rect 17259 38191 17301 38200
rect 17347 38240 17405 38241
rect 17347 38200 17356 38240
rect 17396 38200 17405 38240
rect 17347 38199 17405 38200
rect 17635 38240 17693 38241
rect 17635 38200 17644 38240
rect 17684 38200 17693 38240
rect 17635 38199 17693 38200
rect 18883 38240 18941 38241
rect 18883 38200 18892 38240
rect 18932 38200 18941 38240
rect 18883 38199 18941 38200
rect 19459 38240 19517 38241
rect 19459 38200 19468 38240
rect 19508 38200 19517 38240
rect 19459 38199 19517 38200
rect 19563 38240 19605 38249
rect 19563 38200 19564 38240
rect 19604 38200 19605 38240
rect 19563 38191 19605 38200
rect 19755 38240 19797 38249
rect 19755 38200 19756 38240
rect 19796 38200 19797 38240
rect 19755 38191 19797 38200
rect 19947 38240 19989 38249
rect 19947 38200 19948 38240
rect 19988 38200 19989 38240
rect 19947 38191 19989 38200
rect 20043 38240 20085 38249
rect 20043 38200 20044 38240
rect 20084 38200 20085 38240
rect 20139 38221 20140 38261
rect 20180 38221 20181 38261
rect 20139 38212 20181 38221
rect 20043 38191 20085 38200
rect 16579 38185 16637 38186
rect 1507 38156 1565 38157
rect 1507 38116 1516 38156
rect 1556 38116 1565 38156
rect 1507 38115 1565 38116
rect 2187 38156 2229 38165
rect 2187 38116 2188 38156
rect 2228 38116 2229 38156
rect 2187 38107 2229 38116
rect 2371 38156 2429 38157
rect 2371 38116 2380 38156
rect 2420 38116 2429 38156
rect 2371 38115 2429 38116
rect 2755 38156 2813 38157
rect 2755 38116 2764 38156
rect 2804 38116 2813 38156
rect 2755 38115 2813 38116
rect 6883 38156 6941 38157
rect 6883 38116 6892 38156
rect 6932 38116 6941 38156
rect 6883 38115 6941 38116
rect 10627 38156 10685 38157
rect 10627 38116 10636 38156
rect 10676 38116 10685 38156
rect 10627 38115 10685 38116
rect 11595 38156 11637 38165
rect 11595 38116 11596 38156
rect 11636 38116 11637 38156
rect 13411 38156 13469 38157
rect 11595 38107 11637 38116
rect 13027 38145 13085 38146
rect 13027 38105 13036 38145
rect 13076 38105 13085 38145
rect 13411 38116 13420 38156
rect 13460 38116 13469 38156
rect 13411 38115 13469 38116
rect 13027 38104 13085 38105
rect 1323 38072 1365 38081
rect 1323 38032 1324 38072
rect 1364 38032 1365 38072
rect 1323 38023 1365 38032
rect 2571 38072 2613 38081
rect 2571 38032 2572 38072
rect 2612 38032 2613 38072
rect 2571 38023 2613 38032
rect 4875 38072 4917 38081
rect 4875 38032 4876 38072
rect 4916 38032 4917 38072
rect 4875 38023 4917 38032
rect 7563 38072 7605 38081
rect 7563 38032 7564 38072
rect 7604 38032 7605 38072
rect 7563 38023 7605 38032
rect 15531 38072 15573 38081
rect 15531 38032 15532 38072
rect 15572 38032 15573 38072
rect 15531 38023 15573 38032
rect 16395 38072 16437 38081
rect 16395 38032 16396 38072
rect 16436 38032 16437 38072
rect 16395 38023 16437 38032
rect 4587 37988 4629 37997
rect 4587 37948 4588 37988
rect 4628 37948 4629 37988
rect 4587 37939 4629 37948
rect 6507 37988 6549 37997
rect 6507 37948 6508 37988
rect 6548 37948 6549 37988
rect 6507 37939 6549 37948
rect 9771 37988 9813 37997
rect 9771 37948 9772 37988
rect 9812 37948 9813 37988
rect 9771 37939 9813 37948
rect 9963 37988 10005 37997
rect 9963 37948 9964 37988
rect 10004 37948 10005 37988
rect 9963 37939 10005 37948
rect 10443 37988 10485 37997
rect 10443 37948 10444 37988
rect 10484 37948 10485 37988
rect 10443 37939 10485 37948
rect 15243 37988 15285 37997
rect 15243 37948 15244 37988
rect 15284 37948 15285 37988
rect 15243 37939 15285 37948
rect 15723 37988 15765 37997
rect 15723 37948 15724 37988
rect 15764 37948 15765 37988
rect 15723 37939 15765 37948
rect 17067 37988 17109 37997
rect 17067 37948 17068 37988
rect 17108 37948 17109 37988
rect 17067 37939 17109 37948
rect 19755 37988 19797 37997
rect 19755 37948 19756 37988
rect 19796 37948 19797 37988
rect 19755 37939 19797 37948
rect 1152 37820 20352 37844
rect 1152 37780 3688 37820
rect 3728 37780 3770 37820
rect 3810 37780 3852 37820
rect 3892 37780 3934 37820
rect 3974 37780 4016 37820
rect 4056 37780 18808 37820
rect 18848 37780 18890 37820
rect 18930 37780 18972 37820
rect 19012 37780 19054 37820
rect 19094 37780 19136 37820
rect 19176 37780 20352 37820
rect 1152 37756 20352 37780
rect 1707 37652 1749 37661
rect 1707 37612 1708 37652
rect 1748 37612 1749 37652
rect 1707 37603 1749 37612
rect 4299 37652 4341 37661
rect 4299 37612 4300 37652
rect 4340 37612 4341 37652
rect 4299 37603 4341 37612
rect 9579 37652 9621 37661
rect 9579 37612 9580 37652
rect 9620 37612 9621 37652
rect 9579 37603 9621 37612
rect 14859 37652 14901 37661
rect 14859 37612 14860 37652
rect 14900 37612 14901 37652
rect 14859 37603 14901 37612
rect 16771 37652 16829 37653
rect 16771 37612 16780 37652
rect 16820 37612 16829 37652
rect 16771 37611 16829 37612
rect 17163 37652 17205 37661
rect 17163 37612 17164 37652
rect 17204 37612 17205 37652
rect 17163 37603 17205 37612
rect 18795 37652 18837 37661
rect 18795 37612 18796 37652
rect 18836 37612 18837 37652
rect 18795 37603 18837 37612
rect 6891 37568 6933 37577
rect 6891 37528 6892 37568
rect 6932 37528 6933 37568
rect 6891 37519 6933 37528
rect 15811 37568 15869 37569
rect 15811 37528 15820 37568
rect 15860 37528 15869 37568
rect 15811 37527 15869 37528
rect 1323 37484 1365 37493
rect 1323 37444 1324 37484
rect 1364 37444 1365 37484
rect 1323 37435 1365 37444
rect 1507 37484 1565 37485
rect 1507 37444 1516 37484
rect 1556 37444 1565 37484
rect 1507 37443 1565 37444
rect 3051 37484 3093 37493
rect 3051 37444 3052 37484
rect 3092 37444 3093 37484
rect 3051 37435 3093 37444
rect 4099 37484 4157 37485
rect 4099 37444 4108 37484
rect 4148 37444 4157 37484
rect 4099 37443 4157 37444
rect 9379 37484 9437 37485
rect 9379 37444 9388 37484
rect 9428 37444 9437 37484
rect 9379 37443 9437 37444
rect 16963 37484 17021 37485
rect 16963 37444 16972 37484
rect 17012 37444 17021 37484
rect 16963 37443 17021 37444
rect 8419 37442 8477 37443
rect 2091 37414 2133 37423
rect 2091 37374 2092 37414
rect 2132 37374 2133 37414
rect 4923 37409 4965 37418
rect 2091 37365 2133 37374
rect 2563 37400 2621 37401
rect 2563 37360 2572 37400
rect 2612 37360 2621 37400
rect 2563 37359 2621 37360
rect 3147 37400 3189 37409
rect 3147 37360 3148 37400
rect 3188 37360 3189 37400
rect 3147 37351 3189 37360
rect 3531 37400 3573 37409
rect 3531 37360 3532 37400
rect 3572 37360 3573 37400
rect 3531 37351 3573 37360
rect 3627 37400 3669 37409
rect 3627 37360 3628 37400
rect 3668 37360 3669 37400
rect 4923 37369 4924 37409
rect 4964 37369 4965 37409
rect 4923 37360 4965 37369
rect 5443 37400 5501 37401
rect 5443 37360 5452 37400
rect 5492 37360 5501 37400
rect 3627 37351 3669 37360
rect 5443 37359 5501 37360
rect 5931 37400 5973 37409
rect 5931 37360 5932 37400
rect 5972 37360 5973 37400
rect 5931 37351 5973 37360
rect 6027 37400 6069 37409
rect 6027 37360 6028 37400
rect 6068 37360 6069 37400
rect 6027 37351 6069 37360
rect 6411 37400 6453 37409
rect 6411 37360 6412 37400
rect 6452 37360 6453 37400
rect 6411 37351 6453 37360
rect 6507 37400 6549 37409
rect 8419 37402 8428 37442
rect 8468 37402 8477 37442
rect 13083 37409 13125 37418
rect 8419 37401 8477 37402
rect 6507 37360 6508 37400
rect 6548 37360 6549 37400
rect 6507 37351 6549 37360
rect 7171 37400 7229 37401
rect 7171 37360 7180 37400
rect 7220 37360 7229 37400
rect 7171 37359 7229 37360
rect 9099 37400 9141 37409
rect 9099 37360 9100 37400
rect 9140 37360 9141 37400
rect 9099 37351 9141 37360
rect 9195 37400 9237 37409
rect 9195 37360 9196 37400
rect 9236 37360 9237 37400
rect 9195 37351 9237 37360
rect 9763 37400 9821 37401
rect 9763 37360 9772 37400
rect 9812 37360 9821 37400
rect 9763 37359 9821 37360
rect 11011 37400 11069 37401
rect 11011 37360 11020 37400
rect 11060 37360 11069 37400
rect 11011 37359 11069 37360
rect 11499 37400 11541 37409
rect 11499 37360 11500 37400
rect 11540 37360 11541 37400
rect 11499 37351 11541 37360
rect 11595 37400 11637 37409
rect 11595 37360 11596 37400
rect 11636 37360 11637 37400
rect 11595 37351 11637 37360
rect 11979 37400 12021 37409
rect 11979 37360 11980 37400
rect 12020 37360 12021 37400
rect 11979 37351 12021 37360
rect 12075 37400 12117 37409
rect 12075 37360 12076 37400
rect 12116 37360 12117 37400
rect 12075 37351 12117 37360
rect 12547 37400 12605 37401
rect 12547 37360 12556 37400
rect 12596 37360 12605 37400
rect 13083 37369 13084 37409
rect 13124 37369 13125 37409
rect 13083 37360 13125 37369
rect 13411 37400 13469 37401
rect 13411 37360 13420 37400
rect 13460 37360 13469 37400
rect 12547 37359 12605 37360
rect 13411 37359 13469 37360
rect 14659 37400 14717 37401
rect 14659 37360 14668 37400
rect 14708 37360 14717 37400
rect 14659 37359 14717 37360
rect 15139 37400 15197 37401
rect 15139 37360 15148 37400
rect 15188 37360 15197 37400
rect 15139 37359 15197 37360
rect 15435 37400 15477 37409
rect 15435 37360 15436 37400
rect 15476 37360 15477 37400
rect 15435 37351 15477 37360
rect 15531 37400 15573 37409
rect 15531 37360 15532 37400
rect 15572 37360 15573 37400
rect 15531 37351 15573 37360
rect 16099 37400 16157 37401
rect 16099 37360 16108 37400
rect 16148 37360 16157 37400
rect 16099 37359 16157 37360
rect 16395 37400 16437 37409
rect 16395 37360 16396 37400
rect 16436 37360 16437 37400
rect 16395 37351 16437 37360
rect 17347 37400 17405 37401
rect 17347 37360 17356 37400
rect 17396 37360 17405 37400
rect 17347 37359 17405 37360
rect 18595 37400 18653 37401
rect 18595 37360 18604 37400
rect 18644 37360 18653 37400
rect 18595 37359 18653 37360
rect 18987 37400 19029 37409
rect 18987 37360 18988 37400
rect 19028 37360 19029 37400
rect 18987 37351 19029 37360
rect 19083 37400 19125 37409
rect 19083 37360 19084 37400
rect 19124 37360 19125 37400
rect 19083 37351 19125 37360
rect 19179 37400 19221 37409
rect 19179 37360 19180 37400
rect 19220 37360 19221 37400
rect 19179 37351 19221 37360
rect 19275 37400 19317 37409
rect 19275 37360 19276 37400
rect 19316 37360 19317 37400
rect 19275 37351 19317 37360
rect 19467 37400 19509 37409
rect 19467 37360 19468 37400
rect 19508 37360 19509 37400
rect 19467 37351 19509 37360
rect 19659 37400 19701 37409
rect 19659 37360 19660 37400
rect 19700 37360 19701 37400
rect 19659 37351 19701 37360
rect 19747 37400 19805 37401
rect 19747 37360 19756 37400
rect 19796 37360 19805 37400
rect 19747 37359 19805 37360
rect 19947 37400 19989 37409
rect 19947 37360 19948 37400
rect 19988 37360 19989 37400
rect 20227 37400 20285 37401
rect 19947 37351 19989 37360
rect 20139 37358 20181 37367
rect 20227 37360 20236 37400
rect 20276 37360 20285 37400
rect 20227 37359 20285 37360
rect 1899 37316 1941 37325
rect 1899 37276 1900 37316
rect 1940 37276 1941 37316
rect 1899 37267 1941 37276
rect 11211 37316 11253 37325
rect 11211 37276 11212 37316
rect 11252 37276 11253 37316
rect 11211 37267 11253 37276
rect 13227 37316 13269 37325
rect 13227 37276 13228 37316
rect 13268 37276 13269 37316
rect 13227 37267 13269 37276
rect 16491 37316 16533 37325
rect 16491 37276 16492 37316
rect 16532 37276 16533 37316
rect 16491 37267 16533 37276
rect 19563 37316 19605 37325
rect 19563 37276 19564 37316
rect 19604 37276 19605 37316
rect 19563 37267 19605 37276
rect 20043 37316 20085 37325
rect 20043 37276 20044 37316
rect 20084 37276 20085 37316
rect 20139 37318 20140 37358
rect 20180 37318 20181 37358
rect 20139 37309 20181 37318
rect 20043 37267 20085 37276
rect 4491 37232 4533 37241
rect 4491 37192 4492 37232
rect 4532 37192 4533 37232
rect 4491 37183 4533 37192
rect 4779 37232 4821 37241
rect 4779 37192 4780 37232
rect 4820 37192 4821 37232
rect 4779 37183 4821 37192
rect 6987 37232 7029 37241
rect 6987 37192 6988 37232
rect 7028 37192 7029 37232
rect 6987 37183 7029 37192
rect 8619 37232 8661 37241
rect 8619 37192 8620 37232
rect 8660 37192 8661 37232
rect 8619 37183 8661 37192
rect 8899 37232 8957 37233
rect 8899 37192 8908 37232
rect 8948 37192 8957 37232
rect 8899 37191 8957 37192
rect 18795 37232 18837 37241
rect 18795 37192 18796 37232
rect 18836 37192 18837 37232
rect 18795 37183 18837 37192
rect 1152 37064 20452 37088
rect 1152 37024 4928 37064
rect 4968 37024 5010 37064
rect 5050 37024 5092 37064
rect 5132 37024 5174 37064
rect 5214 37024 5256 37064
rect 5296 37024 20048 37064
rect 20088 37024 20130 37064
rect 20170 37024 20212 37064
rect 20252 37024 20294 37064
rect 20334 37024 20376 37064
rect 20416 37024 20452 37064
rect 1152 37000 20452 37024
rect 1419 36896 1461 36905
rect 1419 36856 1420 36896
rect 1460 36856 1461 36896
rect 1419 36847 1461 36856
rect 1707 36896 1749 36905
rect 1707 36856 1708 36896
rect 1748 36856 1749 36896
rect 1707 36847 1749 36856
rect 4011 36896 4053 36905
rect 4011 36856 4012 36896
rect 4052 36856 4053 36896
rect 4011 36847 4053 36856
rect 4395 36896 4437 36905
rect 4395 36856 4396 36896
rect 4436 36856 4437 36896
rect 4395 36847 4437 36856
rect 4587 36896 4629 36905
rect 4587 36856 4588 36896
rect 4628 36856 4629 36896
rect 4587 36847 4629 36856
rect 5643 36896 5685 36905
rect 5643 36856 5644 36896
rect 5684 36856 5685 36896
rect 5643 36847 5685 36856
rect 6123 36896 6165 36905
rect 6123 36856 6124 36896
rect 6164 36856 6165 36896
rect 6123 36847 6165 36856
rect 8131 36896 8189 36897
rect 8131 36856 8140 36896
rect 8180 36856 8189 36896
rect 8131 36855 8189 36856
rect 11211 36896 11253 36905
rect 11211 36856 11212 36896
rect 11252 36856 11253 36896
rect 11211 36847 11253 36856
rect 13227 36896 13269 36905
rect 13227 36856 13228 36896
rect 13268 36856 13269 36896
rect 13227 36847 13269 36856
rect 14859 36896 14901 36905
rect 14859 36856 14860 36896
rect 14900 36856 14901 36896
rect 14859 36847 14901 36856
rect 16291 36896 16349 36897
rect 16291 36856 16300 36896
rect 16340 36856 16349 36896
rect 16291 36855 16349 36856
rect 16963 36896 17021 36897
rect 16963 36856 16972 36896
rect 17012 36856 17021 36896
rect 16963 36855 17021 36856
rect 17635 36896 17693 36897
rect 17635 36856 17644 36896
rect 17684 36856 17693 36896
rect 17635 36855 17693 36856
rect 19075 36896 19133 36897
rect 19075 36856 19084 36896
rect 19124 36856 19133 36896
rect 19075 36855 19133 36856
rect 19555 36896 19613 36897
rect 19555 36856 19564 36896
rect 19604 36856 19613 36896
rect 19555 36855 19613 36856
rect 20131 36896 20189 36897
rect 20131 36856 20140 36896
rect 20180 36856 20189 36896
rect 20131 36855 20189 36856
rect 5931 36812 5973 36821
rect 5931 36772 5932 36812
rect 5972 36772 5973 36812
rect 5931 36763 5973 36772
rect 10251 36812 10293 36821
rect 10251 36772 10252 36812
rect 10292 36772 10293 36812
rect 10251 36763 10293 36772
rect 18315 36812 18357 36821
rect 18315 36772 18316 36812
rect 18356 36772 18357 36812
rect 18315 36763 18357 36772
rect 16395 36749 16437 36758
rect 2179 36728 2237 36729
rect 2179 36688 2188 36728
rect 2228 36688 2237 36728
rect 2179 36687 2237 36688
rect 3427 36728 3485 36729
rect 3427 36688 3436 36728
rect 3476 36688 3485 36728
rect 3427 36687 3485 36688
rect 5827 36728 5885 36729
rect 5827 36688 5836 36728
rect 5876 36688 5885 36728
rect 5827 36687 5885 36688
rect 6499 36728 6557 36729
rect 6499 36688 6508 36728
rect 6548 36688 6557 36728
rect 6499 36687 6557 36688
rect 7747 36728 7805 36729
rect 7747 36688 7756 36728
rect 7796 36688 7805 36728
rect 7747 36687 7805 36688
rect 8523 36728 8565 36737
rect 8523 36688 8524 36728
rect 8564 36688 8565 36728
rect 8523 36679 8565 36688
rect 8619 36728 8661 36737
rect 8619 36688 8620 36728
rect 8660 36688 8661 36728
rect 8619 36679 8661 36688
rect 9003 36728 9045 36737
rect 9003 36688 9004 36728
rect 9044 36688 9045 36728
rect 9003 36679 9045 36688
rect 9099 36728 9141 36737
rect 9099 36688 9100 36728
rect 9140 36688 9141 36728
rect 9099 36679 9141 36688
rect 9571 36728 9629 36729
rect 9571 36688 9580 36728
rect 9620 36688 9629 36728
rect 9571 36687 9629 36688
rect 10059 36723 10101 36732
rect 10059 36683 10060 36723
rect 10100 36683 10101 36723
rect 11779 36728 11837 36729
rect 11779 36688 11788 36728
rect 11828 36688 11837 36728
rect 11779 36687 11837 36688
rect 13027 36728 13085 36729
rect 13027 36688 13036 36728
rect 13076 36688 13085 36728
rect 13027 36687 13085 36688
rect 13411 36728 13469 36729
rect 13411 36688 13420 36728
rect 13460 36688 13469 36728
rect 13411 36687 13469 36688
rect 14659 36728 14717 36729
rect 14659 36688 14668 36728
rect 14708 36688 14717 36728
rect 14659 36687 14717 36688
rect 15051 36728 15093 36737
rect 15051 36688 15052 36728
rect 15092 36688 15093 36728
rect 15427 36728 15485 36729
rect 10059 36674 10101 36683
rect 15051 36679 15093 36688
rect 15147 36686 15189 36695
rect 15427 36688 15436 36728
rect 15476 36688 15485 36728
rect 15427 36687 15485 36688
rect 15811 36728 15869 36729
rect 15811 36688 15820 36728
rect 15860 36688 15869 36728
rect 15811 36687 15869 36688
rect 15915 36728 15957 36737
rect 15915 36688 15916 36728
rect 15956 36688 15957 36728
rect 15147 36646 15148 36686
rect 15188 36646 15189 36686
rect 15915 36679 15957 36688
rect 16099 36728 16157 36729
rect 16099 36688 16108 36728
rect 16148 36688 16157 36728
rect 16395 36709 16396 36749
rect 16436 36709 16437 36749
rect 16395 36700 16437 36709
rect 16491 36728 16533 36737
rect 16099 36687 16157 36688
rect 16491 36688 16492 36728
rect 16532 36688 16533 36728
rect 16491 36679 16533 36688
rect 16587 36728 16629 36737
rect 16587 36688 16588 36728
rect 16628 36688 16629 36728
rect 16587 36679 16629 36688
rect 16771 36728 16829 36729
rect 16771 36688 16780 36728
rect 16820 36688 16829 36728
rect 16771 36687 16829 36688
rect 16875 36728 16917 36737
rect 16875 36688 16876 36728
rect 16916 36688 16917 36728
rect 16875 36679 16917 36688
rect 17067 36728 17109 36737
rect 17067 36688 17068 36728
rect 17108 36688 17109 36728
rect 17547 36728 17589 36737
rect 17067 36679 17109 36688
rect 17355 36683 17397 36692
rect 17547 36688 17548 36728
rect 17588 36688 17589 36728
rect 1219 36644 1277 36645
rect 1219 36604 1228 36644
rect 1268 36604 1277 36644
rect 1219 36603 1277 36604
rect 3811 36644 3869 36645
rect 3811 36604 3820 36644
rect 3860 36604 3869 36644
rect 3811 36603 3869 36604
rect 4195 36644 4253 36645
rect 4195 36604 4204 36644
rect 4244 36604 4253 36644
rect 4195 36603 4253 36604
rect 4771 36644 4829 36645
rect 4771 36604 4780 36644
rect 4820 36604 4829 36644
rect 4771 36603 4829 36604
rect 5059 36644 5117 36645
rect 5059 36604 5068 36644
rect 5108 36604 5117 36644
rect 5059 36603 5117 36604
rect 5443 36644 5501 36645
rect 5443 36604 5452 36644
rect 5492 36604 5501 36644
rect 5443 36603 5501 36604
rect 6307 36644 6365 36645
rect 6307 36604 6316 36644
rect 6356 36604 6365 36644
rect 6307 36603 6365 36604
rect 10627 36644 10685 36645
rect 10627 36604 10636 36644
rect 10676 36604 10685 36644
rect 10627 36603 10685 36604
rect 11011 36644 11069 36645
rect 11011 36604 11020 36644
rect 11060 36604 11069 36644
rect 11011 36603 11069 36604
rect 11395 36644 11453 36645
rect 11395 36604 11404 36644
rect 11444 36604 11453 36644
rect 15147 36637 15189 36646
rect 15339 36644 15381 36653
rect 11395 36603 11453 36604
rect 15339 36604 15340 36644
rect 15380 36604 15381 36644
rect 17355 36643 17356 36683
rect 17396 36643 17397 36683
rect 17443 36686 17501 36687
rect 17443 36646 17452 36686
rect 17492 36646 17501 36686
rect 17547 36679 17589 36688
rect 17923 36728 17981 36729
rect 17923 36688 17932 36728
rect 17972 36688 17981 36728
rect 17923 36687 17981 36688
rect 18219 36728 18261 36737
rect 18219 36688 18220 36728
rect 18260 36688 18261 36728
rect 18219 36679 18261 36688
rect 18795 36728 18837 36737
rect 18795 36688 18796 36728
rect 18836 36688 18837 36728
rect 18795 36679 18837 36688
rect 18891 36728 18933 36737
rect 18891 36688 18892 36728
rect 18932 36688 18933 36728
rect 18891 36679 18933 36688
rect 18987 36728 19029 36737
rect 18987 36688 18988 36728
rect 19028 36688 19029 36728
rect 18987 36679 19029 36688
rect 19275 36728 19317 36737
rect 19275 36688 19276 36728
rect 19316 36688 19317 36728
rect 19275 36679 19317 36688
rect 19371 36728 19413 36737
rect 19371 36688 19372 36728
rect 19412 36688 19413 36728
rect 19371 36679 19413 36688
rect 19467 36728 19509 36737
rect 19467 36688 19468 36728
rect 19508 36688 19509 36728
rect 19467 36679 19509 36688
rect 19939 36728 19997 36729
rect 19939 36688 19948 36728
rect 19988 36688 19997 36728
rect 19939 36687 19997 36688
rect 20043 36728 20085 36737
rect 20043 36688 20044 36728
rect 20084 36688 20085 36728
rect 20043 36679 20085 36688
rect 20235 36728 20277 36737
rect 20235 36688 20236 36728
rect 20276 36688 20277 36728
rect 20235 36679 20277 36688
rect 17443 36645 17501 36646
rect 17355 36634 17397 36643
rect 15339 36595 15381 36604
rect 1611 36560 1653 36569
rect 1611 36520 1612 36560
rect 1652 36520 1653 36560
rect 1611 36511 1653 36520
rect 1899 36560 1941 36569
rect 1899 36520 1900 36560
rect 1940 36520 1941 36560
rect 1899 36511 1941 36520
rect 5259 36560 5301 36569
rect 5259 36520 5260 36560
rect 5300 36520 5301 36560
rect 5259 36511 5301 36520
rect 7947 36560 7989 36569
rect 7947 36520 7948 36560
rect 7988 36520 7989 36560
rect 7947 36511 7989 36520
rect 10827 36560 10869 36569
rect 10827 36520 10828 36560
rect 10868 36520 10869 36560
rect 10827 36511 10869 36520
rect 15243 36560 15285 36569
rect 15243 36520 15244 36560
rect 15284 36520 15285 36560
rect 15243 36511 15285 36520
rect 18595 36560 18653 36561
rect 18595 36520 18604 36560
rect 18644 36520 18653 36560
rect 18595 36519 18653 36520
rect 3627 36476 3669 36485
rect 3627 36436 3628 36476
rect 3668 36436 3669 36476
rect 3627 36427 3669 36436
rect 11595 36476 11637 36485
rect 11595 36436 11596 36476
rect 11636 36436 11637 36476
rect 11595 36427 11637 36436
rect 16107 36476 16149 36485
rect 16107 36436 16108 36476
rect 16148 36436 16149 36476
rect 16107 36427 16149 36436
rect 1152 36308 20352 36332
rect 1152 36268 3688 36308
rect 3728 36268 3770 36308
rect 3810 36268 3852 36308
rect 3892 36268 3934 36308
rect 3974 36268 4016 36308
rect 4056 36268 18808 36308
rect 18848 36268 18890 36308
rect 18930 36268 18972 36308
rect 19012 36268 19054 36308
rect 19094 36268 19136 36308
rect 19176 36268 20352 36308
rect 1152 36244 20352 36268
rect 1707 36140 1749 36149
rect 1707 36100 1708 36140
rect 1748 36100 1749 36140
rect 1707 36091 1749 36100
rect 4011 36140 4053 36149
rect 4011 36100 4012 36140
rect 4052 36100 4053 36140
rect 4011 36091 4053 36100
rect 14763 36140 14805 36149
rect 14763 36100 14764 36140
rect 14804 36100 14805 36140
rect 14763 36091 14805 36100
rect 18027 36140 18069 36149
rect 18027 36100 18028 36140
rect 18068 36100 18069 36140
rect 18027 36091 18069 36100
rect 19947 36140 19989 36149
rect 19947 36100 19948 36140
rect 19988 36100 19989 36140
rect 19947 36091 19989 36100
rect 9387 36056 9429 36065
rect 9387 36016 9388 36056
rect 9428 36016 9429 36056
rect 9387 36007 9429 36016
rect 20139 36056 20181 36065
rect 20139 36016 20140 36056
rect 20180 36016 20181 36056
rect 20139 36007 20181 36016
rect 1507 35972 1565 35973
rect 1507 35932 1516 35972
rect 1556 35932 1565 35972
rect 1507 35931 1565 35932
rect 3811 35972 3869 35973
rect 3811 35932 3820 35972
rect 3860 35932 3869 35972
rect 3811 35931 3869 35932
rect 4875 35972 4917 35981
rect 4875 35932 4876 35972
rect 4916 35932 4917 35972
rect 4875 35923 4917 35932
rect 7755 35972 7797 35981
rect 7755 35932 7756 35972
rect 7796 35932 7797 35972
rect 7755 35923 7797 35932
rect 9291 35972 9333 35981
rect 9291 35932 9292 35972
rect 9332 35932 9333 35972
rect 9291 35923 9333 35932
rect 9483 35972 9525 35981
rect 9483 35932 9484 35972
rect 9524 35932 9525 35972
rect 9483 35923 9525 35932
rect 5835 35902 5877 35911
rect 2371 35888 2429 35889
rect 2371 35848 2380 35888
rect 2420 35848 2429 35888
rect 2371 35847 2429 35848
rect 3619 35888 3677 35889
rect 3619 35848 3628 35888
rect 3668 35848 3677 35888
rect 3619 35847 3677 35848
rect 4299 35888 4341 35897
rect 4299 35848 4300 35888
rect 4340 35848 4341 35888
rect 4299 35839 4341 35848
rect 4395 35888 4437 35897
rect 4395 35848 4396 35888
rect 4436 35848 4437 35888
rect 4395 35839 4437 35848
rect 4779 35888 4821 35897
rect 4779 35848 4780 35888
rect 4820 35848 4821 35888
rect 4779 35839 4821 35848
rect 5347 35888 5405 35889
rect 5347 35848 5356 35888
rect 5396 35848 5405 35888
rect 5835 35862 5836 35902
rect 5876 35862 5877 35902
rect 8811 35902 8853 35911
rect 5835 35853 5877 35862
rect 6219 35888 6261 35897
rect 5347 35847 5405 35848
rect 6219 35848 6220 35888
rect 6260 35848 6261 35888
rect 6219 35839 6261 35848
rect 6411 35888 6453 35897
rect 6411 35848 6412 35888
rect 6452 35848 6453 35888
rect 6411 35839 6453 35848
rect 6499 35888 6557 35889
rect 6499 35848 6508 35888
rect 6548 35848 6557 35888
rect 6499 35847 6557 35848
rect 6699 35888 6741 35897
rect 6699 35848 6700 35888
rect 6740 35848 6741 35888
rect 6699 35839 6741 35848
rect 6795 35888 6837 35897
rect 6795 35848 6796 35888
rect 6836 35848 6837 35888
rect 6795 35839 6837 35848
rect 6891 35888 6933 35897
rect 6891 35848 6892 35888
rect 6932 35848 6933 35888
rect 6891 35839 6933 35848
rect 7275 35888 7317 35897
rect 7275 35848 7276 35888
rect 7316 35848 7317 35888
rect 7275 35839 7317 35848
rect 7371 35888 7413 35897
rect 7371 35848 7372 35888
rect 7412 35848 7413 35888
rect 7371 35839 7413 35848
rect 7851 35888 7893 35897
rect 7851 35848 7852 35888
rect 7892 35848 7893 35888
rect 7851 35839 7893 35848
rect 8323 35888 8381 35889
rect 8323 35848 8332 35888
rect 8372 35848 8381 35888
rect 8811 35862 8812 35902
rect 8852 35862 8853 35902
rect 8811 35853 8853 35862
rect 9187 35888 9245 35889
rect 8323 35847 8381 35848
rect 9187 35848 9196 35888
rect 9236 35848 9245 35888
rect 9187 35847 9245 35848
rect 9579 35888 9621 35897
rect 9579 35848 9580 35888
rect 9620 35848 9621 35888
rect 9579 35839 9621 35848
rect 9955 35888 10013 35889
rect 9955 35848 9964 35888
rect 10004 35848 10013 35888
rect 9955 35847 10013 35848
rect 11203 35888 11261 35889
rect 11203 35848 11212 35888
rect 11252 35848 11261 35888
rect 11203 35847 11261 35848
rect 11587 35888 11645 35889
rect 11587 35848 11596 35888
rect 11636 35848 11645 35888
rect 11587 35847 11645 35848
rect 12835 35888 12893 35889
rect 12835 35848 12844 35888
rect 12884 35848 12893 35888
rect 12835 35847 12893 35848
rect 13315 35888 13373 35889
rect 13315 35848 13324 35888
rect 13364 35848 13373 35888
rect 13315 35847 13373 35848
rect 14563 35888 14621 35889
rect 14563 35848 14572 35888
rect 14612 35848 14621 35888
rect 14563 35847 14621 35848
rect 14947 35888 15005 35889
rect 14947 35848 14956 35888
rect 14996 35848 15005 35888
rect 14947 35847 15005 35848
rect 16195 35888 16253 35889
rect 16195 35848 16204 35888
rect 16244 35848 16253 35888
rect 16195 35847 16253 35848
rect 16579 35888 16637 35889
rect 16579 35848 16588 35888
rect 16628 35848 16637 35888
rect 16579 35847 16637 35848
rect 17827 35888 17885 35889
rect 17827 35848 17836 35888
rect 17876 35848 17885 35888
rect 17827 35847 17885 35848
rect 18211 35888 18269 35889
rect 18211 35848 18220 35888
rect 18260 35848 18269 35888
rect 18211 35847 18269 35848
rect 19171 35888 19229 35889
rect 19171 35848 19180 35888
rect 19220 35848 19229 35888
rect 19171 35847 19229 35848
rect 19459 35888 19517 35889
rect 19459 35848 19468 35888
rect 19508 35848 19517 35888
rect 19459 35847 19517 35848
rect 19659 35888 19701 35897
rect 19659 35848 19660 35888
rect 19700 35848 19701 35888
rect 19659 35839 19701 35848
rect 19747 35888 19805 35889
rect 19747 35848 19756 35888
rect 19796 35848 19805 35888
rect 19747 35847 19805 35848
rect 20139 35880 20181 35889
rect 20139 35840 20140 35880
rect 20180 35840 20181 35880
rect 20139 35831 20181 35840
rect 9003 35804 9045 35813
rect 9003 35764 9004 35804
rect 9044 35764 9045 35804
rect 9003 35755 9045 35764
rect 1315 35720 1373 35721
rect 1315 35680 1324 35720
rect 1364 35680 1373 35720
rect 1315 35679 1373 35680
rect 1891 35720 1949 35721
rect 1891 35680 1900 35720
rect 1940 35680 1949 35720
rect 1891 35679 1949 35680
rect 2187 35720 2229 35729
rect 2187 35680 2188 35720
rect 2228 35680 2229 35720
rect 2187 35671 2229 35680
rect 6027 35720 6069 35729
rect 6027 35680 6028 35720
rect 6068 35680 6069 35720
rect 6027 35671 6069 35680
rect 6307 35720 6365 35721
rect 6307 35680 6316 35720
rect 6356 35680 6365 35720
rect 6307 35679 6365 35680
rect 6979 35720 7037 35721
rect 6979 35680 6988 35720
rect 7028 35680 7037 35720
rect 6979 35679 7037 35680
rect 11403 35720 11445 35729
rect 11403 35680 11404 35720
rect 11444 35680 11445 35720
rect 11403 35671 11445 35680
rect 13035 35720 13077 35729
rect 13035 35680 13036 35720
rect 13076 35680 13077 35720
rect 13035 35671 13077 35680
rect 14763 35720 14805 35729
rect 14763 35680 14764 35720
rect 14804 35680 14805 35720
rect 14763 35671 14805 35680
rect 16395 35720 16437 35729
rect 16395 35680 16396 35720
rect 16436 35680 16437 35720
rect 16395 35671 16437 35680
rect 18027 35720 18069 35729
rect 18027 35680 18028 35720
rect 18068 35680 18069 35720
rect 18027 35671 18069 35680
rect 19467 35720 19509 35729
rect 19467 35680 19468 35720
rect 19508 35680 19509 35720
rect 19467 35671 19509 35680
rect 1152 35552 20452 35576
rect 1152 35512 4928 35552
rect 4968 35512 5010 35552
rect 5050 35512 5092 35552
rect 5132 35512 5174 35552
rect 5214 35512 5256 35552
rect 5296 35512 20048 35552
rect 20088 35512 20130 35552
rect 20170 35512 20212 35552
rect 20252 35512 20294 35552
rect 20334 35512 20376 35552
rect 20416 35512 20452 35552
rect 1152 35488 20452 35512
rect 13227 35426 13269 35435
rect 13227 35386 13228 35426
rect 13268 35386 13269 35426
rect 13227 35377 13269 35386
rect 17059 35384 17117 35385
rect 17059 35344 17068 35384
rect 17108 35344 17117 35384
rect 17059 35343 17117 35344
rect 3051 35300 3093 35309
rect 3051 35260 3052 35300
rect 3092 35260 3093 35300
rect 3051 35251 3093 35260
rect 4587 35300 4629 35309
rect 4587 35260 4588 35300
rect 4628 35260 4629 35300
rect 4587 35251 4629 35260
rect 9771 35300 9813 35309
rect 9771 35260 9772 35300
rect 9812 35260 9813 35300
rect 9771 35251 9813 35260
rect 17835 35258 17877 35267
rect 1323 35216 1365 35225
rect 1323 35176 1324 35216
rect 1364 35176 1365 35216
rect 1323 35167 1365 35176
rect 1419 35216 1461 35225
rect 1419 35176 1420 35216
rect 1460 35176 1461 35216
rect 1419 35167 1461 35176
rect 1899 35216 1941 35225
rect 1899 35176 1900 35216
rect 1940 35176 1941 35216
rect 4011 35216 4053 35225
rect 1899 35167 1941 35176
rect 2366 35189 2408 35198
rect 2366 35149 2367 35189
rect 2407 35149 2408 35189
rect 1803 35132 1845 35141
rect 2366 35140 2408 35149
rect 2907 35174 2949 35183
rect 1803 35092 1804 35132
rect 1844 35092 1845 35132
rect 2907 35134 2908 35174
rect 2948 35134 2949 35174
rect 4011 35176 4012 35216
rect 4052 35176 4053 35216
rect 4011 35167 4053 35176
rect 4203 35216 4245 35225
rect 4203 35176 4204 35216
rect 4244 35176 4245 35216
rect 4203 35167 4245 35176
rect 4387 35216 4445 35217
rect 4387 35176 4396 35216
rect 4436 35176 4445 35216
rect 4387 35175 4445 35176
rect 4491 35216 4533 35225
rect 4491 35176 4492 35216
rect 4532 35176 4533 35216
rect 4491 35167 4533 35176
rect 4683 35216 4725 35225
rect 4683 35176 4684 35216
rect 4724 35176 4725 35216
rect 4683 35167 4725 35176
rect 4867 35216 4925 35217
rect 4867 35176 4876 35216
rect 4916 35176 4925 35216
rect 4867 35175 4925 35176
rect 6115 35216 6173 35217
rect 6115 35176 6124 35216
rect 6164 35176 6173 35216
rect 6115 35175 6173 35176
rect 6499 35216 6557 35217
rect 6499 35176 6508 35216
rect 6548 35176 6557 35216
rect 6499 35175 6557 35176
rect 7747 35216 7805 35217
rect 7747 35176 7756 35216
rect 7796 35176 7805 35216
rect 7747 35175 7805 35176
rect 8323 35216 8381 35217
rect 8323 35176 8332 35216
rect 8372 35176 8381 35216
rect 8323 35175 8381 35176
rect 9571 35216 9629 35217
rect 9571 35176 9580 35216
rect 9620 35176 9629 35216
rect 9571 35175 9629 35176
rect 11203 35216 11261 35217
rect 11203 35176 11212 35216
rect 11252 35176 11261 35216
rect 11203 35175 11261 35176
rect 11499 35216 11541 35225
rect 11499 35176 11500 35216
rect 11540 35176 11541 35216
rect 9955 35174 10013 35175
rect 2907 35125 2949 35134
rect 9955 35134 9964 35174
rect 10004 35134 10013 35174
rect 11499 35167 11541 35176
rect 11595 35216 11637 35225
rect 11595 35176 11596 35216
rect 11636 35176 11637 35216
rect 11595 35167 11637 35176
rect 12547 35216 12605 35217
rect 12547 35176 12556 35216
rect 12596 35176 12605 35216
rect 12547 35175 12605 35176
rect 13035 35211 13077 35220
rect 13035 35171 13036 35211
rect 13076 35171 13077 35211
rect 15043 35216 15101 35217
rect 15043 35176 15052 35216
rect 15092 35176 15101 35216
rect 15043 35175 15101 35176
rect 15339 35216 15381 35225
rect 15339 35176 15340 35216
rect 15380 35176 15381 35216
rect 13035 35162 13077 35171
rect 15339 35167 15381 35176
rect 15435 35216 15477 35225
rect 15435 35176 15436 35216
rect 15476 35176 15477 35216
rect 15435 35167 15477 35176
rect 16203 35216 16245 35225
rect 16203 35176 16204 35216
rect 16244 35176 16245 35216
rect 16203 35167 16245 35176
rect 16299 35216 16341 35225
rect 16299 35176 16300 35216
rect 16340 35176 16341 35216
rect 16299 35167 16341 35176
rect 16579 35216 16637 35217
rect 16579 35176 16588 35216
rect 16628 35176 16637 35216
rect 17067 35216 17109 35225
rect 16579 35175 16637 35176
rect 16909 35201 16951 35210
rect 16909 35161 16910 35201
rect 16950 35161 16951 35201
rect 17067 35176 17068 35216
rect 17108 35176 17109 35216
rect 17067 35167 17109 35176
rect 17163 35216 17205 35225
rect 17163 35176 17164 35216
rect 17204 35176 17205 35216
rect 17163 35167 17205 35176
rect 17347 35216 17405 35217
rect 17347 35176 17356 35216
rect 17396 35176 17405 35216
rect 17347 35175 17405 35176
rect 17443 35216 17501 35217
rect 17443 35176 17452 35216
rect 17492 35176 17501 35216
rect 17443 35175 17501 35176
rect 17643 35216 17685 35225
rect 17643 35176 17644 35216
rect 17684 35176 17685 35216
rect 17835 35218 17836 35258
rect 17876 35218 17877 35258
rect 17835 35209 17877 35218
rect 18019 35216 18077 35217
rect 17643 35167 17685 35176
rect 17739 35174 17781 35183
rect 18019 35176 18028 35216
rect 18068 35176 18077 35216
rect 18019 35175 18077 35176
rect 18211 35216 18269 35217
rect 18211 35176 18220 35216
rect 18260 35176 18269 35216
rect 18211 35175 18269 35176
rect 18499 35216 18557 35217
rect 18499 35176 18508 35216
rect 18548 35176 18557 35216
rect 18499 35175 18557 35176
rect 19747 35216 19805 35217
rect 19747 35176 19756 35216
rect 19796 35176 19805 35216
rect 19747 35175 19805 35176
rect 16909 35152 16951 35161
rect 13411 35145 13469 35146
rect 9955 35133 10013 35134
rect 3715 35132 3773 35133
rect 1803 35083 1845 35092
rect 3715 35092 3724 35132
rect 3764 35092 3773 35132
rect 3715 35091 3773 35092
rect 11979 35132 12021 35141
rect 11979 35092 11980 35132
rect 12020 35092 12021 35132
rect 11979 35083 12021 35092
rect 12075 35132 12117 35141
rect 12075 35092 12076 35132
rect 12116 35092 12117 35132
rect 13411 35105 13420 35145
rect 13460 35105 13469 35145
rect 17739 35134 17740 35174
rect 17780 35134 17781 35174
rect 13411 35104 13469 35105
rect 13795 35132 13853 35133
rect 12075 35083 12117 35092
rect 13795 35092 13804 35132
rect 13844 35092 13853 35132
rect 13795 35091 13853 35092
rect 14179 35132 14237 35133
rect 14179 35092 14188 35132
rect 14228 35092 14237 35132
rect 14179 35091 14237 35092
rect 14563 35132 14621 35133
rect 14563 35092 14572 35132
rect 14612 35092 14621 35132
rect 17739 35125 17781 35134
rect 17931 35132 17973 35141
rect 14563 35091 14621 35092
rect 17931 35092 17932 35132
rect 17972 35092 17973 35132
rect 17931 35083 17973 35092
rect 3243 35048 3285 35057
rect 3243 35008 3244 35048
rect 3284 35008 3285 35048
rect 3243 34999 3285 35008
rect 7947 35048 7989 35057
rect 7947 35008 7948 35048
rect 7988 35008 7989 35048
rect 7947 34999 7989 35008
rect 8139 35048 8181 35057
rect 8139 35008 8140 35048
rect 8180 35008 8181 35048
rect 8139 34999 8181 35008
rect 13995 35048 14037 35057
rect 13995 35008 13996 35048
rect 14036 35008 14037 35048
rect 13995 34999 14037 35008
rect 14379 35048 14421 35057
rect 14379 35008 14380 35048
rect 14420 35008 14421 35048
rect 14379 34999 14421 35008
rect 15715 35048 15773 35049
rect 15715 35008 15724 35048
rect 15764 35008 15773 35048
rect 15715 35007 15773 35008
rect 15907 35048 15965 35049
rect 15907 35008 15916 35048
rect 15956 35008 15965 35048
rect 15907 35007 15965 35008
rect 20235 35048 20277 35057
rect 20235 35008 20236 35048
rect 20276 35008 20277 35048
rect 20235 34999 20277 35008
rect 3531 34964 3573 34973
rect 3531 34924 3532 34964
rect 3572 34924 3573 34964
rect 3531 34915 3573 34924
rect 4011 34964 4053 34973
rect 4011 34924 4012 34964
rect 4052 34924 4053 34964
rect 4011 34915 4053 34924
rect 6315 34964 6357 34973
rect 6315 34924 6316 34964
rect 6356 34924 6357 34964
rect 6315 34915 6357 34924
rect 13611 34964 13653 34973
rect 13611 34924 13612 34964
rect 13652 34924 13653 34964
rect 13611 34915 13653 34924
rect 14763 34964 14805 34973
rect 14763 34924 14764 34964
rect 14804 34924 14805 34964
rect 14763 34915 14805 34924
rect 18315 34964 18357 34973
rect 18315 34924 18316 34964
rect 18356 34924 18357 34964
rect 18315 34915 18357 34924
rect 19947 34964 19989 34973
rect 19947 34924 19948 34964
rect 19988 34924 19989 34964
rect 19947 34915 19989 34924
rect 1152 34796 20352 34820
rect 1152 34756 3688 34796
rect 3728 34756 3770 34796
rect 3810 34756 3852 34796
rect 3892 34756 3934 34796
rect 3974 34756 4016 34796
rect 4056 34756 18808 34796
rect 18848 34756 18890 34796
rect 18930 34756 18972 34796
rect 19012 34756 19054 34796
rect 19094 34756 19136 34796
rect 19176 34756 20352 34796
rect 1152 34732 20352 34756
rect 1611 34628 1653 34637
rect 1611 34588 1612 34628
rect 1652 34588 1653 34628
rect 1611 34579 1653 34588
rect 1995 34628 2037 34637
rect 1995 34588 1996 34628
rect 2036 34588 2037 34628
rect 1995 34579 2037 34588
rect 5643 34628 5685 34637
rect 5643 34588 5644 34628
rect 5684 34588 5685 34628
rect 5643 34579 5685 34588
rect 13035 34628 13077 34637
rect 13035 34588 13036 34628
rect 13076 34588 13077 34628
rect 13035 34579 13077 34588
rect 17643 34628 17685 34637
rect 17643 34588 17644 34628
rect 17684 34588 17685 34628
rect 17643 34579 17685 34588
rect 8811 34544 8853 34553
rect 8811 34504 8812 34544
rect 8852 34504 8853 34544
rect 8811 34495 8853 34504
rect 13803 34544 13845 34553
rect 13803 34504 13804 34544
rect 13844 34504 13845 34544
rect 13803 34495 13845 34504
rect 18691 34544 18749 34545
rect 18691 34504 18700 34544
rect 18740 34504 18749 34544
rect 18691 34503 18749 34504
rect 19851 34544 19893 34553
rect 19851 34504 19852 34544
rect 19892 34504 19893 34544
rect 19851 34495 19893 34504
rect 1411 34460 1469 34461
rect 1411 34420 1420 34460
rect 1460 34420 1469 34460
rect 1411 34419 1469 34420
rect 1795 34460 1853 34461
rect 1795 34420 1804 34460
rect 1844 34420 1853 34460
rect 1795 34419 1853 34420
rect 8715 34460 8757 34469
rect 8715 34420 8716 34460
rect 8756 34420 8757 34460
rect 8715 34411 8757 34420
rect 8907 34460 8949 34469
rect 8907 34420 8908 34460
rect 8948 34420 8949 34460
rect 8907 34411 8949 34420
rect 12451 34460 12509 34461
rect 12451 34420 12460 34460
rect 12500 34420 12509 34460
rect 12451 34419 12509 34420
rect 12835 34460 12893 34461
rect 12835 34420 12844 34460
rect 12884 34420 12893 34460
rect 12835 34419 12893 34420
rect 13411 34460 13469 34461
rect 13411 34420 13420 34460
rect 13460 34420 13469 34460
rect 13411 34419 13469 34420
rect 19755 34460 19797 34469
rect 19755 34420 19756 34460
rect 19796 34420 19797 34460
rect 19755 34411 19797 34420
rect 19947 34460 19989 34469
rect 19947 34420 19948 34460
rect 19988 34420 19989 34460
rect 19947 34411 19989 34420
rect 2379 34381 2421 34390
rect 2379 34341 2380 34381
rect 2420 34341 2421 34381
rect 2379 34332 2421 34341
rect 2851 34376 2909 34377
rect 2851 34336 2860 34376
rect 2900 34336 2909 34376
rect 2851 34335 2909 34336
rect 3339 34376 3381 34385
rect 3339 34336 3340 34376
rect 3380 34336 3381 34376
rect 3339 34327 3381 34336
rect 3435 34376 3477 34385
rect 3435 34336 3436 34376
rect 3476 34336 3477 34376
rect 3435 34327 3477 34336
rect 3819 34376 3861 34385
rect 3819 34336 3820 34376
rect 3860 34336 3861 34376
rect 3819 34327 3861 34336
rect 3915 34376 3957 34385
rect 6219 34381 6261 34390
rect 3915 34336 3916 34376
rect 3956 34336 3957 34376
rect 3915 34327 3957 34336
rect 4195 34376 4253 34377
rect 4195 34336 4204 34376
rect 4244 34336 4253 34376
rect 4195 34335 4253 34336
rect 5443 34376 5501 34377
rect 5443 34336 5452 34376
rect 5492 34336 5501 34376
rect 5443 34335 5501 34336
rect 6219 34341 6220 34381
rect 6260 34341 6261 34381
rect 6219 34332 6261 34341
rect 6691 34376 6749 34377
rect 6691 34336 6700 34376
rect 6740 34336 6749 34376
rect 6691 34335 6749 34336
rect 7179 34376 7221 34385
rect 7179 34336 7180 34376
rect 7220 34336 7221 34376
rect 7179 34327 7221 34336
rect 7275 34376 7317 34385
rect 7275 34336 7276 34376
rect 7316 34336 7317 34376
rect 7275 34327 7317 34336
rect 7659 34376 7701 34385
rect 7659 34336 7660 34376
rect 7700 34336 7701 34376
rect 7659 34327 7701 34336
rect 7755 34376 7797 34385
rect 7755 34336 7756 34376
rect 7796 34336 7797 34376
rect 7755 34327 7797 34336
rect 8139 34376 8181 34385
rect 8139 34336 8140 34376
rect 8180 34336 8181 34376
rect 8139 34327 8181 34336
rect 8235 34376 8277 34385
rect 8235 34336 8236 34376
rect 8276 34336 8277 34376
rect 8235 34327 8277 34336
rect 8331 34376 8373 34385
rect 8331 34336 8332 34376
rect 8372 34336 8373 34376
rect 8331 34327 8373 34336
rect 8611 34376 8669 34377
rect 8611 34336 8620 34376
rect 8660 34336 8669 34376
rect 8611 34335 8669 34336
rect 9003 34376 9045 34385
rect 9003 34336 9004 34376
rect 9044 34336 9045 34376
rect 9003 34327 9045 34336
rect 9187 34376 9245 34377
rect 9187 34336 9196 34376
rect 9236 34336 9245 34376
rect 9187 34335 9245 34336
rect 10435 34376 10493 34377
rect 10435 34336 10444 34376
rect 10484 34336 10493 34376
rect 10435 34335 10493 34336
rect 10819 34376 10877 34377
rect 10819 34336 10828 34376
rect 10868 34336 10877 34376
rect 10819 34335 10877 34336
rect 12067 34376 12125 34377
rect 12067 34336 12076 34376
rect 12116 34336 12125 34376
rect 12067 34335 12125 34336
rect 14659 34376 14717 34377
rect 14659 34336 14668 34376
rect 14708 34336 14717 34376
rect 14659 34335 14717 34336
rect 15907 34376 15965 34377
rect 15907 34336 15916 34376
rect 15956 34336 15965 34376
rect 15907 34335 15965 34336
rect 16195 34376 16253 34377
rect 16195 34336 16204 34376
rect 16244 34336 16253 34376
rect 16195 34335 16253 34336
rect 17443 34376 17501 34377
rect 17443 34336 17452 34376
rect 17492 34336 17501 34376
rect 17443 34335 17501 34336
rect 18019 34376 18077 34377
rect 18019 34336 18028 34376
rect 18068 34336 18077 34376
rect 18019 34335 18077 34336
rect 18315 34376 18357 34385
rect 18315 34336 18316 34376
rect 18356 34336 18357 34376
rect 18315 34327 18357 34336
rect 18974 34376 19032 34377
rect 18974 34336 18983 34376
rect 19023 34336 19032 34376
rect 18974 34335 19032 34336
rect 19083 34376 19125 34385
rect 19083 34336 19084 34376
rect 19124 34336 19125 34376
rect 19083 34327 19125 34336
rect 19179 34376 19221 34385
rect 19179 34336 19180 34376
rect 19220 34336 19221 34376
rect 19179 34327 19221 34336
rect 19363 34376 19421 34377
rect 19363 34336 19372 34376
rect 19412 34336 19421 34376
rect 19363 34335 19421 34336
rect 19459 34376 19517 34377
rect 19459 34336 19468 34376
rect 19508 34336 19517 34376
rect 19459 34335 19517 34336
rect 19659 34376 19701 34385
rect 19659 34336 19660 34376
rect 19700 34336 19701 34376
rect 19659 34327 19701 34336
rect 20035 34376 20093 34377
rect 20035 34336 20044 34376
rect 20084 34336 20093 34376
rect 20035 34335 20093 34336
rect 2187 34292 2229 34301
rect 2187 34252 2188 34292
rect 2228 34252 2229 34292
rect 2187 34243 2229 34252
rect 6027 34292 6069 34301
rect 6027 34252 6028 34292
rect 6068 34252 6069 34292
rect 6027 34243 6069 34252
rect 18411 34292 18453 34301
rect 18411 34252 18412 34292
rect 18452 34252 18453 34292
rect 18411 34243 18453 34252
rect 8419 34208 8477 34209
rect 8419 34168 8428 34208
rect 8468 34168 8477 34208
rect 8419 34167 8477 34168
rect 10635 34208 10677 34217
rect 10635 34168 10636 34208
rect 10676 34168 10677 34208
rect 10635 34159 10677 34168
rect 12267 34208 12309 34217
rect 12267 34168 12268 34208
rect 12308 34168 12309 34208
rect 12267 34159 12309 34168
rect 12651 34208 12693 34217
rect 12651 34168 12652 34208
rect 12692 34168 12693 34208
rect 12651 34159 12693 34168
rect 13611 34208 13653 34217
rect 13611 34168 13612 34208
rect 13652 34168 13653 34208
rect 13611 34159 13653 34168
rect 13899 34208 13941 34217
rect 13899 34168 13900 34208
rect 13940 34168 13941 34208
rect 13899 34159 13941 34168
rect 14179 34208 14237 34209
rect 14179 34168 14188 34208
rect 14228 34168 14237 34208
rect 14179 34167 14237 34168
rect 14475 34208 14517 34217
rect 14475 34168 14476 34208
rect 14516 34168 14517 34208
rect 14475 34159 14517 34168
rect 19267 34208 19325 34209
rect 19267 34168 19276 34208
rect 19316 34168 19325 34208
rect 19267 34167 19325 34168
rect 1152 34040 20452 34064
rect 1152 34000 4928 34040
rect 4968 34000 5010 34040
rect 5050 34000 5092 34040
rect 5132 34000 5174 34040
rect 5214 34000 5256 34040
rect 5296 34000 20048 34040
rect 20088 34000 20130 34040
rect 20170 34000 20212 34040
rect 20252 34000 20294 34040
rect 20334 34000 20376 34040
rect 20416 34000 20452 34040
rect 1152 33976 20452 34000
rect 1419 33872 1461 33881
rect 1419 33832 1420 33872
rect 1460 33832 1461 33872
rect 1419 33823 1461 33832
rect 3627 33872 3669 33881
rect 3627 33832 3628 33872
rect 3668 33832 3669 33872
rect 3627 33823 3669 33832
rect 4107 33872 4149 33881
rect 4107 33832 4108 33872
rect 4148 33832 4149 33872
rect 4107 33823 4149 33832
rect 7947 33872 7989 33881
rect 7947 33832 7948 33872
rect 7988 33832 7989 33872
rect 7947 33823 7989 33832
rect 12363 33872 12405 33881
rect 12363 33832 12364 33872
rect 12404 33832 12405 33872
rect 12363 33823 12405 33832
rect 14659 33872 14717 33873
rect 14659 33832 14668 33872
rect 14708 33832 14717 33872
rect 14659 33831 14717 33832
rect 16683 33872 16725 33881
rect 16683 33832 16684 33872
rect 16724 33832 16725 33872
rect 16683 33823 16725 33832
rect 8427 33788 8469 33797
rect 8427 33748 8428 33788
rect 8468 33748 8469 33788
rect 8427 33739 8469 33748
rect 1603 33704 1661 33705
rect 1603 33664 1612 33704
rect 1652 33664 1661 33704
rect 1603 33663 1661 33664
rect 2851 33704 2909 33705
rect 2851 33664 2860 33704
rect 2900 33664 2909 33704
rect 4771 33704 4829 33705
rect 2851 33663 2909 33664
rect 4299 33690 4341 33699
rect 4299 33650 4300 33690
rect 4340 33650 4341 33690
rect 4771 33664 4780 33704
rect 4820 33664 4829 33704
rect 4771 33663 4829 33664
rect 5259 33704 5301 33713
rect 5259 33664 5260 33704
rect 5300 33664 5301 33704
rect 5259 33655 5301 33664
rect 5739 33704 5781 33713
rect 5739 33664 5740 33704
rect 5780 33664 5781 33704
rect 5739 33655 5781 33664
rect 5835 33704 5877 33713
rect 5835 33664 5836 33704
rect 5876 33664 5877 33704
rect 5835 33655 5877 33664
rect 6219 33704 6261 33713
rect 6219 33664 6220 33704
rect 6260 33664 6261 33704
rect 6219 33655 6261 33664
rect 6315 33704 6357 33713
rect 6315 33664 6316 33704
rect 6356 33664 6357 33704
rect 6315 33655 6357 33664
rect 7267 33704 7325 33705
rect 7267 33664 7276 33704
rect 7316 33664 7325 33704
rect 7267 33663 7325 33664
rect 7755 33699 7797 33708
rect 7755 33659 7756 33699
rect 7796 33659 7797 33699
rect 8611 33704 8669 33705
rect 8611 33664 8620 33704
rect 8660 33664 8669 33704
rect 8611 33663 8669 33664
rect 9859 33704 9917 33705
rect 9859 33664 9868 33704
rect 9908 33664 9917 33704
rect 9859 33663 9917 33664
rect 10051 33704 10109 33705
rect 10051 33664 10060 33704
rect 10100 33664 10109 33704
rect 10051 33663 10109 33664
rect 10251 33704 10293 33713
rect 10251 33664 10252 33704
rect 10292 33664 10293 33704
rect 7755 33650 7797 33659
rect 10251 33655 10293 33664
rect 10339 33704 10397 33705
rect 10339 33664 10348 33704
rect 10388 33664 10397 33704
rect 10339 33663 10397 33664
rect 10635 33704 10677 33713
rect 10635 33664 10636 33704
rect 10676 33664 10677 33704
rect 10635 33655 10677 33664
rect 10731 33704 10773 33713
rect 10731 33664 10732 33704
rect 10772 33664 10773 33704
rect 10731 33655 10773 33664
rect 11683 33704 11741 33705
rect 11683 33664 11692 33704
rect 11732 33664 11741 33704
rect 13795 33704 13853 33705
rect 11683 33663 11741 33664
rect 12219 33694 12261 33703
rect 12219 33654 12220 33694
rect 12260 33654 12261 33694
rect 13795 33664 13804 33704
rect 13844 33664 13853 33704
rect 13795 33663 13853 33664
rect 14179 33704 14237 33705
rect 14179 33664 14188 33704
rect 14228 33664 14237 33704
rect 14179 33663 14237 33664
rect 14275 33704 14333 33705
rect 14275 33664 14284 33704
rect 14324 33664 14333 33704
rect 14275 33663 14333 33664
rect 14475 33704 14517 33713
rect 14475 33664 14476 33704
rect 14516 33664 14517 33704
rect 4299 33641 4341 33650
rect 12219 33645 12261 33654
rect 12547 33662 12605 33663
rect 1219 33620 1277 33621
rect 1219 33580 1228 33620
rect 1268 33580 1277 33620
rect 1219 33579 1277 33580
rect 3235 33620 3293 33621
rect 3235 33580 3244 33620
rect 3284 33580 3293 33620
rect 3235 33579 3293 33580
rect 3811 33620 3869 33621
rect 3811 33580 3820 33620
rect 3860 33580 3869 33620
rect 3811 33579 3869 33580
rect 5355 33620 5397 33629
rect 5355 33580 5356 33620
rect 5396 33580 5397 33620
rect 5355 33571 5397 33580
rect 6699 33620 6741 33629
rect 6699 33580 6700 33620
rect 6740 33580 6741 33620
rect 6699 33571 6741 33580
rect 6795 33620 6837 33629
rect 6795 33580 6796 33620
rect 6836 33580 6837 33620
rect 6795 33571 6837 33580
rect 11115 33620 11157 33629
rect 11115 33580 11116 33620
rect 11156 33580 11157 33620
rect 11115 33571 11157 33580
rect 11211 33620 11253 33629
rect 12547 33622 12556 33662
rect 12596 33622 12605 33662
rect 14475 33655 14517 33664
rect 14571 33704 14613 33713
rect 14571 33664 14572 33704
rect 14612 33664 14613 33704
rect 14571 33655 14613 33664
rect 14664 33704 14722 33705
rect 14664 33664 14673 33704
rect 14713 33664 14722 33704
rect 14664 33663 14722 33664
rect 15531 33704 15573 33713
rect 15531 33664 15532 33704
rect 15572 33664 15573 33704
rect 15531 33655 15573 33664
rect 15627 33704 15669 33713
rect 15627 33664 15628 33704
rect 15668 33664 15669 33704
rect 15627 33655 15669 33664
rect 15907 33704 15965 33705
rect 15907 33664 15916 33704
rect 15956 33664 15965 33704
rect 16395 33704 16437 33713
rect 15907 33663 15965 33664
rect 16195 33691 16253 33692
rect 16195 33651 16204 33691
rect 16244 33651 16253 33691
rect 16395 33664 16396 33704
rect 16436 33664 16437 33704
rect 16395 33655 16437 33664
rect 16483 33704 16541 33705
rect 16483 33664 16492 33704
rect 16532 33664 16541 33704
rect 16483 33663 16541 33664
rect 16867 33704 16925 33705
rect 16867 33664 16876 33704
rect 16916 33664 16925 33704
rect 16867 33663 16925 33664
rect 18115 33704 18173 33705
rect 18115 33664 18124 33704
rect 18164 33664 18173 33704
rect 18115 33663 18173 33664
rect 18403 33704 18461 33705
rect 18403 33664 18412 33704
rect 18452 33664 18461 33704
rect 18403 33663 18461 33664
rect 18699 33704 18741 33713
rect 18699 33664 18700 33704
rect 18740 33664 18741 33704
rect 18699 33655 18741 33664
rect 18795 33704 18837 33713
rect 18795 33664 18796 33704
rect 18836 33664 18837 33704
rect 18795 33655 18837 33664
rect 19275 33704 19317 33713
rect 19275 33664 19276 33704
rect 19316 33664 19317 33704
rect 19275 33655 19317 33664
rect 19651 33704 19709 33705
rect 19651 33664 19660 33704
rect 19700 33664 19709 33704
rect 19651 33663 19709 33664
rect 16195 33650 16253 33651
rect 12547 33621 12605 33622
rect 11211 33580 11212 33620
rect 11252 33580 11253 33620
rect 11211 33571 11253 33580
rect 19371 33620 19413 33629
rect 19371 33580 19372 33620
rect 19412 33580 19413 33620
rect 19371 33571 19413 33580
rect 19563 33620 19605 33629
rect 19563 33580 19564 33620
rect 19604 33580 19605 33620
rect 19563 33571 19605 33580
rect 19843 33620 19901 33621
rect 19843 33580 19852 33620
rect 19892 33580 19901 33620
rect 19843 33579 19901 33580
rect 8139 33536 8181 33545
rect 8139 33496 8140 33536
rect 8180 33496 8181 33536
rect 8139 33487 8181 33496
rect 14955 33536 14997 33545
rect 14955 33496 14956 33536
rect 14996 33496 14997 33536
rect 14955 33487 14997 33496
rect 19075 33536 19133 33537
rect 19075 33496 19084 33536
rect 19124 33496 19133 33536
rect 19075 33495 19133 33496
rect 19467 33536 19509 33545
rect 19467 33496 19468 33536
rect 19508 33496 19509 33536
rect 19467 33487 19509 33496
rect 3051 33452 3093 33461
rect 3051 33412 3052 33452
rect 3092 33412 3093 33452
rect 3051 33403 3093 33412
rect 3435 33452 3477 33461
rect 3435 33412 3436 33452
rect 3476 33412 3477 33452
rect 3435 33403 3477 33412
rect 10059 33452 10101 33461
rect 10059 33412 10060 33452
rect 10100 33412 10101 33452
rect 10059 33403 10101 33412
rect 13995 33452 14037 33461
rect 13995 33412 13996 33452
rect 14036 33412 14037 33452
rect 13995 33403 14037 33412
rect 15235 33452 15293 33453
rect 15235 33412 15244 33452
rect 15284 33412 15293 33452
rect 15235 33411 15293 33412
rect 16203 33452 16245 33461
rect 16203 33412 16204 33452
rect 16244 33412 16245 33452
rect 16203 33403 16245 33412
rect 20043 33452 20085 33461
rect 20043 33412 20044 33452
rect 20084 33412 20085 33452
rect 20043 33403 20085 33412
rect 1152 33284 20352 33308
rect 1152 33244 3688 33284
rect 3728 33244 3770 33284
rect 3810 33244 3852 33284
rect 3892 33244 3934 33284
rect 3974 33244 4016 33284
rect 4056 33244 18808 33284
rect 18848 33244 18890 33284
rect 18930 33244 18972 33284
rect 19012 33244 19054 33284
rect 19094 33244 19136 33284
rect 19176 33244 20352 33284
rect 1152 33220 20352 33244
rect 3435 33116 3477 33125
rect 3435 33076 3436 33116
rect 3476 33076 3477 33116
rect 3435 33067 3477 33076
rect 3819 33116 3861 33125
rect 3819 33076 3820 33116
rect 3860 33076 3861 33116
rect 3819 33067 3861 33076
rect 6123 33116 6165 33125
rect 6123 33076 6124 33116
rect 6164 33076 6165 33116
rect 6123 33067 6165 33076
rect 7755 33116 7797 33125
rect 7755 33076 7756 33116
rect 7796 33076 7797 33116
rect 7755 33067 7797 33076
rect 12651 33116 12693 33125
rect 12651 33076 12652 33116
rect 12692 33076 12693 33116
rect 12651 33067 12693 33076
rect 15051 33116 15093 33125
rect 15051 33076 15052 33116
rect 15092 33076 15093 33116
rect 15051 33067 15093 33076
rect 15435 33116 15477 33125
rect 15435 33076 15436 33116
rect 15476 33076 15477 33116
rect 15435 33067 15477 33076
rect 19275 33116 19317 33125
rect 19275 33076 19276 33116
rect 19316 33076 19317 33116
rect 19275 33067 19317 33076
rect 5931 33032 5973 33041
rect 5931 32992 5932 33032
rect 5972 32992 5973 33032
rect 5931 32983 5973 32992
rect 14667 33032 14709 33041
rect 14667 32992 14668 33032
rect 14708 32992 14709 33032
rect 14667 32983 14709 32992
rect 17259 33032 17301 33041
rect 17259 32992 17260 33032
rect 17300 32992 17301 33032
rect 17259 32983 17301 32992
rect 18307 33032 18365 33033
rect 18307 32992 18316 33032
rect 18356 32992 18365 33032
rect 18307 32991 18365 32992
rect 19947 33032 19989 33041
rect 19947 32992 19948 33032
rect 19988 32992 19989 33032
rect 19947 32983 19989 32992
rect 14467 32948 14525 32949
rect 14467 32908 14476 32948
rect 14516 32908 14525 32948
rect 14467 32907 14525 32908
rect 14851 32948 14909 32949
rect 14851 32908 14860 32948
rect 14900 32908 14909 32948
rect 14851 32907 14909 32908
rect 19851 32948 19893 32957
rect 19851 32908 19852 32948
rect 19892 32908 19893 32948
rect 19851 32899 19893 32908
rect 20043 32948 20085 32957
rect 20043 32908 20044 32948
rect 20084 32908 20085 32948
rect 20043 32899 20085 32908
rect 20139 32906 20181 32915
rect 1315 32864 1373 32865
rect 1315 32824 1324 32864
rect 1364 32824 1373 32864
rect 1315 32823 1373 32824
rect 2563 32864 2621 32865
rect 2563 32824 2572 32864
rect 2612 32824 2621 32864
rect 2563 32823 2621 32824
rect 3043 32864 3101 32865
rect 3043 32824 3052 32864
rect 3092 32824 3101 32864
rect 3043 32823 3101 32824
rect 3243 32864 3285 32873
rect 3243 32824 3244 32864
rect 3284 32824 3285 32864
rect 3243 32815 3285 32824
rect 3435 32864 3477 32873
rect 3435 32824 3436 32864
rect 3476 32824 3477 32864
rect 3435 32815 3477 32824
rect 3627 32864 3669 32873
rect 3627 32824 3628 32864
rect 3668 32824 3669 32864
rect 3627 32815 3669 32824
rect 3819 32864 3861 32873
rect 3819 32824 3820 32864
rect 3860 32824 3861 32864
rect 3819 32815 3861 32824
rect 4011 32864 4053 32873
rect 4011 32824 4012 32864
rect 4052 32824 4053 32864
rect 4011 32815 4053 32824
rect 4107 32864 4149 32873
rect 4107 32824 4108 32864
rect 4148 32824 4149 32864
rect 4107 32815 4149 32824
rect 4203 32864 4245 32873
rect 4203 32824 4204 32864
rect 4244 32824 4245 32864
rect 4203 32815 4245 32824
rect 4299 32864 4341 32873
rect 4299 32824 4300 32864
rect 4340 32824 4341 32864
rect 4299 32815 4341 32824
rect 4483 32864 4541 32865
rect 4483 32824 4492 32864
rect 4532 32824 4541 32864
rect 4483 32823 4541 32824
rect 5731 32864 5789 32865
rect 5731 32824 5740 32864
rect 5780 32824 5789 32864
rect 5731 32823 5789 32824
rect 6307 32864 6365 32865
rect 6307 32824 6316 32864
rect 6356 32824 6365 32864
rect 6307 32823 6365 32824
rect 7555 32864 7613 32865
rect 7555 32824 7564 32864
rect 7604 32824 7613 32864
rect 7555 32823 7613 32824
rect 7939 32864 7997 32865
rect 7939 32824 7948 32864
rect 7988 32824 7997 32864
rect 7939 32823 7997 32824
rect 9187 32864 9245 32865
rect 9187 32824 9196 32864
rect 9236 32824 9245 32864
rect 9187 32823 9245 32824
rect 9579 32864 9621 32873
rect 9579 32824 9580 32864
rect 9620 32824 9621 32864
rect 9579 32815 9621 32824
rect 9675 32864 9717 32873
rect 9675 32824 9676 32864
rect 9716 32824 9717 32864
rect 9675 32815 9717 32824
rect 10059 32864 10101 32873
rect 10059 32824 10060 32864
rect 10100 32824 10101 32864
rect 10251 32864 10293 32873
rect 10059 32815 10101 32824
rect 10155 32843 10197 32852
rect 10155 32803 10156 32843
rect 10196 32803 10197 32843
rect 10251 32824 10252 32864
rect 10292 32824 10293 32864
rect 10251 32815 10293 32824
rect 10347 32864 10389 32873
rect 10347 32824 10348 32864
rect 10388 32824 10389 32864
rect 10347 32815 10389 32824
rect 10627 32864 10685 32865
rect 10627 32824 10636 32864
rect 10676 32824 10685 32864
rect 10627 32823 10685 32824
rect 11875 32864 11933 32865
rect 11875 32824 11884 32864
rect 11924 32824 11933 32864
rect 11875 32823 11933 32824
rect 12835 32864 12893 32865
rect 12835 32824 12844 32864
rect 12884 32824 12893 32864
rect 12835 32823 12893 32824
rect 14083 32864 14141 32865
rect 14083 32824 14092 32864
rect 14132 32824 14141 32864
rect 14083 32823 14141 32824
rect 15243 32864 15285 32873
rect 15243 32824 15244 32864
rect 15284 32824 15285 32864
rect 15243 32815 15285 32824
rect 15435 32864 15477 32873
rect 15435 32824 15436 32864
rect 15476 32824 15477 32864
rect 15435 32815 15477 32824
rect 15811 32864 15869 32865
rect 15811 32824 15820 32864
rect 15860 32824 15869 32864
rect 15811 32823 15869 32824
rect 17059 32864 17117 32865
rect 17059 32824 17068 32864
rect 17108 32824 17117 32864
rect 17059 32823 17117 32824
rect 17635 32864 17693 32865
rect 17635 32824 17644 32864
rect 17684 32824 17693 32864
rect 17635 32823 17693 32824
rect 17931 32864 17973 32873
rect 17931 32824 17932 32864
rect 17972 32824 17973 32864
rect 17931 32815 17973 32824
rect 18027 32864 18069 32873
rect 20139 32866 20140 32906
rect 20180 32866 20181 32906
rect 18027 32824 18028 32864
rect 18068 32824 18069 32864
rect 18027 32815 18069 32824
rect 18595 32864 18653 32865
rect 18595 32824 18604 32864
rect 18644 32824 18653 32864
rect 18595 32823 18653 32824
rect 19747 32864 19805 32865
rect 19747 32824 19756 32864
rect 19796 32824 19805 32864
rect 20139 32857 20181 32866
rect 19747 32823 19805 32824
rect 10155 32794 10197 32803
rect 12459 32780 12501 32789
rect 12459 32740 12460 32780
rect 12500 32740 12501 32780
rect 12459 32731 12501 32740
rect 19459 32780 19517 32781
rect 19459 32740 19468 32780
rect 19508 32740 19517 32780
rect 19459 32739 19517 32740
rect 2763 32696 2805 32705
rect 2763 32656 2764 32696
rect 2804 32656 2805 32696
rect 2763 32647 2805 32656
rect 2955 32696 2997 32705
rect 2955 32656 2956 32696
rect 2996 32656 2997 32696
rect 2955 32647 2997 32656
rect 9859 32696 9917 32697
rect 9859 32656 9868 32696
rect 9908 32656 9917 32696
rect 9859 32655 9917 32656
rect 12075 32696 12117 32705
rect 12075 32656 12076 32696
rect 12116 32656 12117 32696
rect 12075 32647 12117 32656
rect 15339 32696 15381 32705
rect 15339 32656 15340 32696
rect 15380 32656 15381 32696
rect 15339 32647 15381 32656
rect 15627 32696 15669 32705
rect 15627 32656 15628 32696
rect 15668 32656 15669 32696
rect 15627 32647 15669 32656
rect 1152 32528 20452 32552
rect 1152 32488 4928 32528
rect 4968 32488 5010 32528
rect 5050 32488 5092 32528
rect 5132 32488 5174 32528
rect 5214 32488 5256 32528
rect 5296 32488 20048 32528
rect 20088 32488 20130 32528
rect 20170 32488 20212 32528
rect 20252 32488 20294 32528
rect 20334 32488 20376 32528
rect 20416 32488 20452 32528
rect 1152 32464 20452 32488
rect 1323 32360 1365 32369
rect 1323 32320 1324 32360
rect 1364 32320 1365 32360
rect 1323 32311 1365 32320
rect 1707 32360 1749 32369
rect 1707 32320 1708 32360
rect 1748 32320 1749 32360
rect 1707 32311 1749 32320
rect 3723 32360 3765 32369
rect 3723 32320 3724 32360
rect 3764 32320 3765 32360
rect 3723 32311 3765 32320
rect 4387 32360 4445 32361
rect 4387 32320 4396 32360
rect 4436 32320 4445 32360
rect 4387 32319 4445 32320
rect 6219 32360 6261 32369
rect 6219 32320 6220 32360
rect 6260 32320 6261 32360
rect 6219 32311 6261 32320
rect 8139 32360 8181 32369
rect 8139 32320 8140 32360
rect 8180 32320 8181 32360
rect 8139 32311 8181 32320
rect 12451 32360 12509 32361
rect 12451 32320 12460 32360
rect 12500 32320 12509 32360
rect 12451 32319 12509 32320
rect 15907 32360 15965 32361
rect 15907 32320 15916 32360
rect 15956 32320 15965 32360
rect 15907 32319 15965 32320
rect 17643 32360 17685 32369
rect 17643 32320 17644 32360
rect 17684 32320 17685 32360
rect 17643 32311 17685 32320
rect 10251 32276 10293 32285
rect 10251 32236 10252 32276
rect 10292 32236 10293 32276
rect 10251 32227 10293 32236
rect 12267 32276 12309 32285
rect 12267 32236 12268 32276
rect 12308 32236 12309 32276
rect 12267 32227 12309 32236
rect 1219 32192 1277 32193
rect 1219 32152 1228 32192
rect 1268 32152 1277 32192
rect 1219 32151 1277 32152
rect 1995 32192 2037 32201
rect 1995 32152 1996 32192
rect 2036 32152 2037 32192
rect 1995 32143 2037 32152
rect 2091 32192 2133 32201
rect 2091 32152 2092 32192
rect 2132 32152 2133 32192
rect 2091 32143 2133 32152
rect 3043 32192 3101 32193
rect 3043 32152 3052 32192
rect 3092 32152 3101 32192
rect 3907 32192 3965 32193
rect 3043 32151 3101 32152
rect 3531 32178 3573 32187
rect 3531 32138 3532 32178
rect 3572 32138 3573 32178
rect 3907 32152 3916 32192
rect 3956 32152 3965 32192
rect 3907 32151 3965 32152
rect 4003 32192 4061 32193
rect 4003 32152 4012 32192
rect 4052 32152 4061 32192
rect 4003 32151 4061 32152
rect 4203 32192 4245 32201
rect 4203 32152 4204 32192
rect 4244 32152 4245 32192
rect 4203 32143 4245 32152
rect 4299 32192 4341 32201
rect 4299 32152 4300 32192
rect 4340 32152 4341 32192
rect 4299 32143 4341 32152
rect 4392 32192 4450 32193
rect 4392 32152 4401 32192
rect 4441 32152 4450 32192
rect 4392 32151 4450 32152
rect 4771 32192 4829 32193
rect 4771 32152 4780 32192
rect 4820 32152 4829 32192
rect 4771 32151 4829 32152
rect 6019 32192 6077 32193
rect 6019 32152 6028 32192
rect 6068 32152 6077 32192
rect 6019 32151 6077 32152
rect 6403 32192 6461 32193
rect 6403 32152 6412 32192
rect 6452 32152 6461 32192
rect 6403 32151 6461 32152
rect 7651 32192 7709 32193
rect 7651 32152 7660 32192
rect 7700 32152 7709 32192
rect 7651 32151 7709 32152
rect 8331 32192 8373 32201
rect 8331 32152 8332 32192
rect 8372 32152 8373 32192
rect 8331 32143 8373 32152
rect 8523 32192 8565 32201
rect 8523 32152 8524 32192
rect 8564 32152 8565 32192
rect 8523 32143 8565 32152
rect 8619 32192 8661 32201
rect 8619 32152 8620 32192
rect 8660 32152 8661 32192
rect 8619 32143 8661 32152
rect 8803 32192 8861 32193
rect 8803 32152 8812 32192
rect 8852 32152 8861 32192
rect 8803 32151 8861 32152
rect 10051 32192 10109 32193
rect 10051 32152 10060 32192
rect 10100 32152 10109 32192
rect 10051 32151 10109 32152
rect 10539 32192 10581 32201
rect 10539 32152 10540 32192
rect 10580 32152 10581 32192
rect 10539 32143 10581 32152
rect 10635 32192 10677 32201
rect 10635 32152 10636 32192
rect 10676 32152 10677 32192
rect 10635 32143 10677 32152
rect 11019 32192 11061 32201
rect 11019 32152 11020 32192
rect 11060 32152 11061 32192
rect 11019 32143 11061 32152
rect 11587 32192 11645 32193
rect 11587 32152 11596 32192
rect 11636 32152 11645 32192
rect 11587 32151 11645 32152
rect 12075 32187 12117 32196
rect 12075 32147 12076 32187
rect 12116 32147 12117 32187
rect 12739 32192 12797 32193
rect 12739 32152 12748 32192
rect 12788 32152 12797 32192
rect 12739 32151 12797 32152
rect 13987 32192 14045 32193
rect 13987 32152 13996 32192
rect 14036 32152 14045 32192
rect 13987 32151 14045 32152
rect 14667 32192 14709 32201
rect 14667 32152 14668 32192
rect 14708 32152 14709 32192
rect 12075 32138 12117 32147
rect 14667 32143 14709 32152
rect 14763 32192 14805 32201
rect 14763 32152 14764 32192
rect 14804 32152 14805 32192
rect 14763 32143 14805 32152
rect 15043 32192 15101 32193
rect 15043 32152 15052 32192
rect 15092 32152 15101 32192
rect 15043 32151 15101 32152
rect 15339 32192 15381 32201
rect 15339 32152 15340 32192
rect 15380 32152 15381 32192
rect 15339 32143 15381 32152
rect 15715 32192 15773 32193
rect 15715 32152 15724 32192
rect 15764 32152 15773 32192
rect 15715 32151 15773 32152
rect 16195 32192 16253 32193
rect 16195 32152 16204 32192
rect 16244 32152 16253 32192
rect 16195 32151 16253 32152
rect 17443 32192 17501 32193
rect 17443 32152 17452 32192
rect 17492 32152 17501 32192
rect 17443 32151 17501 32152
rect 17835 32192 17877 32201
rect 17835 32152 17836 32192
rect 17876 32152 17877 32192
rect 17835 32143 17877 32152
rect 18027 32192 18069 32201
rect 18027 32152 18028 32192
rect 18068 32152 18069 32192
rect 18027 32143 18069 32152
rect 18211 32192 18269 32193
rect 18211 32152 18220 32192
rect 18260 32152 18269 32192
rect 18211 32151 18269 32152
rect 19459 32192 19517 32193
rect 19459 32152 19468 32192
rect 19508 32152 19517 32192
rect 19459 32151 19517 32152
rect 3531 32129 3573 32138
rect 1507 32108 1565 32109
rect 1507 32068 1516 32108
rect 1556 32068 1565 32108
rect 1507 32067 1565 32068
rect 2475 32108 2517 32117
rect 2475 32068 2476 32108
rect 2516 32068 2517 32108
rect 2475 32059 2517 32068
rect 2571 32108 2613 32117
rect 2571 32068 2572 32108
rect 2612 32068 2613 32108
rect 2571 32059 2613 32068
rect 11115 32108 11157 32117
rect 11115 32068 11116 32108
rect 11156 32068 11157 32108
rect 11115 32059 11157 32068
rect 15435 32108 15477 32117
rect 15435 32068 15436 32108
rect 15476 32068 15477 32108
rect 15435 32059 15477 32068
rect 15627 32108 15669 32117
rect 15627 32068 15628 32108
rect 15668 32068 15669 32108
rect 15627 32059 15669 32068
rect 19843 32108 19901 32109
rect 19843 32068 19852 32108
rect 19892 32068 19901 32108
rect 19843 32067 19901 32068
rect 8043 32024 8085 32033
rect 8043 31984 8044 32024
rect 8084 31984 8085 32024
rect 8043 31975 8085 31984
rect 8611 32024 8669 32025
rect 8611 31984 8620 32024
rect 8660 31984 8669 32024
rect 8611 31983 8669 31984
rect 14371 32024 14429 32025
rect 14371 31984 14380 32024
rect 14420 31984 14429 32024
rect 14371 31983 14429 31984
rect 15531 32024 15573 32033
rect 15531 31984 15532 32024
rect 15572 31984 15573 32024
rect 15531 31975 15573 31984
rect 7851 31940 7893 31949
rect 7851 31900 7852 31940
rect 7892 31900 7893 31940
rect 7851 31891 7893 31900
rect 14187 31940 14229 31949
rect 14187 31900 14188 31940
rect 14228 31900 14229 31940
rect 14187 31891 14229 31900
rect 17643 31940 17685 31949
rect 17643 31900 17644 31940
rect 17684 31900 17685 31940
rect 17643 31891 17685 31900
rect 17835 31940 17877 31949
rect 17835 31900 17836 31940
rect 17876 31900 17877 31940
rect 17835 31891 17877 31900
rect 19659 31940 19701 31949
rect 19659 31900 19660 31940
rect 19700 31900 19701 31940
rect 19659 31891 19701 31900
rect 20043 31940 20085 31949
rect 20043 31900 20044 31940
rect 20084 31900 20085 31940
rect 20043 31891 20085 31900
rect 1152 31772 20352 31796
rect 1152 31732 3688 31772
rect 3728 31732 3770 31772
rect 3810 31732 3852 31772
rect 3892 31732 3934 31772
rect 3974 31732 4016 31772
rect 4056 31732 18808 31772
rect 18848 31732 18890 31772
rect 18930 31732 18972 31772
rect 19012 31732 19054 31772
rect 19094 31732 19136 31772
rect 19176 31732 20352 31772
rect 1152 31708 20352 31732
rect 9867 31604 9909 31613
rect 9867 31564 9868 31604
rect 9908 31564 9909 31604
rect 9867 31555 9909 31564
rect 2179 31520 2237 31521
rect 2179 31480 2188 31520
rect 2228 31480 2237 31520
rect 2179 31479 2237 31480
rect 16675 31520 16733 31521
rect 16675 31480 16684 31520
rect 16724 31480 16733 31520
rect 16675 31479 16733 31480
rect 18403 31520 18461 31521
rect 18403 31480 18412 31520
rect 18452 31480 18461 31520
rect 18403 31479 18461 31480
rect 19659 31520 19701 31529
rect 19659 31480 19660 31520
rect 19700 31480 19701 31520
rect 19659 31471 19701 31480
rect 6699 31436 6741 31445
rect 6699 31396 6700 31436
rect 6740 31396 6741 31436
rect 2083 31394 2141 31395
rect 2083 31354 2092 31394
rect 2132 31354 2141 31394
rect 6699 31387 6741 31396
rect 8139 31436 8181 31445
rect 8139 31396 8140 31436
rect 8180 31396 8181 31436
rect 14763 31436 14805 31445
rect 8139 31387 8181 31396
rect 13515 31392 13557 31401
rect 7659 31366 7701 31375
rect 2083 31353 2141 31354
rect 1891 31352 1949 31353
rect 1891 31312 1900 31352
rect 1940 31312 1949 31352
rect 1891 31311 1949 31312
rect 2187 31352 2229 31361
rect 2187 31312 2188 31352
rect 2228 31312 2229 31352
rect 2187 31303 2229 31312
rect 2371 31352 2429 31353
rect 2371 31312 2380 31352
rect 2420 31312 2429 31352
rect 2371 31311 2429 31312
rect 2563 31352 2621 31353
rect 2563 31312 2572 31352
rect 2612 31312 2621 31352
rect 2563 31311 2621 31312
rect 3811 31352 3869 31353
rect 3811 31312 3820 31352
rect 3860 31312 3869 31352
rect 3811 31311 3869 31312
rect 4195 31352 4253 31353
rect 4195 31312 4204 31352
rect 4244 31312 4253 31352
rect 4195 31311 4253 31312
rect 5443 31352 5501 31353
rect 5443 31312 5452 31352
rect 5492 31312 5501 31352
rect 5443 31311 5501 31312
rect 6123 31352 6165 31361
rect 6123 31312 6124 31352
rect 6164 31312 6165 31352
rect 6123 31303 6165 31312
rect 6219 31352 6261 31361
rect 6219 31312 6220 31352
rect 6260 31312 6261 31352
rect 6219 31303 6261 31312
rect 6603 31352 6645 31361
rect 6603 31312 6604 31352
rect 6644 31312 6645 31352
rect 6603 31303 6645 31312
rect 7171 31352 7229 31353
rect 7171 31312 7180 31352
rect 7220 31312 7229 31352
rect 7659 31326 7660 31366
rect 7700 31326 7701 31366
rect 7659 31317 7701 31326
rect 8035 31352 8093 31353
rect 7171 31311 7229 31312
rect 8035 31312 8044 31352
rect 8084 31312 8093 31352
rect 8035 31311 8093 31312
rect 8235 31352 8277 31361
rect 8235 31312 8236 31352
rect 8276 31312 8277 31352
rect 8235 31303 8277 31312
rect 8419 31352 8477 31353
rect 8419 31312 8428 31352
rect 8468 31312 8477 31352
rect 8419 31311 8477 31312
rect 9667 31352 9725 31353
rect 9667 31312 9676 31352
rect 9716 31312 9725 31352
rect 9667 31311 9725 31312
rect 10051 31352 10109 31353
rect 10051 31312 10060 31352
rect 10100 31312 10109 31352
rect 10051 31311 10109 31312
rect 11299 31352 11357 31353
rect 11299 31312 11308 31352
rect 11348 31312 11357 31352
rect 11299 31311 11357 31312
rect 11683 31352 11741 31353
rect 11683 31312 11692 31352
rect 11732 31312 11741 31352
rect 11683 31311 11741 31312
rect 12931 31352 12989 31353
rect 12931 31312 12940 31352
rect 12980 31312 12989 31352
rect 13515 31352 13516 31392
rect 13556 31352 13557 31392
rect 14763 31396 14764 31436
rect 14804 31396 14805 31436
rect 14763 31387 14805 31396
rect 19563 31436 19605 31445
rect 19563 31396 19564 31436
rect 19604 31396 19605 31436
rect 19563 31387 19605 31396
rect 19755 31436 19797 31445
rect 19755 31396 19756 31436
rect 19796 31396 19797 31436
rect 19755 31387 19797 31396
rect 20035 31436 20093 31437
rect 20035 31396 20044 31436
rect 20084 31396 20093 31436
rect 20035 31395 20093 31396
rect 18733 31367 18775 31376
rect 13515 31343 13557 31352
rect 13611 31352 13653 31361
rect 12931 31311 12989 31312
rect 13611 31312 13612 31352
rect 13652 31312 13653 31352
rect 13611 31303 13653 31312
rect 13707 31352 13749 31361
rect 13707 31312 13708 31352
rect 13748 31312 13749 31352
rect 13707 31303 13749 31312
rect 13899 31352 13941 31361
rect 13899 31312 13900 31352
rect 13940 31312 13941 31352
rect 13899 31303 13941 31312
rect 14091 31352 14133 31361
rect 14091 31312 14092 31352
rect 14132 31312 14133 31352
rect 14091 31303 14133 31312
rect 14179 31352 14237 31353
rect 14179 31312 14188 31352
rect 14228 31312 14237 31352
rect 14179 31311 14237 31312
rect 14659 31352 14717 31353
rect 14659 31312 14668 31352
rect 14708 31312 14717 31352
rect 14659 31311 14717 31312
rect 15139 31352 15197 31353
rect 15139 31312 15148 31352
rect 15188 31312 15197 31352
rect 15139 31311 15197 31312
rect 16387 31352 16445 31353
rect 16387 31312 16396 31352
rect 16436 31312 16445 31352
rect 16387 31311 16445 31312
rect 17067 31352 17109 31361
rect 17067 31312 17068 31352
rect 17108 31312 17109 31352
rect 17067 31303 17109 31312
rect 17347 31352 17405 31353
rect 17347 31312 17356 31352
rect 17396 31312 17405 31352
rect 17347 31311 17405 31312
rect 17731 31352 17789 31353
rect 17731 31312 17740 31352
rect 17780 31312 17789 31352
rect 17731 31311 17789 31312
rect 18027 31352 18069 31361
rect 18027 31312 18028 31352
rect 18068 31312 18069 31352
rect 18733 31327 18734 31367
rect 18774 31327 18775 31367
rect 18733 31318 18775 31327
rect 18891 31352 18933 31361
rect 18027 31303 18069 31312
rect 18891 31312 18892 31352
rect 18932 31312 18933 31352
rect 18891 31303 18933 31312
rect 18987 31352 19029 31361
rect 18987 31312 18988 31352
rect 19028 31312 19029 31352
rect 18987 31303 19029 31312
rect 19171 31352 19229 31353
rect 19171 31312 19180 31352
rect 19220 31312 19229 31352
rect 19171 31311 19229 31312
rect 19267 31352 19325 31353
rect 19267 31312 19276 31352
rect 19316 31312 19325 31352
rect 19267 31311 19325 31312
rect 19467 31352 19509 31361
rect 19467 31312 19468 31352
rect 19508 31312 19509 31352
rect 19467 31303 19509 31312
rect 19843 31352 19901 31353
rect 19843 31312 19852 31352
rect 19892 31312 19901 31352
rect 19843 31311 19901 31312
rect 1611 31268 1653 31277
rect 1611 31228 1612 31268
rect 1652 31228 1653 31268
rect 1611 31219 1653 31228
rect 5643 31268 5685 31277
rect 5643 31228 5644 31268
rect 5684 31228 5685 31268
rect 5643 31219 5685 31228
rect 7851 31268 7893 31277
rect 7851 31228 7852 31268
rect 7892 31228 7893 31268
rect 7851 31219 7893 31228
rect 13995 31268 14037 31277
rect 13995 31228 13996 31268
rect 14036 31228 14037 31268
rect 13995 31219 14037 31228
rect 16971 31268 17013 31277
rect 16971 31228 16972 31268
rect 17012 31228 17013 31268
rect 16971 31219 17013 31228
rect 18123 31268 18165 31277
rect 18123 31228 18124 31268
rect 18164 31228 18165 31268
rect 18123 31219 18165 31228
rect 1315 31184 1373 31185
rect 1315 31144 1324 31184
rect 1364 31144 1373 31184
rect 1315 31143 1373 31144
rect 1803 31184 1845 31193
rect 1803 31144 1804 31184
rect 1844 31144 1845 31184
rect 1803 31135 1845 31144
rect 4011 31184 4053 31193
rect 4011 31144 4012 31184
rect 4052 31144 4053 31184
rect 4011 31135 4053 31144
rect 9867 31184 9909 31193
rect 9867 31144 9868 31184
rect 9908 31144 9909 31184
rect 9867 31135 9909 31144
rect 11499 31184 11541 31193
rect 11499 31144 11500 31184
rect 11540 31144 11541 31184
rect 11499 31135 11541 31144
rect 13131 31184 13173 31193
rect 13131 31144 13132 31184
rect 13172 31144 13173 31184
rect 13131 31135 13173 31144
rect 13411 31184 13469 31185
rect 13411 31144 13420 31184
rect 13460 31144 13469 31184
rect 13411 31143 13469 31144
rect 14371 31184 14429 31185
rect 14371 31144 14380 31184
rect 14420 31144 14429 31184
rect 14371 31143 14429 31144
rect 14955 31184 14997 31193
rect 14955 31144 14956 31184
rect 14996 31144 14997 31184
rect 14955 31135 14997 31144
rect 19075 31184 19133 31185
rect 19075 31144 19084 31184
rect 19124 31144 19133 31184
rect 19075 31143 19133 31144
rect 20235 31184 20277 31193
rect 20235 31144 20236 31184
rect 20276 31144 20277 31184
rect 20235 31135 20277 31144
rect 1152 31016 20452 31040
rect 1152 30976 4928 31016
rect 4968 30976 5010 31016
rect 5050 30976 5092 31016
rect 5132 30976 5174 31016
rect 5214 30976 5256 31016
rect 5296 30976 20048 31016
rect 20088 30976 20130 31016
rect 20170 30976 20212 31016
rect 20252 30976 20294 31016
rect 20334 30976 20376 31016
rect 20416 30976 20452 31016
rect 1152 30952 20452 30976
rect 5835 30848 5877 30857
rect 5835 30808 5836 30848
rect 5876 30808 5877 30848
rect 5835 30799 5877 30808
rect 9387 30848 9429 30857
rect 9387 30808 9388 30848
rect 9428 30808 9429 30848
rect 9387 30799 9429 30808
rect 9859 30848 9917 30849
rect 9859 30808 9868 30848
rect 9908 30808 9917 30848
rect 9859 30807 9917 30808
rect 14371 30848 14429 30849
rect 14371 30808 14380 30848
rect 14420 30808 14429 30848
rect 14371 30807 14429 30808
rect 17643 30848 17685 30857
rect 17643 30808 17644 30848
rect 17684 30808 17685 30848
rect 17643 30799 17685 30808
rect 20043 30848 20085 30857
rect 20043 30808 20044 30848
rect 20084 30808 20085 30848
rect 20043 30799 20085 30808
rect 2667 30764 2709 30773
rect 2667 30724 2668 30764
rect 2708 30724 2709 30764
rect 2667 30715 2709 30724
rect 11883 30764 11925 30773
rect 11883 30724 11884 30764
rect 11924 30724 11925 30764
rect 11883 30715 11925 30724
rect 13899 30764 13941 30773
rect 13899 30724 13900 30764
rect 13940 30724 13941 30764
rect 13899 30715 13941 30724
rect 17451 30764 17493 30773
rect 17451 30724 17452 30764
rect 17492 30724 17493 30764
rect 17451 30715 17493 30724
rect 19563 30764 19605 30773
rect 19563 30724 19564 30764
rect 19604 30724 19605 30764
rect 19563 30715 19605 30724
rect 14179 30691 14237 30692
rect 1219 30680 1277 30681
rect 1219 30640 1228 30680
rect 1268 30640 1277 30680
rect 1219 30639 1277 30640
rect 2467 30680 2525 30681
rect 2467 30640 2476 30680
rect 2516 30640 2525 30680
rect 2467 30639 2525 30640
rect 2859 30680 2901 30689
rect 2859 30640 2860 30680
rect 2900 30640 2901 30680
rect 2859 30631 2901 30640
rect 3051 30680 3093 30689
rect 3051 30640 3052 30680
rect 3092 30640 3093 30680
rect 3051 30631 3093 30640
rect 3331 30680 3389 30681
rect 3331 30640 3340 30680
rect 3380 30640 3389 30680
rect 3331 30639 3389 30640
rect 3627 30680 3669 30689
rect 3627 30640 3628 30680
rect 3668 30640 3669 30680
rect 3627 30631 3669 30640
rect 3723 30680 3765 30689
rect 3723 30640 3724 30680
rect 3764 30640 3765 30680
rect 3723 30631 3765 30640
rect 4195 30680 4253 30681
rect 4195 30640 4204 30680
rect 4244 30640 4253 30680
rect 4195 30639 4253 30640
rect 5443 30680 5501 30681
rect 5443 30640 5452 30680
rect 5492 30640 5501 30680
rect 5443 30639 5501 30640
rect 6019 30680 6077 30681
rect 6019 30640 6028 30680
rect 6068 30640 6077 30680
rect 6019 30639 6077 30640
rect 7267 30680 7325 30681
rect 7267 30640 7276 30680
rect 7316 30640 7325 30680
rect 7267 30639 7325 30640
rect 7467 30680 7509 30689
rect 7467 30640 7468 30680
rect 7508 30640 7509 30680
rect 7467 30631 7509 30640
rect 7563 30680 7605 30689
rect 7563 30640 7564 30680
rect 7604 30640 7605 30680
rect 7563 30631 7605 30640
rect 7659 30680 7701 30689
rect 7659 30640 7660 30680
rect 7700 30640 7701 30680
rect 7659 30631 7701 30640
rect 7755 30680 7797 30689
rect 7755 30640 7756 30680
rect 7796 30640 7797 30680
rect 7755 30631 7797 30640
rect 7939 30680 7997 30681
rect 7939 30640 7948 30680
rect 7988 30640 7997 30680
rect 7939 30639 7997 30640
rect 9187 30680 9245 30681
rect 9187 30640 9196 30680
rect 9236 30640 9245 30680
rect 9187 30639 9245 30640
rect 9571 30680 9629 30681
rect 9571 30640 9580 30680
rect 9620 30640 9629 30680
rect 9571 30639 9629 30640
rect 9667 30680 9725 30681
rect 9667 30640 9676 30680
rect 9716 30640 9725 30680
rect 9667 30639 9725 30640
rect 9867 30680 9909 30689
rect 9867 30640 9868 30680
rect 9908 30640 9909 30680
rect 9867 30631 9909 30640
rect 9963 30680 10005 30689
rect 9963 30640 9964 30680
rect 10004 30640 10005 30680
rect 9963 30631 10005 30640
rect 10056 30680 10114 30681
rect 10056 30640 10065 30680
rect 10105 30640 10114 30680
rect 10056 30639 10114 30640
rect 10435 30680 10493 30681
rect 10435 30640 10444 30680
rect 10484 30640 10493 30680
rect 10435 30639 10493 30640
rect 11683 30680 11741 30681
rect 11683 30640 11692 30680
rect 11732 30640 11741 30680
rect 11683 30639 11741 30640
rect 12171 30680 12213 30689
rect 12171 30640 12172 30680
rect 12212 30640 12213 30680
rect 12171 30631 12213 30640
rect 12267 30680 12309 30689
rect 12267 30640 12268 30680
rect 12308 30640 12309 30680
rect 12267 30631 12309 30640
rect 12651 30680 12693 30689
rect 12651 30640 12652 30680
rect 12692 30640 12693 30680
rect 12651 30631 12693 30640
rect 13219 30680 13277 30681
rect 13219 30640 13228 30680
rect 13268 30640 13277 30680
rect 13219 30639 13277 30640
rect 13755 30670 13797 30679
rect 13755 30630 13756 30670
rect 13796 30630 13797 30670
rect 14179 30651 14188 30691
rect 14228 30651 14237 30691
rect 14179 30650 14237 30651
rect 14667 30680 14709 30689
rect 14667 30640 14668 30680
rect 14708 30640 14709 30680
rect 14667 30631 14709 30640
rect 14859 30680 14901 30689
rect 14859 30640 14860 30680
rect 14900 30640 14901 30680
rect 14859 30631 14901 30640
rect 15051 30680 15093 30689
rect 15051 30640 15052 30680
rect 15092 30640 15093 30680
rect 15051 30631 15093 30640
rect 15427 30680 15485 30681
rect 15427 30640 15436 30680
rect 15476 30640 15485 30680
rect 15427 30639 15485 30640
rect 15723 30680 15765 30689
rect 15723 30640 15724 30680
rect 15764 30640 15765 30680
rect 15723 30631 15765 30640
rect 15819 30680 15861 30689
rect 15819 30640 15820 30680
rect 15860 30640 15861 30680
rect 15819 30631 15861 30640
rect 16771 30680 16829 30681
rect 16771 30640 16780 30680
rect 16820 30640 16829 30680
rect 17835 30680 17877 30689
rect 16771 30639 16829 30640
rect 17259 30666 17301 30675
rect 13755 30621 13797 30630
rect 17259 30626 17260 30666
rect 17300 30626 17301 30666
rect 17835 30640 17836 30680
rect 17876 30640 17877 30680
rect 17835 30631 17877 30640
rect 18115 30680 18173 30681
rect 18115 30640 18124 30680
rect 18164 30640 18173 30680
rect 18115 30639 18173 30640
rect 19363 30680 19421 30681
rect 19363 30640 19372 30680
rect 19412 30640 19421 30680
rect 19363 30639 19421 30640
rect 19747 30680 19805 30681
rect 19747 30640 19756 30680
rect 19796 30640 19805 30680
rect 19747 30639 19805 30640
rect 19851 30680 19893 30689
rect 19851 30640 19852 30680
rect 19892 30640 19893 30680
rect 19851 30631 19893 30640
rect 20035 30680 20093 30681
rect 20035 30640 20044 30680
rect 20084 30640 20093 30680
rect 20035 30639 20093 30640
rect 17259 30617 17301 30626
rect 12747 30596 12789 30605
rect 12747 30556 12748 30596
rect 12788 30556 12789 30596
rect 12747 30547 12789 30556
rect 15147 30596 15189 30605
rect 15147 30556 15148 30596
rect 15188 30556 15189 30596
rect 15147 30547 15189 30556
rect 15339 30596 15381 30605
rect 15339 30556 15340 30596
rect 15380 30556 15381 30596
rect 15339 30547 15381 30556
rect 16203 30596 16245 30605
rect 16203 30556 16204 30596
rect 16244 30556 16245 30596
rect 16203 30547 16245 30556
rect 16299 30596 16341 30605
rect 16299 30556 16300 30596
rect 16340 30556 16341 30596
rect 16299 30547 16341 30556
rect 15243 30512 15285 30521
rect 15243 30472 15244 30512
rect 15284 30472 15285 30512
rect 15243 30463 15285 30472
rect 17835 30512 17877 30521
rect 17835 30472 17836 30512
rect 17876 30472 17877 30512
rect 17835 30463 17877 30472
rect 3051 30428 3093 30437
rect 3051 30388 3052 30428
rect 3092 30388 3093 30428
rect 3051 30379 3093 30388
rect 4003 30428 4061 30429
rect 4003 30388 4012 30428
rect 4052 30388 4061 30428
rect 4003 30387 4061 30388
rect 5643 30428 5685 30437
rect 5643 30388 5644 30428
rect 5684 30388 5685 30428
rect 5643 30379 5685 30388
rect 14091 30428 14133 30437
rect 14091 30388 14092 30428
rect 14132 30388 14133 30428
rect 14091 30379 14133 30388
rect 14667 30428 14709 30437
rect 14667 30388 14668 30428
rect 14708 30388 14709 30428
rect 14667 30379 14709 30388
rect 1152 30260 20352 30284
rect 1152 30220 3688 30260
rect 3728 30220 3770 30260
rect 3810 30220 3852 30260
rect 3892 30220 3934 30260
rect 3974 30220 4016 30260
rect 4056 30220 18808 30260
rect 18848 30220 18890 30260
rect 18930 30220 18972 30260
rect 19012 30220 19054 30260
rect 19094 30220 19136 30260
rect 19176 30220 20352 30260
rect 1152 30196 20352 30220
rect 2859 30092 2901 30101
rect 2859 30052 2860 30092
rect 2900 30052 2901 30092
rect 2859 30043 2901 30052
rect 10827 30092 10869 30101
rect 10827 30052 10828 30092
rect 10868 30052 10869 30092
rect 10827 30043 10869 30052
rect 17259 30092 17301 30101
rect 17259 30052 17260 30092
rect 17300 30052 17301 30092
rect 17259 30043 17301 30052
rect 7363 30008 7421 30009
rect 7363 29968 7372 30008
rect 7412 29968 7421 30008
rect 7363 29967 7421 29968
rect 11019 30008 11061 30017
rect 11019 29968 11020 30008
rect 11060 29968 11061 30008
rect 11019 29959 11061 29968
rect 20227 30008 20285 30009
rect 20227 29968 20236 30008
rect 20276 29968 20285 30008
rect 20227 29967 20285 29968
rect 5739 29924 5781 29933
rect 5739 29884 5740 29924
rect 5780 29884 5781 29924
rect 5739 29875 5781 29884
rect 12171 29924 12213 29933
rect 12171 29884 12172 29924
rect 12212 29884 12213 29924
rect 12171 29875 12213 29884
rect 17547 29924 17589 29933
rect 17547 29884 17548 29924
rect 17588 29884 17589 29924
rect 17547 29875 17589 29884
rect 4779 29854 4821 29863
rect 1219 29840 1277 29841
rect 1219 29800 1228 29840
rect 1268 29800 1277 29840
rect 1219 29799 1277 29800
rect 2467 29840 2525 29841
rect 2467 29800 2476 29840
rect 2516 29800 2525 29840
rect 2467 29799 2525 29800
rect 3043 29840 3101 29841
rect 3043 29800 3052 29840
rect 3092 29800 3101 29840
rect 3043 29799 3101 29800
rect 4291 29840 4349 29841
rect 4291 29800 4300 29840
rect 4340 29800 4349 29840
rect 4779 29814 4780 29854
rect 4820 29814 4821 29854
rect 4779 29805 4821 29814
rect 5251 29840 5309 29841
rect 4291 29799 4349 29800
rect 5251 29800 5260 29840
rect 5300 29800 5309 29840
rect 5251 29799 5309 29800
rect 5835 29840 5877 29849
rect 5835 29800 5836 29840
rect 5876 29800 5877 29840
rect 5835 29791 5877 29800
rect 6219 29840 6261 29849
rect 6219 29800 6220 29840
rect 6260 29800 6261 29840
rect 6219 29791 6261 29800
rect 6315 29840 6357 29849
rect 6315 29800 6316 29840
rect 6356 29800 6357 29840
rect 6315 29791 6357 29800
rect 6691 29840 6749 29841
rect 6691 29800 6700 29840
rect 6740 29800 6749 29840
rect 6691 29799 6749 29800
rect 6987 29840 7029 29849
rect 6987 29800 6988 29840
rect 7028 29800 7029 29840
rect 6987 29791 7029 29800
rect 7555 29840 7613 29841
rect 7555 29800 7564 29840
rect 7604 29800 7613 29840
rect 7555 29799 7613 29800
rect 8803 29840 8861 29841
rect 8803 29800 8812 29840
rect 8852 29800 8861 29840
rect 8803 29799 8861 29800
rect 9387 29840 9429 29849
rect 9387 29800 9388 29840
rect 9428 29800 9429 29840
rect 9387 29791 9429 29800
rect 9483 29840 9525 29849
rect 9483 29800 9484 29840
rect 9524 29800 9525 29840
rect 9483 29791 9525 29800
rect 9579 29840 9621 29849
rect 9579 29800 9580 29840
rect 9620 29800 9621 29840
rect 9579 29791 9621 29800
rect 9859 29840 9917 29841
rect 9859 29800 9868 29840
rect 9908 29800 9917 29840
rect 9859 29799 9917 29800
rect 9963 29840 10005 29849
rect 9963 29800 9964 29840
rect 10004 29800 10005 29840
rect 9963 29791 10005 29800
rect 10155 29840 10197 29849
rect 10155 29800 10156 29840
rect 10196 29800 10197 29840
rect 10155 29791 10197 29800
rect 10347 29840 10389 29849
rect 10347 29800 10348 29840
rect 10388 29800 10389 29840
rect 10347 29791 10389 29800
rect 10443 29848 10485 29857
rect 13131 29854 13173 29863
rect 10443 29808 10444 29848
rect 10484 29808 10485 29848
rect 10443 29799 10485 29808
rect 10539 29840 10581 29849
rect 10539 29800 10540 29840
rect 10580 29800 10581 29840
rect 10539 29791 10581 29800
rect 11019 29840 11061 29849
rect 11019 29800 11020 29840
rect 11060 29800 11061 29840
rect 11019 29791 11061 29800
rect 11595 29840 11637 29849
rect 11595 29800 11596 29840
rect 11636 29800 11637 29840
rect 11595 29791 11637 29800
rect 11691 29840 11733 29849
rect 11691 29800 11692 29840
rect 11732 29800 11733 29840
rect 11691 29791 11733 29800
rect 12075 29840 12117 29849
rect 12075 29800 12076 29840
rect 12116 29800 12117 29840
rect 12075 29791 12117 29800
rect 12643 29840 12701 29841
rect 12643 29800 12652 29840
rect 12692 29800 12701 29840
rect 13131 29814 13132 29854
rect 13172 29814 13173 29854
rect 13131 29805 13173 29814
rect 13707 29840 13749 29849
rect 12643 29799 12701 29800
rect 13707 29800 13708 29840
rect 13748 29800 13749 29840
rect 13707 29791 13749 29800
rect 13803 29840 13845 29849
rect 13803 29800 13804 29840
rect 13844 29800 13845 29840
rect 13803 29791 13845 29800
rect 13899 29840 13941 29849
rect 13899 29800 13900 29840
rect 13940 29800 13941 29840
rect 13899 29791 13941 29800
rect 13995 29840 14037 29849
rect 13995 29800 13996 29840
rect 14036 29800 14037 29840
rect 13995 29791 14037 29800
rect 14179 29840 14237 29841
rect 14179 29800 14188 29840
rect 14228 29800 14237 29840
rect 14179 29799 14237 29800
rect 15427 29840 15485 29841
rect 15427 29800 15436 29840
rect 15476 29800 15485 29840
rect 15427 29799 15485 29800
rect 15811 29840 15869 29841
rect 15811 29800 15820 29840
rect 15860 29800 15869 29840
rect 15811 29799 15869 29800
rect 17059 29840 17117 29841
rect 17059 29800 17068 29840
rect 17108 29800 17117 29840
rect 17059 29799 17117 29800
rect 17451 29840 17493 29849
rect 17451 29800 17452 29840
rect 17492 29800 17493 29840
rect 17451 29791 17493 29800
rect 17643 29840 17685 29849
rect 17643 29800 17644 29840
rect 17684 29800 17685 29840
rect 17643 29791 17685 29800
rect 17827 29840 17885 29841
rect 17827 29800 17836 29840
rect 17876 29800 17885 29840
rect 17827 29799 17885 29800
rect 19075 29840 19133 29841
rect 19075 29800 19084 29840
rect 19124 29800 19133 29840
rect 19075 29799 19133 29800
rect 19555 29840 19613 29841
rect 19555 29800 19564 29840
rect 19604 29800 19613 29840
rect 19555 29799 19613 29800
rect 19851 29840 19893 29849
rect 19851 29800 19852 29840
rect 19892 29800 19893 29840
rect 19851 29791 19893 29800
rect 4587 29756 4629 29765
rect 4587 29716 4588 29756
rect 4628 29716 4629 29756
rect 4587 29707 4629 29716
rect 7083 29756 7125 29765
rect 7083 29716 7084 29756
rect 7124 29716 7125 29756
rect 7083 29707 7125 29716
rect 13323 29756 13365 29765
rect 13323 29716 13324 29756
rect 13364 29716 13365 29756
rect 13323 29707 13365 29716
rect 19275 29756 19317 29765
rect 19275 29716 19276 29756
rect 19316 29716 19317 29756
rect 19275 29707 19317 29716
rect 19947 29756 19989 29765
rect 19947 29716 19948 29756
rect 19988 29716 19989 29756
rect 19947 29707 19989 29716
rect 2667 29672 2709 29681
rect 2667 29632 2668 29672
rect 2708 29632 2709 29672
rect 2667 29623 2709 29632
rect 9003 29672 9045 29681
rect 9003 29632 9004 29672
rect 9044 29632 9045 29672
rect 9003 29623 9045 29632
rect 9667 29672 9725 29673
rect 9667 29632 9676 29672
rect 9716 29632 9725 29672
rect 9667 29631 9725 29632
rect 10051 29672 10109 29673
rect 10051 29632 10060 29672
rect 10100 29632 10109 29672
rect 10051 29631 10109 29632
rect 10627 29672 10685 29673
rect 10627 29632 10636 29672
rect 10676 29632 10685 29672
rect 10627 29631 10685 29632
rect 15627 29672 15669 29681
rect 15627 29632 15628 29672
rect 15668 29632 15669 29672
rect 15627 29623 15669 29632
rect 1152 29504 20452 29528
rect 1152 29464 4928 29504
rect 4968 29464 5010 29504
rect 5050 29464 5092 29504
rect 5132 29464 5174 29504
rect 5214 29464 5256 29504
rect 5296 29464 20048 29504
rect 20088 29464 20130 29504
rect 20170 29464 20212 29504
rect 20252 29464 20294 29504
rect 20334 29464 20376 29504
rect 20416 29464 20452 29504
rect 1152 29440 20452 29464
rect 3627 29336 3669 29345
rect 3627 29296 3628 29336
rect 3668 29296 3669 29336
rect 3627 29287 3669 29296
rect 8427 29336 8469 29345
rect 8427 29296 8428 29336
rect 8468 29296 8469 29336
rect 8427 29287 8469 29296
rect 8803 29336 8861 29337
rect 8803 29296 8812 29336
rect 8852 29296 8861 29336
rect 8803 29295 8861 29296
rect 9283 29336 9341 29337
rect 9283 29296 9292 29336
rect 9332 29296 9341 29336
rect 9283 29295 9341 29296
rect 15915 29252 15957 29261
rect 15915 29212 15916 29252
rect 15956 29212 15957 29252
rect 15915 29203 15957 29212
rect 1411 29168 1469 29169
rect 1411 29128 1420 29168
rect 1460 29128 1469 29168
rect 1411 29127 1469 29128
rect 1803 29168 1845 29177
rect 1803 29128 1804 29168
rect 1844 29128 1845 29168
rect 1803 29119 1845 29128
rect 1987 29168 2045 29169
rect 1987 29128 1996 29168
rect 2036 29128 2045 29168
rect 1987 29127 2045 29128
rect 3235 29168 3293 29169
rect 3235 29128 3244 29168
rect 3284 29128 3293 29168
rect 3235 29127 3293 29128
rect 3811 29168 3869 29169
rect 3811 29128 3820 29168
rect 3860 29128 3869 29168
rect 3811 29127 3869 29128
rect 5059 29168 5117 29169
rect 5059 29128 5068 29168
rect 5108 29128 5117 29168
rect 5059 29127 5117 29128
rect 5547 29168 5589 29177
rect 5547 29128 5548 29168
rect 5588 29128 5589 29168
rect 5547 29119 5589 29128
rect 5643 29168 5685 29177
rect 5643 29128 5644 29168
rect 5684 29128 5685 29168
rect 5643 29119 5685 29128
rect 5923 29168 5981 29169
rect 5923 29128 5932 29168
rect 5972 29128 5981 29168
rect 5923 29127 5981 29128
rect 6211 29168 6269 29169
rect 6211 29128 6220 29168
rect 6260 29128 6269 29168
rect 6211 29127 6269 29128
rect 6603 29168 6645 29177
rect 6603 29128 6604 29168
rect 6644 29128 6645 29168
rect 6603 29119 6645 29128
rect 6979 29168 7037 29169
rect 6979 29128 6988 29168
rect 7028 29128 7037 29168
rect 6979 29127 7037 29128
rect 8227 29168 8285 29169
rect 8227 29128 8236 29168
rect 8276 29128 8285 29168
rect 8227 29127 8285 29128
rect 8611 29168 8669 29169
rect 8611 29128 8620 29168
rect 8660 29128 8669 29168
rect 8611 29127 8669 29128
rect 8715 29168 8757 29177
rect 8715 29128 8716 29168
rect 8756 29128 8757 29168
rect 8715 29119 8757 29128
rect 8907 29168 8949 29177
rect 8907 29128 8908 29168
rect 8948 29128 8949 29168
rect 8907 29119 8949 29128
rect 9091 29168 9149 29169
rect 9091 29128 9100 29168
rect 9140 29128 9149 29168
rect 9091 29127 9149 29128
rect 9195 29168 9237 29177
rect 9195 29128 9196 29168
rect 9236 29128 9237 29168
rect 9195 29119 9237 29128
rect 9387 29168 9429 29177
rect 9387 29128 9388 29168
rect 9428 29128 9429 29168
rect 9387 29119 9429 29128
rect 9763 29168 9821 29169
rect 9763 29128 9772 29168
rect 9812 29128 9821 29168
rect 9763 29127 9821 29128
rect 11011 29168 11069 29169
rect 11011 29128 11020 29168
rect 11060 29128 11069 29168
rect 11011 29127 11069 29128
rect 11203 29168 11261 29169
rect 11203 29128 11212 29168
rect 11252 29128 11261 29168
rect 11203 29127 11261 29128
rect 12451 29168 12509 29169
rect 12451 29128 12460 29168
rect 12500 29128 12509 29168
rect 12451 29127 12509 29128
rect 12843 29168 12885 29177
rect 12843 29128 12844 29168
rect 12884 29128 12885 29168
rect 12843 29119 12885 29128
rect 13035 29168 13077 29177
rect 13035 29128 13036 29168
rect 13076 29128 13077 29168
rect 13035 29119 13077 29128
rect 13131 29168 13173 29177
rect 13131 29128 13132 29168
rect 13172 29128 13173 29168
rect 13131 29119 13173 29128
rect 13315 29168 13373 29169
rect 13315 29128 13324 29168
rect 13364 29128 13373 29168
rect 13315 29127 13373 29128
rect 13603 29168 13661 29169
rect 13603 29128 13612 29168
rect 13652 29128 13661 29168
rect 13603 29127 13661 29128
rect 14851 29168 14909 29169
rect 14851 29128 14860 29168
rect 14900 29128 14909 29168
rect 14851 29127 14909 29128
rect 15523 29168 15581 29169
rect 15523 29128 15532 29168
rect 15572 29128 15581 29168
rect 15523 29127 15581 29128
rect 15819 29168 15861 29177
rect 15819 29128 15820 29168
rect 15860 29128 15861 29168
rect 15819 29119 15861 29128
rect 16395 29168 16437 29177
rect 16395 29128 16396 29168
rect 16436 29128 16437 29168
rect 16395 29119 16437 29128
rect 16771 29168 16829 29169
rect 16771 29128 16780 29168
rect 16820 29128 16829 29168
rect 16771 29127 16829 29128
rect 17059 29168 17117 29169
rect 17059 29128 17068 29168
rect 17108 29128 17117 29168
rect 17059 29127 17117 29128
rect 18307 29168 18365 29169
rect 18307 29128 18316 29168
rect 18356 29128 18365 29168
rect 18307 29127 18365 29128
rect 19171 29168 19229 29169
rect 19171 29128 19180 29168
rect 19220 29128 19229 29168
rect 19171 29127 19229 29128
rect 1515 29084 1557 29093
rect 1515 29044 1516 29084
rect 1556 29044 1557 29084
rect 1515 29035 1557 29044
rect 1707 29084 1749 29093
rect 1707 29044 1708 29084
rect 1748 29044 1749 29084
rect 1707 29035 1749 29044
rect 16491 29084 16533 29093
rect 16491 29044 16492 29084
rect 16532 29044 16533 29084
rect 16491 29035 16533 29044
rect 16683 29084 16725 29093
rect 16683 29044 16684 29084
rect 16724 29044 16725 29084
rect 16683 29035 16725 29044
rect 18691 29084 18749 29085
rect 18691 29044 18700 29084
rect 18740 29044 18749 29084
rect 18691 29043 18749 29044
rect 1611 29000 1653 29009
rect 1611 28960 1612 29000
rect 1652 28960 1653 29000
rect 1611 28951 1653 28960
rect 6603 29000 6645 29009
rect 6603 28960 6604 29000
rect 6644 28960 6645 29000
rect 6603 28951 6645 28960
rect 9579 29000 9621 29009
rect 9579 28960 9580 29000
rect 9620 28960 9621 29000
rect 9579 28951 9621 28960
rect 13027 29000 13085 29001
rect 13027 28960 13036 29000
rect 13076 28960 13085 29000
rect 13027 28959 13085 28960
rect 16587 29000 16629 29009
rect 16587 28960 16588 29000
rect 16628 28960 16629 29000
rect 16587 28951 16629 28960
rect 18507 29000 18549 29009
rect 18507 28960 18508 29000
rect 18548 28960 18549 29000
rect 18507 28951 18549 28960
rect 18891 29000 18933 29009
rect 18891 28960 18892 29000
rect 18932 28960 18933 29000
rect 18891 28951 18933 28960
rect 19851 29000 19893 29009
rect 19851 28960 19852 29000
rect 19892 28960 19893 29000
rect 19851 28951 19893 28960
rect 3435 28916 3477 28925
rect 3435 28876 3436 28916
rect 3476 28876 3477 28916
rect 3435 28867 3477 28876
rect 5251 28916 5309 28917
rect 5251 28876 5260 28916
rect 5300 28876 5309 28916
rect 5251 28875 5309 28876
rect 6315 28916 6357 28925
rect 6315 28876 6316 28916
rect 6356 28876 6357 28916
rect 6315 28867 6357 28876
rect 6795 28916 6837 28925
rect 6795 28876 6796 28916
rect 6836 28876 6837 28916
rect 6795 28867 6837 28876
rect 12651 28916 12693 28925
rect 12651 28876 12652 28916
rect 12692 28876 12693 28916
rect 12651 28867 12693 28876
rect 13419 28916 13461 28925
rect 13419 28876 13420 28916
rect 13460 28876 13461 28916
rect 13419 28867 13461 28876
rect 15051 28916 15093 28925
rect 15051 28876 15052 28916
rect 15092 28876 15093 28916
rect 15051 28867 15093 28876
rect 16195 28916 16253 28917
rect 16195 28876 16204 28916
rect 16244 28876 16253 28916
rect 16195 28875 16253 28876
rect 1152 28748 20352 28772
rect 1152 28708 3688 28748
rect 3728 28708 3770 28748
rect 3810 28708 3852 28748
rect 3892 28708 3934 28748
rect 3974 28708 4016 28748
rect 4056 28708 18808 28748
rect 18848 28708 18890 28748
rect 18930 28708 18972 28748
rect 19012 28708 19054 28748
rect 19094 28708 19136 28748
rect 19176 28708 20352 28748
rect 1152 28684 20352 28708
rect 9763 28580 9821 28581
rect 9763 28540 9772 28580
rect 9812 28540 9821 28580
rect 9763 28539 9821 28540
rect 10731 28580 10773 28589
rect 10731 28540 10732 28580
rect 10772 28540 10773 28580
rect 10731 28531 10773 28540
rect 12843 28580 12885 28589
rect 12843 28540 12844 28580
rect 12884 28540 12885 28580
rect 12843 28531 12885 28540
rect 15435 28580 15477 28589
rect 15435 28540 15436 28580
rect 15476 28540 15477 28580
rect 15435 28531 15477 28540
rect 4107 28496 4149 28505
rect 4107 28456 4108 28496
rect 4148 28456 4149 28496
rect 4107 28447 4149 28456
rect 5931 28496 5973 28505
rect 5931 28456 5932 28496
rect 5972 28456 5973 28496
rect 5931 28447 5973 28456
rect 6411 28496 6453 28505
rect 6411 28456 6412 28496
rect 6452 28456 6453 28496
rect 6411 28447 6453 28456
rect 2571 28412 2613 28421
rect 2571 28372 2572 28412
rect 2612 28372 2613 28412
rect 2571 28363 2613 28372
rect 4011 28412 4053 28421
rect 4011 28372 4012 28412
rect 4052 28372 4053 28412
rect 4011 28363 4053 28372
rect 4203 28412 4245 28421
rect 4203 28372 4204 28412
rect 4244 28372 4245 28412
rect 4203 28363 4245 28372
rect 6315 28412 6357 28421
rect 6315 28372 6316 28412
rect 6356 28372 6357 28412
rect 6315 28363 6357 28372
rect 6507 28412 6549 28421
rect 6507 28372 6508 28412
rect 6548 28372 6549 28412
rect 6507 28363 6549 28372
rect 19843 28412 19901 28413
rect 19843 28372 19852 28412
rect 19892 28372 19901 28412
rect 19843 28371 19901 28372
rect 3531 28342 3573 28351
rect 1995 28328 2037 28337
rect 1995 28288 1996 28328
rect 2036 28288 2037 28328
rect 1995 28279 2037 28288
rect 2091 28328 2133 28337
rect 2091 28288 2092 28328
rect 2132 28288 2133 28328
rect 2091 28279 2133 28288
rect 2475 28328 2517 28337
rect 2475 28288 2476 28328
rect 2516 28288 2517 28328
rect 2475 28279 2517 28288
rect 3043 28328 3101 28329
rect 3043 28288 3052 28328
rect 3092 28288 3101 28328
rect 3531 28302 3532 28342
rect 3572 28302 3573 28342
rect 10923 28341 10965 28350
rect 3531 28293 3573 28302
rect 3915 28328 3957 28337
rect 3043 28287 3101 28288
rect 3915 28288 3916 28328
rect 3956 28288 3957 28328
rect 3915 28279 3957 28288
rect 4291 28328 4349 28329
rect 4291 28288 4300 28328
rect 4340 28288 4349 28328
rect 4291 28287 4349 28288
rect 4483 28328 4541 28329
rect 4483 28288 4492 28328
rect 4532 28288 4541 28328
rect 4483 28287 4541 28288
rect 5731 28328 5789 28329
rect 5731 28288 5740 28328
rect 5780 28288 5789 28328
rect 5731 28287 5789 28288
rect 6211 28328 6269 28329
rect 6211 28288 6220 28328
rect 6260 28288 6269 28328
rect 6211 28287 6269 28288
rect 6603 28328 6645 28337
rect 6603 28288 6604 28328
rect 6644 28288 6645 28328
rect 6603 28279 6645 28288
rect 6883 28328 6941 28329
rect 6883 28288 6892 28328
rect 6932 28288 6941 28328
rect 6883 28287 6941 28288
rect 8131 28328 8189 28329
rect 8131 28288 8140 28328
rect 8180 28288 8189 28328
rect 8131 28287 8189 28288
rect 8619 28328 8661 28337
rect 8619 28288 8620 28328
rect 8660 28288 8661 28328
rect 8619 28279 8661 28288
rect 8715 28328 8757 28337
rect 8715 28288 8716 28328
rect 8756 28288 8757 28328
rect 8715 28279 8757 28288
rect 8811 28328 8853 28337
rect 8811 28288 8812 28328
rect 8852 28288 8853 28328
rect 8811 28279 8853 28288
rect 9091 28328 9149 28329
rect 9091 28288 9100 28328
rect 9140 28288 9149 28328
rect 9091 28287 9149 28288
rect 9387 28328 9429 28337
rect 9387 28288 9388 28328
rect 9428 28288 9429 28328
rect 9387 28279 9429 28288
rect 9483 28328 9525 28337
rect 9483 28288 9484 28328
rect 9524 28288 9525 28328
rect 9483 28279 9525 28288
rect 9963 28328 10005 28337
rect 9963 28288 9964 28328
rect 10004 28288 10005 28328
rect 9963 28279 10005 28288
rect 10059 28328 10101 28337
rect 10059 28288 10060 28328
rect 10100 28288 10101 28328
rect 10059 28279 10101 28288
rect 10155 28328 10197 28337
rect 10155 28288 10156 28328
rect 10196 28288 10197 28328
rect 10155 28279 10197 28288
rect 10251 28328 10293 28337
rect 10251 28288 10252 28328
rect 10292 28288 10293 28328
rect 10251 28279 10293 28288
rect 10435 28328 10493 28329
rect 10435 28288 10444 28328
rect 10484 28288 10493 28328
rect 10435 28287 10493 28288
rect 10539 28328 10581 28337
rect 10539 28288 10540 28328
rect 10580 28288 10581 28328
rect 10539 28279 10581 28288
rect 10731 28328 10773 28337
rect 10731 28288 10732 28328
rect 10772 28288 10773 28328
rect 10923 28301 10924 28341
rect 10964 28301 10965 28341
rect 15976 28343 16018 28352
rect 10923 28292 10965 28301
rect 11115 28328 11157 28337
rect 10731 28279 10773 28288
rect 11115 28288 11116 28328
rect 11156 28288 11157 28328
rect 11115 28279 11157 28288
rect 11395 28328 11453 28329
rect 11395 28288 11404 28328
rect 11444 28288 11453 28328
rect 11395 28287 11453 28288
rect 12643 28328 12701 28329
rect 12643 28288 12652 28328
rect 12692 28288 12701 28328
rect 12643 28287 12701 28288
rect 13027 28328 13085 28329
rect 13027 28288 13036 28328
rect 13076 28288 13085 28328
rect 13027 28287 13085 28288
rect 13123 28328 13181 28329
rect 13123 28288 13132 28328
rect 13172 28288 13181 28328
rect 13123 28287 13181 28288
rect 13323 28328 13365 28337
rect 13323 28288 13324 28328
rect 13364 28288 13365 28328
rect 13323 28279 13365 28288
rect 13419 28328 13461 28337
rect 13419 28288 13420 28328
rect 13460 28288 13461 28328
rect 13419 28279 13461 28288
rect 13512 28328 13570 28329
rect 13512 28288 13521 28328
rect 13561 28288 13570 28328
rect 13512 28287 13570 28288
rect 13987 28328 14045 28329
rect 13987 28288 13996 28328
rect 14036 28288 14045 28328
rect 13987 28287 14045 28288
rect 15235 28328 15293 28329
rect 15235 28288 15244 28328
rect 15284 28288 15293 28328
rect 15235 28287 15293 28288
rect 15427 28328 15485 28329
rect 15427 28288 15436 28328
rect 15476 28288 15485 28328
rect 15427 28287 15485 28288
rect 15523 28328 15581 28329
rect 15523 28288 15532 28328
rect 15572 28288 15581 28328
rect 15523 28287 15581 28288
rect 15723 28328 15765 28337
rect 15723 28288 15724 28328
rect 15764 28288 15765 28328
rect 15723 28279 15765 28288
rect 15819 28328 15861 28337
rect 15819 28288 15820 28328
rect 15860 28288 15861 28328
rect 15976 28303 15977 28343
rect 16017 28303 16018 28343
rect 15976 28294 16018 28303
rect 16195 28328 16253 28329
rect 15819 28279 15861 28288
rect 16195 28288 16204 28328
rect 16244 28288 16253 28328
rect 16195 28287 16253 28288
rect 17443 28328 17501 28329
rect 17443 28288 17452 28328
rect 17492 28288 17501 28328
rect 17443 28287 17501 28288
rect 17931 28328 17973 28337
rect 17931 28288 17932 28328
rect 17972 28288 17973 28328
rect 17931 28279 17973 28288
rect 18027 28328 18069 28337
rect 18027 28288 18028 28328
rect 18068 28288 18069 28328
rect 18027 28279 18069 28288
rect 18411 28328 18453 28337
rect 18411 28288 18412 28328
rect 18452 28288 18453 28328
rect 18411 28279 18453 28288
rect 18507 28328 18549 28337
rect 19467 28333 19509 28342
rect 18507 28288 18508 28328
rect 18548 28288 18549 28328
rect 18507 28279 18549 28288
rect 18979 28328 19037 28329
rect 18979 28288 18988 28328
rect 19028 28288 19037 28328
rect 18979 28287 19037 28288
rect 19467 28293 19468 28333
rect 19508 28293 19509 28333
rect 19467 28284 19509 28293
rect 3723 28244 3765 28253
rect 3723 28204 3724 28244
rect 3764 28204 3765 28244
rect 3723 28195 3765 28204
rect 8523 28244 8565 28253
rect 8523 28204 8524 28244
rect 8564 28204 8565 28244
rect 8523 28195 8565 28204
rect 19659 28244 19701 28253
rect 19659 28204 19660 28244
rect 19700 28204 19701 28244
rect 19659 28195 19701 28204
rect 1315 28160 1373 28161
rect 1315 28120 1324 28160
rect 1364 28120 1373 28160
rect 1315 28119 1373 28120
rect 1603 28160 1661 28161
rect 1603 28120 1612 28160
rect 1652 28120 1661 28160
rect 1603 28119 1661 28120
rect 8331 28160 8373 28169
rect 8331 28120 8332 28160
rect 8372 28120 8373 28160
rect 8331 28111 8373 28120
rect 11019 28160 11061 28169
rect 11019 28120 11020 28160
rect 11060 28120 11061 28160
rect 11019 28111 11061 28120
rect 13411 28160 13469 28161
rect 13411 28120 13420 28160
rect 13460 28120 13469 28160
rect 13411 28119 13469 28120
rect 13803 28160 13845 28169
rect 13803 28120 13804 28160
rect 13844 28120 13845 28160
rect 13803 28111 13845 28120
rect 17643 28160 17685 28169
rect 17643 28120 17644 28160
rect 17684 28120 17685 28160
rect 17643 28111 17685 28120
rect 20043 28160 20085 28169
rect 20043 28120 20044 28160
rect 20084 28120 20085 28160
rect 20043 28111 20085 28120
rect 1152 27992 20452 28016
rect 1152 27952 4928 27992
rect 4968 27952 5010 27992
rect 5050 27952 5092 27992
rect 5132 27952 5174 27992
rect 5214 27952 5256 27992
rect 5296 27952 20048 27992
rect 20088 27952 20130 27992
rect 20170 27952 20212 27992
rect 20252 27952 20294 27992
rect 20334 27952 20376 27992
rect 20416 27952 20452 27992
rect 1152 27928 20452 27952
rect 9667 27824 9725 27825
rect 9667 27784 9676 27824
rect 9716 27784 9725 27824
rect 9667 27783 9725 27784
rect 9867 27824 9909 27833
rect 9867 27784 9868 27824
rect 9908 27784 9909 27824
rect 9867 27775 9909 27784
rect 13795 27824 13853 27825
rect 13795 27784 13804 27824
rect 13844 27784 13853 27824
rect 13795 27783 13853 27784
rect 14859 27824 14901 27833
rect 14859 27784 14860 27824
rect 14900 27784 14901 27824
rect 14859 27775 14901 27784
rect 3147 27740 3189 27749
rect 3147 27700 3148 27740
rect 3188 27700 3189 27740
rect 3147 27691 3189 27700
rect 7851 27740 7893 27749
rect 7851 27700 7852 27740
rect 7892 27700 7893 27740
rect 7851 27691 7893 27700
rect 19563 27740 19605 27749
rect 19563 27700 19564 27740
rect 19604 27700 19605 27740
rect 19563 27691 19605 27700
rect 1219 27656 1277 27657
rect 1219 27616 1228 27656
rect 1268 27616 1277 27656
rect 1219 27615 1277 27616
rect 2467 27656 2525 27657
rect 2467 27616 2476 27656
rect 2516 27616 2525 27656
rect 2467 27615 2525 27616
rect 3243 27656 3285 27665
rect 3243 27616 3244 27656
rect 3284 27616 3285 27656
rect 3243 27607 3285 27616
rect 3523 27656 3581 27657
rect 3523 27616 3532 27656
rect 3572 27616 3581 27656
rect 3523 27615 3581 27616
rect 3811 27656 3869 27657
rect 3811 27616 3820 27656
rect 3860 27616 3869 27656
rect 3811 27615 3869 27616
rect 3915 27656 3957 27665
rect 3915 27616 3916 27656
rect 3956 27616 3957 27656
rect 3915 27607 3957 27616
rect 4099 27656 4157 27657
rect 4099 27616 4108 27656
rect 4148 27616 4157 27656
rect 4099 27615 4157 27616
rect 4291 27656 4349 27657
rect 4291 27616 4300 27656
rect 4340 27616 4349 27656
rect 4291 27615 4349 27616
rect 5539 27656 5597 27657
rect 5539 27616 5548 27656
rect 5588 27616 5597 27656
rect 5539 27615 5597 27616
rect 6115 27656 6173 27657
rect 6115 27616 6124 27656
rect 6164 27616 6173 27656
rect 6115 27615 6173 27616
rect 7363 27656 7421 27657
rect 7363 27616 7372 27656
rect 7412 27616 7421 27656
rect 7363 27615 7421 27616
rect 7755 27656 7797 27665
rect 7755 27616 7756 27656
rect 7796 27616 7797 27656
rect 7755 27607 7797 27616
rect 7947 27656 7989 27665
rect 7947 27616 7948 27656
rect 7988 27616 7989 27656
rect 7947 27607 7989 27616
rect 8035 27656 8093 27657
rect 8035 27616 8044 27656
rect 8084 27616 8093 27656
rect 8035 27615 8093 27616
rect 8227 27656 8285 27657
rect 8227 27616 8236 27656
rect 8276 27616 8285 27656
rect 8227 27615 8285 27616
rect 8331 27656 8373 27665
rect 8331 27616 8332 27656
rect 8372 27616 8373 27656
rect 8331 27607 8373 27616
rect 8523 27656 8565 27665
rect 8523 27616 8524 27656
rect 8564 27616 8565 27656
rect 8523 27607 8565 27616
rect 8811 27656 8853 27665
rect 8811 27616 8812 27656
rect 8852 27616 8853 27656
rect 8811 27607 8853 27616
rect 8907 27656 8949 27665
rect 8907 27616 8908 27656
rect 8948 27616 8949 27656
rect 8907 27607 8949 27616
rect 9003 27656 9045 27665
rect 9003 27616 9004 27656
rect 9044 27616 9045 27656
rect 9003 27607 9045 27616
rect 9387 27656 9429 27665
rect 9387 27616 9388 27656
rect 9428 27616 9429 27656
rect 9387 27607 9429 27616
rect 9483 27656 9525 27665
rect 9483 27616 9484 27656
rect 9524 27616 9525 27656
rect 9483 27607 9525 27616
rect 9955 27656 10013 27657
rect 9955 27616 9964 27656
rect 10004 27616 10013 27656
rect 9955 27615 10013 27616
rect 10147 27656 10205 27657
rect 10147 27616 10156 27656
rect 10196 27616 10205 27656
rect 10147 27615 10205 27616
rect 11395 27656 11453 27657
rect 11395 27616 11404 27656
rect 11444 27616 11453 27656
rect 11395 27615 11453 27616
rect 11875 27656 11933 27657
rect 11875 27616 11884 27656
rect 11924 27616 11933 27656
rect 11875 27615 11933 27616
rect 13123 27656 13181 27657
rect 13123 27616 13132 27656
rect 13172 27616 13181 27656
rect 13123 27615 13181 27616
rect 13515 27656 13557 27665
rect 13515 27616 13516 27656
rect 13556 27616 13557 27656
rect 13515 27607 13557 27616
rect 13611 27656 13653 27665
rect 13611 27616 13612 27656
rect 13652 27616 13653 27656
rect 13611 27607 13653 27616
rect 14563 27656 14621 27657
rect 14563 27616 14572 27656
rect 14612 27616 14621 27656
rect 14563 27615 14621 27616
rect 14667 27656 14709 27665
rect 14667 27616 14668 27656
rect 14708 27616 14709 27656
rect 14667 27607 14709 27616
rect 14851 27656 14909 27657
rect 14851 27616 14860 27656
rect 14900 27616 14909 27656
rect 15435 27656 15477 27665
rect 14851 27615 14909 27616
rect 15139 27639 15197 27640
rect 15139 27599 15148 27639
rect 15188 27599 15197 27639
rect 15435 27616 15436 27656
rect 15476 27616 15477 27656
rect 15435 27607 15477 27616
rect 15531 27656 15573 27665
rect 15531 27616 15532 27656
rect 15572 27616 15573 27656
rect 15531 27607 15573 27616
rect 16003 27656 16061 27657
rect 16003 27616 16012 27656
rect 16052 27616 16061 27656
rect 16003 27615 16061 27616
rect 16395 27656 16437 27665
rect 16395 27616 16396 27656
rect 16436 27616 16437 27656
rect 16395 27607 16437 27616
rect 16587 27656 16629 27665
rect 16587 27616 16588 27656
rect 16628 27616 16629 27656
rect 16587 27607 16629 27616
rect 16779 27656 16821 27665
rect 16779 27616 16780 27656
rect 16820 27616 16821 27656
rect 16779 27607 16821 27616
rect 17835 27656 17877 27665
rect 17835 27616 17836 27656
rect 17876 27616 17877 27656
rect 17835 27607 17877 27616
rect 17931 27656 17973 27665
rect 17931 27616 17932 27656
rect 17972 27616 17973 27656
rect 17931 27607 17973 27616
rect 18883 27656 18941 27657
rect 18883 27616 18892 27656
rect 18932 27616 18941 27656
rect 18883 27615 18941 27616
rect 19371 27651 19413 27660
rect 19371 27611 19372 27651
rect 19412 27611 19413 27651
rect 19371 27602 19413 27611
rect 20126 27643 20168 27652
rect 20126 27603 20127 27643
rect 20167 27603 20168 27643
rect 15139 27598 15197 27599
rect 20126 27594 20168 27603
rect 14179 27572 14237 27573
rect 14179 27532 14188 27572
rect 14228 27532 14237 27572
rect 14179 27531 14237 27532
rect 16107 27572 16149 27581
rect 16107 27532 16108 27572
rect 16148 27532 16149 27572
rect 16107 27523 16149 27532
rect 16299 27572 16341 27581
rect 16299 27532 16300 27572
rect 16340 27532 16341 27572
rect 16299 27523 16341 27532
rect 16963 27572 17021 27573
rect 16963 27532 16972 27572
rect 17012 27532 17021 27572
rect 16963 27531 17021 27532
rect 17347 27572 17405 27573
rect 17347 27532 17356 27572
rect 17396 27532 17405 27572
rect 17347 27531 17405 27532
rect 18315 27572 18357 27581
rect 18315 27532 18316 27572
rect 18356 27532 18357 27572
rect 18315 27523 18357 27532
rect 18411 27572 18453 27581
rect 18411 27532 18412 27572
rect 18452 27532 18453 27572
rect 18411 27523 18453 27532
rect 19747 27572 19805 27573
rect 19747 27532 19756 27572
rect 19796 27532 19805 27572
rect 19747 27531 19805 27532
rect 2667 27488 2709 27497
rect 2667 27448 2668 27488
rect 2708 27448 2709 27488
rect 2667 27439 2709 27448
rect 8523 27488 8565 27497
rect 8523 27448 8524 27488
rect 8564 27448 8565 27488
rect 8523 27439 8565 27448
rect 15811 27488 15869 27489
rect 15811 27448 15820 27488
rect 15860 27448 15869 27488
rect 15811 27447 15869 27448
rect 16203 27488 16245 27497
rect 16203 27448 16204 27488
rect 16244 27448 16245 27488
rect 16203 27439 16245 27448
rect 16587 27488 16629 27497
rect 16587 27448 16588 27488
rect 16628 27448 16629 27488
rect 16587 27439 16629 27448
rect 17163 27488 17205 27497
rect 17163 27448 17164 27488
rect 17204 27448 17205 27488
rect 17163 27439 17205 27448
rect 17547 27488 17589 27497
rect 17547 27448 17548 27488
rect 17588 27448 17589 27488
rect 17547 27439 17589 27448
rect 2851 27404 2909 27405
rect 2851 27364 2860 27404
rect 2900 27364 2909 27404
rect 2851 27363 2909 27364
rect 4107 27404 4149 27413
rect 4107 27364 4108 27404
rect 4148 27364 4149 27404
rect 4107 27355 4149 27364
rect 5739 27404 5781 27413
rect 5739 27364 5740 27404
rect 5780 27364 5781 27404
rect 5739 27355 5781 27364
rect 7563 27404 7605 27413
rect 7563 27364 7564 27404
rect 7604 27364 7605 27404
rect 7563 27355 7605 27364
rect 9187 27404 9245 27405
rect 9187 27364 9196 27404
rect 9236 27364 9245 27404
rect 9187 27363 9245 27364
rect 11595 27404 11637 27413
rect 11595 27364 11596 27404
rect 11636 27364 11637 27404
rect 11595 27355 11637 27364
rect 13323 27404 13365 27413
rect 13323 27364 13324 27404
rect 13364 27364 13365 27404
rect 13323 27355 13365 27364
rect 13995 27404 14037 27413
rect 13995 27364 13996 27404
rect 14036 27364 14037 27404
rect 13995 27355 14037 27364
rect 19947 27404 19989 27413
rect 19947 27364 19948 27404
rect 19988 27364 19989 27404
rect 19947 27355 19989 27364
rect 20235 27404 20277 27413
rect 20235 27364 20236 27404
rect 20276 27364 20277 27404
rect 20235 27355 20277 27364
rect 1152 27236 20352 27260
rect 1152 27196 3688 27236
rect 3728 27196 3770 27236
rect 3810 27196 3852 27236
rect 3892 27196 3934 27236
rect 3974 27196 4016 27236
rect 4056 27196 18808 27236
rect 18848 27196 18890 27236
rect 18930 27196 18972 27236
rect 19012 27196 19054 27236
rect 19094 27196 19136 27236
rect 19176 27196 20352 27236
rect 1152 27172 20352 27196
rect 2667 27068 2709 27077
rect 2667 27028 2668 27068
rect 2708 27028 2709 27068
rect 2667 27019 2709 27028
rect 8811 27068 8853 27077
rect 8811 27028 8812 27068
rect 8852 27028 8853 27068
rect 8811 27019 8853 27028
rect 13707 27068 13749 27077
rect 13707 27028 13708 27068
rect 13748 27028 13749 27068
rect 13707 27019 13749 27028
rect 17739 27068 17781 27077
rect 17739 27028 17740 27068
rect 17780 27028 17781 27068
rect 17739 27019 17781 27028
rect 18123 27068 18165 27077
rect 18123 27028 18124 27068
rect 18164 27028 18165 27068
rect 18123 27019 18165 27028
rect 3811 26984 3869 26985
rect 3811 26944 3820 26984
rect 3860 26944 3869 26984
rect 3811 26943 3869 26944
rect 4203 26984 4245 26993
rect 4203 26944 4204 26984
rect 4244 26944 4245 26984
rect 4203 26935 4245 26944
rect 6315 26984 6357 26993
rect 6315 26944 6316 26984
rect 6356 26944 6357 26984
rect 6315 26935 6357 26944
rect 9283 26984 9341 26985
rect 9283 26944 9292 26984
rect 9332 26944 9341 26984
rect 9283 26943 9341 26944
rect 11403 26984 11445 26993
rect 11403 26944 11404 26984
rect 11444 26944 11445 26984
rect 11403 26935 11445 26944
rect 13995 26984 14037 26993
rect 13995 26944 13996 26984
rect 14036 26944 14037 26984
rect 13995 26935 14037 26944
rect 16395 26984 16437 26993
rect 16395 26944 16396 26984
rect 16436 26944 16437 26984
rect 16395 26935 16437 26944
rect 18507 26984 18549 26993
rect 18507 26944 18508 26984
rect 18548 26944 18549 26984
rect 18507 26935 18549 26944
rect 18307 26911 18365 26912
rect 6229 26900 6271 26909
rect 6229 26860 6230 26900
rect 6270 26860 6271 26900
rect 6229 26851 6271 26860
rect 6411 26900 6453 26909
rect 6411 26860 6412 26900
rect 6452 26860 6453 26900
rect 6411 26851 6453 26860
rect 12171 26900 12213 26909
rect 12171 26860 12172 26900
rect 12212 26860 12213 26900
rect 12171 26851 12213 26860
rect 14283 26900 14325 26909
rect 14283 26860 14284 26900
rect 14324 26860 14325 26900
rect 14283 26851 14325 26860
rect 16299 26900 16341 26909
rect 16299 26860 16300 26900
rect 16340 26860 16341 26900
rect 16299 26851 16341 26860
rect 16491 26900 16533 26909
rect 16491 26860 16492 26900
rect 16532 26860 16533 26900
rect 16491 26851 16533 26860
rect 17539 26900 17597 26901
rect 17539 26860 17548 26900
rect 17588 26860 17597 26900
rect 17539 26859 17597 26860
rect 17923 26900 17981 26901
rect 17923 26860 17932 26900
rect 17972 26860 17981 26900
rect 18307 26871 18316 26911
rect 18356 26871 18365 26911
rect 18307 26870 18365 26871
rect 19555 26900 19613 26901
rect 17923 26859 17981 26860
rect 19555 26860 19564 26900
rect 19604 26860 19613 26900
rect 19555 26859 19613 26860
rect 19939 26900 19997 26901
rect 19939 26860 19948 26900
rect 19988 26860 19997 26900
rect 19939 26859 19997 26860
rect 16771 26858 16829 26859
rect 8331 26830 8373 26839
rect 1219 26816 1277 26817
rect 1219 26776 1228 26816
rect 1268 26776 1277 26816
rect 1219 26775 1277 26776
rect 2467 26816 2525 26817
rect 2467 26776 2476 26816
rect 2516 26776 2525 26816
rect 2467 26775 2525 26776
rect 3139 26816 3197 26817
rect 3139 26776 3148 26816
rect 3188 26776 3197 26816
rect 3139 26775 3197 26776
rect 3435 26816 3477 26825
rect 3435 26776 3436 26816
rect 3476 26776 3477 26816
rect 3435 26767 3477 26776
rect 4011 26816 4053 26825
rect 4011 26776 4012 26816
rect 4052 26776 4053 26816
rect 4011 26767 4053 26776
rect 4203 26816 4245 26825
rect 4203 26776 4204 26816
rect 4244 26776 4245 26816
rect 4203 26767 4245 26776
rect 4387 26816 4445 26817
rect 4387 26776 4396 26816
rect 4436 26776 4445 26816
rect 4387 26775 4445 26776
rect 5635 26816 5693 26817
rect 5635 26776 5644 26816
rect 5684 26776 5693 26816
rect 5635 26775 5693 26776
rect 6115 26816 6173 26817
rect 6115 26776 6124 26816
rect 6164 26776 6173 26816
rect 6115 26775 6173 26776
rect 6507 26816 6549 26825
rect 6507 26776 6508 26816
rect 6548 26776 6549 26816
rect 6507 26767 6549 26776
rect 6795 26816 6837 26825
rect 6795 26776 6796 26816
rect 6836 26776 6837 26816
rect 6795 26767 6837 26776
rect 6891 26816 6933 26825
rect 6891 26776 6892 26816
rect 6932 26776 6933 26816
rect 6891 26767 6933 26776
rect 7275 26816 7317 26825
rect 7275 26776 7276 26816
rect 7316 26776 7317 26816
rect 7275 26767 7317 26776
rect 7371 26816 7413 26825
rect 7371 26776 7372 26816
rect 7412 26776 7413 26816
rect 7371 26767 7413 26776
rect 7843 26816 7901 26817
rect 7843 26776 7852 26816
rect 7892 26776 7901 26816
rect 8331 26790 8332 26830
rect 8372 26790 8373 26830
rect 11691 26835 11733 26844
rect 8331 26781 8373 26790
rect 8707 26816 8765 26817
rect 7843 26775 7901 26776
rect 8707 26776 8716 26816
rect 8756 26776 8765 26816
rect 8707 26775 8765 26776
rect 9091 26816 9149 26817
rect 9091 26776 9100 26816
rect 9140 26776 9149 26816
rect 9091 26775 9149 26776
rect 9483 26816 9525 26825
rect 9483 26776 9484 26816
rect 9524 26776 9525 26816
rect 9483 26767 9525 26776
rect 9675 26816 9717 26825
rect 9675 26776 9676 26816
rect 9716 26776 9717 26816
rect 9675 26767 9717 26776
rect 9763 26816 9821 26817
rect 9763 26776 9772 26816
rect 9812 26776 9821 26816
rect 9763 26775 9821 26776
rect 9955 26816 10013 26817
rect 9955 26776 9964 26816
rect 10004 26776 10013 26816
rect 9955 26775 10013 26776
rect 11203 26816 11261 26817
rect 11203 26776 11212 26816
rect 11252 26776 11261 26816
rect 11691 26795 11692 26835
rect 11732 26795 11733 26835
rect 13275 26825 13317 26834
rect 12267 26816 12309 26825
rect 11691 26786 11733 26795
rect 11787 26796 11829 26805
rect 11203 26775 11261 26776
rect 11787 26756 11788 26796
rect 11828 26756 11829 26796
rect 12267 26776 12268 26816
rect 12308 26776 12309 26816
rect 12267 26767 12309 26776
rect 12739 26816 12797 26817
rect 12739 26776 12748 26816
rect 12788 26776 12797 26816
rect 13275 26785 13276 26825
rect 13316 26785 13317 26825
rect 13275 26776 13317 26785
rect 13795 26816 13853 26817
rect 13795 26776 13804 26816
rect 13844 26776 13853 26816
rect 12739 26775 12797 26776
rect 13795 26775 13853 26776
rect 14083 26816 14141 26817
rect 14083 26776 14092 26816
rect 14132 26776 14141 26816
rect 14083 26775 14141 26776
rect 14371 26816 14429 26817
rect 14371 26776 14380 26816
rect 14420 26776 14429 26816
rect 14371 26775 14429 26776
rect 14563 26816 14621 26817
rect 14563 26776 14572 26816
rect 14612 26776 14621 26816
rect 14563 26775 14621 26776
rect 15811 26816 15869 26817
rect 15811 26776 15820 26816
rect 15860 26776 15869 26816
rect 15811 26775 15869 26776
rect 16195 26816 16253 26817
rect 16195 26776 16204 26816
rect 16244 26776 16253 26816
rect 16195 26775 16253 26776
rect 16587 26816 16629 26825
rect 16771 26818 16780 26858
rect 16820 26818 16829 26858
rect 16771 26817 16829 26818
rect 16587 26776 16588 26816
rect 16628 26776 16629 26816
rect 16587 26767 16629 26776
rect 16971 26816 17013 26825
rect 16971 26776 16972 26816
rect 17012 26776 17013 26816
rect 16971 26767 17013 26776
rect 17059 26816 17117 26817
rect 17059 26776 17068 26816
rect 17108 26776 17117 26816
rect 17059 26775 17117 26776
rect 17251 26816 17309 26817
rect 17251 26776 17260 26816
rect 17300 26776 17309 26816
rect 17251 26775 17309 26776
rect 18691 26816 18749 26817
rect 18691 26776 18700 26816
rect 18740 26776 18749 26816
rect 18691 26775 18749 26776
rect 18795 26816 18837 26825
rect 18795 26776 18796 26816
rect 18836 26776 18837 26816
rect 18795 26767 18837 26776
rect 18979 26816 19037 26817
rect 18979 26776 18988 26816
rect 19028 26776 19037 26816
rect 18979 26775 19037 26776
rect 19179 26816 19221 26825
rect 19179 26776 19180 26816
rect 19220 26776 19221 26816
rect 19179 26767 19221 26776
rect 19371 26816 19413 26825
rect 19371 26776 19372 26816
rect 19412 26776 19413 26816
rect 19371 26767 19413 26776
rect 11787 26747 11829 26756
rect 3531 26732 3573 26741
rect 3531 26692 3532 26732
rect 3572 26692 3573 26732
rect 3531 26683 3573 26692
rect 5835 26648 5877 26657
rect 5835 26608 5836 26648
rect 5876 26608 5877 26648
rect 5835 26599 5877 26608
rect 8523 26648 8565 26657
rect 8523 26608 8524 26648
rect 8564 26608 8565 26648
rect 8523 26599 8565 26608
rect 8995 26648 9053 26649
rect 8995 26608 9004 26648
rect 9044 26608 9053 26648
rect 8995 26607 9053 26608
rect 9571 26648 9629 26649
rect 9571 26608 9580 26648
rect 9620 26608 9629 26648
rect 9571 26607 9629 26608
rect 13419 26648 13461 26657
rect 13419 26608 13420 26648
rect 13460 26608 13461 26648
rect 13419 26599 13461 26608
rect 16011 26648 16053 26657
rect 16011 26608 16012 26648
rect 16052 26608 16053 26648
rect 16011 26599 16053 26608
rect 16779 26648 16821 26657
rect 16779 26608 16780 26648
rect 16820 26608 16821 26648
rect 16779 26599 16821 26608
rect 17355 26648 17397 26657
rect 17355 26608 17356 26648
rect 17396 26608 17397 26648
rect 17355 26599 17397 26608
rect 18987 26648 19029 26657
rect 18987 26608 18988 26648
rect 19028 26608 19029 26648
rect 18987 26599 19029 26608
rect 19275 26648 19317 26657
rect 19275 26608 19276 26648
rect 19316 26608 19317 26648
rect 19275 26599 19317 26608
rect 19755 26648 19797 26657
rect 19755 26608 19756 26648
rect 19796 26608 19797 26648
rect 19755 26599 19797 26608
rect 20139 26648 20181 26657
rect 20139 26608 20140 26648
rect 20180 26608 20181 26648
rect 20139 26599 20181 26608
rect 1152 26480 20452 26504
rect 1152 26440 4928 26480
rect 4968 26440 5010 26480
rect 5050 26440 5092 26480
rect 5132 26440 5174 26480
rect 5214 26440 5256 26480
rect 5296 26440 20048 26480
rect 20088 26440 20130 26480
rect 20170 26440 20212 26480
rect 20252 26440 20294 26480
rect 20334 26440 20376 26480
rect 20416 26440 20452 26480
rect 1152 26416 20452 26440
rect 3619 26312 3677 26313
rect 3619 26272 3628 26312
rect 3668 26272 3677 26312
rect 3619 26271 3677 26272
rect 6979 26312 7037 26313
rect 6979 26272 6988 26312
rect 7028 26272 7037 26312
rect 6979 26271 7037 26272
rect 11491 26312 11549 26313
rect 11491 26272 11500 26312
rect 11540 26272 11549 26312
rect 11491 26271 11549 26272
rect 11883 26312 11925 26321
rect 11883 26272 11884 26312
rect 11924 26272 11925 26312
rect 11883 26263 11925 26272
rect 15435 26312 15477 26321
rect 15435 26272 15436 26312
rect 15476 26272 15477 26312
rect 15435 26263 15477 26272
rect 16675 26312 16733 26313
rect 16675 26272 16684 26312
rect 16724 26272 16733 26312
rect 16675 26271 16733 26272
rect 17451 26312 17493 26321
rect 17451 26272 17452 26312
rect 17492 26272 17493 26312
rect 17451 26263 17493 26272
rect 12075 26228 12117 26237
rect 12075 26188 12076 26228
rect 12116 26188 12117 26228
rect 12075 26179 12117 26188
rect 3232 26148 3290 26149
rect 1315 26144 1373 26145
rect 1315 26104 1324 26144
rect 1364 26104 1373 26144
rect 1315 26103 1373 26104
rect 1507 26144 1565 26145
rect 1507 26104 1516 26144
rect 1556 26104 1565 26144
rect 1507 26103 1565 26104
rect 2755 26144 2813 26145
rect 2755 26104 2764 26144
rect 2804 26104 2813 26144
rect 3232 26108 3241 26148
rect 3281 26108 3290 26148
rect 3232 26107 3290 26108
rect 3331 26144 3389 26145
rect 2755 26103 2813 26104
rect 3331 26104 3340 26144
rect 3380 26104 3389 26144
rect 3331 26103 3389 26104
rect 3497 26144 3555 26145
rect 3497 26104 3506 26144
rect 3546 26104 3555 26144
rect 3763 26144 3821 26145
rect 3497 26103 3555 26104
rect 3619 26115 3677 26116
rect 3619 26075 3628 26115
rect 3668 26075 3677 26115
rect 3763 26104 3772 26144
rect 3812 26104 3821 26144
rect 3763 26103 3821 26104
rect 4011 26144 4053 26153
rect 4011 26104 4012 26144
rect 4052 26104 4053 26144
rect 4011 26095 4053 26104
rect 4387 26144 4445 26145
rect 4387 26104 4396 26144
rect 4436 26104 4445 26144
rect 4387 26103 4445 26104
rect 4587 26144 4629 26153
rect 4587 26104 4588 26144
rect 4628 26104 4629 26144
rect 4587 26095 4629 26104
rect 4779 26144 4821 26153
rect 4779 26104 4780 26144
rect 4820 26104 4821 26144
rect 4779 26095 4821 26104
rect 5059 26144 5117 26145
rect 5059 26104 5068 26144
rect 5108 26104 5117 26144
rect 5059 26103 5117 26104
rect 5355 26144 5397 26153
rect 5355 26104 5356 26144
rect 5396 26104 5397 26144
rect 5355 26095 5397 26104
rect 5451 26144 5493 26153
rect 5451 26104 5452 26144
rect 5492 26104 5493 26144
rect 5451 26095 5493 26104
rect 6019 26144 6077 26145
rect 6019 26104 6028 26144
rect 6068 26104 6077 26144
rect 6019 26103 6077 26104
rect 6315 26144 6357 26153
rect 6315 26104 6316 26144
rect 6356 26104 6357 26144
rect 6315 26095 6357 26104
rect 6411 26144 6453 26153
rect 6411 26104 6412 26144
rect 6452 26104 6453 26144
rect 7083 26144 7125 26153
rect 6411 26095 6453 26104
rect 6925 26129 6967 26138
rect 6925 26089 6926 26129
rect 6966 26089 6967 26129
rect 7083 26104 7084 26144
rect 7124 26104 7125 26144
rect 7083 26095 7125 26104
rect 7179 26144 7221 26153
rect 7179 26104 7180 26144
rect 7220 26104 7221 26144
rect 7179 26095 7221 26104
rect 7363 26144 7421 26145
rect 7363 26104 7372 26144
rect 7412 26104 7421 26144
rect 7363 26103 7421 26104
rect 7459 26144 7517 26145
rect 7459 26104 7468 26144
rect 7508 26104 7517 26144
rect 7459 26103 7517 26104
rect 7747 26144 7805 26145
rect 7747 26104 7756 26144
rect 7796 26104 7805 26144
rect 7747 26103 7805 26104
rect 7851 26144 7893 26153
rect 7851 26104 7852 26144
rect 7892 26104 7893 26144
rect 7851 26095 7893 26104
rect 8035 26144 8093 26145
rect 8035 26104 8044 26144
rect 8084 26104 8093 26144
rect 8035 26103 8093 26104
rect 8419 26144 8477 26145
rect 8419 26104 8428 26144
rect 8468 26104 8477 26144
rect 8419 26103 8477 26104
rect 9667 26144 9725 26145
rect 9667 26104 9676 26144
rect 9716 26104 9725 26144
rect 9667 26103 9725 26104
rect 9859 26144 9917 26145
rect 9859 26104 9868 26144
rect 9908 26104 9917 26144
rect 9859 26103 9917 26104
rect 11107 26144 11165 26145
rect 11107 26104 11116 26144
rect 11156 26104 11165 26144
rect 11107 26103 11165 26104
rect 11779 26144 11837 26145
rect 11779 26104 11788 26144
rect 11828 26104 11837 26144
rect 11779 26103 11837 26104
rect 12355 26144 12413 26145
rect 12355 26104 12364 26144
rect 12404 26104 12413 26144
rect 12355 26103 12413 26104
rect 13603 26144 13661 26145
rect 13603 26104 13612 26144
rect 13652 26104 13661 26144
rect 13603 26103 13661 26104
rect 13987 26144 14045 26145
rect 13987 26104 13996 26144
rect 14036 26104 14045 26144
rect 13987 26103 14045 26104
rect 15235 26144 15293 26145
rect 15235 26104 15244 26144
rect 15284 26104 15293 26144
rect 15235 26103 15293 26104
rect 15715 26144 15773 26145
rect 15715 26104 15724 26144
rect 15764 26104 15773 26144
rect 15715 26103 15773 26104
rect 16011 26144 16053 26153
rect 16011 26104 16012 26144
rect 16052 26104 16053 26144
rect 16011 26095 16053 26104
rect 16107 26144 16149 26153
rect 16107 26104 16108 26144
rect 16148 26104 16149 26144
rect 16779 26144 16821 26153
rect 16107 26095 16149 26104
rect 16621 26129 16663 26138
rect 6925 26080 6967 26089
rect 16621 26089 16622 26129
rect 16662 26089 16663 26129
rect 16779 26104 16780 26144
rect 16820 26104 16821 26144
rect 16779 26095 16821 26104
rect 16875 26144 16917 26153
rect 16875 26104 16876 26144
rect 16916 26104 16917 26144
rect 16875 26095 16917 26104
rect 17059 26144 17117 26145
rect 17059 26104 17068 26144
rect 17108 26104 17117 26144
rect 17059 26103 17117 26104
rect 17155 26144 17213 26145
rect 17155 26104 17164 26144
rect 17204 26104 17213 26144
rect 17155 26103 17213 26104
rect 17355 26144 17397 26153
rect 17355 26104 17356 26144
rect 17396 26104 17397 26144
rect 17355 26095 17397 26104
rect 17547 26144 17589 26153
rect 17547 26104 17548 26144
rect 17588 26104 17589 26144
rect 17547 26095 17589 26104
rect 17731 26144 17789 26145
rect 17731 26104 17740 26144
rect 17780 26104 17789 26144
rect 17731 26103 17789 26104
rect 18979 26144 19037 26145
rect 18979 26104 18988 26144
rect 19028 26104 19037 26144
rect 18979 26103 19037 26104
rect 19371 26144 19413 26153
rect 19371 26104 19372 26144
rect 19412 26104 19413 26144
rect 19371 26095 19413 26104
rect 19747 26144 19805 26145
rect 19747 26104 19756 26144
rect 19796 26104 19805 26144
rect 19747 26103 19805 26104
rect 16621 26080 16663 26089
rect 3619 26074 3677 26075
rect 1227 26060 1269 26069
rect 1227 26020 1228 26060
rect 1268 26020 1269 26060
rect 1227 26011 1269 26020
rect 4107 26060 4149 26069
rect 4107 26020 4108 26060
rect 4148 26020 4149 26060
rect 4107 26011 4149 26020
rect 4299 26060 4341 26069
rect 4299 26020 4300 26060
rect 4340 26020 4341 26060
rect 4299 26011 4341 26020
rect 19467 26060 19509 26069
rect 19467 26020 19468 26060
rect 19508 26020 19509 26060
rect 19467 26011 19509 26020
rect 19659 26060 19701 26069
rect 19659 26020 19660 26060
rect 19700 26020 19701 26060
rect 19659 26011 19701 26020
rect 19939 26060 19997 26061
rect 19939 26020 19948 26060
rect 19988 26020 19997 26060
rect 19939 26019 19997 26020
rect 2955 25976 2997 25985
rect 2955 25936 2956 25976
rect 2996 25936 2997 25976
rect 2955 25927 2997 25936
rect 4203 25976 4245 25985
rect 4203 25936 4204 25976
rect 4244 25936 4245 25976
rect 4203 25927 4245 25936
rect 5731 25976 5789 25977
rect 5731 25936 5740 25976
rect 5780 25936 5789 25976
rect 5731 25935 5789 25936
rect 6691 25976 6749 25977
rect 6691 25936 6700 25976
rect 6740 25936 6749 25976
rect 6691 25935 6749 25936
rect 16387 25976 16445 25977
rect 16387 25936 16396 25976
rect 16436 25936 16445 25976
rect 16387 25935 16445 25936
rect 19563 25976 19605 25985
rect 19563 25936 19564 25976
rect 19604 25936 19605 25976
rect 19563 25927 19605 25936
rect 4587 25892 4629 25901
rect 4587 25852 4588 25892
rect 4628 25852 4629 25892
rect 4587 25843 4629 25852
rect 7851 25892 7893 25901
rect 7851 25852 7852 25892
rect 7892 25852 7893 25892
rect 7851 25843 7893 25852
rect 8235 25892 8277 25901
rect 8235 25852 8236 25892
rect 8276 25852 8277 25892
rect 8235 25843 8277 25852
rect 11307 25892 11349 25901
rect 11307 25852 11308 25892
rect 11348 25852 11349 25892
rect 11307 25843 11349 25852
rect 13803 25892 13845 25901
rect 13803 25852 13804 25892
rect 13844 25852 13845 25892
rect 13803 25843 13845 25852
rect 19179 25892 19221 25901
rect 19179 25852 19180 25892
rect 19220 25852 19221 25892
rect 19179 25843 19221 25852
rect 20139 25892 20181 25901
rect 20139 25852 20140 25892
rect 20180 25852 20181 25892
rect 20139 25843 20181 25852
rect 1152 25724 20352 25748
rect 1152 25684 3688 25724
rect 3728 25684 3770 25724
rect 3810 25684 3852 25724
rect 3892 25684 3934 25724
rect 3974 25684 4016 25724
rect 4056 25684 18808 25724
rect 18848 25684 18890 25724
rect 18930 25684 18972 25724
rect 19012 25684 19054 25724
rect 19094 25684 19136 25724
rect 19176 25684 20352 25724
rect 1152 25660 20352 25684
rect 5643 25556 5685 25565
rect 5643 25516 5644 25556
rect 5684 25516 5685 25556
rect 5643 25507 5685 25516
rect 6219 25556 6261 25565
rect 6219 25516 6220 25556
rect 6260 25516 6261 25556
rect 6219 25507 6261 25516
rect 8043 25556 8085 25565
rect 8043 25516 8044 25556
rect 8084 25516 8085 25556
rect 8043 25507 8085 25516
rect 15531 25556 15573 25565
rect 15531 25516 15532 25556
rect 15572 25516 15573 25556
rect 15531 25507 15573 25516
rect 16483 25556 16541 25557
rect 16483 25516 16492 25556
rect 16532 25516 16541 25556
rect 16483 25515 16541 25516
rect 19651 25556 19709 25557
rect 19651 25516 19660 25556
rect 19700 25516 19709 25556
rect 19651 25515 19709 25516
rect 3243 25472 3285 25481
rect 3243 25432 3244 25472
rect 3284 25432 3285 25472
rect 3243 25423 3285 25432
rect 8995 25472 9053 25473
rect 8995 25432 9004 25472
rect 9044 25432 9053 25472
rect 8995 25431 9053 25432
rect 9387 25472 9429 25481
rect 9387 25432 9388 25472
rect 9428 25432 9429 25472
rect 9387 25423 9429 25432
rect 16875 25472 16917 25481
rect 16875 25432 16876 25472
rect 16916 25432 16917 25472
rect 16875 25423 16917 25432
rect 20043 25472 20085 25481
rect 20043 25432 20044 25472
rect 20084 25432 20085 25472
rect 20043 25423 20085 25432
rect 3147 25388 3189 25397
rect 3147 25348 3148 25388
rect 3188 25348 3189 25388
rect 3147 25339 3189 25348
rect 3339 25388 3381 25397
rect 3339 25348 3340 25388
rect 3380 25348 3381 25388
rect 3339 25339 3381 25348
rect 9291 25388 9333 25397
rect 9291 25348 9292 25388
rect 9332 25348 9333 25388
rect 9291 25339 9333 25348
rect 9483 25388 9525 25397
rect 9483 25348 9484 25388
rect 9524 25348 9525 25388
rect 9483 25339 9525 25348
rect 11595 25388 11637 25397
rect 11595 25348 11596 25388
rect 11636 25348 11637 25388
rect 11595 25339 11637 25348
rect 12747 25388 12789 25397
rect 12747 25348 12748 25388
rect 12788 25348 12789 25388
rect 12747 25339 12789 25348
rect 16779 25388 16821 25397
rect 16779 25348 16780 25388
rect 16820 25348 16821 25388
rect 16779 25339 16821 25348
rect 16971 25388 17013 25397
rect 16971 25348 16972 25388
rect 17012 25348 17013 25388
rect 16971 25339 17013 25348
rect 19947 25388 19989 25397
rect 19947 25348 19948 25388
rect 19988 25348 19989 25388
rect 19947 25339 19989 25348
rect 20129 25388 20171 25397
rect 20129 25348 20130 25388
rect 20170 25348 20171 25388
rect 20129 25339 20171 25348
rect 13707 25318 13749 25327
rect 1219 25304 1277 25305
rect 1219 25264 1228 25304
rect 1268 25264 1277 25304
rect 1219 25263 1277 25264
rect 2467 25304 2525 25305
rect 2467 25264 2476 25304
rect 2516 25264 2525 25304
rect 2467 25263 2525 25264
rect 3043 25304 3101 25305
rect 3043 25264 3052 25304
rect 3092 25264 3101 25304
rect 3043 25263 3101 25264
rect 3435 25304 3477 25313
rect 3435 25264 3436 25304
rect 3476 25264 3477 25304
rect 3435 25255 3477 25264
rect 3619 25304 3677 25305
rect 3619 25264 3628 25304
rect 3668 25264 3677 25304
rect 3619 25263 3677 25264
rect 4867 25304 4925 25305
rect 4867 25264 4876 25304
rect 4916 25264 4925 25304
rect 4867 25263 4925 25264
rect 5259 25304 5301 25313
rect 5259 25264 5260 25304
rect 5300 25264 5301 25304
rect 5259 25255 5301 25264
rect 5451 25304 5493 25313
rect 5451 25264 5452 25304
rect 5492 25264 5493 25304
rect 5451 25255 5493 25264
rect 5731 25304 5789 25305
rect 5731 25264 5740 25304
rect 5780 25264 5789 25304
rect 5731 25263 5789 25264
rect 5923 25304 5981 25305
rect 5923 25264 5932 25304
rect 5972 25264 5981 25304
rect 5923 25263 5981 25264
rect 6027 25304 6069 25313
rect 6027 25264 6028 25304
rect 6068 25264 6069 25304
rect 6027 25255 6069 25264
rect 6211 25304 6269 25305
rect 6211 25264 6220 25304
rect 6260 25264 6269 25304
rect 6211 25263 6269 25264
rect 6595 25304 6653 25305
rect 6595 25264 6604 25304
rect 6644 25264 6653 25304
rect 6595 25263 6653 25264
rect 7843 25304 7901 25305
rect 7843 25264 7852 25304
rect 7892 25264 7901 25304
rect 7843 25263 7901 25264
rect 8323 25304 8381 25305
rect 8323 25264 8332 25304
rect 8372 25264 8381 25304
rect 8323 25263 8381 25264
rect 8619 25304 8661 25313
rect 8619 25264 8620 25304
rect 8660 25264 8661 25304
rect 8619 25255 8661 25264
rect 8715 25304 8757 25313
rect 8715 25264 8716 25304
rect 8756 25264 8757 25304
rect 8715 25255 8757 25264
rect 9187 25304 9245 25305
rect 9187 25264 9196 25304
rect 9236 25264 9245 25304
rect 9187 25263 9245 25264
rect 9579 25304 9621 25313
rect 9579 25264 9580 25304
rect 9620 25264 9621 25304
rect 9579 25255 9621 25264
rect 9859 25304 9917 25305
rect 9859 25264 9868 25304
rect 9908 25264 9917 25304
rect 9859 25263 9917 25264
rect 11107 25304 11165 25305
rect 11107 25264 11116 25304
rect 11156 25264 11165 25304
rect 11107 25263 11165 25264
rect 12171 25304 12213 25313
rect 12171 25264 12172 25304
rect 12212 25264 12213 25304
rect 12171 25255 12213 25264
rect 12267 25304 12309 25313
rect 12267 25264 12268 25304
rect 12308 25264 12309 25304
rect 12267 25255 12309 25264
rect 12651 25304 12693 25313
rect 12651 25264 12652 25304
rect 12692 25264 12693 25304
rect 12651 25255 12693 25264
rect 13219 25304 13277 25305
rect 13219 25264 13228 25304
rect 13268 25264 13277 25304
rect 13707 25278 13708 25318
rect 13748 25278 13749 25318
rect 13707 25269 13749 25278
rect 14083 25304 14141 25305
rect 13219 25263 13277 25264
rect 14083 25264 14092 25304
rect 14132 25264 14141 25304
rect 14083 25263 14141 25264
rect 15331 25304 15389 25305
rect 15331 25264 15340 25304
rect 15380 25264 15389 25304
rect 15331 25263 15389 25264
rect 15811 25304 15869 25305
rect 15811 25264 15820 25304
rect 15860 25264 15869 25304
rect 15811 25263 15869 25264
rect 16107 25304 16149 25313
rect 16107 25264 16108 25304
rect 16148 25264 16149 25304
rect 16107 25255 16149 25264
rect 16675 25304 16733 25305
rect 16675 25264 16684 25304
rect 16724 25264 16733 25304
rect 16675 25263 16733 25264
rect 17067 25304 17109 25313
rect 17067 25264 17068 25304
rect 17108 25264 17109 25304
rect 17067 25255 17109 25264
rect 17443 25304 17501 25305
rect 17443 25264 17452 25304
rect 17492 25264 17501 25304
rect 17443 25263 17501 25264
rect 18691 25304 18749 25305
rect 18691 25264 18700 25304
rect 18740 25264 18749 25304
rect 18691 25263 18749 25264
rect 18979 25304 19037 25305
rect 18979 25264 18988 25304
rect 19028 25264 19037 25304
rect 18979 25263 19037 25264
rect 19275 25304 19317 25313
rect 19275 25264 19276 25304
rect 19316 25264 19317 25304
rect 19275 25255 19317 25264
rect 19851 25304 19893 25313
rect 19851 25264 19852 25304
rect 19892 25264 19893 25304
rect 19851 25255 19893 25264
rect 20227 25304 20285 25305
rect 20227 25264 20236 25304
rect 20276 25264 20285 25304
rect 20227 25263 20285 25264
rect 5067 25220 5109 25229
rect 5067 25180 5068 25220
rect 5108 25180 5109 25220
rect 5067 25171 5109 25180
rect 13899 25220 13941 25229
rect 13899 25180 13900 25220
rect 13940 25180 13941 25220
rect 13899 25171 13941 25180
rect 16203 25220 16245 25229
rect 16203 25180 16204 25220
rect 16244 25180 16245 25220
rect 16203 25171 16245 25180
rect 17259 25220 17301 25229
rect 17259 25180 17260 25220
rect 17300 25180 17301 25220
rect 17259 25171 17301 25180
rect 19371 25220 19413 25229
rect 19371 25180 19372 25220
rect 19412 25180 19413 25220
rect 19371 25171 19413 25180
rect 2667 25136 2709 25145
rect 2667 25096 2668 25136
rect 2708 25096 2709 25136
rect 2667 25087 2709 25096
rect 5355 25136 5397 25145
rect 5355 25096 5356 25136
rect 5396 25096 5397 25136
rect 5355 25087 5397 25096
rect 8043 25136 8085 25145
rect 8043 25096 8044 25136
rect 8084 25096 8085 25136
rect 8043 25087 8085 25096
rect 11307 25136 11349 25145
rect 11307 25096 11308 25136
rect 11348 25096 11349 25136
rect 11307 25087 11349 25096
rect 1152 24968 20452 24992
rect 1152 24928 4928 24968
rect 4968 24928 5010 24968
rect 5050 24928 5092 24968
rect 5132 24928 5174 24968
rect 5214 24928 5256 24968
rect 5296 24928 20048 24968
rect 20088 24928 20130 24968
rect 20170 24928 20212 24968
rect 20252 24928 20294 24968
rect 20334 24928 20376 24968
rect 20416 24928 20452 24968
rect 1152 24904 20452 24928
rect 6699 24800 6741 24809
rect 6699 24760 6700 24800
rect 6740 24760 6741 24800
rect 6699 24751 6741 24760
rect 9475 24800 9533 24801
rect 9475 24760 9484 24800
rect 9524 24760 9533 24800
rect 9475 24759 9533 24760
rect 19459 24800 19517 24801
rect 19459 24760 19468 24800
rect 19508 24760 19517 24800
rect 19459 24759 19517 24760
rect 3147 24716 3189 24725
rect 3147 24676 3148 24716
rect 3188 24676 3189 24716
rect 3147 24667 3189 24676
rect 4779 24716 4821 24725
rect 4779 24676 4780 24716
rect 4820 24676 4821 24716
rect 4779 24667 4821 24676
rect 12075 24716 12117 24725
rect 12075 24676 12076 24716
rect 12116 24676 12117 24716
rect 12075 24667 12117 24676
rect 17931 24716 17973 24725
rect 17931 24676 17932 24716
rect 17972 24676 17973 24716
rect 17931 24667 17973 24676
rect 18603 24716 18645 24725
rect 18603 24676 18604 24716
rect 18644 24676 18645 24716
rect 18603 24667 18645 24676
rect 4369 24647 4427 24648
rect 1411 24632 1469 24633
rect 1411 24592 1420 24632
rect 1460 24592 1469 24632
rect 1411 24591 1469 24592
rect 2659 24632 2717 24633
rect 2659 24592 2668 24632
rect 2708 24592 2717 24632
rect 2659 24591 2717 24592
rect 3043 24632 3101 24633
rect 3043 24592 3052 24632
rect 3092 24592 3101 24632
rect 3043 24591 3101 24592
rect 3435 24632 3477 24641
rect 3435 24592 3436 24632
rect 3476 24592 3477 24632
rect 3435 24583 3477 24592
rect 3819 24632 3861 24641
rect 3819 24592 3820 24632
rect 3860 24592 3861 24632
rect 3819 24583 3861 24592
rect 3915 24632 3957 24641
rect 3915 24592 3916 24632
rect 3956 24592 3957 24632
rect 3915 24583 3957 24592
rect 4011 24632 4053 24641
rect 4011 24592 4012 24632
rect 4052 24592 4053 24632
rect 4011 24583 4053 24592
rect 4107 24632 4149 24641
rect 4107 24592 4108 24632
rect 4148 24592 4149 24632
rect 4369 24607 4378 24647
rect 4418 24607 4427 24647
rect 18193 24647 18251 24648
rect 4369 24606 4427 24607
rect 4683 24632 4725 24641
rect 4107 24583 4149 24592
rect 4683 24592 4684 24632
rect 4724 24592 4725 24632
rect 4683 24583 4725 24592
rect 5251 24632 5309 24633
rect 5251 24592 5260 24632
rect 5300 24592 5309 24632
rect 5251 24591 5309 24592
rect 5355 24632 5397 24641
rect 5355 24592 5356 24632
rect 5396 24592 5397 24632
rect 5355 24583 5397 24592
rect 5547 24632 5589 24641
rect 5547 24592 5548 24632
rect 5588 24592 5589 24632
rect 5547 24583 5589 24592
rect 5739 24632 5781 24641
rect 5739 24592 5740 24632
rect 5780 24592 5781 24632
rect 5739 24583 5781 24592
rect 5931 24632 5973 24641
rect 5931 24592 5932 24632
rect 5972 24592 5973 24632
rect 5931 24583 5973 24592
rect 6315 24632 6357 24641
rect 6315 24592 6316 24632
rect 6356 24592 6357 24632
rect 6315 24583 6357 24592
rect 6507 24632 6549 24641
rect 6507 24592 6508 24632
rect 6548 24592 6549 24632
rect 6507 24583 6549 24592
rect 6883 24632 6941 24633
rect 6883 24592 6892 24632
rect 6932 24592 6941 24632
rect 6883 24591 6941 24592
rect 8131 24632 8189 24633
rect 8131 24592 8140 24632
rect 8180 24592 8189 24632
rect 8131 24591 8189 24592
rect 8515 24632 8573 24633
rect 8515 24592 8524 24632
rect 8564 24592 8573 24632
rect 8515 24591 8573 24592
rect 8811 24632 8853 24641
rect 8811 24592 8812 24632
rect 8852 24592 8853 24632
rect 8811 24583 8853 24592
rect 8907 24632 8949 24641
rect 8907 24592 8908 24632
rect 8948 24592 8949 24632
rect 9579 24632 9621 24641
rect 8907 24583 8949 24592
rect 9421 24617 9463 24626
rect 9421 24577 9422 24617
rect 9462 24577 9463 24617
rect 9579 24592 9580 24632
rect 9620 24592 9621 24632
rect 9579 24583 9621 24592
rect 9675 24632 9717 24641
rect 9675 24592 9676 24632
rect 9716 24592 9717 24632
rect 9675 24583 9717 24592
rect 9859 24632 9917 24633
rect 9859 24592 9868 24632
rect 9908 24592 9917 24632
rect 9859 24591 9917 24592
rect 9955 24632 10013 24633
rect 9955 24592 9964 24632
rect 10004 24592 10013 24632
rect 9955 24591 10013 24592
rect 10347 24632 10389 24641
rect 10347 24592 10348 24632
rect 10388 24592 10389 24632
rect 10347 24583 10389 24592
rect 10443 24632 10485 24641
rect 10443 24592 10444 24632
rect 10484 24592 10485 24632
rect 10443 24583 10485 24592
rect 10923 24632 10965 24641
rect 10923 24592 10924 24632
rect 10964 24592 10965 24632
rect 10923 24583 10965 24592
rect 11395 24632 11453 24633
rect 11395 24592 11404 24632
rect 11444 24592 11453 24632
rect 13027 24632 13085 24633
rect 11395 24591 11453 24592
rect 11883 24618 11925 24627
rect 9421 24568 9463 24577
rect 11883 24578 11884 24618
rect 11924 24578 11925 24618
rect 13027 24592 13036 24632
rect 13076 24592 13085 24632
rect 13027 24591 13085 24592
rect 14851 24632 14909 24633
rect 14851 24592 14860 24632
rect 14900 24592 14909 24632
rect 14851 24591 14909 24592
rect 16099 24632 16157 24633
rect 16099 24592 16108 24632
rect 16148 24592 16157 24632
rect 16099 24591 16157 24592
rect 16483 24632 16541 24633
rect 16483 24592 16492 24632
rect 16532 24592 16541 24632
rect 16483 24591 16541 24592
rect 17731 24632 17789 24633
rect 17731 24592 17740 24632
rect 17780 24592 17789 24632
rect 18193 24607 18202 24647
rect 18242 24607 18251 24647
rect 18193 24606 18251 24607
rect 18507 24632 18549 24641
rect 17731 24591 17789 24592
rect 18507 24592 18508 24632
rect 18548 24592 18549 24632
rect 19275 24632 19317 24641
rect 11883 24569 11925 24578
rect 14275 24590 14333 24591
rect 5835 24548 5877 24557
rect 5835 24508 5836 24548
rect 5876 24508 5877 24548
rect 5835 24499 5877 24508
rect 10827 24548 10869 24557
rect 14275 24550 14284 24590
rect 14324 24550 14333 24590
rect 18507 24583 18549 24592
rect 19117 24617 19159 24626
rect 19117 24577 19118 24617
rect 19158 24577 19159 24617
rect 19275 24592 19276 24632
rect 19316 24592 19317 24632
rect 19275 24583 19317 24592
rect 19371 24632 19413 24641
rect 19371 24592 19372 24632
rect 19412 24592 19413 24632
rect 19371 24583 19413 24592
rect 19555 24632 19613 24633
rect 19555 24592 19564 24632
rect 19604 24592 19613 24632
rect 19555 24591 19613 24592
rect 19651 24632 19709 24633
rect 19651 24592 19660 24632
rect 19700 24592 19709 24632
rect 19651 24591 19709 24592
rect 19117 24568 19159 24577
rect 14275 24549 14333 24550
rect 10827 24508 10828 24548
rect 10868 24508 10869 24548
rect 10827 24499 10869 24508
rect 19843 24548 19901 24549
rect 19843 24508 19852 24548
rect 19892 24508 19901 24548
rect 19843 24507 19901 24508
rect 2859 24464 2901 24473
rect 2859 24424 2860 24464
rect 2900 24424 2901 24464
rect 2859 24415 2901 24424
rect 3435 24464 3477 24473
rect 3435 24424 3436 24464
rect 3476 24424 3477 24464
rect 3435 24415 3477 24424
rect 5059 24464 5117 24465
rect 5059 24424 5068 24464
rect 5108 24424 5117 24464
rect 5059 24423 5117 24424
rect 6507 24464 6549 24473
rect 6507 24424 6508 24464
rect 6548 24424 6549 24464
rect 6507 24415 6549 24424
rect 9187 24464 9245 24465
rect 9187 24424 9196 24464
rect 9236 24424 9245 24464
rect 9187 24423 9245 24424
rect 18883 24464 18941 24465
rect 18883 24424 18892 24464
rect 18932 24424 18941 24464
rect 18883 24423 18941 24424
rect 20043 24464 20085 24473
rect 20043 24424 20044 24464
rect 20084 24424 20085 24464
rect 20043 24415 20085 24424
rect 3627 24380 3669 24389
rect 3627 24340 3628 24380
rect 3668 24340 3669 24380
rect 3627 24331 3669 24340
rect 5547 24380 5589 24389
rect 5547 24340 5548 24380
rect 5588 24340 5589 24380
rect 5547 24331 5589 24340
rect 6699 24380 6741 24389
rect 6699 24340 6700 24380
rect 6740 24340 6741 24380
rect 6699 24331 6741 24340
rect 14475 24380 14517 24389
rect 14475 24340 14476 24380
rect 14516 24340 14517 24380
rect 14475 24331 14517 24340
rect 16299 24380 16341 24389
rect 16299 24340 16300 24380
rect 16340 24340 16341 24380
rect 16299 24331 16341 24340
rect 1152 24212 20352 24236
rect 1152 24172 3688 24212
rect 3728 24172 3770 24212
rect 3810 24172 3852 24212
rect 3892 24172 3934 24212
rect 3974 24172 4016 24212
rect 4056 24172 18808 24212
rect 18848 24172 18890 24212
rect 18930 24172 18972 24212
rect 19012 24172 19054 24212
rect 19094 24172 19136 24212
rect 19176 24172 20352 24212
rect 1152 24148 20352 24172
rect 8331 23960 8373 23969
rect 8331 23920 8332 23960
rect 8372 23920 8373 23960
rect 8331 23911 8373 23920
rect 8715 23960 8757 23969
rect 8715 23920 8716 23960
rect 8756 23920 8757 23960
rect 8715 23911 8757 23920
rect 8899 23960 8957 23961
rect 8899 23920 8908 23960
rect 8948 23920 8957 23960
rect 8899 23919 8957 23920
rect 12363 23960 12405 23969
rect 12363 23920 12364 23960
rect 12404 23920 12405 23960
rect 12363 23911 12405 23920
rect 18787 23960 18845 23961
rect 18787 23920 18796 23960
rect 18836 23920 18845 23960
rect 18787 23919 18845 23920
rect 20235 23960 20277 23969
rect 20235 23920 20236 23960
rect 20276 23920 20277 23960
rect 20235 23911 20277 23920
rect 1603 23876 1661 23877
rect 1603 23836 1612 23876
rect 1652 23836 1661 23876
rect 1603 23835 1661 23836
rect 6411 23876 6453 23885
rect 6411 23836 6412 23876
rect 6452 23836 6453 23876
rect 6411 23827 6453 23836
rect 10923 23876 10965 23885
rect 10923 23836 10924 23876
rect 10964 23836 10965 23876
rect 19747 23876 19805 23877
rect 10923 23827 10965 23836
rect 16059 23834 16101 23843
rect 19747 23836 19756 23876
rect 19796 23836 19805 23876
rect 19747 23835 19805 23836
rect 4011 23806 4053 23815
rect 1899 23792 1941 23801
rect 1899 23752 1900 23792
rect 1940 23752 1941 23792
rect 1899 23743 1941 23752
rect 2475 23792 2517 23801
rect 2475 23752 2476 23792
rect 2516 23752 2517 23792
rect 2475 23743 2517 23752
rect 2571 23792 2613 23801
rect 2571 23752 2572 23792
rect 2612 23752 2613 23792
rect 2571 23743 2613 23752
rect 2955 23792 2997 23801
rect 2955 23752 2956 23792
rect 2996 23752 2997 23792
rect 2955 23743 2997 23752
rect 3051 23792 3093 23801
rect 3051 23752 3052 23792
rect 3092 23752 3093 23792
rect 3051 23743 3093 23752
rect 3523 23792 3581 23793
rect 3523 23752 3532 23792
rect 3572 23752 3581 23792
rect 4011 23766 4012 23806
rect 4052 23766 4053 23806
rect 6075 23801 6117 23810
rect 11979 23806 12021 23815
rect 4011 23757 4053 23766
rect 4491 23792 4533 23801
rect 3523 23751 3581 23752
rect 4491 23752 4492 23792
rect 4532 23752 4533 23792
rect 4491 23743 4533 23752
rect 4587 23792 4629 23801
rect 4587 23752 4588 23792
rect 4628 23752 4629 23792
rect 4587 23743 4629 23752
rect 4971 23792 5013 23801
rect 4971 23752 4972 23792
rect 5012 23752 5013 23792
rect 4971 23743 5013 23752
rect 5067 23792 5109 23801
rect 5067 23752 5068 23792
rect 5108 23752 5109 23792
rect 5067 23743 5109 23752
rect 5539 23792 5597 23793
rect 5539 23752 5548 23792
rect 5588 23752 5597 23792
rect 6075 23761 6076 23801
rect 6116 23761 6117 23801
rect 6075 23752 6117 23761
rect 6499 23792 6557 23793
rect 6499 23752 6508 23792
rect 6548 23752 6557 23792
rect 5539 23751 5597 23752
rect 6499 23751 6557 23752
rect 6883 23792 6941 23793
rect 6883 23752 6892 23792
rect 6932 23752 6941 23792
rect 6883 23751 6941 23752
rect 8131 23792 8189 23793
rect 8131 23752 8140 23792
rect 8180 23752 8189 23792
rect 8131 23751 8189 23752
rect 8523 23792 8565 23801
rect 8523 23752 8524 23792
rect 8564 23752 8565 23792
rect 8523 23743 8565 23752
rect 8715 23792 8757 23801
rect 8715 23752 8716 23792
rect 8756 23752 8757 23792
rect 8715 23743 8757 23752
rect 9195 23792 9237 23801
rect 9195 23752 9196 23792
rect 9236 23752 9237 23792
rect 9195 23743 9237 23752
rect 9291 23792 9333 23801
rect 9291 23752 9292 23792
rect 9332 23752 9333 23792
rect 9291 23743 9333 23752
rect 9571 23792 9629 23793
rect 9571 23752 9580 23792
rect 9620 23752 9629 23792
rect 9571 23751 9629 23752
rect 9859 23792 9917 23793
rect 9859 23752 9868 23792
rect 9908 23752 9917 23792
rect 9859 23751 9917 23752
rect 9963 23792 10005 23801
rect 9963 23752 9964 23792
rect 10004 23752 10005 23792
rect 9963 23743 10005 23752
rect 10147 23792 10205 23793
rect 10147 23752 10156 23792
rect 10196 23752 10205 23792
rect 10147 23751 10205 23752
rect 10443 23792 10485 23801
rect 10443 23752 10444 23792
rect 10484 23752 10485 23792
rect 10443 23743 10485 23752
rect 10539 23792 10581 23801
rect 10539 23752 10540 23792
rect 10580 23752 10581 23792
rect 10539 23743 10581 23752
rect 11019 23792 11061 23801
rect 11019 23752 11020 23792
rect 11060 23752 11061 23792
rect 11019 23743 11061 23752
rect 11491 23792 11549 23793
rect 11491 23752 11500 23792
rect 11540 23752 11549 23792
rect 11979 23766 11980 23806
rect 12020 23766 12021 23806
rect 11979 23757 12021 23766
rect 12547 23792 12605 23793
rect 11491 23751 11549 23752
rect 12547 23752 12556 23792
rect 12596 23752 12605 23792
rect 12547 23751 12605 23752
rect 13795 23792 13853 23793
rect 13795 23752 13804 23792
rect 13844 23752 13853 23792
rect 13795 23751 13853 23752
rect 14475 23792 14517 23801
rect 14475 23752 14476 23792
rect 14516 23752 14517 23792
rect 14475 23743 14517 23752
rect 14571 23792 14613 23801
rect 14571 23752 14572 23792
rect 14612 23752 14613 23792
rect 14571 23743 14613 23752
rect 14955 23792 14997 23801
rect 14955 23752 14956 23792
rect 14996 23752 14997 23792
rect 14955 23743 14997 23752
rect 15051 23792 15093 23801
rect 16059 23794 16060 23834
rect 16100 23794 16101 23834
rect 19021 23807 19063 23816
rect 15051 23752 15052 23792
rect 15092 23752 15093 23792
rect 15051 23743 15093 23752
rect 15523 23792 15581 23793
rect 15523 23752 15532 23792
rect 15572 23752 15581 23792
rect 16059 23785 16101 23794
rect 16579 23792 16637 23793
rect 15523 23751 15581 23752
rect 16579 23752 16588 23792
rect 16628 23752 16637 23792
rect 16579 23751 16637 23752
rect 17827 23792 17885 23793
rect 17827 23752 17836 23792
rect 17876 23752 17885 23792
rect 17827 23751 17885 23752
rect 18115 23792 18173 23793
rect 18115 23752 18124 23792
rect 18164 23752 18173 23792
rect 18115 23751 18173 23752
rect 18411 23792 18453 23801
rect 18411 23752 18412 23792
rect 18452 23752 18453 23792
rect 19021 23767 19022 23807
rect 19062 23767 19063 23807
rect 20131 23805 20189 23806
rect 19021 23758 19063 23767
rect 19179 23792 19221 23801
rect 18411 23743 18453 23752
rect 19179 23752 19180 23792
rect 19220 23752 19221 23792
rect 19179 23743 19221 23752
rect 19275 23792 19317 23801
rect 19275 23752 19276 23792
rect 19316 23752 19317 23792
rect 19275 23743 19317 23752
rect 19459 23792 19517 23793
rect 19459 23752 19468 23792
rect 19508 23752 19517 23792
rect 19459 23751 19517 23752
rect 19555 23792 19613 23793
rect 19555 23752 19564 23792
rect 19604 23752 19613 23792
rect 20131 23765 20140 23805
rect 20180 23765 20189 23805
rect 20131 23764 20189 23765
rect 19555 23751 19613 23752
rect 4203 23708 4245 23717
rect 4203 23668 4204 23708
rect 4244 23668 4245 23708
rect 4203 23659 4245 23668
rect 18507 23708 18549 23717
rect 18507 23668 18508 23708
rect 18548 23668 18549 23708
rect 18507 23659 18549 23668
rect 1419 23624 1461 23633
rect 1419 23584 1420 23624
rect 1460 23584 1461 23624
rect 1419 23575 1461 23584
rect 2179 23624 2237 23625
rect 2179 23584 2188 23624
rect 2228 23584 2237 23624
rect 2179 23583 2237 23584
rect 6219 23624 6261 23633
rect 6219 23584 6220 23624
rect 6260 23584 6261 23624
rect 6219 23575 6261 23584
rect 10155 23624 10197 23633
rect 10155 23584 10156 23624
rect 10196 23584 10197 23624
rect 10155 23575 10197 23584
rect 12171 23624 12213 23633
rect 12171 23584 12172 23624
rect 12212 23584 12213 23624
rect 12171 23575 12213 23584
rect 16203 23624 16245 23633
rect 16203 23584 16204 23624
rect 16244 23584 16245 23624
rect 16203 23575 16245 23584
rect 16395 23624 16437 23633
rect 16395 23584 16396 23624
rect 16436 23584 16437 23624
rect 16395 23575 16437 23584
rect 19363 23624 19421 23625
rect 19363 23584 19372 23624
rect 19412 23584 19421 23624
rect 19363 23583 19421 23584
rect 19947 23624 19989 23633
rect 19947 23584 19948 23624
rect 19988 23584 19989 23624
rect 19947 23575 19989 23584
rect 1152 23456 20452 23480
rect 1152 23416 4928 23456
rect 4968 23416 5010 23456
rect 5050 23416 5092 23456
rect 5132 23416 5174 23456
rect 5214 23416 5256 23456
rect 5296 23416 20048 23456
rect 20088 23416 20130 23456
rect 20170 23416 20212 23456
rect 20252 23416 20294 23456
rect 20334 23416 20376 23456
rect 20416 23416 20452 23456
rect 1152 23392 20452 23416
rect 1315 23288 1373 23289
rect 1315 23248 1324 23288
rect 1364 23248 1373 23288
rect 1315 23247 1373 23248
rect 3339 23288 3381 23297
rect 3339 23248 3340 23288
rect 3380 23248 3381 23288
rect 3339 23239 3381 23248
rect 3627 23288 3669 23297
rect 3627 23248 3628 23288
rect 3668 23248 3669 23288
rect 3627 23239 3669 23248
rect 4291 23288 4349 23289
rect 4291 23248 4300 23288
rect 4340 23248 4349 23288
rect 4291 23247 4349 23248
rect 6315 23288 6357 23297
rect 6315 23248 6316 23288
rect 6356 23248 6357 23288
rect 6315 23239 6357 23248
rect 10539 23288 10581 23297
rect 10539 23248 10540 23288
rect 10580 23248 10581 23288
rect 10539 23239 10581 23248
rect 10915 23288 10973 23289
rect 10915 23248 10924 23288
rect 10964 23248 10973 23288
rect 10915 23247 10973 23248
rect 18027 23288 18069 23297
rect 18027 23248 18028 23288
rect 18068 23248 18069 23288
rect 18027 23239 18069 23248
rect 11595 23204 11637 23213
rect 11595 23164 11596 23204
rect 11636 23164 11637 23204
rect 11595 23155 11637 23164
rect 12363 23204 12405 23213
rect 12363 23164 12364 23204
rect 12404 23164 12405 23204
rect 12363 23155 12405 23164
rect 14283 23204 14325 23213
rect 14283 23164 14284 23204
rect 14324 23164 14325 23204
rect 14283 23155 14325 23164
rect 16299 23204 16341 23213
rect 16299 23164 16300 23204
rect 16340 23164 16341 23204
rect 16299 23155 16341 23164
rect 1891 23120 1949 23121
rect 1891 23080 1900 23120
rect 1940 23080 1949 23120
rect 1891 23079 1949 23080
rect 3139 23120 3197 23121
rect 3139 23080 3148 23120
rect 3188 23080 3197 23120
rect 3139 23079 3197 23080
rect 3811 23120 3869 23121
rect 3811 23080 3820 23120
rect 3860 23080 3869 23120
rect 3811 23079 3869 23080
rect 4011 23120 4053 23129
rect 4011 23080 4012 23120
rect 4052 23080 4053 23120
rect 4011 23071 4053 23080
rect 4099 23120 4157 23121
rect 4099 23080 4108 23120
rect 4148 23080 4157 23120
rect 4099 23079 4157 23080
rect 4395 23120 4437 23129
rect 4395 23080 4396 23120
rect 4436 23080 4437 23120
rect 4395 23071 4437 23080
rect 4491 23120 4533 23129
rect 4491 23080 4492 23120
rect 4532 23080 4533 23120
rect 4491 23071 4533 23080
rect 4587 23120 4629 23129
rect 4587 23080 4588 23120
rect 4628 23080 4629 23120
rect 4587 23071 4629 23080
rect 4867 23120 4925 23121
rect 4867 23080 4876 23120
rect 4916 23080 4925 23120
rect 4867 23079 4925 23080
rect 6115 23120 6173 23121
rect 6115 23080 6124 23120
rect 6164 23080 6173 23120
rect 6115 23079 6173 23080
rect 6691 23120 6749 23121
rect 6691 23080 6700 23120
rect 6740 23080 6749 23120
rect 6691 23079 6749 23080
rect 7939 23120 7997 23121
rect 7939 23080 7948 23120
rect 7988 23080 7997 23120
rect 7939 23079 7997 23080
rect 8515 23120 8573 23121
rect 8515 23080 8524 23120
rect 8564 23080 8573 23120
rect 8515 23079 8573 23080
rect 8907 23120 8949 23129
rect 8907 23080 8908 23120
rect 8948 23080 8949 23120
rect 8907 23071 8949 23080
rect 9091 23120 9149 23121
rect 9091 23080 9100 23120
rect 9140 23080 9149 23120
rect 9091 23079 9149 23080
rect 10339 23120 10397 23121
rect 10339 23080 10348 23120
rect 10388 23080 10397 23120
rect 10339 23079 10397 23080
rect 10723 23120 10781 23121
rect 10723 23080 10732 23120
rect 10772 23080 10781 23120
rect 11019 23120 11061 23129
rect 10723 23079 10781 23080
rect 10867 23110 10925 23111
rect 10867 23070 10876 23110
rect 10916 23070 10925 23110
rect 11019 23080 11020 23120
rect 11060 23080 11061 23120
rect 11019 23071 11061 23080
rect 11115 23120 11157 23129
rect 11115 23080 11116 23120
rect 11156 23080 11157 23120
rect 11491 23120 11549 23121
rect 11115 23071 11157 23080
rect 11272 23105 11314 23114
rect 10867 23069 10925 23070
rect 11272 23065 11273 23105
rect 11313 23065 11314 23105
rect 11491 23080 11500 23120
rect 11540 23080 11549 23120
rect 11491 23079 11549 23080
rect 11971 23120 12029 23121
rect 11971 23080 11980 23120
rect 12020 23080 12029 23120
rect 11971 23079 12029 23080
rect 12267 23120 12309 23129
rect 12267 23080 12268 23120
rect 12308 23080 12309 23120
rect 12267 23071 12309 23080
rect 12835 23120 12893 23121
rect 12835 23080 12844 23120
rect 12884 23080 12893 23120
rect 12835 23079 12893 23080
rect 14083 23120 14141 23121
rect 14083 23080 14092 23120
rect 14132 23080 14141 23120
rect 14083 23079 14141 23080
rect 14571 23120 14613 23129
rect 14571 23080 14572 23120
rect 14612 23080 14613 23120
rect 14571 23071 14613 23080
rect 14667 23120 14709 23129
rect 14667 23080 14668 23120
rect 14708 23080 14709 23120
rect 14667 23071 14709 23080
rect 15619 23120 15677 23121
rect 15619 23080 15628 23120
rect 15668 23080 15677 23120
rect 16579 23120 16637 23121
rect 15619 23079 15677 23080
rect 16155 23110 16197 23119
rect 11272 23056 11314 23065
rect 16155 23070 16156 23110
rect 16196 23070 16197 23110
rect 16579 23080 16588 23120
rect 16628 23080 16637 23120
rect 16579 23079 16637 23080
rect 17827 23120 17885 23121
rect 17827 23080 17836 23120
rect 17876 23080 17885 23120
rect 17827 23079 17885 23080
rect 18403 23120 18461 23121
rect 18403 23080 18412 23120
rect 18452 23080 18461 23120
rect 18403 23079 18461 23080
rect 19651 23120 19709 23121
rect 19651 23080 19660 23120
rect 19700 23080 19709 23120
rect 19651 23079 19709 23080
rect 20043 23120 20085 23129
rect 20043 23080 20044 23120
rect 20084 23080 20085 23120
rect 20043 23071 20085 23080
rect 20235 23120 20277 23129
rect 20235 23080 20236 23120
rect 20276 23080 20277 23120
rect 20235 23071 20277 23080
rect 16155 23061 16197 23070
rect 1699 23036 1757 23037
rect 1699 22996 1708 23036
rect 1748 22996 1757 23036
rect 1699 22995 1757 22996
rect 8619 23036 8661 23045
rect 8619 22996 8620 23036
rect 8660 22996 8661 23036
rect 8619 22987 8661 22996
rect 8811 23036 8853 23045
rect 8811 22996 8812 23036
rect 8852 22996 8853 23036
rect 8811 22987 8853 22996
rect 15051 23036 15093 23045
rect 15051 22996 15052 23036
rect 15092 22996 15093 23036
rect 15051 22987 15093 22996
rect 15147 23036 15189 23045
rect 15147 22996 15148 23036
rect 15188 22996 15189 23036
rect 15147 22987 15189 22996
rect 20139 23036 20181 23045
rect 20139 22996 20140 23036
rect 20180 22996 20181 23036
rect 20139 22987 20181 22996
rect 3627 22952 3669 22961
rect 3627 22912 3628 22952
rect 3668 22912 3669 22952
rect 3627 22903 3669 22912
rect 8715 22952 8757 22961
rect 8715 22912 8716 22952
rect 8756 22912 8757 22952
rect 8715 22903 8757 22912
rect 19851 22952 19893 22961
rect 19851 22912 19852 22952
rect 19892 22912 19893 22952
rect 19851 22903 19893 22912
rect 1515 22868 1557 22877
rect 1515 22828 1516 22868
rect 1556 22828 1557 22868
rect 1515 22819 1557 22828
rect 3819 22868 3861 22877
rect 3819 22828 3820 22868
rect 3860 22828 3861 22868
rect 3819 22819 3861 22828
rect 8139 22868 8181 22877
rect 8139 22828 8140 22868
rect 8180 22828 8181 22868
rect 8139 22819 8181 22828
rect 12643 22868 12701 22869
rect 12643 22828 12652 22868
rect 12692 22828 12701 22868
rect 12643 22827 12701 22828
rect 18027 22868 18069 22877
rect 18027 22828 18028 22868
rect 18068 22828 18069 22868
rect 18027 22819 18069 22828
rect 1152 22700 20352 22724
rect 1152 22660 3688 22700
rect 3728 22660 3770 22700
rect 3810 22660 3852 22700
rect 3892 22660 3934 22700
rect 3974 22660 4016 22700
rect 4056 22660 18808 22700
rect 18848 22660 18890 22700
rect 18930 22660 18972 22700
rect 19012 22660 19054 22700
rect 19094 22660 19136 22700
rect 19176 22660 20352 22700
rect 1152 22636 20352 22660
rect 10731 22532 10773 22541
rect 10731 22492 10732 22532
rect 10772 22492 10773 22532
rect 10731 22483 10773 22492
rect 11683 22532 11741 22533
rect 11683 22492 11692 22532
rect 11732 22492 11741 22532
rect 11683 22491 11741 22492
rect 20235 22532 20277 22541
rect 20235 22492 20236 22532
rect 20276 22492 20277 22532
rect 20235 22483 20277 22492
rect 3147 22448 3189 22457
rect 3147 22408 3148 22448
rect 3188 22408 3189 22448
rect 3147 22399 3189 22408
rect 4491 22448 4533 22457
rect 4491 22408 4492 22448
rect 4532 22408 4533 22448
rect 4491 22399 4533 22408
rect 4875 22448 4917 22457
rect 4875 22408 4876 22448
rect 4916 22408 4917 22448
rect 4875 22399 4917 22408
rect 8907 22448 8949 22457
rect 8907 22408 8908 22448
rect 8948 22408 8949 22448
rect 8907 22399 8949 22408
rect 18307 22448 18365 22449
rect 18307 22408 18316 22448
rect 18356 22408 18365 22448
rect 18307 22407 18365 22408
rect 3051 22364 3093 22373
rect 3051 22324 3052 22364
rect 3092 22324 3093 22364
rect 3051 22315 3093 22324
rect 3243 22364 3285 22373
rect 3243 22324 3244 22364
rect 3284 22324 3285 22364
rect 3243 22315 3285 22324
rect 4395 22364 4437 22373
rect 4395 22324 4396 22364
rect 4436 22324 4437 22364
rect 4395 22315 4437 22324
rect 4587 22364 4629 22373
rect 4587 22324 4588 22364
rect 4628 22324 4629 22364
rect 4587 22315 4629 22324
rect 5451 22364 5493 22373
rect 5451 22324 5452 22364
rect 5492 22324 5493 22364
rect 5451 22315 5493 22324
rect 6987 22364 7029 22373
rect 6987 22324 6988 22364
rect 7028 22324 7029 22364
rect 6987 22315 7029 22324
rect 7083 22364 7125 22373
rect 7083 22324 7084 22364
rect 7124 22324 7125 22364
rect 7083 22315 7125 22324
rect 8811 22364 8853 22373
rect 8811 22324 8812 22364
rect 8852 22324 8853 22364
rect 8811 22315 8853 22324
rect 9003 22364 9045 22373
rect 9003 22324 9004 22364
rect 9044 22324 9045 22364
rect 9003 22315 9045 22324
rect 11979 22364 12021 22373
rect 11979 22324 11980 22364
rect 12020 22324 12021 22364
rect 11979 22315 12021 22324
rect 13507 22322 13565 22323
rect 8043 22294 8085 22303
rect 1219 22280 1277 22281
rect 1219 22240 1228 22280
rect 1268 22240 1277 22280
rect 1219 22239 1277 22240
rect 2467 22280 2525 22281
rect 2467 22240 2476 22280
rect 2516 22240 2525 22280
rect 2467 22239 2525 22240
rect 2947 22280 3005 22281
rect 2947 22240 2956 22280
rect 2996 22240 3005 22280
rect 2947 22239 3005 22240
rect 3339 22280 3381 22289
rect 3339 22240 3340 22280
rect 3380 22240 3381 22280
rect 3339 22231 3381 22240
rect 3523 22280 3581 22281
rect 3523 22240 3532 22280
rect 3572 22240 3581 22280
rect 3523 22239 3581 22240
rect 3619 22280 3677 22281
rect 3619 22240 3628 22280
rect 3668 22240 3677 22280
rect 3619 22239 3677 22240
rect 3819 22280 3861 22289
rect 3819 22240 3820 22280
rect 3860 22240 3861 22280
rect 3819 22231 3861 22240
rect 3915 22280 3957 22289
rect 3915 22240 3916 22280
rect 3956 22240 3957 22280
rect 3915 22231 3957 22240
rect 4062 22280 4120 22281
rect 4062 22240 4071 22280
rect 4111 22240 4120 22280
rect 4062 22239 4120 22240
rect 4291 22280 4349 22281
rect 4291 22240 4300 22280
rect 4340 22240 4349 22280
rect 4291 22239 4349 22240
rect 4683 22280 4725 22289
rect 4683 22240 4684 22280
rect 4724 22240 4725 22280
rect 4683 22231 4725 22240
rect 6507 22280 6549 22289
rect 6507 22240 6508 22280
rect 6548 22240 6549 22280
rect 6507 22231 6549 22240
rect 6603 22280 6645 22289
rect 6603 22240 6604 22280
rect 6644 22240 6645 22280
rect 6603 22231 6645 22240
rect 7555 22280 7613 22281
rect 7555 22240 7564 22280
rect 7604 22240 7613 22280
rect 8043 22254 8044 22294
rect 8084 22254 8085 22294
rect 8043 22245 8085 22254
rect 8707 22280 8765 22281
rect 7555 22239 7613 22240
rect 8707 22240 8716 22280
rect 8756 22240 8765 22280
rect 8707 22239 8765 22240
rect 9099 22280 9141 22289
rect 9099 22240 9100 22280
rect 9140 22240 9141 22280
rect 9099 22231 9141 22240
rect 9283 22280 9341 22281
rect 9283 22240 9292 22280
rect 9332 22240 9341 22280
rect 9283 22239 9341 22240
rect 10531 22280 10589 22281
rect 10531 22240 10540 22280
rect 10580 22240 10589 22280
rect 10531 22239 10589 22240
rect 11011 22280 11069 22281
rect 11011 22240 11020 22280
rect 11060 22240 11069 22280
rect 11011 22239 11069 22240
rect 11307 22280 11349 22289
rect 11307 22240 11308 22280
rect 11348 22240 11349 22280
rect 11307 22231 11349 22240
rect 11883 22280 11925 22289
rect 11883 22240 11884 22280
rect 11924 22240 11925 22280
rect 11883 22231 11925 22240
rect 12075 22280 12117 22289
rect 13507 22282 13516 22322
rect 13556 22282 13565 22322
rect 13507 22281 13565 22282
rect 12075 22240 12076 22280
rect 12116 22240 12117 22280
rect 12075 22231 12117 22240
rect 12259 22280 12317 22281
rect 12259 22240 12268 22280
rect 12308 22240 12317 22280
rect 12259 22239 12317 22240
rect 14851 22280 14909 22281
rect 14851 22240 14860 22280
rect 14900 22240 14909 22280
rect 14851 22239 14909 22240
rect 16099 22280 16157 22281
rect 16099 22240 16108 22280
rect 16148 22240 16157 22280
rect 16099 22239 16157 22240
rect 16683 22280 16725 22289
rect 16683 22240 16684 22280
rect 16724 22240 16725 22280
rect 16683 22231 16725 22240
rect 16875 22280 16917 22289
rect 16875 22240 16876 22280
rect 16916 22240 16917 22280
rect 16875 22231 16917 22240
rect 17067 22280 17109 22289
rect 17067 22240 17068 22280
rect 17108 22240 17109 22280
rect 17067 22231 17109 22240
rect 17163 22280 17205 22289
rect 17163 22240 17164 22280
rect 17204 22240 17205 22280
rect 17163 22231 17205 22240
rect 17635 22280 17693 22281
rect 17635 22240 17644 22280
rect 17684 22240 17693 22280
rect 17635 22239 17693 22240
rect 17931 22280 17973 22289
rect 17931 22240 17932 22280
rect 17972 22240 17973 22280
rect 17931 22231 17973 22240
rect 18027 22280 18069 22289
rect 18027 22240 18028 22280
rect 18068 22240 18069 22280
rect 18027 22231 18069 22240
rect 18499 22280 18557 22281
rect 18499 22240 18508 22280
rect 18548 22240 18557 22280
rect 18499 22239 18557 22240
rect 19747 22280 19805 22281
rect 19747 22240 19756 22280
rect 19796 22240 19805 22280
rect 19747 22239 19805 22240
rect 20126 22269 20168 22278
rect 20126 22229 20127 22269
rect 20167 22229 20168 22269
rect 20126 22220 20168 22229
rect 5739 22196 5781 22205
rect 5739 22156 5740 22196
rect 5780 22156 5781 22196
rect 5739 22147 5781 22156
rect 11403 22196 11445 22205
rect 11403 22156 11404 22196
rect 11444 22156 11445 22196
rect 11403 22147 11445 22156
rect 19947 22196 19989 22205
rect 19947 22156 19948 22196
rect 19988 22156 19989 22196
rect 19947 22147 19989 22156
rect 2667 22112 2709 22121
rect 2667 22072 2668 22112
rect 2708 22072 2709 22112
rect 2667 22063 2709 22072
rect 3715 22112 3773 22113
rect 3715 22072 3724 22112
rect 3764 22072 3773 22112
rect 3715 22071 3773 22072
rect 5259 22112 5301 22121
rect 5259 22072 5260 22112
rect 5300 22072 5301 22112
rect 5259 22063 5301 22072
rect 6123 22112 6165 22121
rect 6123 22072 6124 22112
rect 6164 22072 6165 22112
rect 6123 22063 6165 22072
rect 8235 22112 8277 22121
rect 8235 22072 8236 22112
rect 8276 22072 8277 22112
rect 8235 22063 8277 22072
rect 8419 22112 8477 22113
rect 8419 22072 8428 22112
rect 8468 22072 8477 22112
rect 8419 22071 8477 22072
rect 10731 22112 10773 22121
rect 10731 22072 10732 22112
rect 10772 22072 10773 22112
rect 10731 22063 10773 22072
rect 13707 22112 13749 22121
rect 13707 22072 13708 22112
rect 13748 22072 13749 22112
rect 13707 22063 13749 22072
rect 16299 22112 16341 22121
rect 16299 22072 16300 22112
rect 16340 22072 16341 22112
rect 16299 22063 16341 22072
rect 16779 22112 16821 22121
rect 16779 22072 16780 22112
rect 16820 22072 16821 22112
rect 16779 22063 16821 22072
rect 17347 22112 17405 22113
rect 17347 22072 17356 22112
rect 17396 22072 17405 22112
rect 17347 22071 17405 22072
rect 20235 22112 20277 22121
rect 20235 22072 20236 22112
rect 20276 22072 20277 22112
rect 20235 22063 20277 22072
rect 1152 21944 20452 21968
rect 1152 21904 4928 21944
rect 4968 21904 5010 21944
rect 5050 21904 5092 21944
rect 5132 21904 5174 21944
rect 5214 21904 5256 21944
rect 5296 21904 20048 21944
rect 20088 21904 20130 21944
rect 20170 21904 20212 21944
rect 20252 21904 20294 21944
rect 20334 21904 20376 21944
rect 20416 21904 20452 21944
rect 1152 21880 20452 21904
rect 3051 21776 3093 21785
rect 3051 21736 3052 21776
rect 3092 21736 3093 21776
rect 3051 21727 3093 21736
rect 3627 21776 3669 21785
rect 3627 21736 3628 21776
rect 3668 21736 3669 21776
rect 3627 21727 3669 21736
rect 6027 21776 6069 21785
rect 6027 21736 6028 21776
rect 6068 21736 6069 21776
rect 6027 21727 6069 21736
rect 9675 21776 9717 21785
rect 9675 21736 9676 21776
rect 9716 21736 9717 21776
rect 9675 21727 9717 21736
rect 16395 21776 16437 21785
rect 16395 21736 16396 21776
rect 16436 21736 16437 21776
rect 16395 21727 16437 21736
rect 18499 21776 18557 21777
rect 18499 21736 18508 21776
rect 18548 21736 18557 21776
rect 18499 21735 18557 21736
rect 8043 21692 8085 21701
rect 8043 21652 8044 21692
rect 8084 21652 8085 21692
rect 8043 21643 8085 21652
rect 11979 21692 12021 21701
rect 11979 21652 11980 21692
rect 12020 21652 12021 21692
rect 11979 21643 12021 21652
rect 13995 21692 14037 21701
rect 13995 21652 13996 21692
rect 14036 21652 14037 21692
rect 13995 21643 14037 21652
rect 20131 21622 20189 21623
rect 1603 21608 1661 21609
rect 1603 21568 1612 21608
rect 1652 21568 1661 21608
rect 1603 21567 1661 21568
rect 2851 21608 2909 21609
rect 2851 21568 2860 21608
rect 2900 21568 2909 21608
rect 2851 21567 2909 21568
rect 4203 21608 4245 21617
rect 4203 21568 4204 21608
rect 4244 21568 4245 21608
rect 4203 21559 4245 21568
rect 4395 21608 4437 21617
rect 4395 21568 4396 21608
rect 4436 21568 4437 21608
rect 4395 21559 4437 21568
rect 4579 21608 4637 21609
rect 4579 21568 4588 21608
rect 4628 21568 4637 21608
rect 4579 21567 4637 21568
rect 5827 21608 5885 21609
rect 5827 21568 5836 21608
rect 5876 21568 5885 21608
rect 5827 21567 5885 21568
rect 6315 21608 6357 21617
rect 6315 21568 6316 21608
rect 6356 21568 6357 21608
rect 6315 21559 6357 21568
rect 6411 21608 6453 21617
rect 6411 21568 6412 21608
rect 6452 21568 6453 21608
rect 6411 21559 6453 21568
rect 6795 21608 6837 21617
rect 6795 21568 6796 21608
rect 6836 21568 6837 21608
rect 6795 21559 6837 21568
rect 6891 21608 6933 21617
rect 6891 21568 6892 21608
rect 6932 21568 6933 21608
rect 6891 21559 6933 21568
rect 7363 21608 7421 21609
rect 7363 21568 7372 21608
rect 7412 21568 7421 21608
rect 8227 21608 8285 21609
rect 7363 21567 7421 21568
rect 7851 21594 7893 21603
rect 7851 21554 7852 21594
rect 7892 21554 7893 21594
rect 8227 21568 8236 21608
rect 8276 21568 8285 21608
rect 8227 21567 8285 21568
rect 9475 21608 9533 21609
rect 9475 21568 9484 21608
rect 9524 21568 9533 21608
rect 9475 21567 9533 21568
rect 9955 21608 10013 21609
rect 9955 21568 9964 21608
rect 10004 21568 10013 21608
rect 9955 21567 10013 21568
rect 10347 21608 10389 21617
rect 10347 21568 10348 21608
rect 10388 21568 10389 21608
rect 10347 21559 10389 21568
rect 10531 21608 10589 21609
rect 10531 21568 10540 21608
rect 10580 21568 10589 21608
rect 10531 21567 10589 21568
rect 11779 21608 11837 21609
rect 11779 21568 11788 21608
rect 11828 21568 11837 21608
rect 11779 21567 11837 21568
rect 12267 21608 12309 21617
rect 12267 21568 12268 21608
rect 12308 21568 12309 21608
rect 12267 21559 12309 21568
rect 12363 21608 12405 21617
rect 12363 21568 12364 21608
rect 12404 21568 12405 21608
rect 12363 21559 12405 21568
rect 12747 21608 12789 21617
rect 12747 21568 12748 21608
rect 12788 21568 12789 21608
rect 12747 21559 12789 21568
rect 12843 21608 12885 21617
rect 12843 21568 12844 21608
rect 12884 21568 12885 21608
rect 12843 21559 12885 21568
rect 13315 21608 13373 21609
rect 13315 21568 13324 21608
rect 13364 21568 13373 21608
rect 13315 21567 13373 21568
rect 13803 21603 13845 21612
rect 13803 21563 13804 21603
rect 13844 21563 13845 21603
rect 13803 21554 13845 21563
rect 14667 21608 14709 21617
rect 14667 21568 14668 21608
rect 14708 21568 14709 21608
rect 14667 21559 14709 21568
rect 14763 21608 14805 21617
rect 14763 21568 14764 21608
rect 14804 21568 14805 21608
rect 14763 21559 14805 21568
rect 15715 21608 15773 21609
rect 15715 21568 15724 21608
rect 15764 21568 15773 21608
rect 16579 21608 16637 21609
rect 15715 21567 15773 21568
rect 16251 21598 16293 21607
rect 16251 21558 16252 21598
rect 16292 21558 16293 21598
rect 16579 21568 16588 21608
rect 16628 21568 16637 21608
rect 16579 21567 16637 21568
rect 17827 21608 17885 21609
rect 17827 21568 17836 21608
rect 17876 21568 17885 21608
rect 17827 21567 17885 21568
rect 18219 21608 18261 21617
rect 18219 21568 18220 21608
rect 18260 21568 18261 21608
rect 18219 21559 18261 21568
rect 18315 21608 18357 21617
rect 18315 21568 18316 21608
rect 18356 21568 18357 21608
rect 18315 21559 18357 21568
rect 18411 21608 18453 21617
rect 18411 21568 18412 21608
rect 18452 21568 18453 21608
rect 18411 21559 18453 21568
rect 18691 21608 18749 21609
rect 18691 21568 18700 21608
rect 18740 21568 18749 21608
rect 18691 21567 18749 21568
rect 19083 21608 19125 21617
rect 19083 21568 19084 21608
rect 19124 21568 19125 21608
rect 19083 21559 19125 21568
rect 19275 21608 19317 21617
rect 19275 21568 19276 21608
rect 19316 21568 19317 21608
rect 19275 21559 19317 21568
rect 19651 21608 19709 21609
rect 19651 21568 19660 21608
rect 19700 21568 19709 21608
rect 19651 21567 19709 21568
rect 19843 21608 19901 21609
rect 19843 21568 19852 21608
rect 19892 21568 19901 21608
rect 19843 21567 19901 21568
rect 19947 21608 19989 21617
rect 19947 21568 19948 21608
rect 19988 21568 19989 21608
rect 20131 21582 20140 21622
rect 20180 21582 20189 21622
rect 20131 21581 20189 21582
rect 19947 21559 19989 21568
rect 7851 21545 7893 21554
rect 16251 21549 16293 21558
rect 1411 21524 1469 21525
rect 1411 21484 1420 21524
rect 1460 21484 1469 21524
rect 1411 21483 1469 21484
rect 3339 21524 3381 21533
rect 3339 21484 3340 21524
rect 3380 21484 3381 21524
rect 3339 21475 3381 21484
rect 3915 21524 3957 21533
rect 3915 21484 3916 21524
rect 3956 21484 3957 21524
rect 3915 21475 3957 21484
rect 10059 21524 10101 21533
rect 10059 21484 10060 21524
rect 10100 21484 10101 21524
rect 10059 21475 10101 21484
rect 10251 21524 10293 21533
rect 10251 21484 10252 21524
rect 10292 21484 10293 21524
rect 10251 21475 10293 21484
rect 15147 21524 15189 21533
rect 15147 21484 15148 21524
rect 15188 21484 15189 21524
rect 15147 21475 15189 21484
rect 15243 21524 15285 21533
rect 15243 21484 15244 21524
rect 15284 21484 15285 21524
rect 15243 21475 15285 21484
rect 18795 21524 18837 21533
rect 18795 21484 18796 21524
rect 18836 21484 18837 21524
rect 18795 21475 18837 21484
rect 18987 21524 19029 21533
rect 18987 21484 18988 21524
rect 19028 21484 19029 21524
rect 18987 21475 19029 21484
rect 19371 21524 19413 21533
rect 19371 21484 19372 21524
rect 19412 21484 19413 21524
rect 19371 21475 19413 21484
rect 19563 21524 19605 21533
rect 19563 21484 19564 21524
rect 19604 21484 19605 21524
rect 19563 21475 19605 21484
rect 3531 21440 3573 21449
rect 3531 21400 3532 21440
rect 3572 21400 3573 21440
rect 3531 21391 3573 21400
rect 4395 21440 4437 21449
rect 4395 21400 4396 21440
rect 4436 21400 4437 21440
rect 4395 21391 4437 21400
rect 10155 21440 10197 21449
rect 10155 21400 10156 21440
rect 10196 21400 10197 21440
rect 10155 21391 10197 21400
rect 18891 21440 18933 21449
rect 18891 21400 18892 21440
rect 18932 21400 18933 21440
rect 18891 21391 18933 21400
rect 19467 21440 19509 21449
rect 19467 21400 19468 21440
rect 19508 21400 19509 21440
rect 19467 21391 19509 21400
rect 19939 21440 19997 21441
rect 19939 21400 19948 21440
rect 19988 21400 19997 21440
rect 19939 21399 19997 21400
rect 1227 21356 1269 21365
rect 1227 21316 1228 21356
rect 1268 21316 1269 21356
rect 1227 21307 1269 21316
rect 18027 21356 18069 21365
rect 18027 21316 18028 21356
rect 18068 21316 18069 21356
rect 18027 21307 18069 21316
rect 1152 21188 20352 21212
rect 1152 21148 3688 21188
rect 3728 21148 3770 21188
rect 3810 21148 3852 21188
rect 3892 21148 3934 21188
rect 3974 21148 4016 21188
rect 4056 21148 18808 21188
rect 18848 21148 18890 21188
rect 18930 21148 18972 21188
rect 19012 21148 19054 21188
rect 19094 21148 19136 21188
rect 19176 21148 20352 21188
rect 1152 21124 20352 21148
rect 6123 21020 6165 21029
rect 6123 20980 6124 21020
rect 6164 20980 6165 21020
rect 6123 20971 6165 20980
rect 7755 21020 7797 21029
rect 7755 20980 7756 21020
rect 7796 20980 7797 21020
rect 7755 20971 7797 20980
rect 14859 21020 14901 21029
rect 14859 20980 14860 21020
rect 14900 20980 14901 21020
rect 14859 20971 14901 20980
rect 15627 21020 15669 21029
rect 15627 20980 15628 21020
rect 15668 20980 15669 21020
rect 15627 20971 15669 20980
rect 17259 21020 17301 21029
rect 17259 20980 17260 21020
rect 17300 20980 17301 21020
rect 17259 20971 17301 20980
rect 2859 20936 2901 20945
rect 2859 20896 2860 20936
rect 2900 20896 2901 20936
rect 2859 20887 2901 20896
rect 3147 20936 3189 20945
rect 3147 20896 3148 20936
rect 3188 20896 3189 20936
rect 3147 20887 3189 20896
rect 3531 20936 3573 20945
rect 3531 20896 3532 20936
rect 3572 20896 3573 20936
rect 3531 20887 3573 20896
rect 4011 20936 4053 20945
rect 4011 20896 4012 20936
rect 4052 20896 4053 20936
rect 4011 20887 4053 20896
rect 3915 20852 3957 20861
rect 3915 20812 3916 20852
rect 3956 20812 3957 20852
rect 3915 20803 3957 20812
rect 4107 20852 4149 20861
rect 4107 20812 4108 20852
rect 4148 20812 4149 20852
rect 4107 20803 4149 20812
rect 15427 20852 15485 20853
rect 15427 20812 15436 20852
rect 15476 20812 15485 20852
rect 15427 20811 15485 20812
rect 20131 20810 20189 20811
rect 1219 20768 1277 20769
rect 1219 20728 1228 20768
rect 1268 20728 1277 20768
rect 1219 20727 1277 20728
rect 2467 20768 2525 20769
rect 2467 20728 2476 20768
rect 2516 20728 2525 20768
rect 2467 20727 2525 20728
rect 3811 20768 3869 20769
rect 3811 20728 3820 20768
rect 3860 20728 3869 20768
rect 3811 20727 3869 20728
rect 4203 20768 4245 20777
rect 4203 20728 4204 20768
rect 4244 20728 4245 20768
rect 4203 20719 4245 20728
rect 4387 20768 4445 20769
rect 4387 20728 4396 20768
rect 4436 20728 4445 20768
rect 4387 20727 4445 20728
rect 4675 20768 4733 20769
rect 4675 20728 4684 20768
rect 4724 20728 4733 20768
rect 4675 20727 4733 20728
rect 5923 20768 5981 20769
rect 5923 20728 5932 20768
rect 5972 20728 5981 20768
rect 5923 20727 5981 20728
rect 6307 20768 6365 20769
rect 6307 20728 6316 20768
rect 6356 20728 6365 20768
rect 6307 20727 6365 20728
rect 7555 20768 7613 20769
rect 7555 20728 7564 20768
rect 7604 20728 7613 20768
rect 7555 20727 7613 20728
rect 9379 20768 9437 20769
rect 9379 20728 9388 20768
rect 9428 20728 9437 20768
rect 9379 20727 9437 20728
rect 10627 20768 10685 20769
rect 10627 20728 10636 20768
rect 10676 20728 10685 20768
rect 10627 20727 10685 20728
rect 11011 20768 11069 20769
rect 11011 20728 11020 20768
rect 11060 20728 11069 20768
rect 11011 20727 11069 20728
rect 12259 20768 12317 20769
rect 12259 20728 12268 20768
rect 12308 20728 12317 20768
rect 12259 20727 12317 20728
rect 13411 20768 13469 20769
rect 13411 20728 13420 20768
rect 13460 20728 13469 20768
rect 13411 20727 13469 20728
rect 14659 20768 14717 20769
rect 14659 20728 14668 20768
rect 14708 20728 14717 20768
rect 14659 20727 14717 20728
rect 15811 20768 15869 20769
rect 15811 20728 15820 20768
rect 15860 20728 15869 20768
rect 15811 20727 15869 20728
rect 17059 20768 17117 20769
rect 17059 20728 17068 20768
rect 17108 20728 17117 20768
rect 17059 20727 17117 20728
rect 17451 20768 17493 20777
rect 17451 20728 17452 20768
rect 17492 20728 17493 20768
rect 17451 20719 17493 20728
rect 17547 20768 17589 20777
rect 17547 20728 17548 20768
rect 17588 20728 17589 20768
rect 17547 20719 17589 20728
rect 17643 20768 17685 20777
rect 17643 20728 17644 20768
rect 17684 20728 17685 20768
rect 17643 20719 17685 20728
rect 17739 20768 17781 20777
rect 17739 20728 17740 20768
rect 17780 20728 17781 20768
rect 17739 20719 17781 20728
rect 17931 20768 17973 20777
rect 17931 20728 17932 20768
rect 17972 20728 17973 20768
rect 17931 20719 17973 20728
rect 18123 20768 18165 20777
rect 18123 20728 18124 20768
rect 18164 20728 18165 20768
rect 18123 20719 18165 20728
rect 18307 20768 18365 20769
rect 18307 20728 18316 20768
rect 18356 20728 18365 20768
rect 18307 20727 18365 20728
rect 19555 20768 19613 20769
rect 19555 20728 19564 20768
rect 19604 20728 19613 20768
rect 19555 20727 19613 20728
rect 19947 20768 19989 20777
rect 19947 20728 19948 20768
rect 19988 20728 19989 20768
rect 19947 20719 19989 20728
rect 20043 20768 20085 20777
rect 20131 20770 20140 20810
rect 20180 20770 20189 20810
rect 20131 20769 20189 20770
rect 20043 20728 20044 20768
rect 20084 20728 20085 20768
rect 20043 20719 20085 20728
rect 2667 20684 2709 20693
rect 2667 20644 2668 20684
rect 2708 20644 2709 20684
rect 2667 20635 2709 20644
rect 19755 20684 19797 20693
rect 19755 20644 19756 20684
rect 19796 20644 19797 20684
rect 19755 20635 19797 20644
rect 4491 20600 4533 20609
rect 4491 20560 4492 20600
rect 4532 20560 4533 20600
rect 4491 20551 4533 20560
rect 10827 20600 10869 20609
rect 10827 20560 10828 20600
rect 10868 20560 10869 20600
rect 10827 20551 10869 20560
rect 12459 20600 12501 20609
rect 12459 20560 12460 20600
rect 12500 20560 12501 20600
rect 12459 20551 12501 20560
rect 18027 20600 18069 20609
rect 18027 20560 18028 20600
rect 18068 20560 18069 20600
rect 18027 20551 18069 20560
rect 20227 20600 20285 20601
rect 20227 20560 20236 20600
rect 20276 20560 20285 20600
rect 20227 20559 20285 20560
rect 1152 20432 20452 20456
rect 1152 20392 4928 20432
rect 4968 20392 5010 20432
rect 5050 20392 5092 20432
rect 5132 20392 5174 20432
rect 5214 20392 5256 20432
rect 5296 20392 20048 20432
rect 20088 20392 20130 20432
rect 20170 20392 20212 20432
rect 20252 20392 20294 20432
rect 20334 20392 20376 20432
rect 20416 20392 20452 20432
rect 1152 20368 20452 20392
rect 19939 20264 19997 20265
rect 19939 20224 19948 20264
rect 19988 20224 19997 20264
rect 19939 20223 19997 20224
rect 3723 20180 3765 20189
rect 3723 20140 3724 20180
rect 3764 20140 3765 20180
rect 3723 20131 3765 20140
rect 8043 20180 8085 20189
rect 8043 20140 8044 20180
rect 8084 20140 8085 20180
rect 8043 20131 8085 20140
rect 11019 20180 11061 20189
rect 11019 20140 11020 20180
rect 11060 20140 11061 20180
rect 11019 20131 11061 20140
rect 13995 20180 14037 20189
rect 13995 20140 13996 20180
rect 14036 20140 14037 20180
rect 13995 20131 14037 20140
rect 19747 20111 19805 20112
rect 1219 20096 1277 20097
rect 1219 20056 1228 20096
rect 1268 20056 1277 20096
rect 1219 20055 1277 20056
rect 2467 20096 2525 20097
rect 2467 20056 2476 20096
rect 2516 20056 2525 20096
rect 2467 20055 2525 20056
rect 2851 20096 2909 20097
rect 2851 20056 2860 20096
rect 2900 20056 2909 20096
rect 2851 20055 2909 20056
rect 3331 20096 3389 20097
rect 3331 20056 3340 20096
rect 3380 20056 3389 20096
rect 3331 20055 3389 20056
rect 3627 20096 3669 20105
rect 3627 20056 3628 20096
rect 3668 20056 3669 20096
rect 3627 20047 3669 20056
rect 4579 20096 4637 20097
rect 4579 20056 4588 20096
rect 4628 20056 4637 20096
rect 4579 20055 4637 20056
rect 5827 20096 5885 20097
rect 5827 20056 5836 20096
rect 5876 20056 5885 20096
rect 5827 20055 5885 20056
rect 6315 20096 6357 20105
rect 6315 20056 6316 20096
rect 6356 20056 6357 20096
rect 6315 20047 6357 20056
rect 6411 20096 6453 20105
rect 6411 20056 6412 20096
rect 6452 20056 6453 20096
rect 6411 20047 6453 20056
rect 7363 20096 7421 20097
rect 7363 20056 7372 20096
rect 7412 20056 7421 20096
rect 9291 20096 9333 20105
rect 7363 20055 7421 20056
rect 7899 20054 7941 20063
rect 4387 20012 4445 20013
rect 4387 19972 4396 20012
rect 4436 19972 4445 20012
rect 4387 19971 4445 19972
rect 6795 20012 6837 20021
rect 6795 19972 6796 20012
rect 6836 19972 6837 20012
rect 6795 19963 6837 19972
rect 6891 20012 6933 20021
rect 6891 19972 6892 20012
rect 6932 19972 6933 20012
rect 7899 20014 7900 20054
rect 7940 20014 7941 20054
rect 9291 20056 9292 20096
rect 9332 20056 9333 20096
rect 9291 20047 9333 20056
rect 9387 20096 9429 20105
rect 9387 20056 9388 20096
rect 9428 20056 9429 20096
rect 9387 20047 9429 20056
rect 10339 20096 10397 20097
rect 10339 20056 10348 20096
rect 10388 20056 10397 20096
rect 10339 20055 10397 20056
rect 10827 20091 10869 20100
rect 10827 20051 10828 20091
rect 10868 20051 10869 20091
rect 10827 20042 10869 20051
rect 12267 20096 12309 20105
rect 12267 20056 12268 20096
rect 12308 20056 12309 20096
rect 12267 20047 12309 20056
rect 12363 20096 12405 20105
rect 12363 20056 12364 20096
rect 12404 20056 12405 20096
rect 12363 20047 12405 20056
rect 13315 20096 13373 20097
rect 13315 20056 13324 20096
rect 13364 20056 13373 20096
rect 14371 20096 14429 20097
rect 13315 20055 13373 20056
rect 13803 20082 13845 20091
rect 13803 20042 13804 20082
rect 13844 20042 13845 20082
rect 14371 20056 14380 20096
rect 14420 20056 14429 20096
rect 14371 20055 14429 20056
rect 15619 20096 15677 20097
rect 15619 20056 15628 20096
rect 15668 20056 15677 20096
rect 15619 20055 15677 20056
rect 15811 20096 15869 20097
rect 15811 20056 15820 20096
rect 15860 20056 15869 20096
rect 17635 20096 17693 20097
rect 15811 20055 15869 20056
rect 17059 20075 17117 20076
rect 13803 20033 13845 20042
rect 17059 20035 17068 20075
rect 17108 20035 17117 20075
rect 17635 20056 17644 20096
rect 17684 20056 17693 20096
rect 17635 20055 17693 20056
rect 18883 20096 18941 20097
rect 18883 20056 18892 20096
rect 18932 20056 18941 20096
rect 18883 20055 18941 20056
rect 19275 20096 19317 20105
rect 19275 20056 19276 20096
rect 19316 20056 19317 20096
rect 19275 20047 19317 20056
rect 19371 20096 19413 20105
rect 19371 20056 19372 20096
rect 19412 20056 19413 20096
rect 19371 20047 19413 20056
rect 19467 20096 19509 20105
rect 19467 20056 19468 20096
rect 19508 20056 19509 20096
rect 19467 20047 19509 20056
rect 19563 20096 19605 20105
rect 19563 20056 19564 20096
rect 19604 20056 19605 20096
rect 19747 20071 19756 20111
rect 19796 20071 19805 20111
rect 19747 20070 19805 20071
rect 19851 20096 19893 20105
rect 19563 20047 19605 20056
rect 19851 20056 19852 20096
rect 19892 20056 19893 20096
rect 19851 20047 19893 20056
rect 20043 20096 20085 20105
rect 20043 20056 20044 20096
rect 20084 20056 20085 20096
rect 20043 20047 20085 20056
rect 17059 20034 17117 20035
rect 7899 20005 7941 20014
rect 9771 20012 9813 20021
rect 6891 19963 6933 19972
rect 9771 19972 9772 20012
rect 9812 19972 9813 20012
rect 9771 19963 9813 19972
rect 9867 20012 9909 20021
rect 9867 19972 9868 20012
rect 9908 19972 9909 20012
rect 9867 19963 9909 19972
rect 12747 20012 12789 20021
rect 12747 19972 12748 20012
rect 12788 19972 12789 20012
rect 12747 19963 12789 19972
rect 12843 20012 12885 20021
rect 12843 19972 12844 20012
rect 12884 19972 12885 20012
rect 12843 19963 12885 19972
rect 4003 19928 4061 19929
rect 4003 19888 4012 19928
rect 4052 19888 4061 19928
rect 4003 19887 4061 19888
rect 2667 19844 2709 19853
rect 2667 19804 2668 19844
rect 2708 19804 2709 19844
rect 2667 19795 2709 19804
rect 2955 19844 2997 19853
rect 2955 19804 2956 19844
rect 2996 19804 2997 19844
rect 2955 19795 2997 19804
rect 4203 19844 4245 19853
rect 4203 19804 4204 19844
rect 4244 19804 4245 19844
rect 4203 19795 4245 19804
rect 6027 19844 6069 19853
rect 6027 19804 6028 19844
rect 6068 19804 6069 19844
rect 6027 19795 6069 19804
rect 14187 19844 14229 19853
rect 14187 19804 14188 19844
rect 14228 19804 14229 19844
rect 14187 19795 14229 19804
rect 17259 19844 17301 19853
rect 17259 19804 17260 19844
rect 17300 19804 17301 19844
rect 17259 19795 17301 19804
rect 19083 19844 19125 19853
rect 19083 19804 19084 19844
rect 19124 19804 19125 19844
rect 19083 19795 19125 19804
rect 1152 19676 20352 19700
rect 1152 19636 3688 19676
rect 3728 19636 3770 19676
rect 3810 19636 3852 19676
rect 3892 19636 3934 19676
rect 3974 19636 4016 19676
rect 4056 19636 18808 19676
rect 18848 19636 18890 19676
rect 18930 19636 18972 19676
rect 19012 19636 19054 19676
rect 19094 19636 19136 19676
rect 19176 19636 20352 19676
rect 1152 19612 20352 19636
rect 5259 19508 5301 19517
rect 5259 19468 5260 19508
rect 5300 19468 5301 19508
rect 5259 19459 5301 19468
rect 19659 19508 19701 19517
rect 19659 19468 19660 19508
rect 19700 19468 19701 19508
rect 19659 19459 19701 19468
rect 3627 19424 3669 19433
rect 3627 19384 3628 19424
rect 3668 19384 3669 19424
rect 3627 19375 3669 19384
rect 7659 19424 7701 19433
rect 7659 19384 7660 19424
rect 7700 19384 7701 19424
rect 7659 19375 7701 19384
rect 16683 19424 16725 19433
rect 16683 19384 16684 19424
rect 16724 19384 16725 19424
rect 16683 19375 16725 19384
rect 17451 19424 17493 19433
rect 17451 19384 17452 19424
rect 17492 19384 17493 19424
rect 17451 19375 17493 19384
rect 1507 19340 1565 19341
rect 1507 19300 1516 19340
rect 1556 19300 1565 19340
rect 1507 19299 1565 19300
rect 7563 19340 7605 19349
rect 7563 19300 7564 19340
rect 7604 19300 7605 19340
rect 7563 19291 7605 19300
rect 7755 19340 7797 19349
rect 7755 19300 7756 19340
rect 7796 19300 7797 19340
rect 7755 19291 7797 19300
rect 13899 19340 13941 19349
rect 13899 19300 13900 19340
rect 13940 19300 13941 19340
rect 13899 19291 13941 19300
rect 7083 19270 7125 19279
rect 1699 19256 1757 19257
rect 1699 19216 1708 19256
rect 1748 19216 1757 19256
rect 1699 19215 1757 19216
rect 2947 19256 3005 19257
rect 2947 19216 2956 19256
rect 2996 19216 3005 19256
rect 2947 19215 3005 19216
rect 3331 19256 3389 19257
rect 3331 19216 3340 19256
rect 3380 19216 3389 19256
rect 3331 19215 3389 19216
rect 3435 19256 3477 19265
rect 3435 19216 3436 19256
rect 3476 19216 3477 19256
rect 3435 19207 3477 19216
rect 3619 19256 3677 19257
rect 3619 19216 3628 19256
rect 3668 19216 3677 19256
rect 3619 19215 3677 19216
rect 3811 19256 3869 19257
rect 3811 19216 3820 19256
rect 3860 19216 3869 19256
rect 3811 19215 3869 19216
rect 5059 19256 5117 19257
rect 5059 19216 5068 19256
rect 5108 19216 5117 19256
rect 5059 19215 5117 19216
rect 5547 19256 5589 19265
rect 5547 19216 5548 19256
rect 5588 19216 5589 19256
rect 5547 19207 5589 19216
rect 5643 19256 5685 19265
rect 5643 19216 5644 19256
rect 5684 19216 5685 19256
rect 5643 19207 5685 19216
rect 6027 19256 6069 19265
rect 6027 19216 6028 19256
rect 6068 19216 6069 19256
rect 6027 19207 6069 19216
rect 6123 19256 6165 19265
rect 6123 19216 6124 19256
rect 6164 19216 6165 19256
rect 6123 19207 6165 19216
rect 6595 19256 6653 19257
rect 6595 19216 6604 19256
rect 6644 19216 6653 19256
rect 7083 19230 7084 19270
rect 7124 19230 7125 19270
rect 10683 19265 10725 19274
rect 14859 19270 14901 19279
rect 7083 19221 7125 19230
rect 7467 19256 7509 19265
rect 6595 19215 6653 19216
rect 7467 19216 7468 19256
rect 7508 19216 7509 19256
rect 7467 19207 7509 19216
rect 7843 19256 7901 19257
rect 7843 19216 7852 19256
rect 7892 19216 7901 19256
rect 7843 19215 7901 19216
rect 9099 19256 9141 19265
rect 9099 19216 9100 19256
rect 9140 19216 9141 19256
rect 9099 19207 9141 19216
rect 9195 19256 9237 19265
rect 9195 19216 9196 19256
rect 9236 19216 9237 19256
rect 9195 19207 9237 19216
rect 9579 19256 9621 19265
rect 9579 19216 9580 19256
rect 9620 19216 9621 19256
rect 9579 19207 9621 19216
rect 9675 19256 9717 19265
rect 9675 19216 9676 19256
rect 9716 19216 9717 19256
rect 9675 19207 9717 19216
rect 10147 19256 10205 19257
rect 10147 19216 10156 19256
rect 10196 19216 10205 19256
rect 10683 19225 10684 19265
rect 10724 19225 10725 19265
rect 10683 19216 10725 19225
rect 11587 19256 11645 19257
rect 11587 19216 11596 19256
rect 11636 19216 11645 19256
rect 10147 19215 10205 19216
rect 11587 19215 11645 19216
rect 12835 19256 12893 19257
rect 12835 19216 12844 19256
rect 12884 19216 12893 19256
rect 12835 19215 12893 19216
rect 13323 19256 13365 19265
rect 13323 19216 13324 19256
rect 13364 19216 13365 19256
rect 13323 19207 13365 19216
rect 13419 19256 13461 19265
rect 13419 19216 13420 19256
rect 13460 19216 13461 19256
rect 13419 19207 13461 19216
rect 13803 19256 13845 19265
rect 13803 19216 13804 19256
rect 13844 19216 13845 19256
rect 13803 19207 13845 19216
rect 14371 19256 14429 19257
rect 14371 19216 14380 19256
rect 14420 19216 14429 19256
rect 14859 19230 14860 19270
rect 14900 19230 14901 19270
rect 14859 19221 14901 19230
rect 15235 19256 15293 19257
rect 14371 19215 14429 19216
rect 15235 19216 15244 19256
rect 15284 19216 15293 19256
rect 15235 19215 15293 19216
rect 16483 19256 16541 19257
rect 16483 19216 16492 19256
rect 16532 19216 16541 19256
rect 16483 19215 16541 19216
rect 17067 19256 17109 19265
rect 17067 19216 17068 19256
rect 17108 19216 17109 19256
rect 17067 19207 17109 19216
rect 17163 19264 17205 19273
rect 20139 19267 20181 19276
rect 17163 19224 17164 19264
rect 17204 19224 17205 19264
rect 17163 19215 17205 19224
rect 17259 19256 17301 19265
rect 17259 19216 17260 19256
rect 17300 19216 17301 19256
rect 17259 19207 17301 19216
rect 17451 19256 17493 19265
rect 17451 19216 17452 19256
rect 17492 19216 17493 19256
rect 17451 19207 17493 19216
rect 17643 19256 17685 19265
rect 17643 19216 17644 19256
rect 17684 19216 17685 19256
rect 17643 19207 17685 19216
rect 17731 19256 17789 19257
rect 17731 19216 17740 19256
rect 17780 19216 17789 19256
rect 17731 19215 17789 19216
rect 18211 19256 18269 19257
rect 18211 19216 18220 19256
rect 18260 19216 18269 19256
rect 18211 19215 18269 19216
rect 19459 19256 19517 19257
rect 19459 19216 19468 19256
rect 19508 19216 19517 19256
rect 19459 19215 19517 19216
rect 19843 19256 19901 19257
rect 19843 19216 19852 19256
rect 19892 19216 19901 19256
rect 19843 19215 19901 19216
rect 19947 19256 19989 19265
rect 19947 19216 19948 19256
rect 19988 19216 19989 19256
rect 20139 19227 20140 19267
rect 20180 19227 20181 19267
rect 20139 19218 20181 19227
rect 19947 19207 19989 19216
rect 3147 19172 3189 19181
rect 3147 19132 3148 19172
rect 3188 19132 3189 19172
rect 3147 19123 3189 19132
rect 10827 19172 10869 19181
rect 10827 19132 10828 19172
rect 10868 19132 10869 19172
rect 10827 19123 10869 19132
rect 13035 19172 13077 19181
rect 13035 19132 13036 19172
rect 13076 19132 13077 19172
rect 13035 19123 13077 19132
rect 1323 19088 1365 19097
rect 1323 19048 1324 19088
rect 1364 19048 1365 19088
rect 1323 19039 1365 19048
rect 7275 19088 7317 19097
rect 7275 19048 7276 19088
rect 7316 19048 7317 19088
rect 7275 19039 7317 19048
rect 15051 19088 15093 19097
rect 15051 19048 15052 19088
rect 15092 19048 15093 19088
rect 15051 19039 15093 19048
rect 16963 19088 17021 19089
rect 16963 19048 16972 19088
rect 17012 19048 17021 19088
rect 16963 19047 17021 19048
rect 20035 19088 20093 19089
rect 20035 19048 20044 19088
rect 20084 19048 20093 19088
rect 20035 19047 20093 19048
rect 1152 18920 20452 18944
rect 1152 18880 4928 18920
rect 4968 18880 5010 18920
rect 5050 18880 5092 18920
rect 5132 18880 5174 18920
rect 5214 18880 5256 18920
rect 5296 18880 20048 18920
rect 20088 18880 20130 18920
rect 20170 18880 20212 18920
rect 20252 18880 20294 18920
rect 20334 18880 20376 18920
rect 20416 18880 20452 18920
rect 1152 18856 20452 18880
rect 3915 18752 3957 18761
rect 3915 18712 3916 18752
rect 3956 18712 3957 18752
rect 3915 18703 3957 18712
rect 5643 18752 5685 18761
rect 5643 18712 5644 18752
rect 5684 18712 5685 18752
rect 5643 18703 5685 18712
rect 7563 18752 7605 18761
rect 7563 18712 7564 18752
rect 7604 18712 7605 18752
rect 7563 18703 7605 18712
rect 9195 18752 9237 18761
rect 9195 18712 9196 18752
rect 9236 18712 9237 18752
rect 9195 18703 9237 18712
rect 10827 18752 10869 18761
rect 10827 18712 10828 18752
rect 10868 18712 10869 18752
rect 10827 18703 10869 18712
rect 14091 18752 14133 18761
rect 14091 18712 14092 18752
rect 14132 18712 14133 18752
rect 14091 18703 14133 18712
rect 14955 18752 14997 18761
rect 14955 18712 14956 18752
rect 14996 18712 14997 18752
rect 14955 18703 14997 18712
rect 20043 18752 20085 18761
rect 20043 18712 20044 18752
rect 20084 18712 20085 18752
rect 20043 18703 20085 18712
rect 3339 18668 3381 18677
rect 3339 18628 3340 18668
rect 3380 18628 3381 18668
rect 3339 18619 3381 18628
rect 15531 18668 15573 18677
rect 15531 18628 15532 18668
rect 15572 18628 15573 18668
rect 15531 18619 15573 18628
rect 1219 18584 1277 18585
rect 1219 18544 1228 18584
rect 1268 18544 1277 18584
rect 1219 18543 1277 18544
rect 2467 18584 2525 18585
rect 2467 18544 2476 18584
rect 2516 18544 2525 18584
rect 2467 18543 2525 18544
rect 2947 18584 3005 18585
rect 2947 18544 2956 18584
rect 2996 18544 3005 18584
rect 2947 18543 3005 18544
rect 3243 18584 3285 18593
rect 3243 18544 3244 18584
rect 3284 18544 3285 18584
rect 3243 18535 3285 18544
rect 3819 18584 3861 18593
rect 3819 18544 3820 18584
rect 3860 18544 3861 18584
rect 3819 18535 3861 18544
rect 4011 18584 4053 18593
rect 4011 18544 4012 18584
rect 4052 18544 4053 18584
rect 4011 18535 4053 18544
rect 4195 18584 4253 18585
rect 4195 18544 4204 18584
rect 4244 18544 4253 18584
rect 4195 18543 4253 18544
rect 5443 18584 5501 18585
rect 5443 18544 5452 18584
rect 5492 18544 5501 18584
rect 5443 18543 5501 18544
rect 6115 18584 6173 18585
rect 6115 18544 6124 18584
rect 6164 18544 6173 18584
rect 6115 18543 6173 18544
rect 7363 18584 7421 18585
rect 7363 18544 7372 18584
rect 7412 18544 7421 18584
rect 7363 18543 7421 18544
rect 7747 18584 7805 18585
rect 7747 18544 7756 18584
rect 7796 18544 7805 18584
rect 7747 18543 7805 18544
rect 8995 18584 9053 18585
rect 8995 18544 9004 18584
rect 9044 18544 9053 18584
rect 8995 18543 9053 18544
rect 9379 18584 9437 18585
rect 9379 18544 9388 18584
rect 9428 18544 9437 18584
rect 9379 18543 9437 18544
rect 10627 18584 10685 18585
rect 10627 18544 10636 18584
rect 10676 18544 10685 18584
rect 10627 18543 10685 18544
rect 11011 18584 11069 18585
rect 11011 18544 11020 18584
rect 11060 18544 11069 18584
rect 11011 18543 11069 18544
rect 12259 18584 12317 18585
rect 12259 18544 12268 18584
rect 12308 18544 12317 18584
rect 12259 18543 12317 18544
rect 12643 18584 12701 18585
rect 12643 18544 12652 18584
rect 12692 18544 12701 18584
rect 12643 18543 12701 18544
rect 15147 18584 15189 18593
rect 15147 18544 15148 18584
rect 15188 18544 15189 18584
rect 13891 18542 13949 18543
rect 13891 18502 13900 18542
rect 13940 18502 13949 18542
rect 15147 18535 15189 18544
rect 15339 18584 15381 18593
rect 15339 18544 15340 18584
rect 15380 18544 15381 18584
rect 15339 18535 15381 18544
rect 15723 18579 15765 18588
rect 15723 18539 15724 18579
rect 15764 18539 15765 18579
rect 16195 18584 16253 18585
rect 16195 18544 16204 18584
rect 16244 18544 16253 18584
rect 16195 18543 16253 18544
rect 17163 18584 17205 18593
rect 17163 18544 17164 18584
rect 17204 18544 17205 18584
rect 15723 18530 15765 18539
rect 17163 18535 17205 18544
rect 17259 18584 17301 18593
rect 17259 18544 17260 18584
rect 17300 18544 17301 18584
rect 17259 18535 17301 18544
rect 17547 18584 17589 18593
rect 17547 18544 17548 18584
rect 17588 18544 17589 18584
rect 17547 18535 17589 18544
rect 17643 18584 17685 18593
rect 17643 18544 17644 18584
rect 17684 18544 17685 18584
rect 17643 18535 17685 18544
rect 17739 18584 17781 18593
rect 17739 18544 17740 18584
rect 17780 18544 17781 18584
rect 17739 18535 17781 18544
rect 17835 18584 17877 18593
rect 17835 18544 17836 18584
rect 17876 18544 17877 18584
rect 17835 18535 17877 18544
rect 18315 18584 18357 18593
rect 18315 18544 18316 18584
rect 18356 18544 18357 18584
rect 18315 18535 18357 18544
rect 18411 18584 18453 18593
rect 18411 18544 18412 18584
rect 18452 18544 18453 18584
rect 18411 18535 18453 18544
rect 19363 18584 19421 18585
rect 19363 18544 19372 18584
rect 19412 18544 19421 18584
rect 19363 18543 19421 18544
rect 19851 18579 19893 18588
rect 19851 18539 19852 18579
rect 19892 18539 19893 18579
rect 19851 18530 19893 18539
rect 13891 18501 13949 18502
rect 14755 18500 14813 18501
rect 14755 18460 14764 18500
rect 14804 18460 14813 18500
rect 14755 18459 14813 18460
rect 16683 18500 16725 18509
rect 16683 18460 16684 18500
rect 16724 18460 16725 18500
rect 16683 18451 16725 18460
rect 16779 18500 16821 18509
rect 16779 18460 16780 18500
rect 16820 18460 16821 18500
rect 16779 18451 16821 18460
rect 18795 18500 18837 18509
rect 18795 18460 18796 18500
rect 18836 18460 18837 18500
rect 18795 18451 18837 18460
rect 18891 18500 18933 18509
rect 18891 18460 18892 18500
rect 18932 18460 18933 18500
rect 18891 18451 18933 18460
rect 3619 18416 3677 18417
rect 3619 18376 3628 18416
rect 3668 18376 3677 18416
rect 3619 18375 3677 18376
rect 2667 18332 2709 18341
rect 2667 18292 2668 18332
rect 2708 18292 2709 18332
rect 2667 18283 2709 18292
rect 12459 18332 12501 18341
rect 12459 18292 12460 18332
rect 12500 18292 12501 18332
rect 12459 18283 12501 18292
rect 15339 18332 15381 18341
rect 15339 18292 15340 18332
rect 15380 18292 15381 18332
rect 15339 18283 15381 18292
rect 1152 18164 20352 18188
rect 1152 18124 3688 18164
rect 3728 18124 3770 18164
rect 3810 18124 3852 18164
rect 3892 18124 3934 18164
rect 3974 18124 4016 18164
rect 4056 18124 18808 18164
rect 18848 18124 18890 18164
rect 18930 18124 18972 18164
rect 19012 18124 19054 18164
rect 19094 18124 19136 18164
rect 19176 18124 20352 18164
rect 1152 18100 20352 18124
rect 14955 17996 14997 18005
rect 14955 17956 14956 17996
rect 14996 17956 14997 17996
rect 14955 17947 14997 17956
rect 15627 17996 15669 18005
rect 15627 17956 15628 17996
rect 15668 17956 15669 17996
rect 15627 17947 15669 17956
rect 20235 17996 20277 18005
rect 20235 17956 20236 17996
rect 20276 17956 20277 17996
rect 20235 17947 20277 17956
rect 3907 17912 3965 17913
rect 3907 17872 3916 17912
rect 3956 17872 3965 17912
rect 3907 17871 3965 17872
rect 7755 17912 7797 17921
rect 7755 17872 7756 17912
rect 7796 17872 7797 17912
rect 7755 17863 7797 17872
rect 1227 17828 1269 17837
rect 1227 17788 1228 17828
rect 1268 17788 1269 17828
rect 1227 17779 1269 17788
rect 6315 17828 6357 17837
rect 6315 17788 6316 17828
rect 6356 17788 6357 17828
rect 6315 17779 6357 17788
rect 6411 17828 6453 17837
rect 6411 17788 6412 17828
rect 6452 17788 6453 17828
rect 6411 17779 6453 17788
rect 7939 17828 7997 17829
rect 7939 17788 7948 17828
rect 7988 17788 7997 17828
rect 7939 17787 7997 17788
rect 11307 17828 11349 17837
rect 11307 17788 11308 17828
rect 11348 17788 11349 17828
rect 11307 17779 11349 17788
rect 11403 17828 11445 17837
rect 11403 17788 11404 17828
rect 11444 17788 11445 17828
rect 13611 17828 13653 17837
rect 11403 17779 11445 17788
rect 12411 17786 12453 17795
rect 1507 17744 1565 17745
rect 1507 17704 1516 17744
rect 1556 17704 1565 17744
rect 1507 17703 1565 17704
rect 2755 17744 2813 17745
rect 2755 17704 2764 17744
rect 2804 17704 2813 17744
rect 2755 17703 2813 17704
rect 3235 17744 3293 17745
rect 3235 17704 3244 17744
rect 3284 17704 3293 17744
rect 3235 17703 3293 17704
rect 3531 17744 3573 17753
rect 3531 17704 3532 17744
rect 3572 17704 3573 17744
rect 3531 17695 3573 17704
rect 3627 17744 3669 17753
rect 3627 17704 3628 17744
rect 3668 17704 3669 17744
rect 3627 17695 3669 17704
rect 4099 17744 4157 17745
rect 4099 17704 4108 17744
rect 4148 17704 4157 17744
rect 4099 17703 4157 17704
rect 5347 17744 5405 17745
rect 5347 17704 5356 17744
rect 5396 17704 5405 17744
rect 5347 17703 5405 17704
rect 5835 17744 5877 17753
rect 5835 17704 5836 17744
rect 5876 17704 5877 17744
rect 5835 17695 5877 17704
rect 5931 17744 5973 17753
rect 7371 17749 7413 17758
rect 5931 17704 5932 17744
rect 5972 17704 5973 17744
rect 5931 17695 5973 17704
rect 6883 17744 6941 17745
rect 6883 17704 6892 17744
rect 6932 17704 6941 17744
rect 6883 17703 6941 17704
rect 7371 17709 7372 17749
rect 7412 17709 7413 17749
rect 7371 17700 7413 17709
rect 8331 17744 8373 17753
rect 8331 17704 8332 17744
rect 8372 17704 8373 17744
rect 8331 17695 8373 17704
rect 8427 17744 8469 17753
rect 8427 17704 8428 17744
rect 8468 17704 8469 17744
rect 8427 17695 8469 17704
rect 8811 17744 8853 17753
rect 8811 17704 8812 17744
rect 8852 17704 8853 17744
rect 8811 17695 8853 17704
rect 8907 17744 8949 17753
rect 9867 17749 9909 17758
rect 8907 17704 8908 17744
rect 8948 17704 8949 17744
rect 8907 17695 8949 17704
rect 9379 17744 9437 17745
rect 9379 17704 9388 17744
rect 9428 17704 9437 17744
rect 9379 17703 9437 17704
rect 9867 17709 9868 17749
rect 9908 17709 9909 17749
rect 9867 17700 9909 17709
rect 10827 17744 10869 17753
rect 10827 17704 10828 17744
rect 10868 17704 10869 17744
rect 10827 17695 10869 17704
rect 10923 17744 10965 17753
rect 12411 17746 12412 17786
rect 12452 17746 12453 17786
rect 13611 17788 13612 17828
rect 13652 17788 13653 17828
rect 13611 17779 13653 17788
rect 15139 17828 15197 17829
rect 15139 17788 15148 17828
rect 15188 17788 15197 17828
rect 15139 17787 15197 17788
rect 18123 17828 18165 17837
rect 18123 17788 18124 17828
rect 18164 17788 18165 17828
rect 18123 17779 18165 17788
rect 14619 17753 14661 17762
rect 10923 17704 10924 17744
rect 10964 17704 10965 17744
rect 10923 17695 10965 17704
rect 11875 17744 11933 17745
rect 11875 17704 11884 17744
rect 11924 17704 11933 17744
rect 12411 17737 12453 17746
rect 13035 17744 13077 17753
rect 11875 17703 11933 17704
rect 13035 17704 13036 17744
rect 13076 17704 13077 17744
rect 13035 17695 13077 17704
rect 13131 17744 13173 17753
rect 13131 17704 13132 17744
rect 13172 17704 13173 17744
rect 13131 17695 13173 17704
rect 13515 17744 13557 17753
rect 13515 17704 13516 17744
rect 13556 17704 13557 17744
rect 13515 17695 13557 17704
rect 14083 17744 14141 17745
rect 14083 17704 14092 17744
rect 14132 17704 14141 17744
rect 14619 17713 14620 17753
rect 14660 17713 14661 17753
rect 14619 17704 14661 17713
rect 15811 17744 15869 17745
rect 15811 17704 15820 17744
rect 15860 17704 15869 17744
rect 14083 17703 14141 17704
rect 15811 17703 15869 17704
rect 17059 17744 17117 17745
rect 17059 17704 17068 17744
rect 17108 17704 17117 17744
rect 17059 17703 17117 17704
rect 17251 17744 17309 17745
rect 17251 17704 17260 17744
rect 17300 17704 17309 17744
rect 17251 17703 17309 17704
rect 17355 17744 17397 17753
rect 17355 17704 17356 17744
rect 17396 17704 17397 17744
rect 17355 17695 17397 17704
rect 17547 17744 17589 17753
rect 17547 17704 17548 17744
rect 17588 17704 17589 17744
rect 17547 17695 17589 17704
rect 17931 17744 17973 17753
rect 17931 17704 17932 17744
rect 17972 17704 17973 17744
rect 17931 17695 17973 17704
rect 18219 17744 18261 17753
rect 18219 17704 18220 17744
rect 18260 17704 18261 17744
rect 18219 17695 18261 17704
rect 18403 17744 18461 17745
rect 18403 17704 18412 17744
rect 18452 17704 18461 17744
rect 18403 17703 18461 17704
rect 19651 17744 19709 17745
rect 19651 17704 19660 17744
rect 19700 17704 19709 17744
rect 19651 17703 19709 17704
rect 20043 17744 20085 17753
rect 20043 17704 20044 17744
rect 20084 17704 20085 17744
rect 20043 17695 20085 17704
rect 20235 17744 20277 17753
rect 20235 17704 20236 17744
rect 20276 17704 20277 17744
rect 20235 17695 20277 17704
rect 5547 17660 5589 17669
rect 5547 17620 5548 17660
rect 5588 17620 5589 17660
rect 5547 17611 5589 17620
rect 7563 17660 7605 17669
rect 7563 17620 7564 17660
rect 7604 17620 7605 17660
rect 7563 17611 7605 17620
rect 10059 17660 10101 17669
rect 10059 17620 10060 17660
rect 10100 17620 10101 17660
rect 10059 17611 10101 17620
rect 14763 17660 14805 17669
rect 14763 17620 14764 17660
rect 14804 17620 14805 17660
rect 14763 17611 14805 17620
rect 2955 17576 2997 17585
rect 2955 17536 2956 17576
rect 2996 17536 2997 17576
rect 2955 17527 2997 17536
rect 12555 17576 12597 17585
rect 12555 17536 12556 17576
rect 12596 17536 12597 17576
rect 12555 17527 12597 17536
rect 17443 17576 17501 17577
rect 17443 17536 17452 17576
rect 17492 17536 17501 17576
rect 17443 17535 17501 17536
rect 19851 17576 19893 17585
rect 19851 17536 19852 17576
rect 19892 17536 19893 17576
rect 19851 17527 19893 17536
rect 1152 17408 20452 17432
rect 1152 17368 4928 17408
rect 4968 17368 5010 17408
rect 5050 17368 5092 17408
rect 5132 17368 5174 17408
rect 5214 17368 5256 17408
rect 5296 17368 20048 17408
rect 20088 17368 20130 17408
rect 20170 17368 20212 17408
rect 20252 17368 20294 17408
rect 20334 17368 20376 17408
rect 20416 17368 20452 17408
rect 1152 17344 20452 17368
rect 5827 17240 5885 17241
rect 5827 17200 5836 17240
rect 5876 17200 5885 17240
rect 5827 17199 5885 17200
rect 8043 17240 8085 17249
rect 8043 17200 8044 17240
rect 8084 17200 8085 17240
rect 8043 17191 8085 17200
rect 9675 17240 9717 17249
rect 9675 17200 9676 17240
rect 9716 17200 9717 17240
rect 9675 17191 9717 17200
rect 9963 17240 10005 17249
rect 9963 17200 9964 17240
rect 10004 17200 10005 17240
rect 9963 17191 10005 17200
rect 13131 17240 13173 17249
rect 13131 17200 13132 17240
rect 13172 17200 13173 17240
rect 13131 17191 13173 17200
rect 14763 17240 14805 17249
rect 14763 17200 14764 17240
rect 14804 17200 14805 17240
rect 14763 17191 14805 17200
rect 3435 17156 3477 17165
rect 3435 17116 3436 17156
rect 3476 17116 3477 17156
rect 3435 17107 3477 17116
rect 17355 17156 17397 17165
rect 17355 17116 17356 17156
rect 17396 17116 17397 17156
rect 17355 17107 17397 17116
rect 1795 17072 1853 17073
rect 1795 17032 1804 17072
rect 1844 17032 1853 17072
rect 1795 17031 1853 17032
rect 3043 17072 3101 17073
rect 3043 17032 3052 17072
rect 3092 17032 3101 17072
rect 4099 17072 4157 17073
rect 3043 17031 3101 17032
rect 3627 17058 3669 17067
rect 3627 17018 3628 17058
rect 3668 17018 3669 17058
rect 4099 17032 4108 17072
rect 4148 17032 4157 17072
rect 4099 17031 4157 17032
rect 4587 17072 4629 17081
rect 4587 17032 4588 17072
rect 4628 17032 4629 17072
rect 4587 17023 4629 17032
rect 5067 17072 5109 17081
rect 5067 17032 5068 17072
rect 5108 17032 5109 17072
rect 5067 17023 5109 17032
rect 5163 17072 5205 17081
rect 5163 17032 5164 17072
rect 5204 17032 5205 17072
rect 5163 17023 5205 17032
rect 5480 17072 5538 17073
rect 5480 17032 5489 17072
rect 5529 17032 5538 17072
rect 5480 17031 5538 17032
rect 5643 17072 5685 17081
rect 5643 17032 5644 17072
rect 5684 17032 5685 17072
rect 5643 17023 5685 17032
rect 5739 17072 5781 17081
rect 5739 17032 5740 17072
rect 5780 17032 5781 17072
rect 5739 17023 5781 17032
rect 5923 17072 5981 17073
rect 5923 17032 5932 17072
rect 5972 17032 5981 17072
rect 5923 17031 5981 17032
rect 6019 17072 6077 17073
rect 6019 17032 6028 17072
rect 6068 17032 6077 17072
rect 6019 17031 6077 17032
rect 6219 17072 6261 17081
rect 6219 17032 6220 17072
rect 6260 17032 6261 17072
rect 6219 17023 6261 17032
rect 6411 17072 6453 17081
rect 6411 17032 6412 17072
rect 6452 17032 6453 17072
rect 6411 17023 6453 17032
rect 6595 17072 6653 17073
rect 6595 17032 6604 17072
rect 6644 17032 6653 17072
rect 6595 17031 6653 17032
rect 7843 17072 7901 17073
rect 7843 17032 7852 17072
rect 7892 17032 7901 17072
rect 7843 17031 7901 17032
rect 8227 17072 8285 17073
rect 8227 17032 8236 17072
rect 8276 17032 8285 17072
rect 8227 17031 8285 17032
rect 9475 17072 9533 17073
rect 9475 17032 9484 17072
rect 9524 17032 9533 17072
rect 9475 17031 9533 17032
rect 11683 17072 11741 17073
rect 11683 17032 11692 17072
rect 11732 17032 11741 17072
rect 11683 17031 11741 17032
rect 12931 17072 12989 17073
rect 12931 17032 12940 17072
rect 12980 17032 12989 17072
rect 12931 17031 12989 17032
rect 13315 17072 13373 17073
rect 13315 17032 13324 17072
rect 13364 17032 13373 17072
rect 13315 17031 13373 17032
rect 14563 17072 14621 17073
rect 14563 17032 14572 17072
rect 14612 17032 14621 17072
rect 14563 17031 14621 17032
rect 14947 17072 15005 17073
rect 14947 17032 14956 17072
rect 14996 17032 15005 17072
rect 14947 17031 15005 17032
rect 16195 17072 16253 17073
rect 16195 17032 16204 17072
rect 16244 17032 16253 17072
rect 16195 17031 16253 17032
rect 16779 17072 16821 17081
rect 16779 17032 16780 17072
rect 16820 17032 16821 17072
rect 16779 17023 16821 17032
rect 17067 17072 17109 17081
rect 17067 17032 17068 17072
rect 17108 17032 17109 17072
rect 17067 17023 17109 17032
rect 17259 17072 17301 17081
rect 17259 17032 17260 17072
rect 17300 17032 17301 17072
rect 17259 17023 17301 17032
rect 17451 17072 17493 17081
rect 17451 17032 17452 17072
rect 17492 17032 17493 17072
rect 17451 17023 17493 17032
rect 17643 17072 17685 17081
rect 17643 17032 17644 17072
rect 17684 17032 17685 17072
rect 17643 17023 17685 17032
rect 17835 17072 17877 17081
rect 17835 17032 17836 17072
rect 17876 17032 17877 17072
rect 17835 17023 17877 17032
rect 18115 17072 18173 17073
rect 18115 17032 18124 17072
rect 18164 17032 18173 17072
rect 18115 17031 18173 17032
rect 19363 17072 19421 17073
rect 19363 17032 19372 17072
rect 19412 17032 19421 17072
rect 19363 17031 19421 17032
rect 19755 17072 19797 17081
rect 19755 17032 19756 17072
rect 19796 17032 19797 17072
rect 19755 17023 19797 17032
rect 20043 17072 20085 17081
rect 20043 17032 20044 17072
rect 20084 17032 20085 17072
rect 20043 17023 20085 17032
rect 3627 17009 3669 17018
rect 1603 16988 1661 16989
rect 1603 16948 1612 16988
rect 1652 16948 1661 16988
rect 1603 16947 1661 16948
rect 4683 16988 4725 16997
rect 4683 16948 4684 16988
rect 4724 16948 4725 16988
rect 4683 16939 4725 16948
rect 9867 16904 9909 16913
rect 9867 16864 9868 16904
rect 9908 16864 9909 16904
rect 9867 16855 9909 16864
rect 17067 16904 17109 16913
rect 17067 16864 17068 16904
rect 17108 16864 17109 16904
rect 17067 16855 17109 16864
rect 1419 16820 1461 16829
rect 1419 16780 1420 16820
rect 1460 16780 1461 16820
rect 1419 16771 1461 16780
rect 3243 16820 3285 16829
rect 3243 16780 3244 16820
rect 3284 16780 3285 16820
rect 3243 16771 3285 16780
rect 6411 16820 6453 16829
rect 6411 16780 6412 16820
rect 6452 16780 6453 16820
rect 6411 16771 6453 16780
rect 16395 16820 16437 16829
rect 16395 16780 16396 16820
rect 16436 16780 16437 16820
rect 16395 16771 16437 16780
rect 17643 16820 17685 16829
rect 17643 16780 17644 16820
rect 17684 16780 17685 16820
rect 17643 16771 17685 16780
rect 19563 16820 19605 16829
rect 19563 16780 19564 16820
rect 19604 16780 19605 16820
rect 19563 16771 19605 16780
rect 19755 16820 19797 16829
rect 19755 16780 19756 16820
rect 19796 16780 19797 16820
rect 19755 16771 19797 16780
rect 1152 16652 20352 16676
rect 1152 16612 3688 16652
rect 3728 16612 3770 16652
rect 3810 16612 3852 16652
rect 3892 16612 3934 16652
rect 3974 16612 4016 16652
rect 4056 16612 18808 16652
rect 18848 16612 18890 16652
rect 18930 16612 18972 16652
rect 19012 16612 19054 16652
rect 19094 16612 19136 16652
rect 19176 16612 20352 16652
rect 1152 16588 20352 16612
rect 2371 16484 2429 16485
rect 2371 16444 2380 16484
rect 2420 16444 2429 16484
rect 2371 16443 2429 16444
rect 1411 16316 1469 16317
rect 1411 16276 1420 16316
rect 1460 16276 1469 16316
rect 1411 16275 1469 16276
rect 4771 16316 4829 16317
rect 4771 16276 4780 16316
rect 4820 16276 4829 16316
rect 4771 16275 4829 16276
rect 8043 16316 8085 16325
rect 8043 16276 8044 16316
rect 8084 16276 8085 16316
rect 8043 16267 8085 16276
rect 9091 16316 9149 16317
rect 9091 16276 9100 16316
rect 9140 16276 9149 16316
rect 9091 16275 9149 16276
rect 9475 16316 9533 16317
rect 9475 16276 9484 16316
rect 9524 16276 9533 16316
rect 9475 16275 9533 16276
rect 10539 16316 10581 16325
rect 10539 16276 10540 16316
rect 10580 16276 10581 16316
rect 13995 16316 14037 16325
rect 10539 16267 10581 16276
rect 11547 16274 11589 16283
rect 2763 16246 2805 16255
rect 1699 16232 1757 16233
rect 1699 16192 1708 16232
rect 1748 16192 1757 16232
rect 1699 16191 1757 16192
rect 1995 16232 2037 16241
rect 1995 16192 1996 16232
rect 2036 16192 2037 16232
rect 1995 16183 2037 16192
rect 2091 16232 2133 16241
rect 2091 16192 2092 16232
rect 2132 16192 2133 16232
rect 2763 16206 2764 16246
rect 2804 16206 2805 16246
rect 2763 16197 2805 16206
rect 3235 16232 3293 16233
rect 2091 16183 2133 16192
rect 3235 16192 3244 16232
rect 3284 16192 3293 16232
rect 3235 16191 3293 16192
rect 3723 16232 3765 16241
rect 3723 16192 3724 16232
rect 3764 16192 3765 16232
rect 3723 16183 3765 16192
rect 3819 16232 3861 16241
rect 3819 16192 3820 16232
rect 3860 16192 3861 16232
rect 3819 16183 3861 16192
rect 4203 16232 4245 16241
rect 4203 16192 4204 16232
rect 4244 16192 4245 16232
rect 4203 16183 4245 16192
rect 4299 16232 4341 16241
rect 7083 16237 7125 16246
rect 4299 16192 4300 16232
rect 4340 16192 4341 16232
rect 4299 16183 4341 16192
rect 5059 16232 5117 16233
rect 5059 16192 5068 16232
rect 5108 16192 5117 16232
rect 5059 16191 5117 16192
rect 5251 16232 5309 16233
rect 5251 16192 5260 16232
rect 5300 16192 5309 16232
rect 5251 16191 5309 16192
rect 6499 16232 6557 16233
rect 6499 16192 6508 16232
rect 6548 16192 6557 16232
rect 6499 16191 6557 16192
rect 7083 16197 7084 16237
rect 7124 16197 7125 16237
rect 7083 16188 7125 16197
rect 7555 16232 7613 16233
rect 7555 16192 7564 16232
rect 7604 16192 7613 16232
rect 7555 16191 7613 16192
rect 8139 16232 8181 16241
rect 8139 16192 8140 16232
rect 8180 16192 8181 16232
rect 8139 16183 8181 16192
rect 8523 16232 8565 16241
rect 8523 16192 8524 16232
rect 8564 16192 8565 16232
rect 8523 16183 8565 16192
rect 8619 16232 8661 16241
rect 8619 16192 8620 16232
rect 8660 16192 8661 16232
rect 8619 16183 8661 16192
rect 9963 16232 10005 16241
rect 9963 16192 9964 16232
rect 10004 16192 10005 16232
rect 9963 16183 10005 16192
rect 10059 16232 10101 16241
rect 10059 16192 10060 16232
rect 10100 16192 10101 16232
rect 10059 16183 10101 16192
rect 10443 16232 10485 16241
rect 11547 16234 11548 16274
rect 11588 16234 11589 16274
rect 13995 16276 13996 16316
rect 14036 16276 14037 16316
rect 13995 16267 14037 16276
rect 16683 16316 16725 16325
rect 16683 16276 16684 16316
rect 16724 16276 16725 16316
rect 16683 16267 16725 16276
rect 15099 16241 15141 16250
rect 10443 16192 10444 16232
rect 10484 16192 10485 16232
rect 10443 16183 10485 16192
rect 11011 16232 11069 16233
rect 11011 16192 11020 16232
rect 11060 16192 11069 16232
rect 11547 16225 11589 16234
rect 13515 16232 13557 16241
rect 11011 16191 11069 16192
rect 13515 16192 13516 16232
rect 13556 16192 13557 16232
rect 13515 16183 13557 16192
rect 13611 16232 13653 16241
rect 13611 16192 13612 16232
rect 13652 16192 13653 16232
rect 13611 16183 13653 16192
rect 14091 16232 14133 16241
rect 14091 16192 14092 16232
rect 14132 16192 14133 16232
rect 14091 16183 14133 16192
rect 14563 16232 14621 16233
rect 14563 16192 14572 16232
rect 14612 16192 14621 16232
rect 15099 16201 15100 16241
rect 15140 16201 15141 16241
rect 15099 16192 15141 16201
rect 15675 16241 15717 16250
rect 15675 16201 15676 16241
rect 15716 16201 15717 16241
rect 15675 16192 15717 16201
rect 16195 16232 16253 16233
rect 16195 16192 16204 16232
rect 16244 16192 16253 16232
rect 14563 16191 14621 16192
rect 16195 16191 16253 16192
rect 16779 16232 16821 16241
rect 16779 16192 16780 16232
rect 16820 16192 16821 16232
rect 16779 16183 16821 16192
rect 17163 16232 17205 16241
rect 17163 16192 17164 16232
rect 17204 16192 17205 16232
rect 17163 16183 17205 16192
rect 17259 16232 17301 16241
rect 17259 16192 17260 16232
rect 17300 16192 17301 16232
rect 17259 16183 17301 16192
rect 17539 16232 17597 16233
rect 17539 16192 17548 16232
rect 17588 16192 17597 16232
rect 17539 16191 17597 16192
rect 18787 16232 18845 16233
rect 18787 16192 18796 16232
rect 18836 16192 18845 16232
rect 18787 16191 18845 16192
rect 19179 16232 19221 16241
rect 19179 16192 19180 16232
rect 19220 16192 19221 16232
rect 19179 16183 19221 16192
rect 19275 16232 19317 16241
rect 19275 16192 19276 16232
rect 19316 16192 19317 16232
rect 19275 16183 19317 16192
rect 19659 16232 19701 16241
rect 19659 16192 19660 16232
rect 19700 16192 19701 16232
rect 19659 16183 19701 16192
rect 19851 16232 19893 16241
rect 19851 16192 19852 16232
rect 19892 16192 19893 16232
rect 19851 16183 19893 16192
rect 19939 16232 19997 16233
rect 19939 16192 19948 16232
rect 19988 16192 19997 16232
rect 19939 16191 19997 16192
rect 6699 16148 6741 16157
rect 6699 16108 6700 16148
rect 6740 16108 6741 16148
rect 6699 16099 6741 16108
rect 1227 16064 1269 16073
rect 1227 16024 1228 16064
rect 1268 16024 1269 16064
rect 1227 16015 1269 16024
rect 2571 16064 2613 16073
rect 2571 16024 2572 16064
rect 2612 16024 2613 16064
rect 2571 16015 2613 16024
rect 4587 16064 4629 16073
rect 4587 16024 4588 16064
rect 4628 16024 4629 16064
rect 4587 16015 4629 16024
rect 4971 16064 5013 16073
rect 4971 16024 4972 16064
rect 5012 16024 5013 16064
rect 4971 16015 5013 16024
rect 6891 16064 6933 16073
rect 6891 16024 6892 16064
rect 6932 16024 6933 16064
rect 6891 16015 6933 16024
rect 8907 16064 8949 16073
rect 8907 16024 8908 16064
rect 8948 16024 8949 16064
rect 8907 16015 8949 16024
rect 9291 16064 9333 16073
rect 9291 16024 9292 16064
rect 9332 16024 9333 16064
rect 9291 16015 9333 16024
rect 11691 16064 11733 16073
rect 11691 16024 11692 16064
rect 11732 16024 11733 16064
rect 11691 16015 11733 16024
rect 15243 16064 15285 16073
rect 15243 16024 15244 16064
rect 15284 16024 15285 16064
rect 15243 16015 15285 16024
rect 15531 16064 15573 16073
rect 15531 16024 15532 16064
rect 15572 16024 15573 16064
rect 15531 16015 15573 16024
rect 18987 16064 19029 16073
rect 18987 16024 18988 16064
rect 19028 16024 19029 16064
rect 18987 16015 19029 16024
rect 19459 16064 19517 16065
rect 19459 16024 19468 16064
rect 19508 16024 19517 16064
rect 19459 16023 19517 16024
rect 19747 16064 19805 16065
rect 19747 16024 19756 16064
rect 19796 16024 19805 16064
rect 19747 16023 19805 16024
rect 1152 15896 20452 15920
rect 1152 15856 4928 15896
rect 4968 15856 5010 15896
rect 5050 15856 5092 15896
rect 5132 15856 5174 15896
rect 5214 15856 5256 15896
rect 5296 15856 20048 15896
rect 20088 15856 20130 15896
rect 20170 15856 20212 15896
rect 20252 15856 20294 15896
rect 20334 15856 20376 15896
rect 20416 15856 20452 15896
rect 1152 15832 20452 15856
rect 4203 15728 4245 15737
rect 4203 15688 4204 15728
rect 4244 15688 4245 15728
rect 4203 15679 4245 15688
rect 5835 15728 5877 15737
rect 5835 15688 5836 15728
rect 5876 15688 5877 15728
rect 5835 15679 5877 15688
rect 7467 15728 7509 15737
rect 7467 15688 7468 15728
rect 7508 15688 7509 15728
rect 7467 15679 7509 15688
rect 9675 15728 9717 15737
rect 9675 15688 9676 15728
rect 9716 15688 9717 15728
rect 9675 15679 9717 15688
rect 9859 15728 9917 15729
rect 9859 15688 9868 15728
rect 9908 15688 9917 15728
rect 9859 15687 9917 15688
rect 11691 15728 11733 15737
rect 11691 15688 11692 15728
rect 11732 15688 11733 15728
rect 11691 15679 11733 15688
rect 15147 15728 15189 15737
rect 15147 15688 15148 15728
rect 15188 15688 15189 15728
rect 15147 15679 15189 15688
rect 15627 15728 15669 15737
rect 15627 15688 15628 15728
rect 15668 15688 15669 15728
rect 15627 15679 15669 15688
rect 18795 15732 18837 15741
rect 18795 15692 18796 15732
rect 18836 15692 18837 15732
rect 18795 15683 18837 15692
rect 20139 15602 20181 15611
rect 2283 15560 2325 15569
rect 2283 15520 2284 15560
rect 2324 15520 2325 15560
rect 2283 15511 2325 15520
rect 2379 15560 2421 15569
rect 2379 15520 2380 15560
rect 2420 15520 2421 15560
rect 2379 15511 2421 15520
rect 2475 15560 2517 15569
rect 2475 15520 2476 15560
rect 2516 15520 2517 15560
rect 2475 15511 2517 15520
rect 2571 15560 2613 15569
rect 2571 15520 2572 15560
rect 2612 15520 2613 15560
rect 2571 15511 2613 15520
rect 2755 15560 2813 15561
rect 2755 15520 2764 15560
rect 2804 15520 2813 15560
rect 2755 15519 2813 15520
rect 4003 15560 4061 15561
rect 4003 15520 4012 15560
rect 4052 15520 4061 15560
rect 4003 15519 4061 15520
rect 4387 15560 4445 15561
rect 4387 15520 4396 15560
rect 4436 15520 4445 15560
rect 4387 15519 4445 15520
rect 5635 15560 5693 15561
rect 5635 15520 5644 15560
rect 5684 15520 5693 15560
rect 5635 15519 5693 15520
rect 6019 15560 6077 15561
rect 6019 15520 6028 15560
rect 6068 15520 6077 15560
rect 6019 15519 6077 15520
rect 7267 15560 7325 15561
rect 7267 15520 7276 15560
rect 7316 15520 7325 15560
rect 7267 15519 7325 15520
rect 7659 15560 7701 15569
rect 7659 15520 7660 15560
rect 7700 15520 7701 15560
rect 7659 15511 7701 15520
rect 7947 15560 7989 15569
rect 7947 15520 7948 15560
rect 7988 15520 7989 15560
rect 7947 15511 7989 15520
rect 8227 15560 8285 15561
rect 8227 15520 8236 15560
rect 8276 15520 8285 15560
rect 8227 15519 8285 15520
rect 9475 15560 9533 15561
rect 9475 15520 9484 15560
rect 9524 15520 9533 15560
rect 9475 15519 9533 15520
rect 10243 15560 10301 15561
rect 10243 15520 10252 15560
rect 10292 15520 10301 15560
rect 10243 15519 10301 15520
rect 11491 15560 11549 15561
rect 11491 15520 11500 15560
rect 11540 15520 11549 15560
rect 11491 15519 11549 15520
rect 11971 15560 12029 15561
rect 11971 15520 11980 15560
rect 12020 15520 12029 15560
rect 11971 15519 12029 15520
rect 13219 15560 13277 15561
rect 13219 15520 13228 15560
rect 13268 15520 13277 15560
rect 13219 15519 13277 15520
rect 13699 15560 13757 15561
rect 13699 15520 13708 15560
rect 13748 15520 13757 15560
rect 13699 15519 13757 15520
rect 14947 15560 15005 15561
rect 14947 15520 14956 15560
rect 14996 15520 15005 15560
rect 14947 15519 15005 15520
rect 15811 15560 15869 15561
rect 15811 15520 15820 15560
rect 15860 15520 15869 15560
rect 15811 15519 15869 15520
rect 17059 15560 17117 15561
rect 17059 15520 17068 15560
rect 17108 15520 17117 15560
rect 17059 15519 17117 15520
rect 17355 15560 17397 15569
rect 17355 15520 17356 15560
rect 17396 15520 17397 15560
rect 17355 15511 17397 15520
rect 17451 15560 17493 15569
rect 17451 15520 17452 15560
rect 17492 15520 17493 15560
rect 17451 15511 17493 15520
rect 17547 15560 17589 15569
rect 17547 15520 17548 15560
rect 17588 15520 17589 15560
rect 17547 15511 17589 15520
rect 17643 15560 17685 15569
rect 17643 15520 17644 15560
rect 17684 15520 17685 15560
rect 17643 15511 17685 15520
rect 17835 15560 17877 15569
rect 17835 15520 17836 15560
rect 17876 15520 17877 15560
rect 17835 15511 17877 15520
rect 18123 15560 18165 15569
rect 18123 15520 18124 15560
rect 18164 15520 18165 15560
rect 18123 15511 18165 15520
rect 18603 15560 18645 15569
rect 18603 15520 18604 15560
rect 18644 15520 18645 15560
rect 18603 15511 18645 15520
rect 18691 15560 18749 15561
rect 18691 15520 18700 15560
rect 18740 15520 18749 15560
rect 18691 15519 18749 15520
rect 19075 15560 19133 15561
rect 19075 15520 19084 15560
rect 19124 15520 19133 15560
rect 19075 15519 19133 15520
rect 19371 15560 19413 15569
rect 19371 15520 19372 15560
rect 19412 15520 19413 15560
rect 19371 15511 19413 15520
rect 19467 15560 19509 15569
rect 19467 15520 19468 15560
rect 19508 15520 19509 15560
rect 19467 15511 19509 15520
rect 19947 15560 19989 15569
rect 19947 15520 19948 15560
rect 19988 15520 19989 15560
rect 20139 15562 20140 15602
rect 20180 15562 20181 15602
rect 20139 15553 20181 15562
rect 20227 15560 20285 15561
rect 19947 15511 19989 15520
rect 20227 15520 20236 15560
rect 20276 15520 20285 15560
rect 20227 15519 20285 15520
rect 1699 15476 1757 15477
rect 1699 15436 1708 15476
rect 1748 15436 1757 15476
rect 1699 15435 1757 15436
rect 2083 15476 2141 15477
rect 2083 15436 2092 15476
rect 2132 15436 2141 15476
rect 2083 15435 2141 15436
rect 1323 15392 1365 15401
rect 1323 15352 1324 15392
rect 1364 15352 1365 15392
rect 1323 15343 1365 15352
rect 1515 15392 1557 15401
rect 1515 15352 1516 15392
rect 1556 15352 1557 15392
rect 1515 15343 1557 15352
rect 13419 15392 13461 15401
rect 13419 15352 13420 15392
rect 13460 15352 13461 15392
rect 13419 15343 13461 15352
rect 19747 15392 19805 15393
rect 19747 15352 19756 15392
rect 19796 15352 19805 15392
rect 19747 15351 19805 15352
rect 1899 15308 1941 15317
rect 1899 15268 1900 15308
rect 1940 15268 1941 15308
rect 1899 15259 1941 15268
rect 7659 15308 7701 15317
rect 7659 15268 7660 15308
rect 7700 15268 7701 15308
rect 7659 15259 7701 15268
rect 18123 15308 18165 15317
rect 18123 15268 18124 15308
rect 18164 15268 18165 15308
rect 18123 15259 18165 15268
rect 18315 15308 18357 15317
rect 18315 15268 18316 15308
rect 18356 15268 18357 15308
rect 18315 15259 18357 15268
rect 19947 15308 19989 15317
rect 19947 15268 19948 15308
rect 19988 15268 19989 15308
rect 19947 15259 19989 15268
rect 1152 15140 20352 15164
rect 1152 15100 3688 15140
rect 3728 15100 3770 15140
rect 3810 15100 3852 15140
rect 3892 15100 3934 15140
rect 3974 15100 4016 15140
rect 4056 15100 18808 15140
rect 18848 15100 18890 15140
rect 18930 15100 18972 15140
rect 19012 15100 19054 15140
rect 19094 15100 19136 15140
rect 19176 15100 20352 15140
rect 1152 15076 20352 15100
rect 2667 14972 2709 14981
rect 2667 14932 2668 14972
rect 2708 14932 2709 14972
rect 2667 14923 2709 14932
rect 6027 14972 6069 14981
rect 6027 14932 6028 14972
rect 6068 14932 6069 14972
rect 6027 14923 6069 14932
rect 7659 14972 7701 14981
rect 7659 14932 7660 14972
rect 7700 14932 7701 14972
rect 7659 14923 7701 14932
rect 9867 14888 9909 14897
rect 9867 14848 9868 14888
rect 9908 14848 9909 14888
rect 9867 14839 9909 14848
rect 18891 14888 18933 14897
rect 18891 14848 18892 14888
rect 18932 14848 18933 14888
rect 18891 14839 18933 14848
rect 19755 14888 19797 14897
rect 19755 14848 19756 14888
rect 19796 14848 19797 14888
rect 19755 14839 19797 14848
rect 3043 14804 3101 14805
rect 3043 14764 3052 14804
rect 3092 14764 3101 14804
rect 3043 14763 3101 14764
rect 3915 14804 3957 14813
rect 3915 14764 3916 14804
rect 3956 14764 3957 14804
rect 3915 14755 3957 14764
rect 4011 14804 4053 14813
rect 4011 14764 4012 14804
rect 4052 14764 4053 14804
rect 4011 14755 4053 14764
rect 12555 14804 12597 14813
rect 12555 14764 12556 14804
rect 12596 14764 12597 14804
rect 12555 14755 12597 14764
rect 12651 14804 12693 14813
rect 12651 14764 12652 14804
rect 12692 14764 12693 14804
rect 12651 14755 12693 14764
rect 18795 14804 18837 14813
rect 18795 14764 18796 14804
rect 18836 14764 18837 14804
rect 18795 14755 18837 14764
rect 18987 14804 19029 14813
rect 18987 14764 18988 14804
rect 19028 14764 19029 14804
rect 18987 14755 19029 14764
rect 1219 14720 1277 14721
rect 1219 14680 1228 14720
rect 1268 14680 1277 14720
rect 1219 14679 1277 14680
rect 2467 14720 2525 14721
rect 2467 14680 2476 14720
rect 2516 14680 2525 14720
rect 2467 14679 2525 14680
rect 3435 14720 3477 14729
rect 3435 14680 3436 14720
rect 3476 14680 3477 14720
rect 3435 14671 3477 14680
rect 3531 14720 3573 14729
rect 4971 14725 5013 14734
rect 3531 14680 3532 14720
rect 3572 14680 3573 14720
rect 3531 14671 3573 14680
rect 4483 14720 4541 14721
rect 4483 14680 4492 14720
rect 4532 14680 4541 14720
rect 4483 14679 4541 14680
rect 4971 14685 4972 14725
rect 5012 14685 5013 14725
rect 4971 14676 5013 14685
rect 5547 14720 5589 14729
rect 5547 14680 5548 14720
rect 5588 14680 5589 14720
rect 5547 14671 5589 14680
rect 5643 14720 5685 14729
rect 5643 14680 5644 14720
rect 5684 14680 5685 14720
rect 5643 14671 5685 14680
rect 5739 14720 5781 14729
rect 5739 14680 5740 14720
rect 5780 14680 5781 14720
rect 5739 14671 5781 14680
rect 5923 14720 5981 14721
rect 5923 14680 5932 14720
rect 5972 14680 5981 14720
rect 5923 14679 5981 14680
rect 6211 14720 6269 14721
rect 6211 14680 6220 14720
rect 6260 14680 6269 14720
rect 6211 14679 6269 14680
rect 7459 14720 7517 14721
rect 7459 14680 7468 14720
rect 7508 14680 7517 14720
rect 7459 14679 7517 14680
rect 7947 14720 7989 14729
rect 7947 14680 7948 14720
rect 7988 14680 7989 14720
rect 7947 14671 7989 14680
rect 8043 14720 8085 14729
rect 8043 14680 8044 14720
rect 8084 14680 8085 14720
rect 8043 14671 8085 14680
rect 8427 14720 8469 14729
rect 8427 14680 8428 14720
rect 8468 14680 8469 14720
rect 8427 14671 8469 14680
rect 8523 14720 8565 14729
rect 9483 14725 9525 14734
rect 8523 14680 8524 14720
rect 8564 14680 8565 14720
rect 8523 14671 8565 14680
rect 8995 14720 9053 14721
rect 8995 14680 9004 14720
rect 9044 14680 9053 14720
rect 8995 14679 9053 14680
rect 9483 14685 9484 14725
rect 9524 14685 9525 14725
rect 9483 14676 9525 14685
rect 10339 14720 10397 14721
rect 10339 14680 10348 14720
rect 10388 14680 10397 14720
rect 10339 14679 10397 14680
rect 11587 14720 11645 14721
rect 11587 14680 11596 14720
rect 11636 14680 11645 14720
rect 11587 14679 11645 14680
rect 12075 14720 12117 14729
rect 12075 14680 12076 14720
rect 12116 14680 12117 14720
rect 12075 14671 12117 14680
rect 12171 14720 12213 14729
rect 13611 14725 13653 14734
rect 12171 14680 12172 14720
rect 12212 14680 12213 14720
rect 12171 14671 12213 14680
rect 13123 14720 13181 14721
rect 13123 14680 13132 14720
rect 13172 14680 13181 14720
rect 13123 14679 13181 14680
rect 13611 14685 13612 14725
rect 13652 14685 13653 14725
rect 13611 14676 13653 14685
rect 15627 14725 15669 14734
rect 15627 14685 15628 14725
rect 15668 14685 15669 14725
rect 15627 14676 15669 14685
rect 16099 14720 16157 14721
rect 16099 14680 16108 14720
rect 16148 14680 16157 14720
rect 16099 14679 16157 14680
rect 16587 14720 16629 14729
rect 16587 14680 16588 14720
rect 16628 14680 16629 14720
rect 16587 14671 16629 14680
rect 16683 14720 16725 14729
rect 16683 14680 16684 14720
rect 16724 14680 16725 14720
rect 16683 14671 16725 14680
rect 17067 14720 17109 14729
rect 17067 14680 17068 14720
rect 17108 14680 17109 14720
rect 17067 14671 17109 14680
rect 17163 14720 17205 14729
rect 17163 14680 17164 14720
rect 17204 14680 17205 14720
rect 17163 14671 17205 14680
rect 17739 14720 17781 14729
rect 17739 14680 17740 14720
rect 17780 14680 17781 14720
rect 17739 14671 17781 14680
rect 17835 14720 17877 14729
rect 17835 14680 17836 14720
rect 17876 14680 17877 14720
rect 17835 14671 17877 14680
rect 17931 14720 17973 14729
rect 17931 14680 17932 14720
rect 17972 14680 17973 14720
rect 17931 14671 17973 14680
rect 18219 14720 18261 14729
rect 18219 14680 18220 14720
rect 18260 14680 18261 14720
rect 18219 14671 18261 14680
rect 18315 14720 18357 14729
rect 18315 14680 18316 14720
rect 18356 14680 18357 14720
rect 18315 14671 18357 14680
rect 18411 14720 18453 14729
rect 18411 14680 18412 14720
rect 18452 14680 18453 14720
rect 18411 14671 18453 14680
rect 18691 14720 18749 14721
rect 18691 14680 18700 14720
rect 18740 14680 18749 14720
rect 18691 14679 18749 14680
rect 19083 14720 19125 14729
rect 19083 14680 19084 14720
rect 19124 14680 19125 14720
rect 19083 14671 19125 14680
rect 19275 14720 19317 14729
rect 19275 14680 19276 14720
rect 19316 14680 19317 14720
rect 19275 14671 19317 14680
rect 19371 14720 19413 14729
rect 19371 14680 19372 14720
rect 19412 14680 19413 14720
rect 19371 14671 19413 14680
rect 19467 14720 19509 14729
rect 19467 14680 19468 14720
rect 19508 14680 19509 14720
rect 19467 14671 19509 14680
rect 19563 14720 19605 14729
rect 19563 14680 19564 14720
rect 19604 14680 19605 14720
rect 19947 14720 19989 14729
rect 19563 14671 19605 14680
rect 19755 14678 19797 14687
rect 5163 14636 5205 14645
rect 5163 14596 5164 14636
rect 5204 14596 5205 14636
rect 19755 14638 19756 14678
rect 19796 14638 19797 14678
rect 19947 14680 19948 14720
rect 19988 14680 19989 14720
rect 19947 14671 19989 14680
rect 20035 14720 20093 14721
rect 20035 14680 20044 14720
rect 20084 14680 20093 14720
rect 20035 14679 20093 14680
rect 19755 14629 19797 14638
rect 5163 14587 5205 14596
rect 2859 14552 2901 14561
rect 2859 14512 2860 14552
rect 2900 14512 2901 14552
rect 2859 14503 2901 14512
rect 5443 14552 5501 14553
rect 5443 14512 5452 14552
rect 5492 14512 5501 14552
rect 5443 14511 5501 14512
rect 9675 14552 9717 14561
rect 9675 14512 9676 14552
rect 9716 14512 9717 14552
rect 9675 14503 9717 14512
rect 11787 14552 11829 14561
rect 11787 14512 11788 14552
rect 11828 14512 11829 14552
rect 11787 14503 11829 14512
rect 13803 14552 13845 14561
rect 13803 14512 13804 14552
rect 13844 14512 13845 14552
rect 13803 14503 13845 14512
rect 15435 14552 15477 14561
rect 15435 14512 15436 14552
rect 15476 14512 15477 14552
rect 15435 14503 15477 14512
rect 18019 14552 18077 14553
rect 18019 14512 18028 14552
rect 18068 14512 18077 14552
rect 18019 14511 18077 14512
rect 18499 14552 18557 14553
rect 18499 14512 18508 14552
rect 18548 14512 18557 14552
rect 18499 14511 18557 14512
rect 1152 14384 20452 14408
rect 1152 14344 4928 14384
rect 4968 14344 5010 14384
rect 5050 14344 5092 14384
rect 5132 14344 5174 14384
rect 5214 14344 5256 14384
rect 5296 14344 20048 14384
rect 20088 14344 20130 14384
rect 20170 14344 20212 14384
rect 20252 14344 20294 14384
rect 20334 14344 20376 14384
rect 20416 14344 20452 14384
rect 1152 14320 20452 14344
rect 1227 14216 1269 14225
rect 1227 14176 1228 14216
rect 1268 14176 1269 14216
rect 1227 14167 1269 14176
rect 9195 14216 9237 14225
rect 9195 14176 9196 14216
rect 9236 14176 9237 14216
rect 9195 14167 9237 14176
rect 11211 14216 11253 14225
rect 11211 14176 11212 14216
rect 11252 14176 11253 14216
rect 11211 14167 11253 14176
rect 11403 14216 11445 14225
rect 11403 14176 11404 14216
rect 11444 14176 11445 14216
rect 11403 14167 11445 14176
rect 16203 14216 16245 14225
rect 16203 14176 16204 14216
rect 16244 14176 16245 14216
rect 16203 14167 16245 14176
rect 1707 14132 1749 14141
rect 1707 14092 1708 14132
rect 1748 14092 1749 14132
rect 1707 14083 1749 14092
rect 2379 14132 2421 14141
rect 2379 14092 2380 14132
rect 2420 14092 2421 14132
rect 2379 14083 2421 14092
rect 2571 14132 2613 14141
rect 2571 14092 2572 14132
rect 2612 14092 2613 14132
rect 2571 14083 2613 14092
rect 7467 14132 7509 14141
rect 7467 14092 7468 14132
rect 7508 14092 7509 14132
rect 7467 14083 7509 14092
rect 14379 14132 14421 14141
rect 14379 14092 14380 14132
rect 14420 14092 14421 14132
rect 14379 14083 14421 14092
rect 16011 14132 16053 14141
rect 16011 14092 16012 14132
rect 16052 14092 16053 14132
rect 16011 14083 16053 14092
rect 20139 14132 20181 14141
rect 20139 14092 20140 14132
rect 20180 14092 20181 14132
rect 20139 14083 20181 14092
rect 1611 14048 1653 14057
rect 1611 14008 1612 14048
rect 1652 14008 1653 14048
rect 1611 13999 1653 14008
rect 1803 14048 1845 14057
rect 1803 14008 1804 14048
rect 1844 14008 1845 14048
rect 1803 13999 1845 14008
rect 1891 14048 1949 14049
rect 1891 14008 1900 14048
rect 1940 14008 1949 14048
rect 1891 14007 1949 14008
rect 2091 14048 2133 14057
rect 2091 14008 2092 14048
rect 2132 14008 2133 14048
rect 2091 13999 2133 14008
rect 2283 14040 2325 14049
rect 3235 14048 3293 14049
rect 2179 14006 2237 14007
rect 2179 13966 2188 14006
rect 2228 13966 2237 14006
rect 2283 14000 2284 14040
rect 2324 14000 2325 14040
rect 2283 13991 2325 14000
rect 2763 14034 2805 14043
rect 2763 13994 2764 14034
rect 2804 13994 2805 14034
rect 3235 14008 3244 14048
rect 3284 14008 3293 14048
rect 3235 14007 3293 14008
rect 3819 14048 3861 14057
rect 3819 14008 3820 14048
rect 3860 14008 3861 14048
rect 3819 13999 3861 14008
rect 4203 14048 4245 14057
rect 4203 14008 4204 14048
rect 4244 14008 4245 14048
rect 4203 13999 4245 14008
rect 4299 14048 4341 14057
rect 4299 14008 4300 14048
rect 4340 14008 4341 14048
rect 4299 13999 4341 14008
rect 4675 14048 4733 14049
rect 4675 14008 4684 14048
rect 4724 14008 4733 14048
rect 4675 14007 4733 14008
rect 4779 14048 4821 14057
rect 4779 14008 4780 14048
rect 4820 14008 4821 14048
rect 4779 13999 4821 14008
rect 4971 14048 5013 14057
rect 4971 14008 4972 14048
rect 5012 14008 5013 14048
rect 4971 13999 5013 14008
rect 5163 14048 5205 14057
rect 5163 14008 5164 14048
rect 5204 14008 5205 14048
rect 5163 13999 5205 14008
rect 5259 14048 5301 14057
rect 5259 14008 5260 14048
rect 5300 14008 5301 14048
rect 5259 13999 5301 14008
rect 5355 14048 5397 14057
rect 5355 14008 5356 14048
rect 5396 14008 5397 14048
rect 5355 13999 5397 14008
rect 5451 14048 5493 14057
rect 5451 14008 5452 14048
rect 5492 14008 5493 14048
rect 5451 13999 5493 14008
rect 5739 14048 5781 14057
rect 5739 14008 5740 14048
rect 5780 14008 5781 14048
rect 5739 13999 5781 14008
rect 5835 14048 5877 14057
rect 5835 14008 5836 14048
rect 5876 14008 5877 14048
rect 5835 13999 5877 14008
rect 6787 14048 6845 14049
rect 6787 14008 6796 14048
rect 6836 14008 6845 14048
rect 6787 14007 6845 14008
rect 7275 14043 7317 14052
rect 7275 14003 7276 14043
rect 7316 14003 7317 14043
rect 7747 14048 7805 14049
rect 7747 14008 7756 14048
rect 7796 14008 7805 14048
rect 7747 14007 7805 14008
rect 8995 14048 9053 14049
rect 8995 14008 9004 14048
rect 9044 14008 9053 14048
rect 8995 14007 9053 14008
rect 9483 14048 9525 14057
rect 9483 14008 9484 14048
rect 9524 14008 9525 14048
rect 7275 13994 7317 14003
rect 9483 13999 9525 14008
rect 9579 14048 9621 14057
rect 9579 14008 9580 14048
rect 9620 14008 9621 14048
rect 9579 13999 9621 14008
rect 9963 14048 10005 14057
rect 9963 14008 9964 14048
rect 10004 14008 10005 14048
rect 9963 13999 10005 14008
rect 10059 14048 10101 14057
rect 10059 14008 10060 14048
rect 10100 14008 10101 14048
rect 10059 13999 10101 14008
rect 10531 14048 10589 14049
rect 10531 14008 10540 14048
rect 10580 14008 10589 14048
rect 12651 14048 12693 14057
rect 10531 14007 10589 14008
rect 11067 14038 11109 14047
rect 11067 13998 11068 14038
rect 11108 13998 11109 14038
rect 12651 14008 12652 14048
rect 12692 14008 12693 14048
rect 12651 13999 12693 14008
rect 12747 14048 12789 14057
rect 12747 14008 12748 14048
rect 12788 14008 12789 14048
rect 12747 13999 12789 14008
rect 13131 14048 13173 14057
rect 13131 14008 13132 14048
rect 13172 14008 13173 14048
rect 13131 13999 13173 14008
rect 13699 14048 13757 14049
rect 13699 14008 13708 14048
rect 13748 14008 13757 14048
rect 14563 14048 14621 14049
rect 13699 14007 13757 14008
rect 14187 14034 14229 14043
rect 2763 13985 2805 13994
rect 11067 13989 11109 13998
rect 14187 13994 14188 14034
rect 14228 13994 14229 14034
rect 14563 14008 14572 14048
rect 14612 14008 14621 14048
rect 14563 14007 14621 14008
rect 15811 14048 15869 14049
rect 15811 14008 15820 14048
rect 15860 14008 15869 14048
rect 15811 14007 15869 14008
rect 16387 14048 16445 14049
rect 16387 14008 16396 14048
rect 16436 14008 16445 14048
rect 16387 14007 16445 14008
rect 17635 14048 17693 14049
rect 17635 14008 17644 14048
rect 17684 14008 17693 14048
rect 17635 14007 17693 14008
rect 17827 14048 17885 14049
rect 17827 14008 17836 14048
rect 17876 14008 17885 14048
rect 17827 14007 17885 14008
rect 19075 14048 19133 14049
rect 19075 14008 19084 14048
rect 19124 14008 19133 14048
rect 19075 14007 19133 14008
rect 19459 14048 19517 14049
rect 19459 14008 19468 14048
rect 19508 14008 19517 14048
rect 19459 14007 19517 14008
rect 19851 14048 19893 14057
rect 19851 14008 19852 14048
rect 19892 14008 19893 14048
rect 19851 13999 19893 14008
rect 20035 14048 20093 14049
rect 20035 14008 20044 14048
rect 20084 14008 20093 14048
rect 20035 14007 20093 14008
rect 20235 14048 20277 14057
rect 20235 14008 20236 14048
rect 20276 14008 20277 14048
rect 20235 13999 20277 14008
rect 14187 13985 14229 13994
rect 2179 13965 2237 13966
rect 1411 13964 1469 13965
rect 1411 13924 1420 13964
rect 1460 13924 1469 13964
rect 1411 13923 1469 13924
rect 3723 13964 3765 13973
rect 3723 13924 3724 13964
rect 3764 13924 3765 13964
rect 3723 13915 3765 13924
rect 6219 13964 6261 13973
rect 6219 13924 6220 13964
rect 6260 13924 6261 13964
rect 6219 13915 6261 13924
rect 6315 13964 6357 13973
rect 6315 13924 6316 13964
rect 6356 13924 6357 13964
rect 6315 13915 6357 13924
rect 11587 13964 11645 13965
rect 11587 13924 11596 13964
rect 11636 13924 11645 13964
rect 11587 13923 11645 13924
rect 11971 13964 12029 13965
rect 11971 13924 11980 13964
rect 12020 13924 12029 13964
rect 11971 13923 12029 13924
rect 12355 13964 12413 13965
rect 12355 13924 12364 13964
rect 12404 13924 12413 13964
rect 12355 13923 12413 13924
rect 13227 13964 13269 13973
rect 13227 13924 13228 13964
rect 13268 13924 13269 13964
rect 13227 13915 13269 13924
rect 19563 13964 19605 13973
rect 19563 13924 19564 13964
rect 19604 13924 19605 13964
rect 19563 13915 19605 13924
rect 19755 13964 19797 13973
rect 19755 13924 19756 13964
rect 19796 13924 19797 13964
rect 19755 13915 19797 13924
rect 11787 13880 11829 13889
rect 11787 13840 11788 13880
rect 11828 13840 11829 13880
rect 11787 13831 11829 13840
rect 12171 13880 12213 13889
rect 12171 13840 12172 13880
rect 12212 13840 12213 13880
rect 12171 13831 12213 13840
rect 19275 13880 19317 13889
rect 19275 13840 19276 13880
rect 19316 13840 19317 13880
rect 19275 13831 19317 13840
rect 19659 13880 19701 13889
rect 19659 13840 19660 13880
rect 19700 13840 19701 13880
rect 19659 13831 19701 13840
rect 4971 13796 5013 13805
rect 4971 13756 4972 13796
rect 5012 13756 5013 13796
rect 4971 13747 5013 13756
rect 1152 13628 20352 13652
rect 1152 13588 3688 13628
rect 3728 13588 3770 13628
rect 3810 13588 3852 13628
rect 3892 13588 3934 13628
rect 3974 13588 4016 13628
rect 4056 13588 18808 13628
rect 18848 13588 18890 13628
rect 18930 13588 18972 13628
rect 19012 13588 19054 13628
rect 19094 13588 19136 13628
rect 19176 13588 20352 13628
rect 1152 13564 20352 13588
rect 1227 13460 1269 13469
rect 1227 13420 1228 13460
rect 1268 13420 1269 13460
rect 1227 13411 1269 13420
rect 3147 13460 3189 13469
rect 3147 13420 3148 13460
rect 3188 13420 3189 13460
rect 3147 13411 3189 13420
rect 5739 13460 5781 13469
rect 5739 13420 5740 13460
rect 5780 13420 5781 13460
rect 5739 13411 5781 13420
rect 7371 13460 7413 13469
rect 7371 13420 7372 13460
rect 7412 13420 7413 13460
rect 7371 13411 7413 13420
rect 9579 13460 9621 13469
rect 9579 13420 9580 13460
rect 9620 13420 9621 13460
rect 9579 13411 9621 13420
rect 11307 13460 11349 13469
rect 11307 13420 11308 13460
rect 11348 13420 11349 13460
rect 11307 13411 11349 13420
rect 13419 13460 13461 13469
rect 13419 13420 13420 13460
rect 13460 13420 13461 13460
rect 13419 13411 13461 13420
rect 18603 13460 18645 13469
rect 18603 13420 18604 13460
rect 18644 13420 18645 13460
rect 18603 13411 18645 13420
rect 19843 13376 19901 13377
rect 19843 13336 19852 13376
rect 19892 13336 19901 13376
rect 19843 13335 19901 13336
rect 3523 13303 3581 13304
rect 1411 13292 1469 13293
rect 1411 13252 1420 13292
rect 1460 13252 1469 13292
rect 3523 13263 3532 13303
rect 3572 13263 3581 13303
rect 3523 13262 3581 13263
rect 3907 13292 3965 13293
rect 1411 13251 1469 13252
rect 3907 13252 3916 13292
rect 3956 13252 3965 13292
rect 3907 13251 3965 13252
rect 11683 13292 11741 13293
rect 11683 13252 11692 13292
rect 11732 13252 11741 13292
rect 11683 13251 11741 13252
rect 13219 13250 13277 13251
rect 1699 13208 1757 13209
rect 1699 13168 1708 13208
rect 1748 13168 1757 13208
rect 1699 13167 1757 13168
rect 2947 13208 3005 13209
rect 2947 13168 2956 13208
rect 2996 13168 3005 13208
rect 2947 13167 3005 13168
rect 4291 13208 4349 13209
rect 4291 13168 4300 13208
rect 4340 13168 4349 13208
rect 4291 13167 4349 13168
rect 5539 13208 5597 13209
rect 5539 13168 5548 13208
rect 5588 13168 5597 13208
rect 5539 13167 5597 13168
rect 5923 13208 5981 13209
rect 5923 13168 5932 13208
rect 5972 13168 5981 13208
rect 5923 13167 5981 13168
rect 7171 13208 7229 13209
rect 7171 13168 7180 13208
rect 7220 13168 7229 13208
rect 7171 13167 7229 13168
rect 7563 13208 7605 13217
rect 7563 13168 7564 13208
rect 7604 13168 7605 13208
rect 7563 13159 7605 13168
rect 7755 13208 7797 13217
rect 13219 13210 13228 13250
rect 13268 13210 13277 13250
rect 13219 13209 13277 13210
rect 7755 13168 7756 13208
rect 7796 13168 7797 13208
rect 7755 13159 7797 13168
rect 7843 13208 7901 13209
rect 7843 13168 7852 13208
rect 7892 13168 7901 13208
rect 7843 13167 7901 13168
rect 8131 13208 8189 13209
rect 8131 13168 8140 13208
rect 8180 13168 8189 13208
rect 8131 13167 8189 13168
rect 9379 13208 9437 13209
rect 9379 13168 9388 13208
rect 9428 13168 9437 13208
rect 9379 13167 9437 13168
rect 9859 13208 9917 13209
rect 9859 13168 9868 13208
rect 9908 13168 9917 13208
rect 9859 13167 9917 13168
rect 11107 13208 11165 13209
rect 11107 13168 11116 13208
rect 11156 13168 11165 13208
rect 11107 13167 11165 13168
rect 11971 13208 12029 13209
rect 11971 13168 11980 13208
rect 12020 13168 12029 13208
rect 11971 13167 12029 13168
rect 13795 13208 13853 13209
rect 13795 13168 13804 13208
rect 13844 13168 13853 13208
rect 13795 13167 13853 13168
rect 15043 13208 15101 13209
rect 15043 13168 15052 13208
rect 15092 13168 15101 13208
rect 15043 13167 15101 13168
rect 15235 13208 15293 13209
rect 15235 13168 15244 13208
rect 15284 13168 15293 13208
rect 15235 13167 15293 13168
rect 16483 13208 16541 13209
rect 16483 13168 16492 13208
rect 16532 13168 16541 13208
rect 16483 13167 16541 13168
rect 17155 13208 17213 13209
rect 17155 13168 17164 13208
rect 17204 13168 17213 13208
rect 17155 13167 17213 13168
rect 18403 13208 18461 13209
rect 18403 13168 18412 13208
rect 18452 13168 18461 13208
rect 18403 13167 18461 13168
rect 19171 13208 19229 13209
rect 19171 13168 19180 13208
rect 19220 13168 19229 13208
rect 19171 13167 19229 13168
rect 19467 13208 19509 13217
rect 19467 13168 19468 13208
rect 19508 13168 19509 13208
rect 19467 13159 19509 13168
rect 19563 13208 19605 13217
rect 19563 13168 19564 13208
rect 19604 13168 19605 13208
rect 19563 13159 19605 13168
rect 20035 13208 20093 13209
rect 20035 13168 20044 13208
rect 20084 13168 20093 13208
rect 20035 13167 20093 13168
rect 20235 13208 20277 13217
rect 20235 13168 20236 13208
rect 20276 13168 20277 13208
rect 20235 13159 20277 13168
rect 13611 13124 13653 13133
rect 13611 13084 13612 13124
rect 13652 13084 13653 13124
rect 13611 13075 13653 13084
rect 20139 13124 20181 13133
rect 20139 13084 20140 13124
rect 20180 13084 20181 13124
rect 20139 13075 20181 13084
rect 3339 13040 3381 13049
rect 3339 13000 3340 13040
rect 3380 13000 3381 13040
rect 3339 12991 3381 13000
rect 3723 13040 3765 13049
rect 3723 13000 3724 13040
rect 3764 13000 3765 13040
rect 3723 12991 3765 13000
rect 7651 13040 7709 13041
rect 7651 13000 7660 13040
rect 7700 13000 7709 13040
rect 7651 12999 7709 13000
rect 11499 13040 11541 13049
rect 11499 13000 11500 13040
rect 11540 13000 11541 13040
rect 11499 12991 11541 13000
rect 16683 13040 16725 13049
rect 16683 13000 16684 13040
rect 16724 13000 16725 13040
rect 16683 12991 16725 13000
rect 1152 12872 20452 12896
rect 1152 12832 4928 12872
rect 4968 12832 5010 12872
rect 5050 12832 5092 12872
rect 5132 12832 5174 12872
rect 5214 12832 5256 12872
rect 5296 12832 20048 12872
rect 20088 12832 20130 12872
rect 20170 12832 20212 12872
rect 20252 12832 20294 12872
rect 20334 12832 20376 12872
rect 20416 12832 20452 12872
rect 1152 12808 20452 12832
rect 18891 12762 18933 12771
rect 18891 12722 18892 12762
rect 18932 12722 18933 12762
rect 18891 12713 18933 12722
rect 2667 12704 2709 12713
rect 2667 12664 2668 12704
rect 2708 12664 2709 12704
rect 2667 12655 2709 12664
rect 19555 12704 19613 12705
rect 19555 12664 19564 12704
rect 19604 12664 19613 12704
rect 19555 12663 19613 12664
rect 2859 12620 2901 12629
rect 2859 12580 2860 12620
rect 2900 12580 2901 12620
rect 2859 12571 2901 12580
rect 5451 12620 5493 12629
rect 5451 12580 5452 12620
rect 5492 12580 5493 12620
rect 5451 12571 5493 12580
rect 9771 12620 9813 12629
rect 9771 12580 9772 12620
rect 9812 12580 9813 12620
rect 9771 12571 9813 12580
rect 12555 12620 12597 12629
rect 12555 12580 12556 12620
rect 12596 12580 12597 12620
rect 12555 12571 12597 12580
rect 15243 12620 15285 12629
rect 15243 12580 15244 12620
rect 15284 12580 15285 12620
rect 15243 12571 15285 12580
rect 17259 12620 17301 12629
rect 17259 12580 17260 12620
rect 17300 12580 17301 12620
rect 17259 12571 17301 12580
rect 5067 12547 5109 12556
rect 1219 12536 1277 12537
rect 1219 12496 1228 12536
rect 1268 12496 1277 12536
rect 1219 12495 1277 12496
rect 2467 12536 2525 12537
rect 2467 12496 2476 12536
rect 2516 12496 2525 12536
rect 3523 12536 3581 12537
rect 2467 12495 2525 12496
rect 3051 12522 3093 12531
rect 3051 12482 3052 12522
rect 3092 12482 3093 12522
rect 3523 12496 3532 12536
rect 3572 12496 3581 12536
rect 3523 12495 3581 12496
rect 4011 12536 4053 12545
rect 4011 12496 4012 12536
rect 4052 12496 4053 12536
rect 4011 12487 4053 12496
rect 4107 12536 4149 12545
rect 4107 12496 4108 12536
rect 4148 12496 4149 12536
rect 4107 12487 4149 12496
rect 4491 12536 4533 12545
rect 4491 12496 4492 12536
rect 4532 12496 4533 12536
rect 4491 12487 4533 12496
rect 4587 12536 4629 12545
rect 4587 12496 4588 12536
rect 4628 12496 4629 12536
rect 4587 12487 4629 12496
rect 4875 12536 4917 12545
rect 4875 12496 4876 12536
rect 4916 12496 4917 12536
rect 5067 12507 5068 12547
rect 5108 12507 5109 12547
rect 5067 12498 5109 12507
rect 5251 12536 5309 12537
rect 4875 12487 4917 12496
rect 5251 12496 5260 12536
rect 5300 12496 5309 12536
rect 5251 12495 5309 12496
rect 5355 12536 5397 12545
rect 5355 12496 5356 12536
rect 5396 12496 5397 12536
rect 5355 12487 5397 12496
rect 5547 12536 5589 12545
rect 5547 12496 5548 12536
rect 5588 12496 5589 12536
rect 5547 12487 5589 12496
rect 6211 12536 6269 12537
rect 6211 12496 6220 12536
rect 6260 12496 6269 12536
rect 6211 12495 6269 12496
rect 7459 12536 7517 12537
rect 7459 12496 7468 12536
rect 7508 12496 7517 12536
rect 7459 12495 7517 12496
rect 8035 12536 8093 12537
rect 8035 12496 8044 12536
rect 8084 12496 8093 12536
rect 8035 12495 8093 12496
rect 9283 12536 9341 12537
rect 9283 12496 9292 12536
rect 9332 12496 9341 12536
rect 9283 12495 9341 12496
rect 9867 12536 9909 12545
rect 9867 12496 9868 12536
rect 9908 12496 9909 12536
rect 10443 12536 10485 12545
rect 9867 12487 9909 12496
rect 10147 12527 10205 12528
rect 10147 12487 10156 12527
rect 10196 12487 10205 12527
rect 10443 12496 10444 12536
rect 10484 12496 10485 12536
rect 10443 12487 10485 12496
rect 10635 12536 10677 12545
rect 10635 12496 10636 12536
rect 10676 12496 10677 12536
rect 10635 12487 10677 12496
rect 10723 12536 10781 12537
rect 10723 12496 10732 12536
rect 10772 12496 10781 12536
rect 10723 12495 10781 12496
rect 11107 12536 11165 12537
rect 11107 12496 11116 12536
rect 11156 12496 11165 12536
rect 11107 12495 11165 12496
rect 12355 12536 12413 12537
rect 12355 12496 12364 12536
rect 12404 12496 12413 12536
rect 12355 12495 12413 12496
rect 12739 12536 12797 12537
rect 12739 12496 12748 12536
rect 12788 12496 12797 12536
rect 12739 12495 12797 12496
rect 13987 12536 14045 12537
rect 13987 12496 13996 12536
rect 14036 12496 14045 12536
rect 13987 12495 14045 12496
rect 14859 12536 14901 12545
rect 14859 12496 14860 12536
rect 14900 12496 14901 12536
rect 14859 12487 14901 12496
rect 15051 12536 15093 12545
rect 15051 12496 15052 12536
rect 15092 12496 15093 12536
rect 15051 12487 15093 12496
rect 15435 12531 15477 12540
rect 15435 12491 15436 12531
rect 15476 12491 15477 12531
rect 15907 12536 15965 12537
rect 15907 12496 15916 12536
rect 15956 12496 15965 12536
rect 15907 12495 15965 12496
rect 16875 12536 16917 12545
rect 16875 12496 16876 12536
rect 16916 12496 16917 12536
rect 10147 12486 10205 12487
rect 15435 12482 15477 12491
rect 16875 12487 16917 12496
rect 16971 12536 17013 12545
rect 16971 12496 16972 12536
rect 17012 12496 17013 12536
rect 16971 12487 17013 12496
rect 17443 12536 17501 12537
rect 17443 12496 17452 12536
rect 17492 12496 17501 12536
rect 17443 12495 17501 12496
rect 18691 12536 18749 12537
rect 18691 12496 18700 12536
rect 18740 12496 18749 12536
rect 18691 12495 18749 12496
rect 18979 12536 19037 12537
rect 18979 12496 18988 12536
rect 19028 12496 19037 12536
rect 18979 12495 19037 12496
rect 19083 12536 19125 12545
rect 19083 12496 19084 12536
rect 19124 12496 19125 12536
rect 19083 12487 19125 12496
rect 19755 12536 19797 12545
rect 19755 12496 19756 12536
rect 19796 12496 19797 12536
rect 19755 12487 19797 12496
rect 19851 12536 19893 12545
rect 19851 12496 19852 12536
rect 19892 12496 19893 12536
rect 19851 12487 19893 12496
rect 3051 12473 3093 12482
rect 5923 12452 5981 12453
rect 5923 12412 5932 12452
rect 5972 12412 5981 12452
rect 5923 12411 5981 12412
rect 14659 12452 14717 12453
rect 14659 12412 14668 12452
rect 14708 12412 14717 12452
rect 14659 12411 14717 12412
rect 16395 12452 16437 12461
rect 16395 12412 16396 12452
rect 16436 12412 16437 12452
rect 16395 12403 16437 12412
rect 16491 12452 16533 12461
rect 16491 12412 16492 12452
rect 16532 12412 16533 12452
rect 16491 12403 16533 12412
rect 20227 12452 20285 12453
rect 20227 12412 20236 12452
rect 20276 12412 20285 12452
rect 20227 12411 20285 12412
rect 7851 12368 7893 12377
rect 7851 12328 7852 12368
rect 7892 12328 7893 12368
rect 7851 12319 7893 12328
rect 9475 12368 9533 12369
rect 9475 12328 9484 12368
rect 9524 12328 9533 12368
rect 9475 12327 9533 12328
rect 19371 12368 19413 12377
rect 19371 12328 19372 12368
rect 19412 12328 19413 12368
rect 19371 12319 19413 12328
rect 5067 12284 5109 12293
rect 5067 12244 5068 12284
rect 5108 12244 5109 12284
rect 5067 12235 5109 12244
rect 5739 12284 5781 12293
rect 5739 12244 5740 12284
rect 5780 12244 5781 12284
rect 5739 12235 5781 12244
rect 7659 12284 7701 12293
rect 7659 12244 7660 12284
rect 7700 12244 7701 12284
rect 7659 12235 7701 12244
rect 10443 12284 10485 12293
rect 10443 12244 10444 12284
rect 10484 12244 10485 12284
rect 10443 12235 10485 12244
rect 14187 12284 14229 12293
rect 14187 12244 14188 12284
rect 14228 12244 14229 12284
rect 14187 12235 14229 12244
rect 14475 12284 14517 12293
rect 14475 12244 14476 12284
rect 14516 12244 14517 12284
rect 14475 12235 14517 12244
rect 14859 12284 14901 12293
rect 14859 12244 14860 12284
rect 14900 12244 14901 12284
rect 14859 12235 14901 12244
rect 20043 12284 20085 12293
rect 20043 12244 20044 12284
rect 20084 12244 20085 12284
rect 20043 12235 20085 12244
rect 1152 12116 20352 12140
rect 1152 12076 3688 12116
rect 3728 12076 3770 12116
rect 3810 12076 3852 12116
rect 3892 12076 3934 12116
rect 3974 12076 4016 12116
rect 4056 12076 18808 12116
rect 18848 12076 18890 12116
rect 18930 12076 18972 12116
rect 19012 12076 19054 12116
rect 19094 12076 19136 12116
rect 19176 12076 20352 12116
rect 1152 12052 20352 12076
rect 2667 11948 2709 11957
rect 2667 11908 2668 11948
rect 2708 11908 2709 11948
rect 2667 11899 2709 11908
rect 7467 11948 7509 11957
rect 7467 11908 7468 11948
rect 7508 11908 7509 11948
rect 7467 11899 7509 11908
rect 7659 11948 7701 11957
rect 7659 11908 7660 11948
rect 7700 11908 7701 11948
rect 7659 11899 7701 11908
rect 4587 11864 4629 11873
rect 4587 11824 4588 11864
rect 4628 11824 4629 11864
rect 4587 11815 4629 11824
rect 10243 11864 10301 11865
rect 10243 11824 10252 11864
rect 10292 11824 10301 11864
rect 10243 11823 10301 11824
rect 19075 11864 19133 11865
rect 19075 11824 19084 11864
rect 19124 11824 19133 11864
rect 19075 11823 19133 11824
rect 5835 11780 5877 11789
rect 5835 11740 5836 11780
rect 5876 11740 5877 11780
rect 5835 11731 5877 11740
rect 5931 11780 5973 11789
rect 5931 11740 5932 11780
rect 5972 11740 5973 11780
rect 5931 11731 5973 11740
rect 12651 11780 12693 11789
rect 12651 11740 12652 11780
rect 12692 11740 12693 11780
rect 12651 11731 12693 11740
rect 12747 11780 12789 11789
rect 12747 11740 12748 11780
rect 12788 11740 12789 11780
rect 12747 11731 12789 11740
rect 14275 11780 14333 11781
rect 14275 11740 14284 11780
rect 14324 11740 14333 11780
rect 14275 11739 14333 11740
rect 14755 11780 14813 11781
rect 14755 11740 14764 11780
rect 14804 11740 14813 11780
rect 14755 11739 14813 11740
rect 15627 11780 15669 11789
rect 15627 11740 15628 11780
rect 15668 11740 15669 11780
rect 17155 11780 17213 11781
rect 15627 11731 15669 11740
rect 16635 11738 16677 11747
rect 17155 11740 17164 11780
rect 17204 11740 17213 11780
rect 17155 11739 17213 11740
rect 20227 11780 20285 11781
rect 20227 11740 20236 11780
rect 20276 11740 20285 11780
rect 20227 11739 20285 11740
rect 13707 11710 13749 11719
rect 1219 11696 1277 11697
rect 1219 11656 1228 11696
rect 1268 11656 1277 11696
rect 1219 11655 1277 11656
rect 2467 11696 2525 11697
rect 2467 11656 2476 11696
rect 2516 11656 2525 11696
rect 2467 11655 2525 11656
rect 2859 11696 2901 11705
rect 2859 11656 2860 11696
rect 2900 11656 2901 11696
rect 2859 11647 2901 11656
rect 2947 11696 3005 11697
rect 2947 11656 2956 11696
rect 2996 11656 3005 11696
rect 2947 11655 3005 11656
rect 3139 11696 3197 11697
rect 3139 11656 3148 11696
rect 3188 11656 3197 11696
rect 3139 11655 3197 11656
rect 4387 11696 4445 11697
rect 4387 11656 4396 11696
rect 4436 11656 4445 11696
rect 4387 11655 4445 11656
rect 4779 11696 4821 11705
rect 4779 11656 4780 11696
rect 4820 11656 4821 11696
rect 4779 11647 4821 11656
rect 4971 11696 5013 11705
rect 4971 11656 4972 11696
rect 5012 11656 5013 11696
rect 4971 11647 5013 11656
rect 5059 11696 5117 11697
rect 5059 11656 5068 11696
rect 5108 11656 5117 11696
rect 5059 11655 5117 11656
rect 5355 11696 5397 11705
rect 5355 11656 5356 11696
rect 5396 11656 5397 11696
rect 5355 11647 5397 11656
rect 5451 11696 5493 11705
rect 6891 11701 6933 11710
rect 5451 11656 5452 11696
rect 5492 11656 5493 11696
rect 5451 11647 5493 11656
rect 6403 11696 6461 11697
rect 6403 11656 6412 11696
rect 6452 11656 6461 11696
rect 6403 11655 6461 11656
rect 6891 11661 6892 11701
rect 6932 11661 6933 11701
rect 6891 11652 6933 11661
rect 7275 11696 7317 11705
rect 7275 11656 7276 11696
rect 7316 11656 7317 11696
rect 7275 11647 7317 11656
rect 7467 11696 7509 11705
rect 7467 11656 7468 11696
rect 7508 11656 7509 11696
rect 7467 11647 7509 11656
rect 7843 11696 7901 11697
rect 7843 11656 7852 11696
rect 7892 11656 7901 11696
rect 7843 11655 7901 11656
rect 9091 11696 9149 11697
rect 9091 11656 9100 11696
rect 9140 11656 9149 11696
rect 9091 11655 9149 11656
rect 9571 11696 9629 11697
rect 9571 11656 9580 11696
rect 9620 11656 9629 11696
rect 9571 11655 9629 11656
rect 9867 11696 9909 11705
rect 9867 11656 9868 11696
rect 9908 11656 9909 11696
rect 9867 11647 9909 11656
rect 10435 11696 10493 11697
rect 10435 11656 10444 11696
rect 10484 11656 10493 11696
rect 10435 11655 10493 11656
rect 11683 11696 11741 11697
rect 11683 11656 11692 11696
rect 11732 11656 11741 11696
rect 11683 11655 11741 11656
rect 12171 11696 12213 11705
rect 12171 11656 12172 11696
rect 12212 11656 12213 11696
rect 12171 11647 12213 11656
rect 12267 11696 12309 11705
rect 12267 11656 12268 11696
rect 12308 11656 12309 11696
rect 12267 11647 12309 11656
rect 13219 11696 13277 11697
rect 13219 11656 13228 11696
rect 13268 11656 13277 11696
rect 13707 11670 13708 11710
rect 13748 11670 13749 11710
rect 13707 11661 13749 11670
rect 15051 11696 15093 11705
rect 13219 11655 13277 11656
rect 15051 11656 15052 11696
rect 15092 11656 15093 11696
rect 15051 11647 15093 11656
rect 15147 11696 15189 11705
rect 15147 11656 15148 11696
rect 15188 11656 15189 11696
rect 15147 11647 15189 11656
rect 15531 11696 15573 11705
rect 16635 11698 16636 11738
rect 16676 11698 16677 11738
rect 15531 11656 15532 11696
rect 15572 11656 15573 11696
rect 15531 11647 15573 11656
rect 16099 11696 16157 11697
rect 16099 11656 16108 11696
rect 16148 11656 16157 11696
rect 16635 11689 16677 11698
rect 17347 11696 17405 11697
rect 16099 11655 16157 11656
rect 17347 11656 17356 11696
rect 17396 11656 17405 11696
rect 17347 11655 17405 11656
rect 18595 11696 18653 11697
rect 18595 11656 18604 11696
rect 18644 11656 18653 11696
rect 18595 11655 18653 11656
rect 19467 11696 19509 11705
rect 19467 11656 19468 11696
rect 19508 11656 19509 11696
rect 19467 11647 19509 11656
rect 19747 11696 19805 11697
rect 19747 11656 19756 11696
rect 19796 11656 19805 11696
rect 19747 11655 19805 11656
rect 9963 11612 10005 11621
rect 9963 11572 9964 11612
rect 10004 11572 10005 11612
rect 9963 11563 10005 11572
rect 11883 11612 11925 11621
rect 11883 11572 11884 11612
rect 11924 11572 11925 11612
rect 11883 11563 11925 11572
rect 18795 11612 18837 11621
rect 18795 11572 18796 11612
rect 18836 11572 18837 11612
rect 18795 11563 18837 11572
rect 19371 11612 19413 11621
rect 19371 11572 19372 11612
rect 19412 11572 19413 11612
rect 19371 11563 19413 11572
rect 4867 11528 4925 11529
rect 4867 11488 4876 11528
rect 4916 11488 4925 11528
rect 4867 11487 4925 11488
rect 7083 11528 7125 11537
rect 7083 11488 7084 11528
rect 7124 11488 7125 11528
rect 7083 11479 7125 11488
rect 7659 11528 7701 11537
rect 7659 11488 7660 11528
rect 7700 11488 7701 11528
rect 7659 11479 7701 11488
rect 13899 11528 13941 11537
rect 13899 11488 13900 11528
rect 13940 11488 13941 11528
rect 13899 11479 13941 11488
rect 14091 11528 14133 11537
rect 14091 11488 14092 11528
rect 14132 11488 14133 11528
rect 14091 11479 14133 11488
rect 14571 11528 14613 11537
rect 14571 11488 14572 11528
rect 14612 11488 14613 11528
rect 14571 11479 14613 11488
rect 16779 11528 16821 11537
rect 16779 11488 16780 11528
rect 16820 11488 16821 11528
rect 16779 11479 16821 11488
rect 16971 11528 17013 11537
rect 16971 11488 16972 11528
rect 17012 11488 17013 11528
rect 16971 11479 17013 11488
rect 20043 11528 20085 11537
rect 20043 11488 20044 11528
rect 20084 11488 20085 11528
rect 20043 11479 20085 11488
rect 1152 11360 20452 11384
rect 1152 11320 4928 11360
rect 4968 11320 5010 11360
rect 5050 11320 5092 11360
rect 5132 11320 5174 11360
rect 5214 11320 5256 11360
rect 5296 11320 20048 11360
rect 20088 11320 20130 11360
rect 20170 11320 20212 11360
rect 20252 11320 20294 11360
rect 20334 11320 20376 11360
rect 20416 11320 20452 11360
rect 1152 11296 20452 11320
rect 1515 11192 1557 11201
rect 1515 11152 1516 11192
rect 1556 11152 1557 11192
rect 1515 11143 1557 11152
rect 5259 11192 5301 11201
rect 5259 11152 5260 11192
rect 5300 11152 5301 11192
rect 5259 11143 5301 11152
rect 5739 11192 5781 11201
rect 5739 11152 5740 11192
rect 5780 11152 5781 11192
rect 5739 11143 5781 11152
rect 16779 11192 16821 11201
rect 16779 11152 16780 11192
rect 16820 11152 16821 11192
rect 16779 11143 16821 11152
rect 18411 11192 18453 11201
rect 18411 11152 18412 11192
rect 18452 11152 18453 11192
rect 18411 11143 18453 11152
rect 9483 11108 9525 11117
rect 9483 11068 9484 11108
rect 9524 11068 9525 11108
rect 9483 11059 9525 11068
rect 13131 11108 13173 11117
rect 13131 11068 13132 11108
rect 13172 11068 13173 11108
rect 13131 11059 13173 11068
rect 13323 11108 13365 11117
rect 13323 11068 13324 11108
rect 13364 11068 13365 11108
rect 13323 11059 13365 11068
rect 1323 11024 1365 11033
rect 1323 10984 1324 11024
rect 1364 10984 1365 11024
rect 1323 10975 1365 10984
rect 1611 11024 1653 11033
rect 1611 10984 1612 11024
rect 1652 10984 1653 11024
rect 1611 10975 1653 10984
rect 2179 11024 2237 11025
rect 2179 10984 2188 11024
rect 2228 10984 2237 11024
rect 2179 10983 2237 10984
rect 3427 11024 3485 11025
rect 3427 10984 3436 11024
rect 3476 10984 3485 11024
rect 3427 10983 3485 10984
rect 3811 11024 3869 11025
rect 3811 10984 3820 11024
rect 3860 10984 3869 11024
rect 3811 10983 3869 10984
rect 5059 11024 5117 11025
rect 5059 10984 5068 11024
rect 5108 10984 5117 11024
rect 5059 10983 5117 10984
rect 5539 11024 5597 11025
rect 5539 10984 5548 11024
rect 5588 10984 5597 11024
rect 5539 10983 5597 10984
rect 5923 11024 5981 11025
rect 5923 10984 5932 11024
rect 5972 10984 5981 11024
rect 5923 10983 5981 10984
rect 7171 11024 7229 11025
rect 7171 10984 7180 11024
rect 7220 10984 7229 11024
rect 7171 10983 7229 10984
rect 7363 11024 7421 11025
rect 7363 10984 7372 11024
rect 7412 10984 7421 11024
rect 7363 10983 7421 10984
rect 8611 11024 8669 11025
rect 8611 10984 8620 11024
rect 8660 10984 8669 11024
rect 8611 10983 8669 10984
rect 9091 11024 9149 11025
rect 9091 10984 9100 11024
rect 9140 10984 9149 11024
rect 9091 10983 9149 10984
rect 9387 11024 9429 11033
rect 9387 10984 9388 11024
rect 9428 10984 9429 11024
rect 9387 10975 9429 10984
rect 10243 11024 10301 11025
rect 10243 10984 10252 11024
rect 10292 10984 10301 11024
rect 10243 10983 10301 10984
rect 11491 11024 11549 11025
rect 11491 10984 11500 11024
rect 11540 10984 11549 11024
rect 11491 10983 11549 10984
rect 11683 11024 11741 11025
rect 11683 10984 11692 11024
rect 11732 10984 11741 11024
rect 11683 10983 11741 10984
rect 12931 11024 12989 11025
rect 12931 10984 12940 11024
rect 12980 10984 12989 11024
rect 13987 11024 14045 11025
rect 12931 10983 12989 10984
rect 13515 11010 13557 11019
rect 13515 10970 13516 11010
rect 13556 10970 13557 11010
rect 13987 10984 13996 11024
rect 14036 10984 14045 11024
rect 13987 10983 14045 10984
rect 14475 11024 14517 11033
rect 14475 10984 14476 11024
rect 14516 10984 14517 11024
rect 14475 10975 14517 10984
rect 14571 11024 14613 11033
rect 14571 10984 14572 11024
rect 14612 10984 14613 11024
rect 14571 10975 14613 10984
rect 14955 11024 14997 11033
rect 14955 10984 14956 11024
rect 14996 10984 14997 11024
rect 14955 10975 14997 10984
rect 15051 11024 15093 11033
rect 15051 10984 15052 11024
rect 15092 10984 15093 11024
rect 15051 10975 15093 10984
rect 15331 11024 15389 11025
rect 15331 10984 15340 11024
rect 15380 10984 15389 11024
rect 15331 10983 15389 10984
rect 16579 11024 16637 11025
rect 16579 10984 16588 11024
rect 16628 10984 16637 11024
rect 16579 10983 16637 10984
rect 18211 11024 18269 11025
rect 18211 10984 18220 11024
rect 18260 10984 18269 11024
rect 18211 10983 18269 10984
rect 18691 11024 18749 11025
rect 18691 10984 18700 11024
rect 18740 10984 18749 11024
rect 18691 10983 18749 10984
rect 18987 11024 19029 11033
rect 18987 10984 18988 11024
rect 19028 10984 19029 11024
rect 16963 10982 17021 10983
rect 13515 10961 13557 10970
rect 16963 10942 16972 10982
rect 17012 10942 17021 10982
rect 18987 10975 19029 10984
rect 19083 11024 19125 11033
rect 19083 10984 19084 11024
rect 19124 10984 19125 11024
rect 19083 10975 19125 10984
rect 19563 11024 19605 11033
rect 19563 10984 19564 11024
rect 19604 10984 19605 11024
rect 19563 10975 19605 10984
rect 19939 11024 19997 11025
rect 19939 10984 19948 11024
rect 19988 10984 19997 11024
rect 19939 10983 19997 10984
rect 20227 11024 20285 11025
rect 20227 10984 20236 11024
rect 20276 10984 20285 11024
rect 20227 10983 20285 10984
rect 16963 10941 17021 10942
rect 1987 10940 2045 10941
rect 1987 10900 1996 10940
rect 2036 10900 2045 10940
rect 1987 10899 2045 10900
rect 19659 10940 19701 10949
rect 19659 10900 19660 10940
rect 19700 10900 19701 10940
rect 19659 10891 19701 10900
rect 19851 10940 19893 10949
rect 19851 10900 19852 10940
rect 19892 10900 19893 10940
rect 19851 10891 19893 10900
rect 5451 10856 5493 10865
rect 5451 10816 5452 10856
rect 5492 10816 5493 10856
rect 5451 10807 5493 10816
rect 9763 10856 9821 10857
rect 9763 10816 9772 10856
rect 9812 10816 9821 10856
rect 9763 10815 9821 10816
rect 19755 10856 19797 10865
rect 19755 10816 19756 10856
rect 19796 10816 19797 10856
rect 19755 10807 19797 10816
rect 1803 10772 1845 10781
rect 1803 10732 1804 10772
rect 1844 10732 1845 10772
rect 1803 10723 1845 10732
rect 3627 10772 3669 10781
rect 3627 10732 3628 10772
rect 3668 10732 3669 10772
rect 3627 10723 3669 10732
rect 8811 10772 8853 10781
rect 8811 10732 8812 10772
rect 8852 10732 8853 10772
rect 8811 10723 8853 10732
rect 10059 10772 10101 10781
rect 10059 10732 10060 10772
rect 10100 10732 10101 10772
rect 10059 10723 10101 10732
rect 19363 10772 19421 10773
rect 19363 10732 19372 10772
rect 19412 10732 19421 10772
rect 19363 10731 19421 10732
rect 20139 10772 20181 10781
rect 20139 10732 20140 10772
rect 20180 10732 20181 10772
rect 20139 10723 20181 10732
rect 1152 10604 20352 10628
rect 1152 10564 3688 10604
rect 3728 10564 3770 10604
rect 3810 10564 3852 10604
rect 3892 10564 3934 10604
rect 3974 10564 4016 10604
rect 4056 10564 18808 10604
rect 18848 10564 18890 10604
rect 18930 10564 18972 10604
rect 19012 10564 19054 10604
rect 19094 10564 19136 10604
rect 19176 10564 20352 10604
rect 1152 10540 20352 10564
rect 2859 10436 2901 10445
rect 2859 10396 2860 10436
rect 2900 10396 2901 10436
rect 2859 10387 2901 10396
rect 3051 10436 3093 10445
rect 3051 10396 3052 10436
rect 3092 10396 3093 10436
rect 3051 10387 3093 10396
rect 5067 10436 5109 10445
rect 5067 10396 5068 10436
rect 5108 10396 5109 10436
rect 5067 10387 5109 10396
rect 6891 10436 6933 10445
rect 6891 10396 6892 10436
rect 6932 10396 6933 10436
rect 6891 10387 6933 10396
rect 11787 10436 11829 10445
rect 11787 10396 11788 10436
rect 11828 10396 11829 10436
rect 11787 10387 11829 10396
rect 14859 10436 14901 10445
rect 14859 10396 14860 10436
rect 14900 10396 14901 10436
rect 14859 10387 14901 10396
rect 18891 10436 18933 10445
rect 18891 10396 18892 10436
rect 18932 10396 18933 10436
rect 18891 10387 18933 10396
rect 4683 10352 4725 10361
rect 4683 10312 4684 10352
rect 4724 10312 4725 10352
rect 4683 10303 4725 10312
rect 9963 10352 10005 10361
rect 9963 10312 9964 10352
rect 10004 10312 10005 10352
rect 9963 10303 10005 10312
rect 12739 10352 12797 10353
rect 12739 10312 12748 10352
rect 12788 10312 12797 10352
rect 12739 10311 12797 10312
rect 19075 10352 19133 10353
rect 19075 10312 19084 10352
rect 19124 10312 19133 10352
rect 19075 10311 19133 10312
rect 20043 10352 20085 10361
rect 20043 10312 20044 10352
rect 20084 10312 20085 10352
rect 20043 10303 20085 10312
rect 5251 10268 5309 10269
rect 5251 10228 5260 10268
rect 5300 10228 5309 10268
rect 5251 10227 5309 10228
rect 9867 10268 9909 10277
rect 9867 10228 9868 10268
rect 9908 10228 9909 10268
rect 9867 10219 9909 10228
rect 10059 10268 10101 10277
rect 10059 10228 10060 10268
rect 10100 10228 10101 10268
rect 10059 10219 10101 10228
rect 20227 10268 20285 10269
rect 20227 10228 20236 10268
rect 20276 10228 20285 10268
rect 20227 10227 20285 10228
rect 1411 10184 1469 10185
rect 1411 10144 1420 10184
rect 1460 10144 1469 10184
rect 1411 10143 1469 10144
rect 2659 10184 2717 10185
rect 2659 10144 2668 10184
rect 2708 10144 2717 10184
rect 2659 10143 2717 10144
rect 3235 10184 3293 10185
rect 3235 10144 3244 10184
rect 3284 10144 3293 10184
rect 3235 10143 3293 10144
rect 4483 10184 4541 10185
rect 4483 10144 4492 10184
rect 4532 10144 4541 10184
rect 4483 10143 4541 10144
rect 4683 10184 4725 10193
rect 4683 10144 4684 10184
rect 4724 10144 4725 10184
rect 4683 10135 4725 10144
rect 4875 10184 4917 10193
rect 4875 10144 4876 10184
rect 4916 10144 4917 10184
rect 4875 10135 4917 10144
rect 5443 10184 5501 10185
rect 5443 10144 5452 10184
rect 5492 10144 5501 10184
rect 5443 10143 5501 10144
rect 6691 10184 6749 10185
rect 6691 10144 6700 10184
rect 6740 10144 6749 10184
rect 6691 10143 6749 10144
rect 7179 10184 7221 10193
rect 7179 10144 7180 10184
rect 7220 10144 7221 10184
rect 7179 10135 7221 10144
rect 7275 10184 7317 10193
rect 7275 10144 7276 10184
rect 7316 10144 7317 10184
rect 7275 10135 7317 10144
rect 7371 10184 7413 10193
rect 7371 10144 7372 10184
rect 7412 10144 7413 10184
rect 7371 10135 7413 10144
rect 7467 10184 7509 10193
rect 7467 10144 7468 10184
rect 7508 10144 7509 10184
rect 7467 10135 7509 10144
rect 7659 10184 7701 10193
rect 7659 10144 7660 10184
rect 7700 10144 7701 10184
rect 7659 10135 7701 10144
rect 7755 10184 7797 10193
rect 7755 10144 7756 10184
rect 7796 10144 7797 10184
rect 7755 10135 7797 10144
rect 8131 10184 8189 10185
rect 8131 10144 8140 10184
rect 8180 10144 8189 10184
rect 8131 10143 8189 10144
rect 9379 10184 9437 10185
rect 9379 10144 9388 10184
rect 9428 10144 9437 10184
rect 9379 10143 9437 10144
rect 9763 10184 9821 10185
rect 9763 10144 9772 10184
rect 9812 10144 9821 10184
rect 9763 10143 9821 10144
rect 10155 10184 10197 10193
rect 10155 10144 10156 10184
rect 10196 10144 10197 10184
rect 10155 10135 10197 10144
rect 10339 10184 10397 10185
rect 10339 10144 10348 10184
rect 10388 10144 10397 10184
rect 10339 10143 10397 10144
rect 11587 10184 11645 10185
rect 11587 10144 11596 10184
rect 11636 10144 11645 10184
rect 11587 10143 11645 10144
rect 12067 10184 12125 10185
rect 12067 10144 12076 10184
rect 12116 10144 12125 10184
rect 12067 10143 12125 10144
rect 12363 10184 12405 10193
rect 12363 10144 12364 10184
rect 12404 10144 12405 10184
rect 12363 10135 12405 10144
rect 12459 10184 12501 10193
rect 12459 10144 12460 10184
rect 12500 10144 12501 10184
rect 12459 10135 12501 10144
rect 12939 10184 12981 10193
rect 12939 10144 12940 10184
rect 12980 10144 12981 10184
rect 12939 10135 12981 10144
rect 13131 10184 13173 10193
rect 13131 10144 13132 10184
rect 13172 10144 13173 10184
rect 13131 10135 13173 10144
rect 13219 10184 13277 10185
rect 13219 10144 13228 10184
rect 13268 10144 13277 10184
rect 13219 10143 13277 10144
rect 13411 10184 13469 10185
rect 13411 10144 13420 10184
rect 13460 10144 13469 10184
rect 13411 10143 13469 10144
rect 14659 10184 14717 10185
rect 14659 10144 14668 10184
rect 14708 10144 14717 10184
rect 14659 10143 14717 10144
rect 15051 10184 15093 10193
rect 15051 10144 15052 10184
rect 15092 10144 15093 10184
rect 15051 10135 15093 10144
rect 15139 10184 15197 10185
rect 15139 10144 15148 10184
rect 15188 10144 15197 10184
rect 15139 10143 15197 10144
rect 15331 10184 15389 10185
rect 15331 10144 15340 10184
rect 15380 10144 15389 10184
rect 15331 10143 15389 10144
rect 16579 10184 16637 10185
rect 16579 10144 16588 10184
rect 16628 10144 16637 10184
rect 16579 10143 16637 10144
rect 16963 10184 17021 10185
rect 16963 10144 16972 10184
rect 17012 10144 17021 10184
rect 16963 10143 17021 10144
rect 17067 10184 17109 10193
rect 17067 10144 17068 10184
rect 17108 10144 17109 10184
rect 17067 10135 17109 10144
rect 17259 10184 17301 10193
rect 17259 10144 17260 10184
rect 17300 10144 17301 10184
rect 17259 10135 17301 10144
rect 17443 10184 17501 10185
rect 17443 10144 17452 10184
rect 17492 10144 17501 10184
rect 17443 10143 17501 10144
rect 18691 10184 18749 10185
rect 18691 10144 18700 10184
rect 18740 10144 18749 10184
rect 18691 10143 18749 10144
rect 19371 10184 19413 10193
rect 19371 10144 19372 10184
rect 19412 10144 19413 10184
rect 19371 10135 19413 10144
rect 19467 10184 19509 10193
rect 19467 10144 19468 10184
rect 19508 10144 19509 10184
rect 19467 10135 19509 10144
rect 19747 10184 19805 10185
rect 19747 10144 19756 10184
rect 19796 10144 19805 10184
rect 19747 10143 19805 10144
rect 7939 10016 7997 10017
rect 7939 9976 7948 10016
rect 7988 9976 7997 10016
rect 7939 9975 7997 9976
rect 9579 10016 9621 10025
rect 9579 9976 9580 10016
rect 9620 9976 9621 10016
rect 9579 9967 9621 9976
rect 13027 10016 13085 10017
rect 13027 9976 13036 10016
rect 13076 9976 13085 10016
rect 13027 9975 13085 9976
rect 16779 10016 16821 10025
rect 16779 9976 16780 10016
rect 16820 9976 16821 10016
rect 16779 9967 16821 9976
rect 17155 10016 17213 10017
rect 17155 9976 17164 10016
rect 17204 9976 17213 10016
rect 17155 9975 17213 9976
rect 1152 9848 20452 9872
rect 1152 9808 4928 9848
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 5296 9808 20048 9848
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20416 9808 20452 9848
rect 1152 9784 20452 9808
rect 3051 9680 3093 9689
rect 3051 9640 3052 9680
rect 3092 9640 3093 9680
rect 3051 9631 3093 9640
rect 13323 9680 13365 9689
rect 13323 9640 13324 9680
rect 13364 9640 13365 9680
rect 13323 9631 13365 9640
rect 16779 9680 16821 9689
rect 16779 9640 16780 9680
rect 16820 9640 16821 9680
rect 16779 9631 16821 9640
rect 17923 9680 17981 9681
rect 17923 9640 17932 9680
rect 17972 9640 17981 9680
rect 17923 9639 17981 9640
rect 3243 9596 3285 9605
rect 3243 9556 3244 9596
rect 3284 9556 3285 9596
rect 3243 9547 3285 9556
rect 7659 9596 7701 9605
rect 7659 9556 7660 9596
rect 7700 9556 7701 9596
rect 7659 9547 7701 9556
rect 1227 9512 1269 9521
rect 1227 9472 1228 9512
rect 1268 9472 1269 9512
rect 1227 9463 1269 9472
rect 1419 9512 1461 9521
rect 1419 9472 1420 9512
rect 1460 9472 1461 9512
rect 1419 9463 1461 9472
rect 1603 9512 1661 9513
rect 1603 9472 1612 9512
rect 1652 9472 1661 9512
rect 3435 9507 3477 9516
rect 1603 9471 1661 9472
rect 2851 9491 2909 9492
rect 2851 9451 2860 9491
rect 2900 9451 2909 9491
rect 3435 9467 3436 9507
rect 3476 9467 3477 9507
rect 3907 9512 3965 9513
rect 3907 9472 3916 9512
rect 3956 9472 3965 9512
rect 3907 9471 3965 9472
rect 4491 9512 4533 9521
rect 4491 9472 4492 9512
rect 4532 9472 4533 9512
rect 3435 9458 3477 9467
rect 4491 9463 4533 9472
rect 4875 9512 4917 9521
rect 4875 9472 4876 9512
rect 4916 9472 4917 9512
rect 4875 9463 4917 9472
rect 4971 9512 5013 9521
rect 4971 9472 4972 9512
rect 5012 9472 5013 9512
rect 4971 9463 5013 9472
rect 5355 9512 5397 9521
rect 5355 9472 5356 9512
rect 5396 9472 5397 9512
rect 5355 9463 5397 9472
rect 5547 9512 5589 9521
rect 5547 9472 5548 9512
rect 5588 9472 5589 9512
rect 5931 9512 5973 9521
rect 5547 9463 5589 9472
rect 5635 9510 5693 9511
rect 5635 9470 5644 9510
rect 5684 9470 5693 9510
rect 5635 9469 5693 9470
rect 5931 9472 5932 9512
rect 5972 9472 5973 9512
rect 5931 9463 5973 9472
rect 6027 9512 6069 9521
rect 6027 9472 6028 9512
rect 6068 9472 6069 9512
rect 6027 9463 6069 9472
rect 6979 9512 7037 9513
rect 6979 9472 6988 9512
rect 7028 9472 7037 9512
rect 7851 9512 7893 9521
rect 6979 9471 7037 9472
rect 7467 9498 7509 9507
rect 7467 9458 7468 9498
rect 7508 9458 7509 9498
rect 7851 9472 7852 9512
rect 7892 9472 7893 9512
rect 7851 9463 7893 9472
rect 8043 9512 8085 9521
rect 8043 9472 8044 9512
rect 8084 9472 8085 9512
rect 8043 9463 8085 9472
rect 8523 9512 8565 9521
rect 8523 9472 8524 9512
rect 8564 9472 8565 9512
rect 8523 9463 8565 9472
rect 8619 9512 8661 9521
rect 8619 9472 8620 9512
rect 8660 9472 8661 9512
rect 8619 9463 8661 9472
rect 8899 9512 8957 9513
rect 8899 9472 8908 9512
rect 8948 9472 8957 9512
rect 8899 9471 8957 9472
rect 9187 9512 9245 9513
rect 9187 9472 9196 9512
rect 9236 9472 9245 9512
rect 9187 9471 9245 9472
rect 10435 9512 10493 9513
rect 10435 9472 10444 9512
rect 10484 9472 10493 9512
rect 10435 9471 10493 9472
rect 10915 9512 10973 9513
rect 10915 9472 10924 9512
rect 10964 9472 10973 9512
rect 10915 9471 10973 9472
rect 11307 9512 11349 9521
rect 11307 9472 11308 9512
rect 11348 9472 11349 9512
rect 11307 9463 11349 9472
rect 11491 9512 11549 9513
rect 11491 9472 11500 9512
rect 11540 9472 11549 9512
rect 11491 9471 11549 9472
rect 12739 9512 12797 9513
rect 12739 9472 12748 9512
rect 12788 9472 12797 9512
rect 12739 9471 12797 9472
rect 13507 9512 13565 9513
rect 13507 9472 13516 9512
rect 13556 9472 13565 9512
rect 13507 9471 13565 9472
rect 14755 9512 14813 9513
rect 14755 9472 14764 9512
rect 14804 9472 14813 9512
rect 14755 9471 14813 9472
rect 15051 9512 15093 9521
rect 15051 9472 15052 9512
rect 15092 9472 15093 9512
rect 15051 9463 15093 9472
rect 15147 9512 15189 9521
rect 15147 9472 15148 9512
rect 15188 9472 15189 9512
rect 15147 9463 15189 9472
rect 16099 9512 16157 9513
rect 16099 9472 16108 9512
rect 16148 9472 16157 9512
rect 16971 9512 17013 9521
rect 16099 9471 16157 9472
rect 16587 9498 16629 9507
rect 2851 9450 2909 9451
rect 7467 9449 7509 9458
rect 16587 9458 16588 9498
rect 16628 9458 16629 9498
rect 16971 9472 16972 9512
rect 17012 9472 17013 9512
rect 16971 9463 17013 9472
rect 17067 9512 17109 9521
rect 17067 9472 17068 9512
rect 17108 9472 17109 9512
rect 17067 9463 17109 9472
rect 17163 9512 17205 9521
rect 17163 9472 17164 9512
rect 17204 9472 17205 9512
rect 17163 9463 17205 9472
rect 17259 9512 17301 9521
rect 17259 9472 17260 9512
rect 17300 9472 17301 9512
rect 17259 9463 17301 9472
rect 17451 9512 17493 9521
rect 17451 9472 17452 9512
rect 17492 9472 17493 9512
rect 17451 9463 17493 9472
rect 17643 9512 17685 9521
rect 17643 9472 17644 9512
rect 17684 9472 17685 9512
rect 17643 9463 17685 9472
rect 17835 9512 17877 9521
rect 17835 9472 17836 9512
rect 17876 9472 17877 9512
rect 17835 9463 17877 9472
rect 18027 9512 18069 9521
rect 18027 9472 18028 9512
rect 18068 9472 18069 9512
rect 18027 9463 18069 9472
rect 18115 9512 18173 9513
rect 18115 9472 18124 9512
rect 18164 9472 18173 9512
rect 18115 9471 18173 9472
rect 18307 9512 18365 9513
rect 18307 9472 18316 9512
rect 18356 9472 18365 9512
rect 18307 9471 18365 9472
rect 19555 9512 19613 9513
rect 19555 9472 19564 9512
rect 19604 9472 19613 9512
rect 19555 9471 19613 9472
rect 19939 9512 19997 9513
rect 19939 9472 19948 9512
rect 19988 9472 19997 9512
rect 19939 9471 19997 9472
rect 20043 9512 20085 9521
rect 20043 9472 20044 9512
rect 20084 9472 20085 9512
rect 20043 9463 20085 9472
rect 20235 9512 20277 9521
rect 20235 9472 20236 9512
rect 20276 9472 20277 9512
rect 20235 9463 20277 9472
rect 16587 9449 16629 9458
rect 4395 9428 4437 9437
rect 4395 9388 4396 9428
rect 4436 9388 4437 9428
rect 4395 9379 4437 9388
rect 6411 9428 6453 9437
rect 6411 9388 6412 9428
rect 6452 9388 6453 9428
rect 6411 9379 6453 9388
rect 6507 9428 6549 9437
rect 6507 9388 6508 9428
rect 6548 9388 6549 9428
rect 6507 9379 6549 9388
rect 11019 9428 11061 9437
rect 11019 9388 11020 9428
rect 11060 9388 11061 9428
rect 15531 9428 15573 9437
rect 11019 9379 11061 9388
rect 11211 9386 11253 9395
rect 8227 9344 8285 9345
rect 8227 9304 8236 9344
rect 8276 9304 8285 9344
rect 8227 9303 8285 9304
rect 11115 9344 11157 9353
rect 11115 9304 11116 9344
rect 11156 9304 11157 9344
rect 11211 9346 11212 9386
rect 11252 9346 11253 9386
rect 15531 9388 15532 9428
rect 15572 9388 15573 9428
rect 15531 9379 15573 9388
rect 15627 9428 15669 9437
rect 15627 9388 15628 9428
rect 15668 9388 15669 9428
rect 15627 9379 15669 9388
rect 11211 9337 11253 9346
rect 11115 9295 11157 9304
rect 1419 9260 1461 9269
rect 1419 9220 1420 9260
rect 1460 9220 1461 9260
rect 1419 9211 1461 9220
rect 5355 9260 5397 9269
rect 5355 9220 5356 9260
rect 5396 9220 5397 9260
rect 5355 9211 5397 9220
rect 7851 9260 7893 9269
rect 7851 9220 7852 9260
rect 7892 9220 7893 9260
rect 7851 9211 7893 9220
rect 10635 9260 10677 9269
rect 10635 9220 10636 9260
rect 10676 9220 10677 9260
rect 10635 9211 10677 9220
rect 12939 9260 12981 9269
rect 12939 9220 12940 9260
rect 12980 9220 12981 9260
rect 12939 9211 12981 9220
rect 17451 9260 17493 9269
rect 17451 9220 17452 9260
rect 17492 9220 17493 9260
rect 17451 9211 17493 9220
rect 19755 9260 19797 9269
rect 19755 9220 19756 9260
rect 19796 9220 19797 9260
rect 19755 9211 19797 9220
rect 20235 9260 20277 9269
rect 20235 9220 20236 9260
rect 20276 9220 20277 9260
rect 20235 9211 20277 9220
rect 1152 9092 20352 9116
rect 1152 9052 3688 9092
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 4056 9052 18808 9092
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 19176 9052 20352 9092
rect 1152 9028 20352 9052
rect 6795 8924 6837 8933
rect 6795 8884 6796 8924
rect 6836 8884 6837 8924
rect 6795 8875 6837 8884
rect 6987 8924 7029 8933
rect 6987 8884 6988 8924
rect 7028 8884 7029 8924
rect 6987 8875 7029 8884
rect 11595 8924 11637 8933
rect 11595 8884 11596 8924
rect 11636 8884 11637 8924
rect 11595 8875 11637 8884
rect 15051 8924 15093 8933
rect 15051 8884 15052 8924
rect 15092 8884 15093 8924
rect 15051 8875 15093 8884
rect 16683 8924 16725 8933
rect 16683 8884 16684 8924
rect 16724 8884 16725 8924
rect 16683 8875 16725 8884
rect 1227 8840 1269 8849
rect 1227 8800 1228 8840
rect 1268 8800 1269 8840
rect 1227 8791 1269 8800
rect 1611 8840 1653 8849
rect 1611 8800 1612 8840
rect 1652 8800 1653 8840
rect 1611 8791 1653 8800
rect 1995 8840 2037 8849
rect 1995 8800 1996 8840
rect 2036 8800 2037 8840
rect 1995 8791 2037 8800
rect 4395 8840 4437 8849
rect 4395 8800 4396 8840
rect 4436 8800 4437 8840
rect 4395 8791 4437 8800
rect 12547 8840 12605 8841
rect 12547 8800 12556 8840
rect 12596 8800 12605 8840
rect 12547 8799 12605 8800
rect 13035 8840 13077 8849
rect 13035 8800 13036 8840
rect 13076 8800 13077 8840
rect 13035 8791 13077 8800
rect 18211 8840 18269 8841
rect 18211 8800 18220 8840
rect 18260 8800 18269 8840
rect 18211 8799 18269 8800
rect 4568 8767 4626 8768
rect 1411 8756 1469 8757
rect 1411 8716 1420 8756
rect 1460 8716 1469 8756
rect 1411 8715 1469 8716
rect 1795 8756 1853 8757
rect 1795 8716 1804 8756
rect 1844 8716 1853 8756
rect 2955 8756 2997 8765
rect 1795 8715 1853 8716
rect 2179 8743 2237 8744
rect 2179 8703 2188 8743
rect 2228 8703 2237 8743
rect 2955 8716 2956 8756
rect 2996 8716 2997 8756
rect 4568 8727 4577 8767
rect 4617 8727 4626 8767
rect 4568 8726 4626 8727
rect 13411 8756 13469 8757
rect 2955 8707 2997 8716
rect 13411 8716 13420 8756
rect 13460 8716 13469 8756
rect 13411 8715 13469 8716
rect 2179 8702 2237 8703
rect 10827 8686 10869 8695
rect 2475 8672 2517 8681
rect 2475 8632 2476 8672
rect 2516 8632 2517 8672
rect 2475 8623 2517 8632
rect 2571 8672 2613 8681
rect 2571 8632 2572 8672
rect 2612 8632 2613 8672
rect 2571 8623 2613 8632
rect 3051 8672 3093 8681
rect 4011 8677 4053 8686
rect 3051 8632 3052 8672
rect 3092 8632 3093 8672
rect 3051 8623 3093 8632
rect 3523 8672 3581 8673
rect 3523 8632 3532 8672
rect 3572 8632 3581 8672
rect 3523 8631 3581 8632
rect 4011 8637 4012 8677
rect 4052 8637 4053 8677
rect 4011 8628 4053 8637
rect 4971 8672 5013 8681
rect 4971 8632 4972 8672
rect 5012 8632 5013 8672
rect 4971 8623 5013 8632
rect 5163 8672 5205 8681
rect 5163 8632 5164 8672
rect 5204 8632 5205 8672
rect 5163 8623 5205 8632
rect 5347 8672 5405 8673
rect 5347 8632 5356 8672
rect 5396 8632 5405 8672
rect 5347 8631 5405 8632
rect 6595 8672 6653 8673
rect 6595 8632 6604 8672
rect 6644 8632 6653 8672
rect 6595 8631 6653 8632
rect 7171 8672 7229 8673
rect 7171 8632 7180 8672
rect 7220 8632 7229 8672
rect 7171 8631 7229 8632
rect 8419 8672 8477 8673
rect 8419 8632 8428 8672
rect 8468 8632 8477 8672
rect 8419 8631 8477 8632
rect 8715 8672 8757 8681
rect 8715 8632 8716 8672
rect 8756 8632 8757 8672
rect 8907 8672 8949 8681
rect 8715 8623 8757 8632
rect 8811 8651 8853 8660
rect 8811 8611 8812 8651
rect 8852 8611 8853 8651
rect 8907 8632 8908 8672
rect 8948 8632 8949 8672
rect 8907 8623 8949 8632
rect 9003 8672 9045 8681
rect 9003 8632 9004 8672
rect 9044 8632 9045 8672
rect 9003 8623 9045 8632
rect 9291 8672 9333 8681
rect 9291 8632 9292 8672
rect 9332 8632 9333 8672
rect 9291 8623 9333 8632
rect 9387 8672 9429 8681
rect 9387 8632 9388 8672
rect 9428 8632 9429 8672
rect 9387 8623 9429 8632
rect 9771 8672 9813 8681
rect 9771 8632 9772 8672
rect 9812 8632 9813 8672
rect 9771 8623 9813 8632
rect 9867 8672 9909 8681
rect 9867 8632 9868 8672
rect 9908 8632 9909 8672
rect 9867 8623 9909 8632
rect 10339 8672 10397 8673
rect 10339 8632 10348 8672
rect 10388 8632 10397 8672
rect 10827 8646 10828 8686
rect 10868 8646 10869 8686
rect 11403 8672 11445 8681
rect 10827 8637 10869 8646
rect 11299 8657 11357 8658
rect 10339 8631 10397 8632
rect 11299 8617 11308 8657
rect 11348 8617 11357 8657
rect 11403 8632 11404 8672
rect 11444 8632 11445 8672
rect 11403 8623 11445 8632
rect 11595 8672 11637 8681
rect 11595 8632 11596 8672
rect 11636 8632 11637 8672
rect 11595 8623 11637 8632
rect 11875 8672 11933 8673
rect 11875 8632 11884 8672
rect 11924 8632 11933 8672
rect 11875 8631 11933 8632
rect 12171 8672 12213 8681
rect 12171 8632 12172 8672
rect 12212 8632 12213 8672
rect 12171 8623 12213 8632
rect 12739 8672 12797 8673
rect 12739 8632 12748 8672
rect 12788 8632 12797 8672
rect 12739 8631 12797 8632
rect 12843 8672 12885 8681
rect 12843 8632 12844 8672
rect 12884 8632 12885 8672
rect 12843 8623 12885 8632
rect 13035 8672 13077 8681
rect 13035 8632 13036 8672
rect 13076 8632 13077 8672
rect 13035 8623 13077 8632
rect 13603 8672 13661 8673
rect 13603 8632 13612 8672
rect 13652 8632 13661 8672
rect 13603 8631 13661 8632
rect 14851 8672 14909 8673
rect 14851 8632 14860 8672
rect 14900 8632 14909 8672
rect 14851 8631 14909 8632
rect 15235 8672 15293 8673
rect 15235 8632 15244 8672
rect 15284 8632 15293 8672
rect 15235 8631 15293 8632
rect 16483 8672 16541 8673
rect 16483 8632 16492 8672
rect 16532 8632 16541 8672
rect 16483 8631 16541 8632
rect 16875 8672 16917 8681
rect 16875 8632 16876 8672
rect 16916 8632 16917 8672
rect 17067 8672 17109 8681
rect 16875 8623 16917 8632
rect 16971 8651 17013 8660
rect 11299 8616 11357 8617
rect 8811 8602 8853 8611
rect 16971 8611 16972 8651
rect 17012 8611 17013 8651
rect 17067 8632 17068 8672
rect 17108 8632 17109 8672
rect 17067 8623 17109 8632
rect 17355 8672 17397 8681
rect 17355 8632 17356 8672
rect 17396 8632 17397 8672
rect 17355 8623 17397 8632
rect 17643 8672 17685 8681
rect 17643 8632 17644 8672
rect 17684 8632 17685 8672
rect 17643 8623 17685 8632
rect 17835 8672 17877 8681
rect 17835 8632 17836 8672
rect 17876 8632 17877 8672
rect 17835 8623 17877 8632
rect 18027 8672 18069 8681
rect 18027 8632 18028 8672
rect 18068 8632 18069 8672
rect 18027 8623 18069 8632
rect 18603 8672 18645 8681
rect 18603 8632 18604 8672
rect 18644 8632 18645 8672
rect 18603 8623 18645 8632
rect 18883 8672 18941 8673
rect 18883 8632 18892 8672
rect 18932 8632 18941 8672
rect 18883 8631 18941 8632
rect 19179 8672 19221 8681
rect 19179 8632 19180 8672
rect 19220 8632 19221 8672
rect 19179 8623 19221 8632
rect 19371 8672 19413 8681
rect 19371 8632 19372 8672
rect 19412 8632 19413 8672
rect 19371 8623 19413 8632
rect 19459 8672 19517 8673
rect 19459 8632 19468 8672
rect 19508 8632 19517 8672
rect 19459 8631 19517 8632
rect 19659 8672 19701 8681
rect 19659 8632 19660 8672
rect 19700 8632 19701 8672
rect 19851 8672 19893 8681
rect 19659 8623 19701 8632
rect 19755 8651 19797 8660
rect 16971 8602 17013 8611
rect 19755 8611 19756 8651
rect 19796 8611 19797 8651
rect 19851 8632 19852 8672
rect 19892 8632 19893 8672
rect 19851 8623 19893 8632
rect 19947 8672 19989 8681
rect 19947 8632 19948 8672
rect 19988 8632 19989 8672
rect 19947 8623 19989 8632
rect 20126 8661 20168 8670
rect 20126 8621 20127 8661
rect 20167 8621 20168 8661
rect 20126 8612 20168 8621
rect 19755 8602 19797 8611
rect 4203 8588 4245 8597
rect 4203 8548 4204 8588
rect 4244 8548 4245 8588
rect 4203 8539 4245 8548
rect 12267 8588 12309 8597
rect 12267 8548 12268 8588
rect 12308 8548 12309 8588
rect 12267 8539 12309 8548
rect 17163 8588 17205 8597
rect 17163 8548 17164 8588
rect 17204 8548 17205 8588
rect 17163 8539 17205 8548
rect 18507 8588 18549 8597
rect 18507 8548 18508 8588
rect 18548 8548 18549 8588
rect 18507 8539 18549 8548
rect 5067 8504 5109 8513
rect 5067 8464 5068 8504
rect 5108 8464 5109 8504
rect 5067 8455 5109 8464
rect 6795 8504 6837 8513
rect 6795 8464 6796 8504
rect 6836 8464 6837 8504
rect 6795 8455 6837 8464
rect 6987 8504 7029 8513
rect 6987 8464 6988 8504
rect 7028 8464 7029 8504
rect 6987 8455 7029 8464
rect 11019 8504 11061 8513
rect 11019 8464 11020 8504
rect 11060 8464 11061 8504
rect 11019 8455 11061 8464
rect 13227 8504 13269 8513
rect 13227 8464 13228 8504
rect 13268 8464 13269 8504
rect 13227 8455 13269 8464
rect 17451 8504 17493 8513
rect 17451 8464 17452 8504
rect 17492 8464 17493 8504
rect 17451 8455 17493 8464
rect 17931 8504 17973 8513
rect 17931 8464 17932 8504
rect 17972 8464 17973 8504
rect 17931 8455 17973 8464
rect 19267 8504 19325 8505
rect 19267 8464 19276 8504
rect 19316 8464 19325 8504
rect 19267 8463 19325 8464
rect 20235 8504 20277 8513
rect 20235 8464 20236 8504
rect 20276 8464 20277 8504
rect 20235 8455 20277 8464
rect 1152 8336 20452 8360
rect 1152 8296 4928 8336
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 5296 8296 20048 8336
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20416 8296 20452 8336
rect 1152 8272 20452 8296
rect 1227 8168 1269 8177
rect 1227 8128 1228 8168
rect 1268 8128 1269 8168
rect 1227 8119 1269 8128
rect 3051 8168 3093 8177
rect 3051 8128 3052 8168
rect 3092 8128 3093 8168
rect 3051 8119 3093 8128
rect 5259 8168 5301 8177
rect 5259 8128 5260 8168
rect 5300 8128 5301 8168
rect 5259 8119 5301 8128
rect 7267 8168 7325 8169
rect 7267 8128 7276 8168
rect 7316 8128 7325 8168
rect 7267 8127 7325 8128
rect 12547 8168 12605 8169
rect 12547 8128 12556 8168
rect 12596 8128 12605 8168
rect 12547 8127 12605 8128
rect 13131 8168 13173 8177
rect 13131 8128 13132 8168
rect 13172 8128 13173 8168
rect 13131 8119 13173 8128
rect 14955 8168 14997 8177
rect 14955 8128 14956 8168
rect 14996 8128 14997 8168
rect 14955 8119 14997 8128
rect 17155 8168 17213 8169
rect 17155 8128 17164 8168
rect 17204 8128 17213 8168
rect 17155 8127 17213 8128
rect 17539 8168 17597 8169
rect 17539 8128 17548 8168
rect 17588 8128 17597 8168
rect 17539 8127 17597 8128
rect 20131 8168 20189 8169
rect 20131 8128 20140 8168
rect 20180 8128 20189 8168
rect 20131 8127 20189 8128
rect 14763 8084 14805 8093
rect 14763 8044 14764 8084
rect 14804 8044 14805 8084
rect 14763 8035 14805 8044
rect 1603 8000 1661 8001
rect 1603 7960 1612 8000
rect 1652 7960 1661 8000
rect 3435 8000 3477 8009
rect 1603 7959 1661 7960
rect 2851 7979 2909 7980
rect 2851 7939 2860 7979
rect 2900 7939 2909 7979
rect 3435 7960 3436 8000
rect 3476 7960 3477 8000
rect 3435 7951 3477 7960
rect 3627 8000 3669 8009
rect 3627 7960 3628 8000
rect 3668 7960 3669 8000
rect 3627 7951 3669 7960
rect 3811 8000 3869 8001
rect 3811 7960 3820 8000
rect 3860 7960 3869 8000
rect 3811 7959 3869 7960
rect 5059 8000 5117 8001
rect 5059 7960 5068 8000
rect 5108 7960 5117 8000
rect 5059 7959 5117 7960
rect 5443 8000 5501 8001
rect 5443 7960 5452 8000
rect 5492 7960 5501 8000
rect 5443 7959 5501 7960
rect 6691 8000 6749 8001
rect 6691 7960 6700 8000
rect 6740 7960 6749 8000
rect 6691 7959 6749 7960
rect 7075 8000 7133 8001
rect 7075 7960 7084 8000
rect 7124 7960 7133 8000
rect 7075 7959 7133 7960
rect 7179 8000 7221 8009
rect 7179 7960 7180 8000
rect 7220 7960 7221 8000
rect 7179 7951 7221 7960
rect 7371 8000 7413 8009
rect 7371 7960 7372 8000
rect 7412 7960 7413 8000
rect 7371 7951 7413 7960
rect 7555 8000 7613 8001
rect 7555 7960 7564 8000
rect 7604 7960 7613 8000
rect 7555 7959 7613 7960
rect 8803 8000 8861 8001
rect 8803 7960 8812 8000
rect 8852 7960 8861 8000
rect 8803 7959 8861 7960
rect 9187 8000 9245 8001
rect 9187 7960 9196 8000
rect 9236 7960 9245 8000
rect 9187 7959 9245 7960
rect 10435 8000 10493 8001
rect 10435 7960 10444 8000
rect 10484 7960 10493 8000
rect 10435 7959 10493 7960
rect 10915 8000 10973 8001
rect 10915 7960 10924 8000
rect 10964 7960 10973 8000
rect 10915 7959 10973 7960
rect 12163 8000 12221 8001
rect 12163 7960 12172 8000
rect 12212 7960 12221 8000
rect 12163 7959 12221 7960
rect 12747 8000 12789 8009
rect 12747 7960 12748 8000
rect 12788 7960 12789 8000
rect 12747 7951 12789 7960
rect 12843 8000 12885 8009
rect 12843 7960 12844 8000
rect 12884 7960 12885 8000
rect 12843 7951 12885 7960
rect 13027 8000 13085 8001
rect 13027 7960 13036 8000
rect 13076 7960 13085 8000
rect 13027 7959 13085 7960
rect 13315 8000 13373 8001
rect 13315 7960 13324 8000
rect 13364 7960 13373 8000
rect 13315 7959 13373 7960
rect 14563 8000 14621 8001
rect 14563 7960 14572 8000
rect 14612 7960 14621 8000
rect 15619 8000 15677 8001
rect 14563 7959 14621 7960
rect 15147 7986 15189 7995
rect 2851 7938 2909 7939
rect 15147 7946 15148 7986
rect 15188 7946 15189 7986
rect 15619 7960 15628 8000
rect 15668 7960 15677 8000
rect 15619 7959 15677 7960
rect 16107 8000 16149 8009
rect 16107 7960 16108 8000
rect 16148 7960 16149 8000
rect 16107 7951 16149 7960
rect 16203 8000 16245 8009
rect 16203 7960 16204 8000
rect 16244 7960 16245 8000
rect 16203 7951 16245 7960
rect 16587 8000 16629 8009
rect 16587 7960 16588 8000
rect 16628 7960 16629 8000
rect 16587 7951 16629 7960
rect 16683 8000 16725 8009
rect 16683 7960 16684 8000
rect 16724 7960 16725 8000
rect 16683 7951 16725 7960
rect 16963 8000 17021 8001
rect 16963 7960 16972 8000
rect 17012 7960 17021 8000
rect 16963 7959 17021 7960
rect 17067 8000 17109 8009
rect 17067 7960 17068 8000
rect 17108 7960 17109 8000
rect 17067 7951 17109 7960
rect 17259 8000 17301 8009
rect 17259 7960 17260 8000
rect 17300 7960 17301 8000
rect 17259 7951 17301 7960
rect 17451 8000 17493 8009
rect 17451 7960 17452 8000
rect 17492 7960 17493 8000
rect 17451 7951 17493 7960
rect 17643 8000 17685 8009
rect 17643 7960 17644 8000
rect 17684 7960 17685 8000
rect 17643 7951 17685 7960
rect 17731 8000 17789 8001
rect 17731 7960 17740 8000
rect 17780 7960 17789 8000
rect 17731 7959 17789 7960
rect 17923 8000 17981 8001
rect 17923 7960 17932 8000
rect 17972 7960 17981 8000
rect 17923 7959 17981 7960
rect 18211 8000 18269 8001
rect 18211 7960 18220 8000
rect 18260 7960 18269 8000
rect 18211 7959 18269 7960
rect 19459 8000 19517 8001
rect 19459 7960 19468 8000
rect 19508 7960 19517 8000
rect 19459 7959 19517 7960
rect 19851 8000 19893 8009
rect 19851 7960 19852 8000
rect 19892 7960 19893 8000
rect 19851 7951 19893 7960
rect 19947 8000 19989 8009
rect 19947 7960 19948 8000
rect 19988 7960 19989 8000
rect 19947 7951 19989 7960
rect 15147 7937 15189 7946
rect 1411 7916 1469 7917
rect 1411 7876 1420 7916
rect 1460 7876 1469 7916
rect 1411 7875 1469 7876
rect 3531 7916 3573 7925
rect 3531 7876 3532 7916
rect 3572 7876 3573 7916
rect 3531 7867 3573 7876
rect 6891 7748 6933 7757
rect 6891 7708 6892 7748
rect 6932 7708 6933 7748
rect 6891 7699 6933 7708
rect 9003 7748 9045 7757
rect 9003 7708 9004 7748
rect 9044 7708 9045 7748
rect 9003 7699 9045 7708
rect 10635 7748 10677 7757
rect 10635 7708 10636 7748
rect 10676 7708 10677 7748
rect 10635 7699 10677 7708
rect 12363 7748 12405 7757
rect 12363 7708 12364 7748
rect 12404 7708 12405 7748
rect 12363 7699 12405 7708
rect 18027 7748 18069 7757
rect 18027 7708 18028 7748
rect 18068 7708 18069 7748
rect 18027 7699 18069 7708
rect 19659 7748 19701 7757
rect 19659 7708 19660 7748
rect 19700 7708 19701 7748
rect 19659 7699 19701 7708
rect 1152 7580 20352 7604
rect 1152 7540 3688 7580
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 4056 7540 18808 7580
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 19176 7540 20352 7580
rect 1152 7516 20352 7540
rect 2763 7412 2805 7421
rect 2763 7372 2764 7412
rect 2804 7372 2805 7412
rect 2763 7363 2805 7372
rect 5163 7412 5205 7421
rect 5163 7372 5164 7412
rect 5204 7372 5205 7412
rect 5163 7363 5205 7372
rect 14763 7412 14805 7421
rect 14763 7372 14764 7412
rect 14804 7372 14805 7412
rect 14763 7363 14805 7372
rect 20139 7412 20181 7421
rect 20139 7372 20140 7412
rect 20180 7372 20181 7412
rect 20139 7363 20181 7372
rect 18595 7328 18653 7329
rect 18595 7288 18604 7328
rect 18644 7288 18653 7328
rect 18595 7287 18653 7288
rect 19755 7328 19797 7337
rect 19755 7288 19756 7328
rect 19796 7288 19797 7328
rect 19755 7279 19797 7288
rect 3531 7244 3573 7253
rect 3531 7204 3532 7244
rect 3572 7204 3573 7244
rect 3531 7195 3573 7204
rect 10635 7244 10677 7253
rect 10635 7204 10636 7244
rect 10676 7204 10677 7244
rect 10635 7195 10677 7204
rect 10731 7244 10773 7253
rect 10731 7204 10732 7244
rect 10772 7204 10773 7244
rect 10731 7195 10773 7204
rect 12747 7244 12789 7253
rect 12747 7204 12748 7244
rect 12788 7204 12789 7244
rect 12747 7195 12789 7204
rect 17067 7244 17109 7253
rect 17067 7204 17068 7244
rect 17108 7204 17109 7244
rect 17067 7195 17109 7204
rect 19659 7244 19701 7253
rect 19659 7204 19660 7244
rect 19700 7204 19701 7244
rect 19659 7195 19701 7204
rect 19851 7244 19893 7253
rect 19851 7204 19852 7244
rect 19892 7204 19893 7244
rect 19851 7195 19893 7204
rect 6987 7174 7029 7183
rect 1315 7160 1373 7161
rect 1315 7120 1324 7160
rect 1364 7120 1373 7160
rect 1315 7119 1373 7120
rect 2563 7160 2621 7161
rect 2563 7120 2572 7160
rect 2612 7120 2621 7160
rect 2563 7119 2621 7120
rect 3051 7160 3093 7169
rect 3051 7120 3052 7160
rect 3092 7120 3093 7160
rect 3051 7111 3093 7120
rect 3147 7160 3189 7169
rect 3147 7120 3148 7160
rect 3188 7120 3189 7160
rect 3147 7111 3189 7120
rect 3627 7160 3669 7169
rect 4587 7165 4629 7174
rect 3627 7120 3628 7160
rect 3668 7120 3669 7160
rect 3627 7111 3669 7120
rect 4099 7160 4157 7161
rect 4099 7120 4108 7160
rect 4148 7120 4157 7160
rect 4099 7119 4157 7120
rect 4587 7125 4588 7165
rect 4628 7125 4629 7165
rect 4587 7116 4629 7125
rect 4971 7160 5013 7169
rect 4971 7120 4972 7160
rect 5012 7120 5013 7160
rect 4971 7111 5013 7120
rect 5163 7160 5205 7169
rect 5163 7120 5164 7160
rect 5204 7120 5205 7160
rect 5163 7111 5205 7120
rect 5451 7160 5493 7169
rect 5451 7120 5452 7160
rect 5492 7120 5493 7160
rect 5451 7111 5493 7120
rect 5547 7160 5589 7169
rect 5547 7120 5548 7160
rect 5588 7120 5589 7160
rect 5547 7111 5589 7120
rect 5931 7160 5973 7169
rect 5931 7120 5932 7160
rect 5972 7120 5973 7160
rect 5931 7111 5973 7120
rect 6027 7160 6069 7169
rect 6027 7120 6028 7160
rect 6068 7120 6069 7160
rect 6027 7111 6069 7120
rect 6499 7160 6557 7161
rect 6499 7120 6508 7160
rect 6548 7120 6557 7160
rect 6987 7134 6988 7174
rect 7028 7134 7029 7174
rect 11739 7169 11781 7178
rect 13851 7169 13893 7178
rect 6987 7125 7029 7134
rect 7555 7160 7613 7161
rect 6499 7119 6557 7120
rect 7555 7120 7564 7160
rect 7604 7120 7613 7160
rect 7555 7119 7613 7120
rect 8803 7160 8861 7161
rect 8803 7120 8812 7160
rect 8852 7120 8861 7160
rect 8803 7119 8861 7120
rect 8995 7160 9053 7161
rect 8995 7120 9004 7160
rect 9044 7120 9053 7160
rect 8995 7119 9053 7120
rect 9099 7160 9141 7169
rect 9099 7120 9100 7160
rect 9140 7120 9141 7160
rect 9099 7111 9141 7120
rect 9291 7160 9333 7169
rect 9291 7120 9292 7160
rect 9332 7120 9333 7160
rect 9291 7111 9333 7120
rect 9475 7160 9533 7161
rect 9475 7120 9484 7160
rect 9524 7120 9533 7160
rect 9475 7119 9533 7120
rect 9579 7160 9621 7169
rect 9579 7120 9580 7160
rect 9620 7120 9621 7160
rect 9579 7111 9621 7120
rect 9771 7160 9813 7169
rect 9771 7120 9772 7160
rect 9812 7120 9813 7160
rect 9771 7111 9813 7120
rect 10155 7160 10197 7169
rect 10155 7120 10156 7160
rect 10196 7120 10197 7160
rect 10155 7111 10197 7120
rect 10251 7160 10293 7169
rect 10251 7120 10252 7160
rect 10292 7120 10293 7160
rect 10251 7111 10293 7120
rect 11203 7160 11261 7161
rect 11203 7120 11212 7160
rect 11252 7120 11261 7160
rect 11739 7129 11740 7169
rect 11780 7129 11781 7169
rect 11739 7120 11781 7129
rect 12267 7160 12309 7169
rect 12267 7120 12268 7160
rect 12308 7120 12309 7160
rect 11203 7119 11261 7120
rect 12267 7111 12309 7120
rect 12363 7160 12405 7169
rect 12363 7120 12364 7160
rect 12404 7120 12405 7160
rect 12363 7111 12405 7120
rect 12843 7160 12885 7169
rect 12843 7120 12844 7160
rect 12884 7120 12885 7160
rect 12843 7111 12885 7120
rect 13315 7160 13373 7161
rect 13315 7120 13324 7160
rect 13364 7120 13373 7160
rect 13851 7129 13852 7169
rect 13892 7129 13893 7169
rect 13851 7120 13893 7129
rect 14276 7162 14334 7163
rect 14276 7122 14285 7162
rect 14325 7122 14334 7162
rect 14276 7121 14334 7122
rect 14379 7160 14421 7169
rect 14379 7120 14380 7160
rect 14420 7120 14421 7160
rect 13315 7119 13373 7120
rect 14379 7111 14421 7120
rect 14571 7160 14613 7169
rect 14571 7120 14572 7160
rect 14612 7120 14613 7160
rect 14571 7111 14613 7120
rect 14947 7160 15005 7161
rect 14947 7120 14956 7160
rect 14996 7120 15005 7160
rect 14947 7119 15005 7120
rect 16195 7160 16253 7161
rect 16195 7120 16204 7160
rect 16244 7120 16253 7160
rect 16195 7119 16253 7120
rect 16491 7160 16533 7169
rect 16491 7120 16492 7160
rect 16532 7120 16533 7160
rect 16491 7111 16533 7120
rect 16587 7160 16629 7169
rect 16587 7120 16588 7160
rect 16628 7120 16629 7160
rect 16587 7111 16629 7120
rect 16971 7160 17013 7169
rect 18027 7165 18069 7174
rect 16971 7120 16972 7160
rect 17012 7120 17013 7160
rect 16971 7111 17013 7120
rect 17539 7160 17597 7161
rect 17539 7120 17548 7160
rect 17588 7120 17597 7160
rect 17539 7119 17597 7120
rect 18027 7125 18028 7165
rect 18068 7125 18069 7165
rect 18027 7116 18069 7125
rect 18891 7160 18933 7169
rect 18891 7120 18892 7160
rect 18932 7120 18933 7160
rect 18891 7111 18933 7120
rect 18987 7160 19029 7169
rect 18987 7120 18988 7160
rect 19028 7120 19029 7160
rect 18987 7111 19029 7120
rect 19267 7160 19325 7161
rect 19267 7120 19276 7160
rect 19316 7120 19325 7160
rect 19267 7119 19325 7120
rect 19563 7160 19605 7169
rect 19563 7120 19564 7160
rect 19604 7120 19605 7160
rect 19563 7111 19605 7120
rect 19939 7160 19997 7161
rect 19939 7120 19948 7160
rect 19988 7120 19997 7160
rect 19939 7119 19997 7120
rect 20227 7160 20285 7161
rect 20227 7120 20236 7160
rect 20276 7120 20285 7160
rect 20227 7119 20285 7120
rect 7179 7076 7221 7085
rect 7179 7036 7180 7076
rect 7220 7036 7221 7076
rect 7179 7027 7221 7036
rect 9675 7076 9717 7085
rect 9675 7036 9676 7076
rect 9716 7036 9717 7076
rect 9675 7027 9717 7036
rect 11883 7076 11925 7085
rect 11883 7036 11884 7076
rect 11924 7036 11925 7076
rect 11883 7027 11925 7036
rect 13995 7076 14037 7085
rect 13995 7036 13996 7076
rect 14036 7036 14037 7076
rect 13995 7027 14037 7036
rect 4779 6992 4821 7001
rect 4779 6952 4780 6992
rect 4820 6952 4821 6992
rect 4779 6943 4821 6952
rect 7371 6992 7413 7001
rect 7371 6952 7372 6992
rect 7412 6952 7413 6992
rect 7371 6943 7413 6952
rect 9187 6992 9245 6993
rect 9187 6952 9196 6992
rect 9236 6952 9245 6992
rect 9187 6951 9245 6952
rect 14467 6992 14525 6993
rect 14467 6952 14476 6992
rect 14516 6952 14525 6992
rect 14467 6951 14525 6952
rect 18219 6992 18261 7001
rect 18219 6952 18220 6992
rect 18260 6952 18261 6992
rect 18219 6943 18261 6952
rect 1152 6824 20452 6848
rect 1152 6784 4928 6824
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 5296 6784 20048 6824
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20416 6784 20452 6824
rect 1152 6760 20452 6784
rect 8427 6714 8469 6723
rect 8427 6674 8428 6714
rect 8468 6674 8469 6714
rect 8427 6665 8469 6674
rect 9387 6698 9429 6707
rect 1227 6656 1269 6665
rect 1227 6616 1228 6656
rect 1268 6616 1269 6656
rect 1227 6607 1269 6616
rect 1611 6656 1653 6665
rect 1611 6616 1612 6656
rect 1652 6616 1653 6656
rect 1611 6607 1653 6616
rect 2091 6656 2133 6665
rect 2091 6616 2092 6656
rect 2132 6616 2133 6656
rect 2091 6607 2133 6616
rect 4203 6656 4245 6665
rect 9387 6658 9388 6698
rect 9428 6658 9429 6698
rect 4203 6616 4204 6656
rect 4244 6616 4245 6656
rect 4203 6607 4245 6616
rect 6499 6656 6557 6657
rect 6499 6616 6508 6656
rect 6548 6616 6557 6656
rect 9387 6649 9429 6658
rect 11883 6656 11925 6665
rect 6499 6615 6557 6616
rect 11883 6616 11884 6656
rect 11924 6616 11925 6656
rect 11883 6607 11925 6616
rect 12075 6656 12117 6665
rect 12075 6616 12076 6656
rect 12116 6616 12117 6656
rect 12075 6607 12117 6616
rect 13899 6656 13941 6665
rect 13899 6616 13900 6656
rect 13940 6616 13941 6656
rect 13899 6607 13941 6616
rect 15819 6656 15861 6665
rect 15819 6616 15820 6656
rect 15860 6616 15861 6656
rect 15819 6607 15861 6616
rect 18499 6656 18557 6657
rect 18499 6616 18508 6656
rect 18548 6616 18557 6656
rect 18499 6615 18557 6616
rect 4395 6572 4437 6581
rect 4395 6532 4396 6572
rect 4436 6532 4437 6572
rect 4395 6523 4437 6532
rect 6891 6572 6933 6581
rect 6891 6532 6892 6572
rect 6932 6532 6933 6572
rect 6891 6523 6933 6532
rect 9099 6572 9141 6581
rect 9099 6532 9100 6572
rect 9140 6532 9141 6572
rect 9099 6523 9141 6532
rect 1995 6488 2037 6497
rect 1995 6448 1996 6488
rect 2036 6448 2037 6488
rect 1995 6439 2037 6448
rect 2187 6488 2229 6497
rect 2187 6448 2188 6488
rect 2228 6448 2229 6488
rect 2187 6439 2229 6448
rect 2379 6488 2421 6497
rect 2379 6448 2380 6488
rect 2420 6448 2421 6488
rect 2379 6439 2421 6448
rect 2571 6488 2613 6497
rect 2571 6448 2572 6488
rect 2612 6448 2613 6488
rect 2571 6439 2613 6448
rect 2755 6488 2813 6489
rect 2755 6448 2764 6488
rect 2804 6448 2813 6488
rect 2755 6447 2813 6448
rect 4003 6488 4061 6489
rect 4003 6448 4012 6488
rect 4052 6448 4061 6488
rect 5059 6488 5117 6489
rect 4003 6447 4061 6448
rect 4587 6474 4629 6483
rect 4587 6434 4588 6474
rect 4628 6434 4629 6474
rect 5059 6448 5068 6488
rect 5108 6448 5117 6488
rect 5059 6447 5117 6448
rect 5547 6488 5589 6497
rect 5547 6448 5548 6488
rect 5588 6448 5589 6488
rect 5547 6439 5589 6448
rect 5643 6488 5685 6497
rect 5643 6448 5644 6488
rect 5684 6448 5685 6488
rect 5643 6439 5685 6448
rect 6027 6488 6069 6497
rect 6027 6448 6028 6488
rect 6068 6448 6069 6488
rect 6027 6439 6069 6448
rect 6123 6488 6165 6497
rect 6123 6448 6124 6488
rect 6164 6448 6165 6488
rect 6123 6439 6165 6448
rect 6411 6488 6453 6497
rect 6411 6448 6412 6488
rect 6452 6448 6453 6488
rect 6411 6439 6453 6448
rect 6603 6488 6645 6497
rect 6603 6448 6604 6488
rect 6644 6448 6645 6488
rect 6603 6439 6645 6448
rect 6691 6488 6749 6489
rect 6691 6448 6700 6488
rect 6740 6448 6749 6488
rect 6691 6447 6749 6448
rect 6987 6488 7029 6497
rect 6987 6448 6988 6488
rect 7028 6448 7029 6488
rect 6987 6439 7029 6448
rect 7083 6488 7125 6497
rect 7083 6448 7084 6488
rect 7124 6448 7125 6488
rect 7083 6439 7125 6448
rect 7179 6488 7221 6497
rect 7179 6448 7180 6488
rect 7220 6448 7221 6488
rect 7179 6439 7221 6448
rect 7363 6488 7421 6489
rect 7363 6448 7372 6488
rect 7412 6448 7421 6488
rect 7363 6447 7421 6448
rect 7755 6488 7797 6497
rect 7755 6448 7756 6488
rect 7796 6448 7797 6488
rect 7755 6439 7797 6448
rect 8235 6488 8277 6497
rect 8235 6448 8236 6488
rect 8276 6448 8277 6488
rect 8235 6439 8277 6448
rect 8323 6488 8381 6489
rect 8323 6448 8332 6488
rect 8372 6448 8381 6488
rect 8323 6447 8381 6448
rect 8707 6488 8765 6489
rect 8707 6448 8716 6488
rect 8756 6448 8765 6488
rect 8707 6447 8765 6448
rect 9003 6488 9045 6497
rect 9003 6448 9004 6488
rect 9044 6448 9045 6488
rect 9003 6439 9045 6448
rect 9579 6488 9621 6497
rect 9579 6448 9580 6488
rect 9620 6448 9621 6488
rect 9579 6439 9621 6448
rect 9867 6488 9909 6497
rect 9867 6448 9868 6488
rect 9908 6448 9909 6488
rect 9867 6439 9909 6448
rect 10059 6488 10101 6497
rect 10059 6448 10060 6488
rect 10100 6448 10101 6488
rect 10059 6439 10101 6448
rect 10251 6487 10293 6496
rect 10251 6447 10252 6487
rect 10292 6447 10293 6487
rect 10435 6488 10493 6489
rect 10435 6448 10444 6488
rect 10484 6448 10493 6488
rect 10435 6447 10493 6448
rect 11683 6488 11741 6489
rect 11683 6448 11692 6488
rect 11732 6448 11741 6488
rect 11683 6447 11741 6448
rect 12451 6488 12509 6489
rect 12451 6448 12460 6488
rect 12500 6448 12509 6488
rect 12451 6447 12509 6448
rect 13699 6488 13757 6489
rect 13699 6448 13708 6488
rect 13748 6448 13757 6488
rect 13699 6447 13757 6448
rect 14083 6488 14141 6489
rect 14083 6448 14092 6488
rect 14132 6448 14141 6488
rect 14083 6447 14141 6448
rect 15331 6488 15389 6489
rect 15331 6448 15340 6488
rect 15380 6448 15389 6488
rect 15331 6447 15389 6448
rect 15723 6488 15765 6497
rect 15723 6448 15724 6488
rect 15764 6448 15765 6488
rect 10251 6438 10293 6447
rect 15723 6439 15765 6448
rect 15915 6488 15957 6497
rect 15915 6448 15916 6488
rect 15956 6448 15957 6488
rect 15915 6439 15957 6448
rect 16107 6488 16149 6497
rect 16107 6448 16108 6488
rect 16148 6448 16149 6488
rect 16107 6439 16149 6448
rect 16299 6488 16341 6497
rect 16299 6448 16300 6488
rect 16340 6448 16341 6488
rect 16299 6439 16341 6448
rect 16387 6488 16445 6489
rect 16387 6448 16396 6488
rect 16436 6448 16445 6488
rect 16387 6447 16445 6448
rect 16963 6488 17021 6489
rect 16963 6448 16972 6488
rect 17012 6448 17021 6488
rect 16963 6447 17021 6448
rect 17259 6488 17301 6497
rect 17259 6448 17260 6488
rect 17300 6448 17301 6488
rect 17259 6439 17301 6448
rect 17355 6488 17397 6497
rect 17355 6448 17356 6488
rect 17396 6448 17397 6488
rect 17355 6439 17397 6448
rect 17835 6488 17877 6497
rect 17835 6448 17836 6488
rect 17876 6448 17877 6488
rect 17835 6439 17877 6448
rect 18027 6488 18069 6497
rect 18027 6448 18028 6488
rect 18068 6448 18069 6488
rect 18027 6439 18069 6448
rect 18115 6488 18173 6489
rect 18115 6448 18124 6488
rect 18164 6448 18173 6488
rect 18115 6447 18173 6448
rect 18307 6488 18365 6489
rect 18307 6448 18316 6488
rect 18356 6448 18365 6488
rect 18307 6447 18365 6448
rect 18411 6488 18453 6497
rect 18411 6448 18412 6488
rect 18452 6448 18453 6488
rect 19187 6488 19229 6497
rect 18411 6439 18453 6448
rect 18603 6477 18645 6486
rect 4587 6425 4629 6434
rect 18603 6437 18604 6477
rect 18644 6437 18645 6477
rect 19187 6448 19188 6488
rect 19228 6448 19229 6488
rect 19187 6439 19229 6448
rect 19467 6488 19509 6497
rect 19467 6448 19468 6488
rect 19508 6448 19509 6488
rect 19467 6439 19509 6448
rect 19563 6488 19605 6497
rect 19563 6448 19564 6488
rect 19604 6448 19605 6488
rect 19563 6439 19605 6448
rect 20043 6488 20085 6497
rect 20043 6448 20044 6488
rect 20084 6448 20085 6488
rect 20043 6439 20085 6448
rect 20235 6488 20277 6497
rect 20235 6448 20236 6488
rect 20276 6448 20277 6488
rect 20235 6439 20277 6448
rect 18603 6428 18645 6437
rect 1411 6404 1469 6405
rect 1411 6364 1420 6404
rect 1460 6364 1469 6404
rect 1411 6363 1469 6364
rect 1795 6404 1853 6405
rect 1795 6364 1804 6404
rect 1844 6364 1853 6404
rect 1795 6363 1853 6364
rect 7467 6404 7509 6413
rect 7467 6364 7468 6404
rect 7508 6364 7509 6404
rect 7467 6355 7509 6364
rect 7659 6404 7701 6413
rect 7659 6364 7660 6404
rect 7700 6364 7701 6404
rect 7659 6355 7701 6364
rect 12259 6404 12317 6405
rect 12259 6364 12268 6404
rect 12308 6364 12317 6404
rect 12259 6363 12317 6364
rect 2379 6320 2421 6329
rect 2379 6280 2380 6320
rect 2420 6280 2421 6320
rect 2379 6271 2421 6280
rect 7563 6320 7605 6329
rect 7563 6280 7564 6320
rect 7604 6280 7605 6320
rect 7563 6271 7605 6280
rect 7947 6320 7989 6329
rect 7947 6280 7948 6320
rect 7988 6280 7989 6320
rect 7947 6271 7989 6280
rect 9579 6320 9621 6329
rect 9579 6280 9580 6320
rect 9620 6280 9621 6320
rect 9579 6271 9621 6280
rect 16587 6320 16629 6329
rect 16587 6280 16588 6320
rect 16628 6280 16629 6320
rect 16587 6271 16629 6280
rect 17635 6320 17693 6321
rect 17635 6280 17644 6320
rect 17684 6280 17693 6320
rect 17635 6279 17693 6280
rect 19843 6320 19901 6321
rect 19843 6280 19852 6320
rect 19892 6280 19901 6320
rect 19843 6279 19901 6280
rect 10059 6236 10101 6245
rect 10059 6196 10060 6236
rect 10100 6196 10101 6236
rect 10059 6187 10101 6196
rect 15531 6236 15573 6245
rect 15531 6196 15532 6236
rect 15572 6196 15573 6236
rect 15531 6187 15573 6196
rect 16107 6236 16149 6245
rect 16107 6196 16108 6236
rect 16148 6196 16149 6236
rect 16107 6187 16149 6196
rect 17835 6236 17877 6245
rect 17835 6196 17836 6236
rect 17876 6196 17877 6236
rect 17835 6187 17877 6196
rect 20043 6236 20085 6245
rect 20043 6196 20044 6236
rect 20084 6196 20085 6236
rect 20043 6187 20085 6196
rect 1152 6068 20352 6092
rect 1152 6028 3688 6068
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 4056 6028 18808 6068
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 19176 6028 20352 6068
rect 1152 6004 20352 6028
rect 3147 5900 3189 5909
rect 3147 5860 3148 5900
rect 3188 5860 3189 5900
rect 3147 5851 3189 5860
rect 5259 5900 5301 5909
rect 5259 5860 5260 5900
rect 5300 5860 5301 5900
rect 5259 5851 5301 5860
rect 6219 5900 6261 5909
rect 6219 5860 6220 5900
rect 6260 5860 6261 5900
rect 6219 5851 6261 5860
rect 9283 5900 9341 5901
rect 9283 5860 9292 5900
rect 9332 5860 9341 5900
rect 9283 5859 9341 5860
rect 20139 5900 20181 5909
rect 20139 5860 20140 5900
rect 20180 5860 20181 5900
rect 20139 5851 20181 5860
rect 2667 5816 2709 5825
rect 2667 5776 2668 5816
rect 2708 5776 2709 5816
rect 2667 5767 2709 5776
rect 9667 5816 9725 5817
rect 9667 5776 9676 5816
rect 9716 5776 9725 5816
rect 9667 5775 9725 5776
rect 15427 5816 15485 5817
rect 15427 5776 15436 5816
rect 15476 5776 15485 5816
rect 15427 5775 15485 5776
rect 13995 5732 14037 5741
rect 13995 5692 13996 5732
rect 14036 5692 14037 5732
rect 13995 5683 14037 5692
rect 15051 5662 15093 5671
rect 1219 5648 1277 5649
rect 1219 5608 1228 5648
rect 1268 5608 1277 5648
rect 1219 5607 1277 5608
rect 2467 5648 2525 5649
rect 2467 5608 2476 5648
rect 2516 5608 2525 5648
rect 2467 5607 2525 5608
rect 2859 5648 2901 5657
rect 2859 5608 2860 5648
rect 2900 5608 2901 5648
rect 2859 5599 2901 5608
rect 3147 5648 3189 5657
rect 3147 5608 3148 5648
rect 3188 5608 3189 5648
rect 3147 5599 3189 5608
rect 3435 5648 3477 5657
rect 3435 5608 3436 5648
rect 3476 5608 3477 5648
rect 3435 5599 3477 5608
rect 3531 5648 3573 5657
rect 3531 5608 3532 5648
rect 3572 5608 3573 5648
rect 3531 5599 3573 5608
rect 3627 5648 3669 5657
rect 3627 5608 3628 5648
rect 3668 5608 3669 5648
rect 3627 5599 3669 5608
rect 3811 5648 3869 5649
rect 3811 5608 3820 5648
rect 3860 5608 3869 5648
rect 3811 5607 3869 5608
rect 5059 5648 5117 5649
rect 5059 5608 5068 5648
rect 5108 5608 5117 5648
rect 5059 5607 5117 5608
rect 5451 5648 5493 5657
rect 5451 5608 5452 5648
rect 5492 5608 5493 5648
rect 5451 5599 5493 5608
rect 5643 5648 5685 5657
rect 5643 5608 5644 5648
rect 5684 5608 5685 5648
rect 5643 5599 5685 5608
rect 5731 5648 5789 5649
rect 5731 5608 5740 5648
rect 5780 5608 5789 5648
rect 5731 5607 5789 5608
rect 5931 5648 5973 5657
rect 5931 5608 5932 5648
rect 5972 5608 5973 5648
rect 5931 5599 5973 5608
rect 6219 5648 6261 5657
rect 6219 5608 6220 5648
rect 6260 5608 6261 5648
rect 6219 5599 6261 5608
rect 6411 5648 6453 5657
rect 6411 5608 6412 5648
rect 6452 5608 6453 5648
rect 6411 5599 6453 5608
rect 6507 5648 6549 5657
rect 6507 5608 6508 5648
rect 6548 5608 6549 5648
rect 6507 5599 6549 5608
rect 6603 5648 6645 5657
rect 6603 5608 6604 5648
rect 6644 5608 6645 5648
rect 6603 5599 6645 5608
rect 6699 5648 6741 5657
rect 6699 5608 6700 5648
rect 6740 5608 6741 5648
rect 6699 5599 6741 5608
rect 6883 5648 6941 5649
rect 6883 5608 6892 5648
rect 6932 5608 6941 5648
rect 6883 5607 6941 5608
rect 8131 5648 8189 5649
rect 8131 5608 8140 5648
rect 8180 5608 8189 5648
rect 8131 5607 8189 5608
rect 8611 5648 8669 5649
rect 8611 5608 8620 5648
rect 8660 5608 8669 5648
rect 8611 5607 8669 5608
rect 8907 5648 8949 5657
rect 8907 5608 8908 5648
rect 8948 5608 8949 5648
rect 8907 5599 8949 5608
rect 9483 5648 9525 5657
rect 9483 5608 9484 5648
rect 9524 5608 9525 5648
rect 9483 5599 9525 5608
rect 9675 5648 9717 5657
rect 9675 5608 9676 5648
rect 9716 5608 9717 5648
rect 9675 5599 9717 5608
rect 9771 5648 9813 5657
rect 9771 5608 9772 5648
rect 9812 5608 9813 5648
rect 9771 5599 9813 5608
rect 10147 5648 10205 5649
rect 10147 5608 10156 5648
rect 10196 5608 10205 5648
rect 10147 5607 10205 5608
rect 11395 5648 11453 5649
rect 11395 5608 11404 5648
rect 11444 5608 11453 5648
rect 11395 5607 11453 5608
rect 11779 5648 11837 5649
rect 11779 5608 11788 5648
rect 11828 5608 11837 5648
rect 11779 5607 11837 5608
rect 13027 5648 13085 5649
rect 13027 5608 13036 5648
rect 13076 5608 13085 5648
rect 13027 5607 13085 5608
rect 13515 5648 13557 5657
rect 13515 5608 13516 5648
rect 13556 5608 13557 5648
rect 13515 5599 13557 5608
rect 13611 5648 13653 5657
rect 13611 5608 13612 5648
rect 13652 5608 13653 5648
rect 13611 5599 13653 5608
rect 14091 5648 14133 5657
rect 14091 5608 14092 5648
rect 14132 5608 14133 5648
rect 14091 5599 14133 5608
rect 14563 5648 14621 5649
rect 14563 5608 14572 5648
rect 14612 5608 14621 5648
rect 15051 5622 15052 5662
rect 15092 5622 15093 5662
rect 15051 5613 15093 5622
rect 15819 5648 15861 5657
rect 14563 5607 14621 5608
rect 15819 5608 15820 5648
rect 15860 5608 15861 5648
rect 15819 5599 15861 5608
rect 16099 5648 16157 5649
rect 16099 5608 16108 5648
rect 16148 5608 16157 5648
rect 16099 5607 16157 5608
rect 16387 5648 16445 5649
rect 16387 5608 16396 5648
rect 16436 5608 16445 5648
rect 16387 5607 16445 5608
rect 17635 5648 17693 5649
rect 17635 5608 17644 5648
rect 17684 5608 17693 5648
rect 17635 5607 17693 5608
rect 18027 5648 18069 5657
rect 18027 5608 18028 5648
rect 18068 5608 18069 5648
rect 18027 5599 18069 5608
rect 18123 5648 18165 5657
rect 18123 5608 18124 5648
rect 18164 5608 18165 5648
rect 18123 5599 18165 5608
rect 18219 5648 18261 5657
rect 18219 5608 18220 5648
rect 18260 5608 18261 5648
rect 18219 5599 18261 5608
rect 18315 5648 18357 5657
rect 18315 5608 18316 5648
rect 18356 5608 18357 5648
rect 18315 5599 18357 5608
rect 18499 5648 18557 5649
rect 18499 5608 18508 5648
rect 18548 5608 18557 5648
rect 18499 5607 18557 5608
rect 19747 5648 19805 5649
rect 19747 5608 19756 5648
rect 19796 5608 19805 5648
rect 19747 5607 19805 5608
rect 20227 5648 20285 5649
rect 20227 5608 20236 5648
rect 20276 5608 20285 5648
rect 20227 5607 20285 5608
rect 9003 5564 9045 5573
rect 9003 5524 9004 5564
rect 9044 5524 9045 5564
rect 9003 5515 9045 5524
rect 13227 5564 13269 5573
rect 13227 5524 13228 5564
rect 13268 5524 13269 5564
rect 13227 5515 13269 5524
rect 15243 5564 15285 5573
rect 15243 5524 15244 5564
rect 15284 5524 15285 5564
rect 15243 5515 15285 5524
rect 15723 5564 15765 5573
rect 15723 5524 15724 5564
rect 15764 5524 15765 5564
rect 15723 5515 15765 5524
rect 19947 5564 19989 5573
rect 19947 5524 19948 5564
rect 19988 5524 19989 5564
rect 19947 5515 19989 5524
rect 3331 5480 3389 5481
rect 3331 5440 3340 5480
rect 3380 5440 3389 5480
rect 3331 5439 3389 5440
rect 5539 5480 5597 5481
rect 5539 5440 5548 5480
rect 5588 5440 5597 5480
rect 5539 5439 5597 5440
rect 8331 5480 8373 5489
rect 8331 5440 8332 5480
rect 8372 5440 8373 5480
rect 8331 5431 8373 5440
rect 11595 5480 11637 5489
rect 11595 5440 11596 5480
rect 11636 5440 11637 5480
rect 11595 5431 11637 5440
rect 17835 5480 17877 5489
rect 17835 5440 17836 5480
rect 17876 5440 17877 5480
rect 17835 5431 17877 5440
rect 1152 5312 20452 5336
rect 1152 5272 4928 5312
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 5296 5272 20048 5312
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20416 5272 20452 5312
rect 1152 5248 20452 5272
rect 4491 5144 4533 5153
rect 4491 5104 4492 5144
rect 4532 5104 4533 5144
rect 4491 5095 4533 5104
rect 15627 5144 15669 5153
rect 15627 5104 15628 5144
rect 15668 5104 15669 5144
rect 15627 5095 15669 5104
rect 4299 5060 4341 5069
rect 4299 5020 4300 5060
rect 4340 5020 4341 5060
rect 4299 5011 4341 5020
rect 6123 5060 6165 5069
rect 6123 5020 6124 5060
rect 6164 5020 6165 5060
rect 6123 5011 6165 5020
rect 11307 5060 11349 5069
rect 11307 5020 11308 5060
rect 11348 5020 11349 5060
rect 11307 5011 11349 5020
rect 11499 5060 11541 5069
rect 11499 5020 11500 5060
rect 11540 5020 11541 5060
rect 11499 5011 11541 5020
rect 13611 5060 13653 5069
rect 13611 5020 13612 5060
rect 13652 5020 13653 5060
rect 13611 5011 13653 5020
rect 17547 5060 17589 5069
rect 17547 5020 17548 5060
rect 17588 5020 17589 5060
rect 17547 5011 17589 5020
rect 2571 4976 2613 4985
rect 2571 4936 2572 4976
rect 2612 4936 2613 4976
rect 2571 4927 2613 4936
rect 2667 4976 2709 4985
rect 2667 4936 2668 4976
rect 2708 4936 2709 4976
rect 2667 4927 2709 4936
rect 3619 4976 3677 4977
rect 3619 4936 3628 4976
rect 3668 4936 3677 4976
rect 4675 4976 4733 4977
rect 3619 4935 3677 4936
rect 4107 4962 4149 4971
rect 4107 4922 4108 4962
rect 4148 4922 4149 4962
rect 4675 4936 4684 4976
rect 4724 4936 4733 4976
rect 4675 4935 4733 4936
rect 5923 4976 5981 4977
rect 5923 4936 5932 4976
rect 5972 4936 5981 4976
rect 5923 4935 5981 4936
rect 6307 4976 6365 4977
rect 6307 4936 6316 4976
rect 6356 4936 6365 4976
rect 6307 4935 6365 4936
rect 7555 4976 7613 4977
rect 7555 4936 7564 4976
rect 7604 4936 7613 4976
rect 7555 4935 7613 4936
rect 7939 4976 7997 4977
rect 7939 4936 7948 4976
rect 7988 4936 7997 4976
rect 7939 4935 7997 4936
rect 9187 4976 9245 4977
rect 9187 4936 9196 4976
rect 9236 4936 9245 4976
rect 9187 4935 9245 4936
rect 9579 4976 9621 4985
rect 9579 4936 9580 4976
rect 9620 4936 9621 4976
rect 9579 4927 9621 4936
rect 9675 4976 9717 4985
rect 9675 4936 9676 4976
rect 9716 4936 9717 4976
rect 9675 4927 9717 4936
rect 10155 4976 10197 4985
rect 10155 4936 10156 4976
rect 10196 4936 10197 4976
rect 10155 4927 10197 4936
rect 10627 4976 10685 4977
rect 10627 4936 10636 4976
rect 10676 4936 10685 4976
rect 10627 4935 10685 4936
rect 11115 4971 11157 4980
rect 11115 4931 11116 4971
rect 11156 4931 11157 4971
rect 11587 4976 11645 4977
rect 11587 4936 11596 4976
rect 11636 4936 11645 4976
rect 11587 4935 11645 4936
rect 11883 4976 11925 4985
rect 11883 4936 11884 4976
rect 11924 4936 11925 4976
rect 11115 4922 11157 4931
rect 11883 4927 11925 4936
rect 11979 4976 12021 4985
rect 11979 4936 11980 4976
rect 12020 4936 12021 4976
rect 11979 4927 12021 4936
rect 12363 4976 12405 4985
rect 12363 4936 12364 4976
rect 12404 4936 12405 4976
rect 12363 4927 12405 4936
rect 12931 4976 12989 4977
rect 12931 4936 12940 4976
rect 12980 4936 12989 4976
rect 13899 4976 13941 4985
rect 12931 4935 12989 4936
rect 13419 4962 13461 4971
rect 13419 4922 13420 4962
rect 13460 4922 13461 4962
rect 13899 4936 13900 4976
rect 13940 4936 13941 4976
rect 13899 4927 13941 4936
rect 13995 4976 14037 4985
rect 13995 4936 13996 4976
rect 14036 4936 14037 4976
rect 13995 4927 14037 4936
rect 14947 4976 15005 4977
rect 14947 4936 14956 4976
rect 14996 4936 15005 4976
rect 14947 4935 15005 4936
rect 15435 4971 15477 4980
rect 15435 4931 15436 4971
rect 15476 4931 15477 4971
rect 16099 4976 16157 4977
rect 16099 4936 16108 4976
rect 16148 4936 16157 4976
rect 16099 4935 16157 4936
rect 17347 4976 17405 4977
rect 17347 4936 17356 4976
rect 17396 4936 17405 4976
rect 17347 4935 17405 4936
rect 17739 4976 17781 4985
rect 17739 4936 17740 4976
rect 17780 4936 17781 4976
rect 15435 4922 15477 4931
rect 17739 4927 17781 4936
rect 18019 4976 18077 4977
rect 18019 4936 18028 4976
rect 18068 4936 18077 4976
rect 18019 4935 18077 4936
rect 18123 4976 18165 4985
rect 18123 4936 18124 4976
rect 18164 4936 18165 4976
rect 18123 4927 18165 4936
rect 18315 4976 18357 4985
rect 18315 4936 18316 4976
rect 18356 4936 18357 4976
rect 18315 4927 18357 4936
rect 18499 4976 18557 4977
rect 18499 4936 18508 4976
rect 18548 4936 18557 4976
rect 18499 4935 18557 4936
rect 19747 4976 19805 4977
rect 19747 4936 19756 4976
rect 19796 4936 19805 4976
rect 19747 4935 19805 4936
rect 4107 4913 4149 4922
rect 13419 4913 13461 4922
rect 1411 4892 1469 4893
rect 1411 4852 1420 4892
rect 1460 4852 1469 4892
rect 1411 4851 1469 4852
rect 1891 4892 1949 4893
rect 1891 4852 1900 4892
rect 1940 4852 1949 4892
rect 1891 4851 1949 4852
rect 2083 4892 2141 4893
rect 2083 4852 2092 4892
rect 2132 4852 2141 4892
rect 2083 4851 2141 4852
rect 3051 4892 3093 4901
rect 3051 4852 3052 4892
rect 3092 4852 3093 4892
rect 3051 4843 3093 4852
rect 3147 4892 3189 4901
rect 3147 4852 3148 4892
rect 3188 4852 3189 4892
rect 3147 4843 3189 4852
rect 10059 4892 10101 4901
rect 10059 4852 10060 4892
rect 10100 4852 10101 4892
rect 10059 4843 10101 4852
rect 12459 4892 12501 4901
rect 12459 4852 12460 4892
rect 12500 4852 12501 4892
rect 12459 4843 12501 4852
rect 14379 4892 14421 4901
rect 14379 4852 14380 4892
rect 14420 4852 14421 4892
rect 14379 4843 14421 4852
rect 14475 4892 14517 4901
rect 14475 4852 14476 4892
rect 14516 4852 14517 4892
rect 14475 4843 14517 4852
rect 1227 4808 1269 4817
rect 1227 4768 1228 4808
rect 1268 4768 1269 4808
rect 1227 4759 1269 4768
rect 1707 4808 1749 4817
rect 1707 4768 1708 4808
rect 1748 4768 1749 4808
rect 1707 4759 1749 4768
rect 15819 4808 15861 4817
rect 15819 4768 15820 4808
rect 15860 4768 15861 4808
rect 15819 4759 15861 4768
rect 18315 4808 18357 4817
rect 18315 4768 18316 4808
rect 18356 4768 18357 4808
rect 18315 4759 18357 4768
rect 2283 4724 2325 4733
rect 2283 4684 2284 4724
rect 2324 4684 2325 4724
rect 2283 4675 2325 4684
rect 7755 4724 7797 4733
rect 7755 4684 7756 4724
rect 7796 4684 7797 4724
rect 7755 4675 7797 4684
rect 19947 4724 19989 4733
rect 19947 4684 19948 4724
rect 19988 4684 19989 4724
rect 19947 4675 19989 4684
rect 1152 4556 20352 4580
rect 1152 4516 3688 4556
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 4056 4516 18808 4556
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 19176 4516 20352 4556
rect 1152 4492 20352 4516
rect 2763 4388 2805 4397
rect 2763 4348 2764 4388
rect 2804 4348 2805 4388
rect 2763 4339 2805 4348
rect 4395 4388 4437 4397
rect 4395 4348 4396 4388
rect 4436 4348 4437 4388
rect 4395 4339 4437 4348
rect 10251 4388 10293 4397
rect 10251 4348 10252 4388
rect 10292 4348 10293 4388
rect 10251 4339 10293 4348
rect 13323 4388 13365 4397
rect 13323 4348 13324 4388
rect 13364 4348 13365 4388
rect 13323 4339 13365 4348
rect 15531 4388 15573 4397
rect 15531 4348 15532 4388
rect 15572 4348 15573 4388
rect 15531 4339 15573 4348
rect 17835 4388 17877 4397
rect 17835 4348 17836 4388
rect 17876 4348 17877 4388
rect 17835 4339 17877 4348
rect 11115 4304 11157 4313
rect 11115 4264 11116 4304
rect 11156 4264 11157 4304
rect 11115 4255 11157 4264
rect 7275 4220 7317 4229
rect 7275 4180 7276 4220
rect 7316 4180 7317 4220
rect 7275 4171 7317 4180
rect 7371 4220 7413 4229
rect 7371 4180 7372 4220
rect 7412 4180 7413 4220
rect 7371 4171 7413 4180
rect 11883 4220 11925 4229
rect 11883 4180 11884 4220
rect 11924 4180 11925 4220
rect 11883 4171 11925 4180
rect 13507 4220 13565 4221
rect 13507 4180 13516 4220
rect 13556 4180 13565 4220
rect 13507 4179 13565 4180
rect 13891 4220 13949 4221
rect 13891 4180 13900 4220
rect 13940 4180 13949 4220
rect 13891 4179 13949 4180
rect 8379 4145 8421 4154
rect 12987 4145 13029 4154
rect 1315 4136 1373 4137
rect 1315 4096 1324 4136
rect 1364 4096 1373 4136
rect 1315 4095 1373 4096
rect 2563 4136 2621 4137
rect 2563 4096 2572 4136
rect 2612 4096 2621 4136
rect 2563 4095 2621 4096
rect 2947 4136 3005 4137
rect 2947 4096 2956 4136
rect 2996 4096 3005 4136
rect 2947 4095 3005 4096
rect 4195 4136 4253 4137
rect 4195 4096 4204 4136
rect 4244 4096 4253 4136
rect 4195 4095 4253 4096
rect 4579 4136 4637 4137
rect 4579 4096 4588 4136
rect 4628 4096 4637 4136
rect 4579 4095 4637 4096
rect 5827 4136 5885 4137
rect 5827 4096 5836 4136
rect 5876 4096 5885 4136
rect 5827 4095 5885 4096
rect 6219 4136 6261 4145
rect 6219 4096 6220 4136
rect 6260 4096 6261 4136
rect 6219 4087 6261 4096
rect 6315 4136 6357 4145
rect 6315 4096 6316 4136
rect 6356 4096 6357 4136
rect 6315 4087 6357 4096
rect 6411 4136 6453 4145
rect 6411 4096 6412 4136
rect 6452 4096 6453 4136
rect 6411 4087 6453 4096
rect 6507 4136 6549 4145
rect 6507 4096 6508 4136
rect 6548 4096 6549 4136
rect 6507 4087 6549 4096
rect 6795 4136 6837 4145
rect 6795 4096 6796 4136
rect 6836 4096 6837 4136
rect 6795 4087 6837 4096
rect 6891 4136 6933 4145
rect 6891 4096 6892 4136
rect 6932 4096 6933 4136
rect 6891 4087 6933 4096
rect 7843 4136 7901 4137
rect 7843 4096 7852 4136
rect 7892 4096 7901 4136
rect 8379 4105 8380 4145
rect 8420 4105 8421 4145
rect 8379 4096 8421 4105
rect 8803 4136 8861 4137
rect 8803 4096 8812 4136
rect 8852 4096 8861 4136
rect 7843 4095 7901 4096
rect 8803 4095 8861 4096
rect 10051 4136 10109 4137
rect 10051 4096 10060 4136
rect 10100 4096 10109 4136
rect 10051 4095 10109 4096
rect 10443 4136 10485 4145
rect 10443 4096 10444 4136
rect 10484 4096 10485 4136
rect 10443 4087 10485 4096
rect 10539 4136 10581 4145
rect 10539 4096 10540 4136
rect 10580 4096 10581 4136
rect 10539 4087 10581 4096
rect 10635 4136 10677 4145
rect 10635 4096 10636 4136
rect 10676 4096 10677 4136
rect 10635 4087 10677 4096
rect 10731 4136 10773 4145
rect 10731 4096 10732 4136
rect 10772 4096 10773 4136
rect 10731 4087 10773 4096
rect 10923 4136 10965 4145
rect 10923 4096 10924 4136
rect 10964 4096 10965 4136
rect 10923 4087 10965 4096
rect 11115 4136 11157 4145
rect 11115 4096 11116 4136
rect 11156 4096 11157 4136
rect 11115 4087 11157 4096
rect 11403 4136 11445 4145
rect 11403 4096 11404 4136
rect 11444 4096 11445 4136
rect 11403 4087 11445 4096
rect 11499 4136 11541 4145
rect 11499 4096 11500 4136
rect 11540 4096 11541 4136
rect 11499 4087 11541 4096
rect 11979 4136 12021 4145
rect 11979 4096 11980 4136
rect 12020 4096 12021 4136
rect 11979 4087 12021 4096
rect 12451 4136 12509 4137
rect 12451 4096 12460 4136
rect 12500 4096 12509 4136
rect 12987 4105 12988 4145
rect 13028 4105 13029 4145
rect 12987 4096 13029 4105
rect 14083 4136 14141 4137
rect 14083 4096 14092 4136
rect 14132 4096 14141 4136
rect 12451 4095 12509 4096
rect 14083 4095 14141 4096
rect 15331 4136 15389 4137
rect 15331 4096 15340 4136
rect 15380 4096 15389 4136
rect 15331 4095 15389 4096
rect 15915 4136 15957 4145
rect 15915 4096 15916 4136
rect 15956 4096 15957 4136
rect 15915 4087 15957 4096
rect 16011 4136 16053 4145
rect 16011 4096 16012 4136
rect 16052 4096 16053 4136
rect 16011 4087 16053 4096
rect 16387 4136 16445 4137
rect 16387 4096 16396 4136
rect 16436 4096 16445 4136
rect 16387 4095 16445 4096
rect 17635 4136 17693 4137
rect 17635 4096 17644 4136
rect 17684 4096 17693 4136
rect 17635 4095 17693 4096
rect 18019 4136 18077 4137
rect 18019 4096 18028 4136
rect 18068 4096 18077 4136
rect 18019 4095 18077 4096
rect 18123 4136 18165 4145
rect 18123 4096 18124 4136
rect 18164 4096 18165 4136
rect 18123 4087 18165 4096
rect 18315 4136 18357 4145
rect 18315 4096 18316 4136
rect 18356 4096 18357 4136
rect 18315 4087 18357 4096
rect 18499 4136 18557 4137
rect 18499 4096 18508 4136
rect 18548 4096 18557 4136
rect 18499 4095 18557 4096
rect 19747 4136 19805 4137
rect 19747 4096 19756 4136
rect 19796 4096 19805 4136
rect 19747 4095 19805 4096
rect 8523 4052 8565 4061
rect 8523 4012 8524 4052
rect 8564 4012 8565 4052
rect 8523 4003 8565 4012
rect 18219 4052 18261 4061
rect 18219 4012 18220 4052
rect 18260 4012 18261 4052
rect 18219 4003 18261 4012
rect 6027 3968 6069 3977
rect 6027 3928 6028 3968
rect 6068 3928 6069 3968
rect 6027 3919 6069 3928
rect 13131 3968 13173 3977
rect 13131 3928 13132 3968
rect 13172 3928 13173 3968
rect 13131 3919 13173 3928
rect 13707 3968 13749 3977
rect 13707 3928 13708 3968
rect 13748 3928 13749 3968
rect 13707 3919 13749 3928
rect 16195 3968 16253 3969
rect 16195 3928 16204 3968
rect 16244 3928 16253 3968
rect 16195 3927 16253 3928
rect 17835 3968 17877 3977
rect 17835 3928 17836 3968
rect 17876 3928 17877 3968
rect 17835 3919 17877 3928
rect 19947 3968 19989 3977
rect 19947 3928 19948 3968
rect 19988 3928 19989 3968
rect 19947 3919 19989 3928
rect 1152 3800 20452 3824
rect 1152 3760 4928 3800
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 5296 3760 20048 3800
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20416 3760 20452 3800
rect 1152 3736 20452 3760
rect 1323 3632 1365 3641
rect 1323 3592 1324 3632
rect 1364 3592 1365 3632
rect 1323 3583 1365 3592
rect 1995 3632 2037 3641
rect 1995 3592 1996 3632
rect 2036 3592 2037 3632
rect 1995 3583 2037 3592
rect 4299 3632 4341 3641
rect 4299 3592 4300 3632
rect 4340 3592 4341 3632
rect 4299 3583 4341 3592
rect 6403 3632 6461 3633
rect 6403 3592 6412 3632
rect 6452 3592 6461 3632
rect 6403 3591 6461 3592
rect 8619 3632 8661 3641
rect 8619 3592 8620 3632
rect 8660 3592 8661 3632
rect 8619 3583 8661 3592
rect 8811 3632 8853 3641
rect 8811 3592 8812 3632
rect 8852 3592 8853 3632
rect 8811 3583 8853 3592
rect 10443 3632 10485 3641
rect 10443 3592 10444 3632
rect 10484 3592 10485 3632
rect 10443 3583 10485 3592
rect 11203 3632 11261 3633
rect 11203 3592 11212 3632
rect 11252 3592 11261 3632
rect 11203 3591 11261 3592
rect 13227 3632 13269 3641
rect 13227 3592 13228 3632
rect 13268 3592 13269 3632
rect 13227 3583 13269 3592
rect 16971 3632 17013 3641
rect 16971 3592 16972 3632
rect 17012 3592 17013 3632
rect 16971 3583 17013 3592
rect 17355 3632 17397 3641
rect 17355 3592 17356 3632
rect 17396 3592 17397 3632
rect 17355 3583 17397 3592
rect 19939 3632 19997 3633
rect 19939 3592 19948 3632
rect 19988 3592 19997 3632
rect 19939 3591 19997 3592
rect 4011 3548 4053 3557
rect 4011 3508 4012 3548
rect 4052 3508 4053 3548
rect 4011 3499 4053 3508
rect 4587 3548 4629 3557
rect 4587 3508 4588 3548
rect 4628 3508 4629 3548
rect 4587 3499 4629 3508
rect 13899 3548 13941 3557
rect 13899 3508 13900 3548
rect 13940 3508 13941 3548
rect 13899 3499 13941 3508
rect 19467 3548 19509 3557
rect 19467 3508 19468 3548
rect 19508 3508 19509 3548
rect 19467 3499 19509 3508
rect 2187 3459 2229 3468
rect 2187 3419 2188 3459
rect 2228 3419 2229 3459
rect 2659 3464 2717 3465
rect 2659 3424 2668 3464
rect 2708 3424 2717 3464
rect 2659 3423 2717 3424
rect 3243 3464 3285 3473
rect 3243 3424 3244 3464
rect 3284 3424 3285 3464
rect 2187 3410 2229 3419
rect 3243 3415 3285 3424
rect 3627 3464 3669 3473
rect 3627 3424 3628 3464
rect 3668 3424 3669 3464
rect 3627 3415 3669 3424
rect 3723 3464 3765 3473
rect 3723 3424 3724 3464
rect 3764 3424 3765 3464
rect 3723 3415 3765 3424
rect 4387 3464 4445 3465
rect 4387 3424 4396 3464
rect 4436 3424 4445 3464
rect 4387 3423 4445 3424
rect 4771 3464 4829 3465
rect 4771 3424 4780 3464
rect 4820 3424 4829 3464
rect 4771 3423 4829 3424
rect 6019 3464 6077 3465
rect 6019 3424 6028 3464
rect 6068 3424 6077 3464
rect 6019 3423 6077 3424
rect 6315 3464 6357 3473
rect 6315 3424 6316 3464
rect 6356 3424 6357 3464
rect 6315 3415 6357 3424
rect 6507 3464 6549 3473
rect 6507 3424 6508 3464
rect 6548 3424 6549 3464
rect 6507 3415 6549 3424
rect 6595 3464 6653 3465
rect 6595 3424 6604 3464
rect 6644 3424 6653 3464
rect 6595 3423 6653 3424
rect 6891 3464 6933 3473
rect 6891 3424 6892 3464
rect 6932 3424 6933 3464
rect 6891 3415 6933 3424
rect 6987 3464 7029 3473
rect 6987 3424 6988 3464
rect 7028 3424 7029 3464
rect 6987 3415 7029 3424
rect 7467 3464 7509 3473
rect 7467 3424 7468 3464
rect 7508 3424 7509 3464
rect 7467 3415 7509 3424
rect 7939 3464 7997 3465
rect 7939 3424 7948 3464
rect 7988 3424 7997 3464
rect 8995 3464 9053 3465
rect 7939 3423 7997 3424
rect 8427 3450 8469 3459
rect 8427 3410 8428 3450
rect 8468 3410 8469 3450
rect 8995 3424 9004 3464
rect 9044 3424 9053 3464
rect 8995 3423 9053 3424
rect 10243 3464 10301 3465
rect 10243 3424 10252 3464
rect 10292 3424 10301 3464
rect 10243 3423 10301 3424
rect 11011 3464 11069 3465
rect 11011 3424 11020 3464
rect 11060 3424 11069 3464
rect 11011 3423 11069 3424
rect 11107 3464 11165 3465
rect 11107 3424 11116 3464
rect 11156 3424 11165 3464
rect 11107 3423 11165 3424
rect 11307 3464 11349 3473
rect 11307 3424 11308 3464
rect 11348 3424 11349 3464
rect 11307 3415 11349 3424
rect 11403 3464 11445 3473
rect 11403 3424 11404 3464
rect 11444 3424 11445 3464
rect 11403 3415 11445 3424
rect 11496 3464 11554 3465
rect 11496 3424 11505 3464
rect 11545 3424 11554 3464
rect 11496 3423 11554 3424
rect 11779 3464 11837 3465
rect 11779 3424 11788 3464
rect 11828 3424 11837 3464
rect 11779 3423 11837 3424
rect 13027 3464 13085 3465
rect 13027 3424 13036 3464
rect 13076 3424 13085 3464
rect 13027 3423 13085 3424
rect 13507 3464 13565 3465
rect 13507 3424 13516 3464
rect 13556 3424 13565 3464
rect 13507 3423 13565 3424
rect 13803 3464 13845 3473
rect 13803 3424 13804 3464
rect 13844 3424 13845 3464
rect 13803 3415 13845 3424
rect 15243 3464 15285 3473
rect 15243 3424 15244 3464
rect 15284 3424 15285 3464
rect 15243 3415 15285 3424
rect 15339 3464 15381 3473
rect 15339 3424 15340 3464
rect 15380 3424 15381 3464
rect 15339 3415 15381 3424
rect 15723 3464 15765 3473
rect 15723 3424 15724 3464
rect 15764 3424 15765 3464
rect 15723 3415 15765 3424
rect 15819 3464 15861 3473
rect 15819 3424 15820 3464
rect 15860 3424 15861 3464
rect 15819 3415 15861 3424
rect 16291 3464 16349 3465
rect 16291 3424 16300 3464
rect 16340 3424 16349 3464
rect 17163 3464 17205 3473
rect 16291 3423 16349 3424
rect 16779 3450 16821 3459
rect 8427 3401 8469 3410
rect 16779 3410 16780 3450
rect 16820 3410 16821 3450
rect 17163 3424 17164 3464
rect 17204 3424 17205 3464
rect 17163 3415 17205 3424
rect 17451 3464 17493 3473
rect 17451 3424 17452 3464
rect 17492 3424 17493 3464
rect 17451 3415 17493 3424
rect 17739 3464 17781 3473
rect 17739 3424 17740 3464
rect 17780 3424 17781 3464
rect 17739 3415 17781 3424
rect 17835 3464 17877 3473
rect 17835 3424 17836 3464
rect 17876 3424 17877 3464
rect 17835 3415 17877 3424
rect 18219 3464 18261 3473
rect 18219 3424 18220 3464
rect 18260 3424 18261 3464
rect 18219 3415 18261 3424
rect 18315 3464 18357 3473
rect 18315 3424 18316 3464
rect 18356 3424 18357 3464
rect 18315 3415 18357 3424
rect 18787 3464 18845 3465
rect 18787 3424 18796 3464
rect 18836 3424 18845 3464
rect 19659 3464 19701 3473
rect 18787 3423 18845 3424
rect 19323 3454 19365 3463
rect 16779 3401 16821 3410
rect 19323 3414 19324 3454
rect 19364 3414 19365 3454
rect 19659 3424 19660 3464
rect 19700 3424 19701 3464
rect 19659 3415 19701 3424
rect 19755 3464 19797 3473
rect 19755 3424 19756 3464
rect 19796 3424 19797 3464
rect 19755 3415 19797 3424
rect 19851 3464 19893 3473
rect 19851 3424 19852 3464
rect 19892 3424 19893 3464
rect 19851 3415 19893 3424
rect 19323 3405 19365 3414
rect 1507 3380 1565 3381
rect 1507 3340 1516 3380
rect 1556 3340 1565 3380
rect 1507 3339 1565 3340
rect 3147 3380 3189 3389
rect 3147 3340 3148 3380
rect 3188 3340 3189 3380
rect 3147 3331 3189 3340
rect 7371 3380 7413 3389
rect 7371 3340 7372 3380
rect 7412 3340 7413 3380
rect 7371 3331 7413 3340
rect 10627 3380 10685 3381
rect 10627 3340 10636 3380
rect 10676 3340 10685 3380
rect 10627 3339 10685 3340
rect 14371 3380 14429 3381
rect 14371 3340 14380 3380
rect 14420 3340 14429 3380
rect 14371 3339 14429 3340
rect 14947 3380 15005 3381
rect 14947 3340 14956 3380
rect 14996 3340 15005 3380
rect 14947 3339 15005 3340
rect 20139 3380 20181 3389
rect 20139 3340 20140 3380
rect 20180 3340 20181 3380
rect 20139 3331 20181 3340
rect 1803 3296 1845 3305
rect 1803 3256 1804 3296
rect 1844 3256 1845 3296
rect 1803 3247 1845 3256
rect 14179 3296 14237 3297
rect 14179 3256 14188 3296
rect 14228 3256 14237 3296
rect 14179 3255 14237 3256
rect 14571 3212 14613 3221
rect 14571 3172 14572 3212
rect 14612 3172 14613 3212
rect 14571 3163 14613 3172
rect 14763 3212 14805 3221
rect 14763 3172 14764 3212
rect 14804 3172 14805 3212
rect 14763 3163 14805 3172
rect 1152 3044 20352 3068
rect 1152 3004 3688 3044
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 4056 3004 18808 3044
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 19176 3004 20352 3044
rect 1152 2980 20352 3004
rect 2859 2876 2901 2885
rect 2859 2836 2860 2876
rect 2900 2836 2901 2876
rect 2859 2827 2901 2836
rect 9195 2876 9237 2885
rect 9195 2836 9196 2876
rect 9236 2836 9237 2876
rect 9195 2827 9237 2836
rect 9963 2876 10005 2885
rect 9963 2836 9964 2876
rect 10004 2836 10005 2876
rect 9963 2827 10005 2836
rect 14187 2876 14229 2885
rect 14187 2836 14188 2876
rect 14228 2836 14229 2876
rect 14187 2827 14229 2836
rect 14379 2876 14421 2885
rect 14379 2836 14380 2876
rect 14420 2836 14421 2876
rect 14379 2827 14421 2836
rect 3819 2792 3861 2801
rect 3819 2752 3820 2792
rect 3860 2752 3861 2792
rect 3819 2743 3861 2752
rect 4395 2792 4437 2801
rect 4395 2752 4396 2792
rect 4436 2752 4437 2792
rect 4395 2743 4437 2752
rect 9667 2792 9725 2793
rect 9667 2752 9676 2792
rect 9716 2752 9725 2792
rect 9667 2751 9725 2752
rect 17643 2792 17685 2801
rect 17643 2752 17644 2792
rect 17684 2752 17685 2792
rect 17643 2743 17685 2752
rect 3147 2708 3189 2717
rect 3147 2668 3148 2708
rect 3188 2668 3189 2708
rect 3147 2659 3189 2668
rect 3619 2708 3677 2709
rect 3619 2668 3628 2708
rect 3668 2668 3677 2708
rect 3619 2667 3677 2668
rect 4195 2708 4253 2709
rect 4195 2668 4204 2708
rect 4244 2668 4253 2708
rect 4195 2667 4253 2668
rect 5643 2708 5685 2717
rect 5643 2668 5644 2708
rect 5684 2668 5685 2708
rect 5643 2659 5685 2668
rect 6979 2708 7037 2709
rect 6979 2668 6988 2708
rect 7028 2668 7037 2708
rect 6979 2667 7037 2668
rect 7363 2708 7421 2709
rect 7363 2668 7372 2708
rect 7412 2668 7421 2708
rect 7363 2667 7421 2668
rect 10147 2708 10205 2709
rect 10147 2668 10156 2708
rect 10196 2668 10205 2708
rect 10147 2667 10205 2668
rect 10531 2708 10589 2709
rect 10531 2668 10540 2708
rect 10580 2668 10589 2708
rect 10531 2667 10589 2668
rect 11403 2708 11445 2717
rect 11403 2668 11404 2708
rect 11444 2668 11445 2708
rect 11403 2659 11445 2668
rect 14563 2708 14621 2709
rect 14563 2668 14572 2708
rect 14612 2668 14621 2708
rect 14563 2667 14621 2668
rect 15435 2708 15477 2717
rect 15435 2668 15436 2708
rect 15476 2668 15477 2708
rect 15435 2659 15477 2668
rect 15531 2708 15573 2717
rect 15531 2668 15532 2708
rect 15572 2668 15573 2708
rect 17059 2708 17117 2709
rect 15531 2659 15573 2668
rect 16539 2666 16581 2675
rect 17059 2668 17068 2708
rect 17108 2668 17117 2708
rect 17059 2667 17117 2668
rect 17443 2708 17501 2709
rect 17443 2668 17452 2708
rect 17492 2668 17501 2708
rect 17443 2667 17501 2668
rect 18507 2708 18549 2717
rect 18507 2668 18508 2708
rect 18548 2668 18549 2708
rect 15051 2643 15093 2652
rect 1411 2624 1469 2625
rect 1411 2584 1420 2624
rect 1460 2584 1469 2624
rect 1411 2583 1469 2584
rect 2659 2624 2717 2625
rect 2659 2584 2668 2624
rect 2708 2584 2717 2624
rect 2659 2583 2717 2584
rect 3051 2624 3093 2633
rect 3051 2584 3052 2624
rect 3092 2584 3093 2624
rect 3051 2575 3093 2584
rect 3243 2624 3285 2633
rect 3243 2584 3244 2624
rect 3284 2584 3285 2624
rect 3243 2575 3285 2584
rect 4683 2624 4725 2633
rect 4683 2584 4684 2624
rect 4724 2584 4725 2624
rect 4683 2575 4725 2584
rect 5067 2624 5109 2633
rect 5067 2584 5068 2624
rect 5108 2584 5109 2624
rect 5067 2575 5109 2584
rect 5163 2624 5205 2633
rect 5163 2584 5164 2624
rect 5204 2584 5205 2624
rect 5163 2575 5205 2584
rect 5547 2624 5589 2633
rect 6603 2629 6645 2638
rect 5547 2584 5548 2624
rect 5588 2584 5589 2624
rect 5547 2575 5589 2584
rect 6115 2624 6173 2625
rect 6115 2584 6124 2624
rect 6164 2584 6173 2624
rect 6115 2583 6173 2584
rect 6603 2589 6604 2629
rect 6644 2589 6645 2629
rect 6603 2580 6645 2589
rect 7747 2624 7805 2625
rect 7747 2584 7756 2624
rect 7796 2584 7805 2624
rect 7747 2583 7805 2584
rect 8995 2624 9053 2625
rect 8995 2584 9004 2624
rect 9044 2584 9053 2624
rect 8995 2583 9053 2584
rect 9387 2624 9429 2633
rect 9387 2584 9388 2624
rect 9428 2584 9429 2624
rect 9387 2575 9429 2584
rect 9579 2624 9621 2633
rect 9579 2584 9580 2624
rect 9620 2584 9621 2624
rect 9579 2575 9621 2584
rect 9675 2624 9717 2633
rect 9675 2584 9676 2624
rect 9716 2584 9717 2624
rect 9675 2575 9717 2584
rect 10827 2624 10869 2633
rect 10827 2584 10828 2624
rect 10868 2584 10869 2624
rect 10827 2575 10869 2584
rect 10923 2624 10965 2633
rect 10923 2584 10924 2624
rect 10964 2584 10965 2624
rect 10923 2575 10965 2584
rect 11307 2624 11349 2633
rect 12363 2629 12405 2638
rect 11307 2584 11308 2624
rect 11348 2584 11349 2624
rect 11307 2575 11349 2584
rect 11875 2624 11933 2625
rect 11875 2584 11884 2624
rect 11924 2584 11933 2624
rect 11875 2583 11933 2584
rect 12363 2589 12364 2629
rect 12404 2589 12405 2629
rect 12363 2580 12405 2589
rect 12739 2624 12797 2625
rect 12739 2584 12748 2624
rect 12788 2584 12797 2624
rect 12739 2583 12797 2584
rect 13987 2624 14045 2625
rect 13987 2584 13996 2624
rect 14036 2584 14045 2624
rect 13987 2583 14045 2584
rect 14955 2604 14997 2613
rect 14955 2564 14956 2604
rect 14996 2564 14997 2604
rect 15051 2603 15052 2643
rect 15092 2603 15093 2643
rect 16539 2626 16540 2666
rect 16580 2626 16581 2666
rect 18507 2659 18549 2668
rect 19563 2638 19605 2647
rect 15051 2594 15093 2603
rect 16003 2624 16061 2625
rect 16003 2584 16012 2624
rect 16052 2584 16061 2624
rect 16539 2617 16581 2626
rect 18027 2624 18069 2633
rect 16003 2583 16061 2584
rect 18027 2584 18028 2624
rect 18068 2584 18069 2624
rect 18027 2575 18069 2584
rect 18123 2624 18165 2633
rect 18123 2584 18124 2624
rect 18164 2584 18165 2624
rect 18123 2575 18165 2584
rect 18603 2624 18645 2633
rect 18603 2584 18604 2624
rect 18644 2584 18645 2624
rect 18603 2575 18645 2584
rect 19075 2624 19133 2625
rect 19075 2584 19084 2624
rect 19124 2584 19133 2624
rect 19563 2598 19564 2638
rect 19604 2598 19605 2638
rect 19563 2589 19605 2598
rect 19947 2624 19989 2633
rect 19075 2583 19133 2584
rect 19947 2584 19948 2624
rect 19988 2584 19989 2624
rect 19947 2575 19989 2584
rect 20043 2624 20085 2633
rect 20043 2584 20044 2624
rect 20084 2584 20085 2624
rect 20043 2575 20085 2584
rect 20139 2624 20181 2633
rect 20139 2584 20140 2624
rect 20180 2584 20181 2624
rect 20139 2575 20181 2584
rect 20235 2624 20277 2633
rect 20235 2584 20236 2624
rect 20276 2584 20277 2624
rect 20235 2575 20277 2584
rect 14955 2555 14997 2564
rect 6795 2540 6837 2549
rect 6795 2500 6796 2540
rect 6836 2500 6837 2540
rect 6795 2491 6837 2500
rect 12555 2540 12597 2549
rect 12555 2500 12556 2540
rect 12596 2500 12597 2540
rect 12555 2491 12597 2500
rect 16683 2540 16725 2549
rect 16683 2500 16684 2540
rect 16724 2500 16725 2540
rect 16683 2491 16725 2500
rect 4011 2456 4053 2465
rect 4011 2416 4012 2456
rect 4052 2416 4053 2456
rect 4011 2407 4053 2416
rect 7179 2456 7221 2465
rect 7179 2416 7180 2456
rect 7220 2416 7221 2456
rect 7179 2407 7221 2416
rect 7563 2456 7605 2465
rect 7563 2416 7564 2456
rect 7604 2416 7605 2456
rect 7563 2407 7605 2416
rect 10347 2456 10389 2465
rect 10347 2416 10348 2456
rect 10388 2416 10389 2456
rect 10347 2407 10389 2416
rect 16875 2456 16917 2465
rect 16875 2416 16876 2456
rect 16916 2416 16917 2456
rect 16875 2407 16917 2416
rect 17259 2456 17301 2465
rect 17259 2416 17260 2456
rect 17300 2416 17301 2456
rect 17259 2407 17301 2416
rect 19755 2456 19797 2465
rect 19755 2416 19756 2456
rect 19796 2416 19797 2456
rect 19755 2407 19797 2416
rect 1152 2288 20452 2312
rect 1152 2248 4928 2288
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 5296 2248 20048 2288
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20416 2248 20452 2288
rect 1152 2224 20452 2248
rect 4291 2120 4349 2121
rect 4291 2080 4300 2120
rect 4340 2080 4349 2120
rect 4291 2079 4349 2080
rect 5443 2120 5501 2121
rect 5443 2080 5452 2120
rect 5492 2080 5501 2120
rect 5443 2079 5501 2080
rect 9003 2120 9045 2129
rect 9003 2080 9004 2120
rect 9044 2080 9045 2120
rect 9003 2071 9045 2080
rect 9291 2120 9333 2129
rect 9291 2080 9292 2120
rect 9332 2080 9333 2120
rect 9291 2071 9333 2080
rect 11691 2120 11733 2129
rect 11691 2080 11692 2120
rect 11732 2080 11733 2120
rect 11691 2071 11733 2080
rect 11979 2120 12021 2129
rect 11979 2080 11980 2120
rect 12020 2080 12021 2120
rect 11979 2071 12021 2080
rect 15243 2120 15285 2129
rect 15243 2080 15244 2120
rect 15284 2080 15285 2120
rect 15243 2071 15285 2080
rect 15427 2120 15485 2121
rect 15427 2080 15436 2120
rect 15476 2080 15485 2120
rect 15427 2079 15485 2080
rect 17163 2120 17205 2129
rect 17163 2080 17164 2120
rect 17204 2080 17205 2120
rect 17163 2071 17205 2080
rect 19659 2120 19701 2129
rect 19659 2080 19660 2120
rect 19700 2080 19701 2120
rect 19659 2071 19701 2080
rect 3819 2036 3861 2045
rect 3819 1996 3820 2036
rect 3860 1996 3861 2036
rect 3819 1987 3861 1996
rect 2371 1952 2429 1953
rect 2371 1912 2380 1952
rect 2420 1912 2429 1952
rect 2371 1911 2429 1912
rect 3619 1952 3677 1953
rect 3619 1912 3628 1952
rect 3668 1912 3677 1952
rect 3619 1911 3677 1912
rect 4011 1952 4053 1961
rect 4011 1912 4012 1952
rect 4052 1912 4053 1952
rect 4011 1903 4053 1912
rect 4107 1952 4149 1961
rect 4107 1912 4108 1952
rect 4148 1912 4149 1952
rect 4107 1903 4149 1912
rect 5547 1952 5589 1961
rect 5547 1912 5548 1952
rect 5588 1912 5589 1952
rect 5547 1903 5589 1912
rect 5643 1952 5685 1961
rect 5643 1912 5644 1952
rect 5684 1912 5685 1952
rect 5643 1903 5685 1912
rect 5739 1952 5781 1961
rect 5739 1912 5740 1952
rect 5780 1912 5781 1952
rect 5739 1903 5781 1912
rect 5923 1952 5981 1953
rect 5923 1912 5932 1952
rect 5972 1912 5981 1952
rect 5923 1911 5981 1912
rect 7171 1952 7229 1953
rect 7171 1912 7180 1952
rect 7220 1912 7229 1952
rect 7171 1911 7229 1912
rect 7555 1952 7613 1953
rect 7555 1912 7564 1952
rect 7604 1912 7613 1952
rect 7555 1911 7613 1912
rect 8803 1952 8861 1953
rect 8803 1912 8812 1952
rect 8852 1912 8861 1952
rect 8803 1911 8861 1912
rect 9963 1952 10005 1961
rect 9963 1912 9964 1952
rect 10004 1912 10005 1952
rect 9963 1903 10005 1912
rect 10059 1952 10101 1961
rect 10059 1912 10060 1952
rect 10100 1912 10101 1952
rect 10059 1903 10101 1912
rect 10539 1952 10581 1961
rect 10539 1912 10540 1952
rect 10580 1912 10581 1952
rect 10539 1903 10581 1912
rect 11011 1952 11069 1953
rect 11011 1912 11020 1952
rect 11060 1912 11069 1952
rect 12163 1952 12221 1953
rect 11011 1911 11069 1912
rect 11499 1938 11541 1947
rect 11499 1898 11500 1938
rect 11540 1898 11541 1938
rect 12163 1912 12172 1952
rect 12212 1912 12221 1952
rect 12163 1911 12221 1912
rect 13411 1952 13469 1953
rect 13411 1912 13420 1952
rect 13460 1912 13469 1952
rect 13411 1911 13469 1912
rect 13795 1952 13853 1953
rect 13795 1912 13804 1952
rect 13844 1912 13853 1952
rect 13795 1911 13853 1912
rect 15043 1952 15101 1953
rect 15043 1912 15052 1952
rect 15092 1912 15101 1952
rect 15043 1911 15101 1912
rect 15715 1952 15773 1953
rect 15715 1912 15724 1952
rect 15764 1912 15773 1952
rect 15715 1911 15773 1912
rect 16963 1952 17021 1953
rect 16963 1912 16972 1952
rect 17012 1912 17021 1952
rect 16963 1911 17021 1912
rect 17923 1952 17981 1953
rect 17923 1912 17932 1952
rect 17972 1912 17981 1952
rect 17923 1911 17981 1912
rect 19171 1952 19229 1953
rect 19171 1912 19180 1952
rect 19220 1912 19229 1952
rect 19171 1911 19229 1912
rect 19563 1952 19605 1961
rect 19563 1912 19564 1952
rect 19604 1912 19605 1952
rect 19563 1903 19605 1912
rect 19755 1952 19797 1961
rect 19755 1912 19756 1952
rect 19796 1912 19797 1952
rect 19755 1903 19797 1912
rect 19939 1952 19997 1953
rect 19939 1912 19948 1952
rect 19988 1912 19997 1952
rect 19939 1911 19997 1912
rect 20043 1952 20085 1961
rect 20043 1912 20044 1952
rect 20084 1912 20085 1952
rect 20043 1903 20085 1912
rect 20235 1952 20277 1961
rect 20235 1912 20236 1952
rect 20276 1912 20277 1952
rect 20235 1903 20277 1912
rect 11499 1889 11541 1898
rect 1219 1868 1277 1869
rect 1219 1828 1228 1868
rect 1268 1828 1277 1868
rect 1219 1827 1277 1828
rect 1603 1868 1661 1869
rect 1603 1828 1612 1868
rect 1652 1828 1661 1868
rect 1603 1827 1661 1828
rect 1987 1868 2045 1869
rect 1987 1828 1996 1868
rect 2036 1828 2045 1868
rect 1987 1827 2045 1828
rect 4675 1868 4733 1869
rect 4675 1828 4684 1868
rect 4724 1828 4733 1868
rect 4675 1827 4733 1828
rect 5059 1868 5117 1869
rect 5059 1828 5068 1868
rect 5108 1828 5117 1868
rect 5059 1827 5117 1828
rect 9475 1868 9533 1869
rect 9475 1828 9484 1868
rect 9524 1828 9533 1868
rect 9475 1827 9533 1828
rect 10443 1868 10485 1877
rect 10443 1828 10444 1868
rect 10484 1828 10485 1868
rect 10443 1819 10485 1828
rect 17539 1868 17597 1869
rect 17539 1828 17548 1868
rect 17588 1828 17597 1868
rect 17539 1827 17597 1828
rect 4875 1784 4917 1793
rect 4875 1744 4876 1784
rect 4916 1744 4917 1784
rect 4875 1735 4917 1744
rect 7371 1784 7413 1793
rect 7371 1744 7372 1784
rect 7412 1744 7413 1784
rect 7371 1735 7413 1744
rect 20235 1784 20277 1793
rect 20235 1744 20236 1784
rect 20276 1744 20277 1784
rect 20235 1735 20277 1744
rect 1419 1700 1461 1709
rect 1419 1660 1420 1700
rect 1460 1660 1461 1700
rect 1419 1651 1461 1660
rect 1803 1700 1845 1709
rect 1803 1660 1804 1700
rect 1844 1660 1845 1700
rect 1803 1651 1845 1660
rect 2187 1700 2229 1709
rect 2187 1660 2188 1700
rect 2228 1660 2229 1700
rect 2187 1651 2229 1660
rect 5259 1700 5301 1709
rect 5259 1660 5260 1700
rect 5300 1660 5301 1700
rect 5259 1651 5301 1660
rect 9675 1700 9717 1709
rect 9675 1660 9676 1700
rect 9716 1660 9717 1700
rect 9675 1651 9717 1660
rect 17355 1700 17397 1709
rect 17355 1660 17356 1700
rect 17396 1660 17397 1700
rect 17355 1651 17397 1660
rect 19371 1700 19413 1709
rect 19371 1660 19372 1700
rect 19412 1660 19413 1700
rect 19371 1651 19413 1660
rect 1152 1532 20352 1556
rect 1152 1492 3688 1532
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 4056 1492 18808 1532
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 19176 1492 20352 1532
rect 1152 1468 20352 1492
rect 20035 1364 20093 1365
rect 20035 1324 20044 1364
rect 20084 1324 20093 1364
rect 20035 1323 20093 1324
rect 2859 1280 2901 1289
rect 2859 1240 2860 1280
rect 2900 1240 2901 1280
rect 2859 1231 2901 1240
rect 4491 1280 4533 1289
rect 4491 1240 4492 1280
rect 4532 1240 4533 1280
rect 4491 1231 4533 1240
rect 5835 1280 5877 1289
rect 5835 1240 5836 1280
rect 5876 1240 5877 1280
rect 5835 1231 5877 1240
rect 7563 1280 7605 1289
rect 7563 1240 7564 1280
rect 7604 1240 7605 1280
rect 7563 1231 7605 1240
rect 11019 1280 11061 1289
rect 11019 1240 11020 1280
rect 11060 1240 11061 1280
rect 11019 1231 11061 1240
rect 12843 1280 12885 1289
rect 12843 1240 12844 1280
rect 12884 1240 12885 1280
rect 12843 1231 12885 1240
rect 14571 1280 14613 1289
rect 14571 1240 14572 1280
rect 14612 1240 14613 1280
rect 14571 1231 14613 1240
rect 16683 1280 16725 1289
rect 16683 1240 16684 1280
rect 16724 1240 16725 1280
rect 16683 1231 16725 1240
rect 17451 1280 17493 1289
rect 17451 1240 17452 1280
rect 17492 1240 17493 1280
rect 17451 1231 17493 1240
rect 17643 1280 17685 1289
rect 17643 1240 17644 1280
rect 17684 1240 17685 1280
rect 17643 1231 17685 1240
rect 5059 1196 5117 1197
rect 5059 1156 5068 1196
rect 5108 1156 5117 1196
rect 5059 1155 5117 1156
rect 5635 1196 5693 1197
rect 5635 1156 5644 1196
rect 5684 1156 5693 1196
rect 5635 1155 5693 1156
rect 14947 1196 15005 1197
rect 14947 1156 14956 1196
rect 14996 1156 15005 1196
rect 14947 1155 15005 1156
rect 17059 1196 17117 1197
rect 17059 1156 17068 1196
rect 17108 1156 17117 1196
rect 17059 1155 17117 1156
rect 1411 1112 1469 1113
rect 1411 1072 1420 1112
rect 1460 1072 1469 1112
rect 1411 1071 1469 1072
rect 2659 1112 2717 1113
rect 2659 1072 2668 1112
rect 2708 1072 2717 1112
rect 2659 1071 2717 1072
rect 3043 1112 3101 1113
rect 3043 1072 3052 1112
rect 3092 1072 3101 1112
rect 3043 1071 3101 1072
rect 4291 1112 4349 1113
rect 4291 1072 4300 1112
rect 4340 1072 4349 1112
rect 4291 1071 4349 1072
rect 6115 1112 6173 1113
rect 6115 1072 6124 1112
rect 6164 1072 6173 1112
rect 6115 1071 6173 1072
rect 7363 1112 7421 1113
rect 7363 1072 7372 1112
rect 7412 1072 7421 1112
rect 7363 1071 7421 1072
rect 7747 1112 7805 1113
rect 7747 1072 7756 1112
rect 7796 1072 7805 1112
rect 7747 1071 7805 1072
rect 8995 1112 9053 1113
rect 8995 1072 9004 1112
rect 9044 1072 9053 1112
rect 8995 1071 9053 1072
rect 9571 1112 9629 1113
rect 9571 1072 9580 1112
rect 9620 1072 9629 1112
rect 9571 1071 9629 1072
rect 10819 1112 10877 1113
rect 10819 1072 10828 1112
rect 10868 1072 10877 1112
rect 10819 1071 10877 1072
rect 11203 1112 11261 1113
rect 11203 1072 11212 1112
rect 11252 1072 11261 1112
rect 11203 1071 11261 1072
rect 12451 1112 12509 1113
rect 12451 1072 12460 1112
rect 12500 1072 12509 1112
rect 12451 1071 12509 1072
rect 13027 1112 13085 1113
rect 13027 1072 13036 1112
rect 13076 1072 13085 1112
rect 13027 1071 13085 1072
rect 14275 1112 14333 1113
rect 14275 1072 14284 1112
rect 14324 1072 14333 1112
rect 14275 1071 14333 1072
rect 15235 1112 15293 1113
rect 15235 1072 15244 1112
rect 15284 1072 15293 1112
rect 15235 1071 15293 1072
rect 16483 1112 16541 1113
rect 16483 1072 16492 1112
rect 16532 1072 16541 1112
rect 16483 1071 16541 1072
rect 17827 1112 17885 1113
rect 17827 1072 17836 1112
rect 17876 1072 17885 1112
rect 17827 1071 17885 1072
rect 19075 1112 19133 1113
rect 19075 1072 19084 1112
rect 19124 1072 19133 1112
rect 19075 1071 19133 1072
rect 19363 1112 19421 1113
rect 19363 1072 19372 1112
rect 19412 1072 19421 1112
rect 19363 1071 19421 1072
rect 19659 1112 19701 1121
rect 19659 1072 19660 1112
rect 19700 1072 19701 1112
rect 19659 1063 19701 1072
rect 19755 1112 19797 1121
rect 19755 1072 19756 1112
rect 19796 1072 19797 1112
rect 19755 1063 19797 1072
rect 4875 1028 4917 1037
rect 4875 988 4876 1028
rect 4916 988 4917 1028
rect 4875 979 4917 988
rect 9195 1028 9237 1037
rect 9195 988 9196 1028
rect 9236 988 9237 1028
rect 9195 979 9237 988
rect 5259 944 5301 953
rect 5259 904 5260 944
rect 5300 904 5301 944
rect 5259 895 5301 904
rect 5451 944 5493 953
rect 5451 904 5452 944
rect 5492 904 5493 944
rect 5451 895 5493 904
rect 9387 944 9429 953
rect 9387 904 9388 944
rect 9428 904 9429 944
rect 9387 895 9429 904
rect 14763 944 14805 953
rect 14763 904 14764 944
rect 14804 904 14805 944
rect 14763 895 14805 904
rect 16875 944 16917 953
rect 16875 904 16876 944
rect 16916 904 16917 944
rect 16875 895 16917 904
rect 1152 776 20452 800
rect 1152 736 4928 776
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 5296 736 20048 776
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20416 736 20452 776
rect 1152 712 20452 736
<< via1 >>
rect 4928 41560 4968 41600
rect 5010 41560 5050 41600
rect 5092 41560 5132 41600
rect 5174 41560 5214 41600
rect 5256 41560 5296 41600
rect 20048 41560 20088 41600
rect 20130 41560 20170 41600
rect 20212 41560 20252 41600
rect 20294 41560 20334 41600
rect 20376 41560 20416 41600
rect 1516 41392 1556 41432
rect 19564 41392 19604 41432
rect 19948 41392 19988 41432
rect 1708 41224 1748 41264
rect 2956 41224 2996 41264
rect 3340 41224 3380 41264
rect 4588 41224 4628 41264
rect 4972 41224 5012 41264
rect 6220 41224 6260 41264
rect 6604 41224 6644 41264
rect 7852 41224 7892 41264
rect 8236 41224 8276 41264
rect 9484 41224 9524 41264
rect 10252 41224 10292 41264
rect 10636 41224 10676 41264
rect 11884 41224 11924 41264
rect 12460 41224 12500 41264
rect 13708 41224 13748 41264
rect 14092 41224 14132 41264
rect 15340 41224 15380 41264
rect 15724 41224 15764 41264
rect 16972 41224 17012 41264
rect 1324 41140 1364 41180
rect 17356 41140 17396 41180
rect 17740 41140 17780 41180
rect 18124 41140 18164 41180
rect 18508 41140 18548 41180
rect 18892 41140 18932 41180
rect 19372 41140 19412 41180
rect 19756 41140 19796 41180
rect 20121 41137 20161 41177
rect 9868 41056 9908 41096
rect 19180 41056 19220 41096
rect 3148 40972 3188 41012
rect 4780 40972 4820 41012
rect 6412 40972 6452 41012
rect 8044 40972 8084 41012
rect 9676 40972 9716 41012
rect 10156 40972 10196 41012
rect 12076 40972 12116 41012
rect 12268 40972 12308 41012
rect 13900 40972 13940 41012
rect 15532 40972 15572 41012
rect 17164 40972 17204 41012
rect 17548 40972 17588 41012
rect 17932 40972 17972 41012
rect 18316 40972 18356 41012
rect 18700 40972 18740 41012
rect 3688 40804 3728 40844
rect 3770 40804 3810 40844
rect 3852 40804 3892 40844
rect 3934 40804 3974 40844
rect 4016 40804 4056 40844
rect 18808 40804 18848 40844
rect 18890 40804 18930 40844
rect 18972 40804 19012 40844
rect 19054 40804 19094 40844
rect 19136 40804 19176 40844
rect 1612 40636 1652 40676
rect 5836 40636 5876 40676
rect 7660 40636 7700 40676
rect 14284 40636 14324 40676
rect 18412 40636 18452 40676
rect 18796 40636 18836 40676
rect 19948 40636 19988 40676
rect 2092 40552 2132 40592
rect 14572 40552 14612 40592
rect 17164 40552 17204 40592
rect 17548 40552 17588 40592
rect 17932 40552 17972 40592
rect 19372 40552 19412 40592
rect 1420 40468 1460 40508
rect 1900 40468 1940 40508
rect 5644 40468 5684 40508
rect 7852 40468 7892 40508
rect 10444 40468 10484 40508
rect 10540 40468 10580 40508
rect 16588 40468 16628 40508
rect 16972 40468 17012 40508
rect 17356 40468 17396 40508
rect 17740 40468 17780 40508
rect 18124 40468 18164 40508
rect 18604 40468 18644 40508
rect 18988 40468 19028 40508
rect 19180 40468 19220 40508
rect 20121 40468 20161 40508
rect 2284 40384 2324 40424
rect 3532 40384 3572 40424
rect 3916 40384 3956 40424
rect 5164 40384 5204 40424
rect 6028 40384 6068 40424
rect 7276 40384 7316 40424
rect 8044 40384 8084 40424
rect 9292 40384 9332 40424
rect 9964 40384 10004 40424
rect 10060 40384 10100 40424
rect 11020 40384 11060 40424
rect 11500 40398 11540 40438
rect 12076 40384 12116 40424
rect 13324 40405 13364 40445
rect 13742 40391 13782 40431
rect 13900 40384 13940 40424
rect 13996 40384 14036 40424
rect 14188 40384 14228 40424
rect 14284 40384 14324 40424
rect 14476 40384 14516 40424
rect 14764 40384 14804 40424
rect 16012 40384 16052 40424
rect 19564 40384 19604 40424
rect 19756 40384 19796 40424
rect 5356 40300 5396 40340
rect 9484 40300 9524 40340
rect 13516 40300 13556 40340
rect 3724 40216 3764 40256
rect 7468 40216 7508 40256
rect 11692 40216 11732 40256
rect 16204 40216 16244 40256
rect 16396 40216 16436 40256
rect 16780 40216 16820 40256
rect 19660 40216 19700 40256
rect 4928 40048 4968 40088
rect 5010 40048 5050 40088
rect 5092 40048 5132 40088
rect 5174 40048 5214 40088
rect 5256 40048 5296 40088
rect 20048 40048 20088 40088
rect 20130 40048 20170 40088
rect 20212 40048 20252 40088
rect 20294 40048 20334 40088
rect 20376 40048 20416 40088
rect 3916 39880 3956 39920
rect 4300 39880 4340 39920
rect 4684 39880 4724 39920
rect 5068 39880 5108 39920
rect 7852 39880 7892 39920
rect 10540 39880 10580 39920
rect 10828 39880 10868 39920
rect 14668 39880 14708 39920
rect 15340 39880 15380 39920
rect 17836 39880 17876 39920
rect 18028 39880 18068 39920
rect 1420 39796 1460 39836
rect 3532 39796 3572 39836
rect 7372 39796 7412 39836
rect 14380 39796 14420 39836
rect 1612 39698 1652 39738
rect 2092 39712 2132 39752
rect 2668 39712 2708 39752
rect 3052 39712 3092 39752
rect 3148 39712 3188 39752
rect 5356 39712 5396 39752
rect 5644 39712 5684 39752
rect 5740 39712 5780 39752
rect 6700 39712 6740 39752
rect 7180 39707 7220 39747
rect 7564 39712 7604 39752
rect 7660 39712 7700 39752
rect 8236 39712 8276 39752
rect 9484 39712 9524 39752
rect 11308 39712 11348 39752
rect 12556 39712 12596 39752
rect 12940 39712 12980 39752
rect 14188 39712 14228 39752
rect 14572 39712 14612 39752
rect 14764 39712 14804 39752
rect 14860 39712 14900 39752
rect 15052 39712 15092 39752
rect 15148 39712 15188 39752
rect 16108 39712 16148 39752
rect 16204 39712 16244 39752
rect 17164 39712 17204 39752
rect 2572 39628 2612 39668
rect 3724 39628 3764 39668
rect 4108 39628 4148 39668
rect 4492 39628 4532 39668
rect 4876 39628 4916 39668
rect 6124 39628 6164 39668
rect 6220 39628 6260 39668
rect 10156 39625 10196 39665
rect 15724 39628 15764 39668
rect 16588 39628 16628 39668
rect 16684 39628 16724 39668
rect 17692 39670 17732 39710
rect 19948 39712 19988 39752
rect 20140 39699 20180 39739
rect 18220 39628 18260 39668
rect 18604 39628 18644 39668
rect 18796 39628 18836 39668
rect 19180 39628 19220 39668
rect 19564 39628 19604 39668
rect 20044 39628 20084 39668
rect 9868 39544 9908 39584
rect 10924 39544 10964 39584
rect 5260 39460 5300 39500
rect 9676 39460 9716 39500
rect 10348 39460 10388 39500
rect 12748 39460 12788 39500
rect 15532 39460 15572 39500
rect 18412 39460 18452 39500
rect 18988 39460 19028 39500
rect 19372 39460 19412 39500
rect 19756 39460 19796 39500
rect 3688 39292 3728 39332
rect 3770 39292 3810 39332
rect 3852 39292 3892 39332
rect 3934 39292 3974 39332
rect 4016 39292 4056 39332
rect 18808 39292 18848 39332
rect 18890 39292 18930 39332
rect 18972 39292 19012 39332
rect 19054 39292 19094 39332
rect 19136 39292 19176 39332
rect 17740 39124 17780 39164
rect 1420 39040 1460 39080
rect 2188 39040 2228 39080
rect 1228 38956 1268 38996
rect 1612 38956 1652 38996
rect 1996 38956 2036 38996
rect 2380 38956 2420 38996
rect 2764 38956 2804 38996
rect 3148 38956 3188 38996
rect 3532 38956 3572 38996
rect 4588 38956 4628 38996
rect 7756 38956 7796 38996
rect 8716 38956 8756 38996
rect 10540 38956 10580 38996
rect 11404 38956 11444 38996
rect 18412 38956 18452 38996
rect 19372 38956 19412 38996
rect 19852 38956 19892 38996
rect 4012 38891 4052 38931
rect 4108 38872 4148 38912
rect 4492 38872 4532 38912
rect 5068 38872 5108 38912
rect 5548 38886 5588 38926
rect 5932 38872 5972 38912
rect 7180 38872 7220 38912
rect 8140 38872 8180 38912
rect 8236 38872 8276 38912
rect 8620 38872 8660 38912
rect 9196 38872 9236 38912
rect 9676 38886 9716 38926
rect 10828 38872 10868 38912
rect 10924 38872 10964 38912
rect 11308 38872 11348 38912
rect 11884 38872 11924 38912
rect 12364 38886 12404 38926
rect 12940 38872 12980 38912
rect 14188 38872 14228 38912
rect 14380 38872 14420 38912
rect 15628 38872 15668 38912
rect 16300 38872 16340 38912
rect 17548 38872 17588 38912
rect 17932 38872 17972 38912
rect 18028 38872 18068 38912
rect 18220 38872 18260 38912
rect 18796 38872 18836 38912
rect 18988 38872 19028 38912
rect 9868 38788 9908 38828
rect 1804 38704 1844 38744
rect 2572 38704 2612 38744
rect 2956 38704 2996 38744
rect 3340 38704 3380 38744
rect 3724 38704 3764 38744
rect 5740 38704 5780 38744
rect 7372 38704 7412 38744
rect 7564 38704 7604 38744
rect 10060 38704 10100 38744
rect 10348 38704 10388 38744
rect 12556 38704 12596 38744
rect 12748 38704 12788 38744
rect 15820 38704 15860 38744
rect 16012 38704 16052 38744
rect 18124 38704 18164 38744
rect 18604 38704 18644 38744
rect 18892 38704 18932 38744
rect 19564 38704 19604 38744
rect 20044 38704 20084 38744
rect 4928 38536 4968 38576
rect 5010 38536 5050 38576
rect 5092 38536 5132 38576
rect 5174 38536 5214 38576
rect 5256 38536 5296 38576
rect 20048 38536 20088 38576
rect 20130 38536 20170 38576
rect 20212 38536 20252 38576
rect 20294 38536 20334 38576
rect 20376 38536 20416 38576
rect 1708 38368 1748 38408
rect 2956 38368 2996 38408
rect 7084 38368 7124 38408
rect 7852 38368 7892 38408
rect 10828 38368 10868 38408
rect 13228 38368 13268 38408
rect 13612 38368 13652 38408
rect 20236 38368 20276 38408
rect 8044 38284 8084 38324
rect 12844 38284 12884 38324
rect 19084 38284 19124 38324
rect 3148 38200 3188 38240
rect 4396 38200 4436 38240
rect 5068 38200 5108 38240
rect 6316 38200 6356 38240
rect 8332 38200 8372 38240
rect 9580 38200 9620 38240
rect 10060 38200 10100 38240
rect 10252 38200 10292 38240
rect 10444 38200 10484 38240
rect 11116 38200 11156 38240
rect 11212 38200 11252 38240
rect 11692 38200 11732 38240
rect 12172 38200 12212 38240
rect 12652 38195 12692 38235
rect 13804 38200 13844 38240
rect 15052 38200 15092 38240
rect 15532 38200 15572 38240
rect 15916 38200 15956 38240
rect 16012 38200 16052 38240
rect 16108 38200 16148 38240
rect 16204 38200 16244 38240
rect 16396 38200 16436 38240
rect 16588 38186 16628 38226
rect 16684 38200 16724 38240
rect 17068 38200 17108 38240
rect 17260 38200 17300 38240
rect 17356 38200 17396 38240
rect 17644 38200 17684 38240
rect 18892 38200 18932 38240
rect 19468 38200 19508 38240
rect 19564 38200 19604 38240
rect 19756 38200 19796 38240
rect 19948 38200 19988 38240
rect 20044 38200 20084 38240
rect 20140 38221 20180 38261
rect 1516 38116 1556 38156
rect 2188 38116 2228 38156
rect 2380 38116 2420 38156
rect 2764 38116 2804 38156
rect 6892 38116 6932 38156
rect 10636 38116 10676 38156
rect 11596 38116 11636 38156
rect 13036 38105 13076 38145
rect 13420 38116 13460 38156
rect 1324 38032 1364 38072
rect 2572 38032 2612 38072
rect 4876 38032 4916 38072
rect 7564 38032 7604 38072
rect 15532 38032 15572 38072
rect 16396 38032 16436 38072
rect 4588 37948 4628 37988
rect 6508 37948 6548 37988
rect 9772 37948 9812 37988
rect 9964 37948 10004 37988
rect 10444 37948 10484 37988
rect 15244 37948 15284 37988
rect 15724 37948 15764 37988
rect 17068 37948 17108 37988
rect 19756 37948 19796 37988
rect 3688 37780 3728 37820
rect 3770 37780 3810 37820
rect 3852 37780 3892 37820
rect 3934 37780 3974 37820
rect 4016 37780 4056 37820
rect 18808 37780 18848 37820
rect 18890 37780 18930 37820
rect 18972 37780 19012 37820
rect 19054 37780 19094 37820
rect 19136 37780 19176 37820
rect 1708 37612 1748 37652
rect 4300 37612 4340 37652
rect 9580 37612 9620 37652
rect 14860 37612 14900 37652
rect 16780 37612 16820 37652
rect 17164 37612 17204 37652
rect 18796 37612 18836 37652
rect 6892 37528 6932 37568
rect 15820 37528 15860 37568
rect 1324 37444 1364 37484
rect 1516 37444 1556 37484
rect 3052 37444 3092 37484
rect 4108 37444 4148 37484
rect 9388 37444 9428 37484
rect 16972 37444 17012 37484
rect 2092 37374 2132 37414
rect 2572 37360 2612 37400
rect 3148 37360 3188 37400
rect 3532 37360 3572 37400
rect 3628 37360 3668 37400
rect 4924 37369 4964 37409
rect 5452 37360 5492 37400
rect 5932 37360 5972 37400
rect 6028 37360 6068 37400
rect 6412 37360 6452 37400
rect 8428 37402 8468 37442
rect 6508 37360 6548 37400
rect 7180 37360 7220 37400
rect 9100 37360 9140 37400
rect 9196 37360 9236 37400
rect 9772 37360 9812 37400
rect 11020 37360 11060 37400
rect 11500 37360 11540 37400
rect 11596 37360 11636 37400
rect 11980 37360 12020 37400
rect 12076 37360 12116 37400
rect 12556 37360 12596 37400
rect 13084 37369 13124 37409
rect 13420 37360 13460 37400
rect 14668 37360 14708 37400
rect 15148 37360 15188 37400
rect 15436 37360 15476 37400
rect 15532 37360 15572 37400
rect 16108 37360 16148 37400
rect 16396 37360 16436 37400
rect 17356 37360 17396 37400
rect 18604 37360 18644 37400
rect 18988 37360 19028 37400
rect 19084 37360 19124 37400
rect 19180 37360 19220 37400
rect 19276 37360 19316 37400
rect 19468 37360 19508 37400
rect 19660 37360 19700 37400
rect 19756 37360 19796 37400
rect 19948 37360 19988 37400
rect 20236 37360 20276 37400
rect 1900 37276 1940 37316
rect 11212 37276 11252 37316
rect 13228 37276 13268 37316
rect 16492 37276 16532 37316
rect 19564 37276 19604 37316
rect 20044 37276 20084 37316
rect 20140 37318 20180 37358
rect 4492 37192 4532 37232
rect 4780 37192 4820 37232
rect 6988 37192 7028 37232
rect 8620 37192 8660 37232
rect 8908 37192 8948 37232
rect 18796 37192 18836 37232
rect 4928 37024 4968 37064
rect 5010 37024 5050 37064
rect 5092 37024 5132 37064
rect 5174 37024 5214 37064
rect 5256 37024 5296 37064
rect 20048 37024 20088 37064
rect 20130 37024 20170 37064
rect 20212 37024 20252 37064
rect 20294 37024 20334 37064
rect 20376 37024 20416 37064
rect 1420 36856 1460 36896
rect 1708 36856 1748 36896
rect 4012 36856 4052 36896
rect 4396 36856 4436 36896
rect 4588 36856 4628 36896
rect 5644 36856 5684 36896
rect 6124 36856 6164 36896
rect 8140 36856 8180 36896
rect 11212 36856 11252 36896
rect 13228 36856 13268 36896
rect 14860 36856 14900 36896
rect 16300 36856 16340 36896
rect 16972 36856 17012 36896
rect 17644 36856 17684 36896
rect 19084 36856 19124 36896
rect 19564 36856 19604 36896
rect 20140 36856 20180 36896
rect 5932 36772 5972 36812
rect 10252 36772 10292 36812
rect 18316 36772 18356 36812
rect 2188 36688 2228 36728
rect 3436 36688 3476 36728
rect 5836 36688 5876 36728
rect 6508 36688 6548 36728
rect 7756 36688 7796 36728
rect 8524 36688 8564 36728
rect 8620 36688 8660 36728
rect 9004 36688 9044 36728
rect 9100 36688 9140 36728
rect 9580 36688 9620 36728
rect 10060 36683 10100 36723
rect 11788 36688 11828 36728
rect 13036 36688 13076 36728
rect 13420 36688 13460 36728
rect 14668 36688 14708 36728
rect 15052 36688 15092 36728
rect 15436 36688 15476 36728
rect 15820 36688 15860 36728
rect 15916 36688 15956 36728
rect 15148 36646 15188 36686
rect 16108 36688 16148 36728
rect 16396 36709 16436 36749
rect 16492 36688 16532 36728
rect 16588 36688 16628 36728
rect 16780 36688 16820 36728
rect 16876 36688 16916 36728
rect 17068 36688 17108 36728
rect 17548 36688 17588 36728
rect 1228 36604 1268 36644
rect 3820 36604 3860 36644
rect 4204 36604 4244 36644
rect 4780 36604 4820 36644
rect 5068 36604 5108 36644
rect 5452 36604 5492 36644
rect 6316 36604 6356 36644
rect 10636 36604 10676 36644
rect 11020 36604 11060 36644
rect 11404 36604 11444 36644
rect 15340 36604 15380 36644
rect 17356 36643 17396 36683
rect 17452 36646 17492 36686
rect 17932 36688 17972 36728
rect 18220 36688 18260 36728
rect 18796 36688 18836 36728
rect 18892 36688 18932 36728
rect 18988 36688 19028 36728
rect 19276 36688 19316 36728
rect 19372 36688 19412 36728
rect 19468 36688 19508 36728
rect 19948 36688 19988 36728
rect 20044 36688 20084 36728
rect 20236 36688 20276 36728
rect 1612 36520 1652 36560
rect 1900 36520 1940 36560
rect 5260 36520 5300 36560
rect 7948 36520 7988 36560
rect 10828 36520 10868 36560
rect 15244 36520 15284 36560
rect 18604 36520 18644 36560
rect 3628 36436 3668 36476
rect 11596 36436 11636 36476
rect 16108 36436 16148 36476
rect 3688 36268 3728 36308
rect 3770 36268 3810 36308
rect 3852 36268 3892 36308
rect 3934 36268 3974 36308
rect 4016 36268 4056 36308
rect 18808 36268 18848 36308
rect 18890 36268 18930 36308
rect 18972 36268 19012 36308
rect 19054 36268 19094 36308
rect 19136 36268 19176 36308
rect 1708 36100 1748 36140
rect 4012 36100 4052 36140
rect 14764 36100 14804 36140
rect 18028 36100 18068 36140
rect 19948 36100 19988 36140
rect 9388 36016 9428 36056
rect 20140 36016 20180 36056
rect 1516 35932 1556 35972
rect 3820 35932 3860 35972
rect 4876 35932 4916 35972
rect 7756 35932 7796 35972
rect 9292 35932 9332 35972
rect 9484 35932 9524 35972
rect 2380 35848 2420 35888
rect 3628 35848 3668 35888
rect 4300 35848 4340 35888
rect 4396 35848 4436 35888
rect 4780 35848 4820 35888
rect 5356 35848 5396 35888
rect 5836 35862 5876 35902
rect 6220 35848 6260 35888
rect 6412 35848 6452 35888
rect 6508 35848 6548 35888
rect 6700 35848 6740 35888
rect 6796 35848 6836 35888
rect 6892 35848 6932 35888
rect 7276 35848 7316 35888
rect 7372 35848 7412 35888
rect 7852 35848 7892 35888
rect 8332 35848 8372 35888
rect 8812 35862 8852 35902
rect 9196 35848 9236 35888
rect 9580 35848 9620 35888
rect 9964 35848 10004 35888
rect 11212 35848 11252 35888
rect 11596 35848 11636 35888
rect 12844 35848 12884 35888
rect 13324 35848 13364 35888
rect 14572 35848 14612 35888
rect 14956 35848 14996 35888
rect 16204 35848 16244 35888
rect 16588 35848 16628 35888
rect 17836 35848 17876 35888
rect 18220 35848 18260 35888
rect 19180 35848 19220 35888
rect 19468 35848 19508 35888
rect 19660 35848 19700 35888
rect 19756 35848 19796 35888
rect 20140 35840 20180 35880
rect 9004 35764 9044 35804
rect 1324 35680 1364 35720
rect 1900 35680 1940 35720
rect 2188 35680 2228 35720
rect 6028 35680 6068 35720
rect 6316 35680 6356 35720
rect 6988 35680 7028 35720
rect 11404 35680 11444 35720
rect 13036 35680 13076 35720
rect 14764 35680 14804 35720
rect 16396 35680 16436 35720
rect 18028 35680 18068 35720
rect 19468 35680 19508 35720
rect 4928 35512 4968 35552
rect 5010 35512 5050 35552
rect 5092 35512 5132 35552
rect 5174 35512 5214 35552
rect 5256 35512 5296 35552
rect 20048 35512 20088 35552
rect 20130 35512 20170 35552
rect 20212 35512 20252 35552
rect 20294 35512 20334 35552
rect 20376 35512 20416 35552
rect 13228 35386 13268 35426
rect 17068 35344 17108 35384
rect 3052 35260 3092 35300
rect 4588 35260 4628 35300
rect 9772 35260 9812 35300
rect 1324 35176 1364 35216
rect 1420 35176 1460 35216
rect 1900 35176 1940 35216
rect 2367 35149 2407 35189
rect 1804 35092 1844 35132
rect 2908 35134 2948 35174
rect 4012 35176 4052 35216
rect 4204 35176 4244 35216
rect 4396 35176 4436 35216
rect 4492 35176 4532 35216
rect 4684 35176 4724 35216
rect 4876 35176 4916 35216
rect 6124 35176 6164 35216
rect 6508 35176 6548 35216
rect 7756 35176 7796 35216
rect 8332 35176 8372 35216
rect 9580 35176 9620 35216
rect 11212 35176 11252 35216
rect 11500 35176 11540 35216
rect 9964 35134 10004 35174
rect 11596 35176 11636 35216
rect 12556 35176 12596 35216
rect 13036 35171 13076 35211
rect 15052 35176 15092 35216
rect 15340 35176 15380 35216
rect 15436 35176 15476 35216
rect 16204 35176 16244 35216
rect 16300 35176 16340 35216
rect 16588 35176 16628 35216
rect 16910 35161 16950 35201
rect 17068 35176 17108 35216
rect 17164 35176 17204 35216
rect 17356 35176 17396 35216
rect 17452 35176 17492 35216
rect 17644 35176 17684 35216
rect 17836 35218 17876 35258
rect 18028 35176 18068 35216
rect 18220 35176 18260 35216
rect 18508 35176 18548 35216
rect 19756 35176 19796 35216
rect 3724 35092 3764 35132
rect 11980 35092 12020 35132
rect 12076 35092 12116 35132
rect 13420 35105 13460 35145
rect 17740 35134 17780 35174
rect 13804 35092 13844 35132
rect 14188 35092 14228 35132
rect 14572 35092 14612 35132
rect 17932 35092 17972 35132
rect 3244 35008 3284 35048
rect 7948 35008 7988 35048
rect 8140 35008 8180 35048
rect 13996 35008 14036 35048
rect 14380 35008 14420 35048
rect 15724 35008 15764 35048
rect 15916 35008 15956 35048
rect 20236 35008 20276 35048
rect 3532 34924 3572 34964
rect 4012 34924 4052 34964
rect 6316 34924 6356 34964
rect 13612 34924 13652 34964
rect 14764 34924 14804 34964
rect 18316 34924 18356 34964
rect 19948 34924 19988 34964
rect 3688 34756 3728 34796
rect 3770 34756 3810 34796
rect 3852 34756 3892 34796
rect 3934 34756 3974 34796
rect 4016 34756 4056 34796
rect 18808 34756 18848 34796
rect 18890 34756 18930 34796
rect 18972 34756 19012 34796
rect 19054 34756 19094 34796
rect 19136 34756 19176 34796
rect 1612 34588 1652 34628
rect 1996 34588 2036 34628
rect 5644 34588 5684 34628
rect 13036 34588 13076 34628
rect 17644 34588 17684 34628
rect 8812 34504 8852 34544
rect 13804 34504 13844 34544
rect 18700 34504 18740 34544
rect 19852 34504 19892 34544
rect 1420 34420 1460 34460
rect 1804 34420 1844 34460
rect 8716 34420 8756 34460
rect 8908 34420 8948 34460
rect 12460 34420 12500 34460
rect 12844 34420 12884 34460
rect 13420 34420 13460 34460
rect 19756 34420 19796 34460
rect 19948 34420 19988 34460
rect 2380 34341 2420 34381
rect 2860 34336 2900 34376
rect 3340 34336 3380 34376
rect 3436 34336 3476 34376
rect 3820 34336 3860 34376
rect 3916 34336 3956 34376
rect 4204 34336 4244 34376
rect 5452 34336 5492 34376
rect 6220 34341 6260 34381
rect 6700 34336 6740 34376
rect 7180 34336 7220 34376
rect 7276 34336 7316 34376
rect 7660 34336 7700 34376
rect 7756 34336 7796 34376
rect 8140 34336 8180 34376
rect 8236 34336 8276 34376
rect 8332 34336 8372 34376
rect 8620 34336 8660 34376
rect 9004 34336 9044 34376
rect 9196 34336 9236 34376
rect 10444 34336 10484 34376
rect 10828 34336 10868 34376
rect 12076 34336 12116 34376
rect 14668 34336 14708 34376
rect 15916 34336 15956 34376
rect 16204 34336 16244 34376
rect 17452 34336 17492 34376
rect 18028 34336 18068 34376
rect 18316 34336 18356 34376
rect 18983 34336 19023 34376
rect 19084 34336 19124 34376
rect 19180 34336 19220 34376
rect 19372 34336 19412 34376
rect 19468 34336 19508 34376
rect 19660 34336 19700 34376
rect 20044 34336 20084 34376
rect 2188 34252 2228 34292
rect 6028 34252 6068 34292
rect 18412 34252 18452 34292
rect 8428 34168 8468 34208
rect 10636 34168 10676 34208
rect 12268 34168 12308 34208
rect 12652 34168 12692 34208
rect 13612 34168 13652 34208
rect 13900 34168 13940 34208
rect 14188 34168 14228 34208
rect 14476 34168 14516 34208
rect 19276 34168 19316 34208
rect 4928 34000 4968 34040
rect 5010 34000 5050 34040
rect 5092 34000 5132 34040
rect 5174 34000 5214 34040
rect 5256 34000 5296 34040
rect 20048 34000 20088 34040
rect 20130 34000 20170 34040
rect 20212 34000 20252 34040
rect 20294 34000 20334 34040
rect 20376 34000 20416 34040
rect 1420 33832 1460 33872
rect 3628 33832 3668 33872
rect 4108 33832 4148 33872
rect 7948 33832 7988 33872
rect 12364 33832 12404 33872
rect 14668 33832 14708 33872
rect 16684 33832 16724 33872
rect 8428 33748 8468 33788
rect 1612 33664 1652 33704
rect 2860 33664 2900 33704
rect 4300 33650 4340 33690
rect 4780 33664 4820 33704
rect 5260 33664 5300 33704
rect 5740 33664 5780 33704
rect 5836 33664 5876 33704
rect 6220 33664 6260 33704
rect 6316 33664 6356 33704
rect 7276 33664 7316 33704
rect 7756 33659 7796 33699
rect 8620 33664 8660 33704
rect 9868 33664 9908 33704
rect 10060 33664 10100 33704
rect 10252 33664 10292 33704
rect 10348 33664 10388 33704
rect 10636 33664 10676 33704
rect 10732 33664 10772 33704
rect 11692 33664 11732 33704
rect 12220 33654 12260 33694
rect 13804 33664 13844 33704
rect 14188 33664 14228 33704
rect 14284 33664 14324 33704
rect 14476 33664 14516 33704
rect 1228 33580 1268 33620
rect 3244 33580 3284 33620
rect 3820 33580 3860 33620
rect 5356 33580 5396 33620
rect 6700 33580 6740 33620
rect 6796 33580 6836 33620
rect 11116 33580 11156 33620
rect 12556 33622 12596 33662
rect 14572 33664 14612 33704
rect 14673 33664 14713 33704
rect 15532 33664 15572 33704
rect 15628 33664 15668 33704
rect 15916 33664 15956 33704
rect 16204 33651 16244 33691
rect 16396 33664 16436 33704
rect 16492 33664 16532 33704
rect 16876 33664 16916 33704
rect 18124 33664 18164 33704
rect 18412 33664 18452 33704
rect 18700 33664 18740 33704
rect 18796 33664 18836 33704
rect 19276 33664 19316 33704
rect 19660 33664 19700 33704
rect 11212 33580 11252 33620
rect 19372 33580 19412 33620
rect 19564 33580 19604 33620
rect 19852 33580 19892 33620
rect 8140 33496 8180 33536
rect 14956 33496 14996 33536
rect 19084 33496 19124 33536
rect 19468 33496 19508 33536
rect 3052 33412 3092 33452
rect 3436 33412 3476 33452
rect 10060 33412 10100 33452
rect 13996 33412 14036 33452
rect 15244 33412 15284 33452
rect 16204 33412 16244 33452
rect 20044 33412 20084 33452
rect 3688 33244 3728 33284
rect 3770 33244 3810 33284
rect 3852 33244 3892 33284
rect 3934 33244 3974 33284
rect 4016 33244 4056 33284
rect 18808 33244 18848 33284
rect 18890 33244 18930 33284
rect 18972 33244 19012 33284
rect 19054 33244 19094 33284
rect 19136 33244 19176 33284
rect 3436 33076 3476 33116
rect 3820 33076 3860 33116
rect 6124 33076 6164 33116
rect 7756 33076 7796 33116
rect 12652 33076 12692 33116
rect 15052 33076 15092 33116
rect 15436 33076 15476 33116
rect 19276 33076 19316 33116
rect 5932 32992 5972 33032
rect 14668 32992 14708 33032
rect 17260 32992 17300 33032
rect 18316 32992 18356 33032
rect 19948 32992 19988 33032
rect 14476 32908 14516 32948
rect 14860 32908 14900 32948
rect 19852 32908 19892 32948
rect 20044 32908 20084 32948
rect 1324 32824 1364 32864
rect 2572 32824 2612 32864
rect 3052 32824 3092 32864
rect 3244 32824 3284 32864
rect 3436 32824 3476 32864
rect 3628 32824 3668 32864
rect 3820 32824 3860 32864
rect 4012 32824 4052 32864
rect 4108 32824 4148 32864
rect 4204 32824 4244 32864
rect 4300 32824 4340 32864
rect 4492 32824 4532 32864
rect 5740 32824 5780 32864
rect 6316 32824 6356 32864
rect 7564 32824 7604 32864
rect 7948 32824 7988 32864
rect 9196 32824 9236 32864
rect 9580 32824 9620 32864
rect 9676 32824 9716 32864
rect 10060 32824 10100 32864
rect 10156 32803 10196 32843
rect 10252 32824 10292 32864
rect 10348 32824 10388 32864
rect 10636 32824 10676 32864
rect 11884 32824 11924 32864
rect 12844 32824 12884 32864
rect 14092 32824 14132 32864
rect 15244 32824 15284 32864
rect 15436 32824 15476 32864
rect 15820 32824 15860 32864
rect 17068 32824 17108 32864
rect 17644 32824 17684 32864
rect 17932 32824 17972 32864
rect 20140 32866 20180 32906
rect 18028 32824 18068 32864
rect 18604 32824 18644 32864
rect 19756 32824 19796 32864
rect 12460 32740 12500 32780
rect 19468 32740 19508 32780
rect 2764 32656 2804 32696
rect 2956 32656 2996 32696
rect 9868 32656 9908 32696
rect 12076 32656 12116 32696
rect 15340 32656 15380 32696
rect 15628 32656 15668 32696
rect 4928 32488 4968 32528
rect 5010 32488 5050 32528
rect 5092 32488 5132 32528
rect 5174 32488 5214 32528
rect 5256 32488 5296 32528
rect 20048 32488 20088 32528
rect 20130 32488 20170 32528
rect 20212 32488 20252 32528
rect 20294 32488 20334 32528
rect 20376 32488 20416 32528
rect 1324 32320 1364 32360
rect 1708 32320 1748 32360
rect 3724 32320 3764 32360
rect 4396 32320 4436 32360
rect 6220 32320 6260 32360
rect 8140 32320 8180 32360
rect 12460 32320 12500 32360
rect 15916 32320 15956 32360
rect 17644 32320 17684 32360
rect 10252 32236 10292 32276
rect 12268 32236 12308 32276
rect 1228 32152 1268 32192
rect 1996 32152 2036 32192
rect 2092 32152 2132 32192
rect 3052 32152 3092 32192
rect 3532 32138 3572 32178
rect 3916 32152 3956 32192
rect 4012 32152 4052 32192
rect 4204 32152 4244 32192
rect 4300 32152 4340 32192
rect 4401 32152 4441 32192
rect 4780 32152 4820 32192
rect 6028 32152 6068 32192
rect 6412 32152 6452 32192
rect 7660 32152 7700 32192
rect 8332 32152 8372 32192
rect 8524 32152 8564 32192
rect 8620 32152 8660 32192
rect 8812 32152 8852 32192
rect 10060 32152 10100 32192
rect 10540 32152 10580 32192
rect 10636 32152 10676 32192
rect 11020 32152 11060 32192
rect 11596 32152 11636 32192
rect 12076 32147 12116 32187
rect 12748 32152 12788 32192
rect 13996 32152 14036 32192
rect 14668 32152 14708 32192
rect 14764 32152 14804 32192
rect 15052 32152 15092 32192
rect 15340 32152 15380 32192
rect 15724 32152 15764 32192
rect 16204 32152 16244 32192
rect 17452 32152 17492 32192
rect 17836 32152 17876 32192
rect 18028 32152 18068 32192
rect 18220 32152 18260 32192
rect 19468 32152 19508 32192
rect 1516 32068 1556 32108
rect 2476 32068 2516 32108
rect 2572 32068 2612 32108
rect 11116 32068 11156 32108
rect 15436 32068 15476 32108
rect 15628 32068 15668 32108
rect 19852 32068 19892 32108
rect 8044 31984 8084 32024
rect 8620 31984 8660 32024
rect 14380 31984 14420 32024
rect 15532 31984 15572 32024
rect 7852 31900 7892 31940
rect 14188 31900 14228 31940
rect 17644 31900 17684 31940
rect 17836 31900 17876 31940
rect 19660 31900 19700 31940
rect 20044 31900 20084 31940
rect 3688 31732 3728 31772
rect 3770 31732 3810 31772
rect 3852 31732 3892 31772
rect 3934 31732 3974 31772
rect 4016 31732 4056 31772
rect 18808 31732 18848 31772
rect 18890 31732 18930 31772
rect 18972 31732 19012 31772
rect 19054 31732 19094 31772
rect 19136 31732 19176 31772
rect 9868 31564 9908 31604
rect 2188 31480 2228 31520
rect 16684 31480 16724 31520
rect 18412 31480 18452 31520
rect 19660 31480 19700 31520
rect 6700 31396 6740 31436
rect 2092 31354 2132 31394
rect 8140 31396 8180 31436
rect 1900 31312 1940 31352
rect 2188 31312 2228 31352
rect 2380 31312 2420 31352
rect 2572 31312 2612 31352
rect 3820 31312 3860 31352
rect 4204 31312 4244 31352
rect 5452 31312 5492 31352
rect 6124 31312 6164 31352
rect 6220 31312 6260 31352
rect 6604 31312 6644 31352
rect 7180 31312 7220 31352
rect 7660 31326 7700 31366
rect 8044 31312 8084 31352
rect 8236 31312 8276 31352
rect 8428 31312 8468 31352
rect 9676 31312 9716 31352
rect 10060 31312 10100 31352
rect 11308 31312 11348 31352
rect 11692 31312 11732 31352
rect 12940 31312 12980 31352
rect 13516 31352 13556 31392
rect 14764 31396 14804 31436
rect 19564 31396 19604 31436
rect 19756 31396 19796 31436
rect 20044 31396 20084 31436
rect 13612 31312 13652 31352
rect 13708 31312 13748 31352
rect 13900 31312 13940 31352
rect 14092 31312 14132 31352
rect 14188 31312 14228 31352
rect 14668 31312 14708 31352
rect 15148 31312 15188 31352
rect 16396 31312 16436 31352
rect 17068 31312 17108 31352
rect 17356 31312 17396 31352
rect 17740 31312 17780 31352
rect 18028 31312 18068 31352
rect 18734 31327 18774 31367
rect 18892 31312 18932 31352
rect 18988 31312 19028 31352
rect 19180 31312 19220 31352
rect 19276 31312 19316 31352
rect 19468 31312 19508 31352
rect 19852 31312 19892 31352
rect 1612 31228 1652 31268
rect 5644 31228 5684 31268
rect 7852 31228 7892 31268
rect 13996 31228 14036 31268
rect 16972 31228 17012 31268
rect 18124 31228 18164 31268
rect 1324 31144 1364 31184
rect 1804 31144 1844 31184
rect 4012 31144 4052 31184
rect 9868 31144 9908 31184
rect 11500 31144 11540 31184
rect 13132 31144 13172 31184
rect 13420 31144 13460 31184
rect 14380 31144 14420 31184
rect 14956 31144 14996 31184
rect 19084 31144 19124 31184
rect 20236 31144 20276 31184
rect 4928 30976 4968 31016
rect 5010 30976 5050 31016
rect 5092 30976 5132 31016
rect 5174 30976 5214 31016
rect 5256 30976 5296 31016
rect 20048 30976 20088 31016
rect 20130 30976 20170 31016
rect 20212 30976 20252 31016
rect 20294 30976 20334 31016
rect 20376 30976 20416 31016
rect 5836 30808 5876 30848
rect 9388 30808 9428 30848
rect 9868 30808 9908 30848
rect 14380 30808 14420 30848
rect 17644 30808 17684 30848
rect 20044 30808 20084 30848
rect 2668 30724 2708 30764
rect 11884 30724 11924 30764
rect 13900 30724 13940 30764
rect 17452 30724 17492 30764
rect 19564 30724 19604 30764
rect 1228 30640 1268 30680
rect 2476 30640 2516 30680
rect 2860 30640 2900 30680
rect 3052 30640 3092 30680
rect 3340 30640 3380 30680
rect 3628 30640 3668 30680
rect 3724 30640 3764 30680
rect 4204 30640 4244 30680
rect 5452 30640 5492 30680
rect 6028 30640 6068 30680
rect 7276 30640 7316 30680
rect 7468 30640 7508 30680
rect 7564 30640 7604 30680
rect 7660 30640 7700 30680
rect 7756 30640 7796 30680
rect 7948 30640 7988 30680
rect 9196 30640 9236 30680
rect 9580 30640 9620 30680
rect 9676 30640 9716 30680
rect 9868 30640 9908 30680
rect 9964 30640 10004 30680
rect 10065 30640 10105 30680
rect 10444 30640 10484 30680
rect 11692 30640 11732 30680
rect 12172 30640 12212 30680
rect 12268 30640 12308 30680
rect 12652 30640 12692 30680
rect 13228 30640 13268 30680
rect 13756 30630 13796 30670
rect 14188 30651 14228 30691
rect 14668 30640 14708 30680
rect 14860 30640 14900 30680
rect 15052 30640 15092 30680
rect 15436 30640 15476 30680
rect 15724 30640 15764 30680
rect 15820 30640 15860 30680
rect 16780 30640 16820 30680
rect 17260 30626 17300 30666
rect 17836 30640 17876 30680
rect 18124 30640 18164 30680
rect 19372 30640 19412 30680
rect 19756 30640 19796 30680
rect 19852 30640 19892 30680
rect 20044 30640 20084 30680
rect 12748 30556 12788 30596
rect 15148 30556 15188 30596
rect 15340 30556 15380 30596
rect 16204 30556 16244 30596
rect 16300 30556 16340 30596
rect 15244 30472 15284 30512
rect 17836 30472 17876 30512
rect 3052 30388 3092 30428
rect 4012 30388 4052 30428
rect 5644 30388 5684 30428
rect 14092 30388 14132 30428
rect 14668 30388 14708 30428
rect 3688 30220 3728 30260
rect 3770 30220 3810 30260
rect 3852 30220 3892 30260
rect 3934 30220 3974 30260
rect 4016 30220 4056 30260
rect 18808 30220 18848 30260
rect 18890 30220 18930 30260
rect 18972 30220 19012 30260
rect 19054 30220 19094 30260
rect 19136 30220 19176 30260
rect 2860 30052 2900 30092
rect 10828 30052 10868 30092
rect 17260 30052 17300 30092
rect 7372 29968 7412 30008
rect 11020 29968 11060 30008
rect 20236 29968 20276 30008
rect 5740 29884 5780 29924
rect 12172 29884 12212 29924
rect 17548 29884 17588 29924
rect 1228 29800 1268 29840
rect 2476 29800 2516 29840
rect 3052 29800 3092 29840
rect 4300 29800 4340 29840
rect 4780 29814 4820 29854
rect 5260 29800 5300 29840
rect 5836 29800 5876 29840
rect 6220 29800 6260 29840
rect 6316 29800 6356 29840
rect 6700 29800 6740 29840
rect 6988 29800 7028 29840
rect 7564 29800 7604 29840
rect 8812 29800 8852 29840
rect 9388 29800 9428 29840
rect 9484 29800 9524 29840
rect 9580 29800 9620 29840
rect 9868 29800 9908 29840
rect 9964 29800 10004 29840
rect 10156 29800 10196 29840
rect 10348 29800 10388 29840
rect 10444 29808 10484 29848
rect 10540 29800 10580 29840
rect 11020 29800 11060 29840
rect 11596 29800 11636 29840
rect 11692 29800 11732 29840
rect 12076 29800 12116 29840
rect 12652 29800 12692 29840
rect 13132 29814 13172 29854
rect 13708 29800 13748 29840
rect 13804 29800 13844 29840
rect 13900 29800 13940 29840
rect 13996 29800 14036 29840
rect 14188 29800 14228 29840
rect 15436 29800 15476 29840
rect 15820 29800 15860 29840
rect 17068 29800 17108 29840
rect 17452 29800 17492 29840
rect 17644 29800 17684 29840
rect 17836 29800 17876 29840
rect 19084 29800 19124 29840
rect 19564 29800 19604 29840
rect 19852 29800 19892 29840
rect 4588 29716 4628 29756
rect 7084 29716 7124 29756
rect 13324 29716 13364 29756
rect 19276 29716 19316 29756
rect 19948 29716 19988 29756
rect 2668 29632 2708 29672
rect 9004 29632 9044 29672
rect 9676 29632 9716 29672
rect 10060 29632 10100 29672
rect 10636 29632 10676 29672
rect 15628 29632 15668 29672
rect 4928 29464 4968 29504
rect 5010 29464 5050 29504
rect 5092 29464 5132 29504
rect 5174 29464 5214 29504
rect 5256 29464 5296 29504
rect 20048 29464 20088 29504
rect 20130 29464 20170 29504
rect 20212 29464 20252 29504
rect 20294 29464 20334 29504
rect 20376 29464 20416 29504
rect 3628 29296 3668 29336
rect 8428 29296 8468 29336
rect 8812 29296 8852 29336
rect 9292 29296 9332 29336
rect 15916 29212 15956 29252
rect 1420 29128 1460 29168
rect 1804 29128 1844 29168
rect 1996 29128 2036 29168
rect 3244 29128 3284 29168
rect 3820 29128 3860 29168
rect 5068 29128 5108 29168
rect 5548 29128 5588 29168
rect 5644 29128 5684 29168
rect 5932 29128 5972 29168
rect 6220 29128 6260 29168
rect 6604 29128 6644 29168
rect 6988 29128 7028 29168
rect 8236 29128 8276 29168
rect 8620 29128 8660 29168
rect 8716 29128 8756 29168
rect 8908 29128 8948 29168
rect 9100 29128 9140 29168
rect 9196 29128 9236 29168
rect 9388 29128 9428 29168
rect 9772 29128 9812 29168
rect 11020 29128 11060 29168
rect 11212 29128 11252 29168
rect 12460 29128 12500 29168
rect 12844 29128 12884 29168
rect 13036 29128 13076 29168
rect 13132 29128 13172 29168
rect 13324 29128 13364 29168
rect 13612 29128 13652 29168
rect 14860 29128 14900 29168
rect 15532 29128 15572 29168
rect 15820 29128 15860 29168
rect 16396 29128 16436 29168
rect 16780 29128 16820 29168
rect 17068 29128 17108 29168
rect 18316 29128 18356 29168
rect 19180 29128 19220 29168
rect 1516 29044 1556 29084
rect 1708 29044 1748 29084
rect 16492 29044 16532 29084
rect 16684 29044 16724 29084
rect 18700 29044 18740 29084
rect 1612 28960 1652 29000
rect 6604 28960 6644 29000
rect 9580 28960 9620 29000
rect 13036 28960 13076 29000
rect 16588 28960 16628 29000
rect 18508 28960 18548 29000
rect 18892 28960 18932 29000
rect 19852 28960 19892 29000
rect 3436 28876 3476 28916
rect 5260 28876 5300 28916
rect 6316 28876 6356 28916
rect 6796 28876 6836 28916
rect 12652 28876 12692 28916
rect 13420 28876 13460 28916
rect 15052 28876 15092 28916
rect 16204 28876 16244 28916
rect 3688 28708 3728 28748
rect 3770 28708 3810 28748
rect 3852 28708 3892 28748
rect 3934 28708 3974 28748
rect 4016 28708 4056 28748
rect 18808 28708 18848 28748
rect 18890 28708 18930 28748
rect 18972 28708 19012 28748
rect 19054 28708 19094 28748
rect 19136 28708 19176 28748
rect 9772 28540 9812 28580
rect 10732 28540 10772 28580
rect 12844 28540 12884 28580
rect 15436 28540 15476 28580
rect 4108 28456 4148 28496
rect 5932 28456 5972 28496
rect 6412 28456 6452 28496
rect 2572 28372 2612 28412
rect 4012 28372 4052 28412
rect 4204 28372 4244 28412
rect 6316 28372 6356 28412
rect 6508 28372 6548 28412
rect 19852 28372 19892 28412
rect 1996 28288 2036 28328
rect 2092 28288 2132 28328
rect 2476 28288 2516 28328
rect 3052 28288 3092 28328
rect 3532 28302 3572 28342
rect 3916 28288 3956 28328
rect 4300 28288 4340 28328
rect 4492 28288 4532 28328
rect 5740 28288 5780 28328
rect 6220 28288 6260 28328
rect 6604 28288 6644 28328
rect 6892 28288 6932 28328
rect 8140 28288 8180 28328
rect 8620 28288 8660 28328
rect 8716 28288 8756 28328
rect 8812 28288 8852 28328
rect 9100 28288 9140 28328
rect 9388 28288 9428 28328
rect 9484 28288 9524 28328
rect 9964 28288 10004 28328
rect 10060 28288 10100 28328
rect 10156 28288 10196 28328
rect 10252 28288 10292 28328
rect 10444 28288 10484 28328
rect 10540 28288 10580 28328
rect 10732 28288 10772 28328
rect 10924 28301 10964 28341
rect 11116 28288 11156 28328
rect 11404 28288 11444 28328
rect 12652 28288 12692 28328
rect 13036 28288 13076 28328
rect 13132 28288 13172 28328
rect 13324 28288 13364 28328
rect 13420 28288 13460 28328
rect 13521 28288 13561 28328
rect 13996 28288 14036 28328
rect 15244 28288 15284 28328
rect 15436 28288 15476 28328
rect 15532 28288 15572 28328
rect 15724 28288 15764 28328
rect 15820 28288 15860 28328
rect 15977 28303 16017 28343
rect 16204 28288 16244 28328
rect 17452 28288 17492 28328
rect 17932 28288 17972 28328
rect 18028 28288 18068 28328
rect 18412 28288 18452 28328
rect 18508 28288 18548 28328
rect 18988 28288 19028 28328
rect 19468 28293 19508 28333
rect 3724 28204 3764 28244
rect 8524 28204 8564 28244
rect 19660 28204 19700 28244
rect 1324 28120 1364 28160
rect 1612 28120 1652 28160
rect 8332 28120 8372 28160
rect 11020 28120 11060 28160
rect 13420 28120 13460 28160
rect 13804 28120 13844 28160
rect 17644 28120 17684 28160
rect 20044 28120 20084 28160
rect 4928 27952 4968 27992
rect 5010 27952 5050 27992
rect 5092 27952 5132 27992
rect 5174 27952 5214 27992
rect 5256 27952 5296 27992
rect 20048 27952 20088 27992
rect 20130 27952 20170 27992
rect 20212 27952 20252 27992
rect 20294 27952 20334 27992
rect 20376 27952 20416 27992
rect 9676 27784 9716 27824
rect 9868 27784 9908 27824
rect 13804 27784 13844 27824
rect 14860 27784 14900 27824
rect 3148 27700 3188 27740
rect 7852 27700 7892 27740
rect 19564 27700 19604 27740
rect 1228 27616 1268 27656
rect 2476 27616 2516 27656
rect 3244 27616 3284 27656
rect 3532 27616 3572 27656
rect 3820 27616 3860 27656
rect 3916 27616 3956 27656
rect 4108 27616 4148 27656
rect 4300 27616 4340 27656
rect 5548 27616 5588 27656
rect 6124 27616 6164 27656
rect 7372 27616 7412 27656
rect 7756 27616 7796 27656
rect 7948 27616 7988 27656
rect 8044 27616 8084 27656
rect 8236 27616 8276 27656
rect 8332 27616 8372 27656
rect 8524 27616 8564 27656
rect 8812 27616 8852 27656
rect 8908 27616 8948 27656
rect 9004 27616 9044 27656
rect 9388 27616 9428 27656
rect 9484 27616 9524 27656
rect 9964 27616 10004 27656
rect 10156 27616 10196 27656
rect 11404 27616 11444 27656
rect 11884 27616 11924 27656
rect 13132 27616 13172 27656
rect 13516 27616 13556 27656
rect 13612 27616 13652 27656
rect 14572 27616 14612 27656
rect 14668 27616 14708 27656
rect 14860 27616 14900 27656
rect 15148 27599 15188 27639
rect 15436 27616 15476 27656
rect 15532 27616 15572 27656
rect 16012 27616 16052 27656
rect 16396 27616 16436 27656
rect 16588 27616 16628 27656
rect 16780 27616 16820 27656
rect 17836 27616 17876 27656
rect 17932 27616 17972 27656
rect 18892 27616 18932 27656
rect 19372 27611 19412 27651
rect 20127 27603 20167 27643
rect 14188 27532 14228 27572
rect 16108 27532 16148 27572
rect 16300 27532 16340 27572
rect 16972 27532 17012 27572
rect 17356 27532 17396 27572
rect 18316 27532 18356 27572
rect 18412 27532 18452 27572
rect 19756 27532 19796 27572
rect 2668 27448 2708 27488
rect 8524 27448 8564 27488
rect 15820 27448 15860 27488
rect 16204 27448 16244 27488
rect 16588 27448 16628 27488
rect 17164 27448 17204 27488
rect 17548 27448 17588 27488
rect 2860 27364 2900 27404
rect 4108 27364 4148 27404
rect 5740 27364 5780 27404
rect 7564 27364 7604 27404
rect 9196 27364 9236 27404
rect 11596 27364 11636 27404
rect 13324 27364 13364 27404
rect 13996 27364 14036 27404
rect 19948 27364 19988 27404
rect 20236 27364 20276 27404
rect 3688 27196 3728 27236
rect 3770 27196 3810 27236
rect 3852 27196 3892 27236
rect 3934 27196 3974 27236
rect 4016 27196 4056 27236
rect 18808 27196 18848 27236
rect 18890 27196 18930 27236
rect 18972 27196 19012 27236
rect 19054 27196 19094 27236
rect 19136 27196 19176 27236
rect 2668 27028 2708 27068
rect 8812 27028 8852 27068
rect 13708 27028 13748 27068
rect 17740 27028 17780 27068
rect 18124 27028 18164 27068
rect 3820 26944 3860 26984
rect 4204 26944 4244 26984
rect 6316 26944 6356 26984
rect 9292 26944 9332 26984
rect 11404 26944 11444 26984
rect 13996 26944 14036 26984
rect 16396 26944 16436 26984
rect 18508 26944 18548 26984
rect 6230 26860 6270 26900
rect 6412 26860 6452 26900
rect 12172 26860 12212 26900
rect 14284 26860 14324 26900
rect 16300 26860 16340 26900
rect 16492 26860 16532 26900
rect 17548 26860 17588 26900
rect 17932 26860 17972 26900
rect 18316 26871 18356 26911
rect 19564 26860 19604 26900
rect 19948 26860 19988 26900
rect 1228 26776 1268 26816
rect 2476 26776 2516 26816
rect 3148 26776 3188 26816
rect 3436 26776 3476 26816
rect 4012 26776 4052 26816
rect 4204 26776 4244 26816
rect 4396 26776 4436 26816
rect 5644 26776 5684 26816
rect 6124 26776 6164 26816
rect 6508 26776 6548 26816
rect 6796 26776 6836 26816
rect 6892 26776 6932 26816
rect 7276 26776 7316 26816
rect 7372 26776 7412 26816
rect 7852 26776 7892 26816
rect 8332 26790 8372 26830
rect 8716 26776 8756 26816
rect 9100 26776 9140 26816
rect 9484 26776 9524 26816
rect 9676 26776 9716 26816
rect 9772 26776 9812 26816
rect 9964 26776 10004 26816
rect 11212 26776 11252 26816
rect 11692 26795 11732 26835
rect 11788 26756 11828 26796
rect 12268 26776 12308 26816
rect 12748 26776 12788 26816
rect 13276 26785 13316 26825
rect 13804 26776 13844 26816
rect 14092 26776 14132 26816
rect 14380 26776 14420 26816
rect 14572 26776 14612 26816
rect 15820 26776 15860 26816
rect 16204 26776 16244 26816
rect 16780 26818 16820 26858
rect 16588 26776 16628 26816
rect 16972 26776 17012 26816
rect 17068 26776 17108 26816
rect 17260 26776 17300 26816
rect 18700 26776 18740 26816
rect 18796 26776 18836 26816
rect 18988 26776 19028 26816
rect 19180 26776 19220 26816
rect 19372 26776 19412 26816
rect 3532 26692 3572 26732
rect 5836 26608 5876 26648
rect 8524 26608 8564 26648
rect 9004 26608 9044 26648
rect 9580 26608 9620 26648
rect 13420 26608 13460 26648
rect 16012 26608 16052 26648
rect 16780 26608 16820 26648
rect 17356 26608 17396 26648
rect 18988 26608 19028 26648
rect 19276 26608 19316 26648
rect 19756 26608 19796 26648
rect 20140 26608 20180 26648
rect 4928 26440 4968 26480
rect 5010 26440 5050 26480
rect 5092 26440 5132 26480
rect 5174 26440 5214 26480
rect 5256 26440 5296 26480
rect 20048 26440 20088 26480
rect 20130 26440 20170 26480
rect 20212 26440 20252 26480
rect 20294 26440 20334 26480
rect 20376 26440 20416 26480
rect 3628 26272 3668 26312
rect 6988 26272 7028 26312
rect 11500 26272 11540 26312
rect 11884 26272 11924 26312
rect 15436 26272 15476 26312
rect 16684 26272 16724 26312
rect 17452 26272 17492 26312
rect 12076 26188 12116 26228
rect 1324 26104 1364 26144
rect 1516 26104 1556 26144
rect 2764 26104 2804 26144
rect 3241 26108 3281 26148
rect 3340 26104 3380 26144
rect 3506 26104 3546 26144
rect 3628 26075 3668 26115
rect 3772 26104 3812 26144
rect 4012 26104 4052 26144
rect 4396 26104 4436 26144
rect 4588 26104 4628 26144
rect 4780 26104 4820 26144
rect 5068 26104 5108 26144
rect 5356 26104 5396 26144
rect 5452 26104 5492 26144
rect 6028 26104 6068 26144
rect 6316 26104 6356 26144
rect 6412 26104 6452 26144
rect 6926 26089 6966 26129
rect 7084 26104 7124 26144
rect 7180 26104 7220 26144
rect 7372 26104 7412 26144
rect 7468 26104 7508 26144
rect 7756 26104 7796 26144
rect 7852 26104 7892 26144
rect 8044 26104 8084 26144
rect 8428 26104 8468 26144
rect 9676 26104 9716 26144
rect 9868 26104 9908 26144
rect 11116 26104 11156 26144
rect 11788 26104 11828 26144
rect 12364 26104 12404 26144
rect 13612 26104 13652 26144
rect 13996 26104 14036 26144
rect 15244 26104 15284 26144
rect 15724 26104 15764 26144
rect 16012 26104 16052 26144
rect 16108 26104 16148 26144
rect 16622 26089 16662 26129
rect 16780 26104 16820 26144
rect 16876 26104 16916 26144
rect 17068 26104 17108 26144
rect 17164 26104 17204 26144
rect 17356 26104 17396 26144
rect 17548 26104 17588 26144
rect 17740 26104 17780 26144
rect 18988 26104 19028 26144
rect 19372 26104 19412 26144
rect 19756 26104 19796 26144
rect 1228 26020 1268 26060
rect 4108 26020 4148 26060
rect 4300 26020 4340 26060
rect 19468 26020 19508 26060
rect 19660 26020 19700 26060
rect 19948 26020 19988 26060
rect 2956 25936 2996 25976
rect 4204 25936 4244 25976
rect 5740 25936 5780 25976
rect 6700 25936 6740 25976
rect 16396 25936 16436 25976
rect 19564 25936 19604 25976
rect 4588 25852 4628 25892
rect 7852 25852 7892 25892
rect 8236 25852 8276 25892
rect 11308 25852 11348 25892
rect 13804 25852 13844 25892
rect 19180 25852 19220 25892
rect 20140 25852 20180 25892
rect 3688 25684 3728 25724
rect 3770 25684 3810 25724
rect 3852 25684 3892 25724
rect 3934 25684 3974 25724
rect 4016 25684 4056 25724
rect 18808 25684 18848 25724
rect 18890 25684 18930 25724
rect 18972 25684 19012 25724
rect 19054 25684 19094 25724
rect 19136 25684 19176 25724
rect 5644 25516 5684 25556
rect 6220 25516 6260 25556
rect 8044 25516 8084 25556
rect 15532 25516 15572 25556
rect 16492 25516 16532 25556
rect 19660 25516 19700 25556
rect 3244 25432 3284 25472
rect 9004 25432 9044 25472
rect 9388 25432 9428 25472
rect 16876 25432 16916 25472
rect 20044 25432 20084 25472
rect 3148 25348 3188 25388
rect 3340 25348 3380 25388
rect 9292 25348 9332 25388
rect 9484 25348 9524 25388
rect 11596 25348 11636 25388
rect 12748 25348 12788 25388
rect 16780 25348 16820 25388
rect 16972 25348 17012 25388
rect 19948 25348 19988 25388
rect 20130 25348 20170 25388
rect 1228 25264 1268 25304
rect 2476 25264 2516 25304
rect 3052 25264 3092 25304
rect 3436 25264 3476 25304
rect 3628 25264 3668 25304
rect 4876 25264 4916 25304
rect 5260 25264 5300 25304
rect 5452 25264 5492 25304
rect 5740 25264 5780 25304
rect 5932 25264 5972 25304
rect 6028 25264 6068 25304
rect 6220 25264 6260 25304
rect 6604 25264 6644 25304
rect 7852 25264 7892 25304
rect 8332 25264 8372 25304
rect 8620 25264 8660 25304
rect 8716 25264 8756 25304
rect 9196 25264 9236 25304
rect 9580 25264 9620 25304
rect 9868 25264 9908 25304
rect 11116 25264 11156 25304
rect 12172 25264 12212 25304
rect 12268 25264 12308 25304
rect 12652 25264 12692 25304
rect 13228 25264 13268 25304
rect 13708 25278 13748 25318
rect 14092 25264 14132 25304
rect 15340 25264 15380 25304
rect 15820 25264 15860 25304
rect 16108 25264 16148 25304
rect 16684 25264 16724 25304
rect 17068 25264 17108 25304
rect 17452 25264 17492 25304
rect 18700 25264 18740 25304
rect 18988 25264 19028 25304
rect 19276 25264 19316 25304
rect 19852 25264 19892 25304
rect 20236 25264 20276 25304
rect 5068 25180 5108 25220
rect 13900 25180 13940 25220
rect 16204 25180 16244 25220
rect 17260 25180 17300 25220
rect 19372 25180 19412 25220
rect 2668 25096 2708 25136
rect 5356 25096 5396 25136
rect 8044 25096 8084 25136
rect 11308 25096 11348 25136
rect 4928 24928 4968 24968
rect 5010 24928 5050 24968
rect 5092 24928 5132 24968
rect 5174 24928 5214 24968
rect 5256 24928 5296 24968
rect 20048 24928 20088 24968
rect 20130 24928 20170 24968
rect 20212 24928 20252 24968
rect 20294 24928 20334 24968
rect 20376 24928 20416 24968
rect 6700 24760 6740 24800
rect 9484 24760 9524 24800
rect 19468 24760 19508 24800
rect 3148 24676 3188 24716
rect 4780 24676 4820 24716
rect 12076 24676 12116 24716
rect 17932 24676 17972 24716
rect 18604 24676 18644 24716
rect 1420 24592 1460 24632
rect 2668 24592 2708 24632
rect 3052 24592 3092 24632
rect 3436 24592 3476 24632
rect 3820 24592 3860 24632
rect 3916 24592 3956 24632
rect 4012 24592 4052 24632
rect 4108 24592 4148 24632
rect 4378 24607 4418 24647
rect 4684 24592 4724 24632
rect 5260 24592 5300 24632
rect 5356 24592 5396 24632
rect 5548 24592 5588 24632
rect 5740 24592 5780 24632
rect 5932 24592 5972 24632
rect 6316 24592 6356 24632
rect 6508 24592 6548 24632
rect 6892 24592 6932 24632
rect 8140 24592 8180 24632
rect 8524 24592 8564 24632
rect 8812 24592 8852 24632
rect 8908 24592 8948 24632
rect 9422 24577 9462 24617
rect 9580 24592 9620 24632
rect 9676 24592 9716 24632
rect 9868 24592 9908 24632
rect 9964 24592 10004 24632
rect 10348 24592 10388 24632
rect 10444 24592 10484 24632
rect 10924 24592 10964 24632
rect 11404 24592 11444 24632
rect 11884 24578 11924 24618
rect 13036 24592 13076 24632
rect 14860 24592 14900 24632
rect 16108 24592 16148 24632
rect 16492 24592 16532 24632
rect 17740 24592 17780 24632
rect 18202 24607 18242 24647
rect 18508 24592 18548 24632
rect 5836 24508 5876 24548
rect 14284 24550 14324 24590
rect 19118 24577 19158 24617
rect 19276 24592 19316 24632
rect 19372 24592 19412 24632
rect 19564 24592 19604 24632
rect 19660 24592 19700 24632
rect 10828 24508 10868 24548
rect 19852 24508 19892 24548
rect 2860 24424 2900 24464
rect 3436 24424 3476 24464
rect 5068 24424 5108 24464
rect 6508 24424 6548 24464
rect 9196 24424 9236 24464
rect 18892 24424 18932 24464
rect 20044 24424 20084 24464
rect 3628 24340 3668 24380
rect 5548 24340 5588 24380
rect 6700 24340 6740 24380
rect 14476 24340 14516 24380
rect 16300 24340 16340 24380
rect 3688 24172 3728 24212
rect 3770 24172 3810 24212
rect 3852 24172 3892 24212
rect 3934 24172 3974 24212
rect 4016 24172 4056 24212
rect 18808 24172 18848 24212
rect 18890 24172 18930 24212
rect 18972 24172 19012 24212
rect 19054 24172 19094 24212
rect 19136 24172 19176 24212
rect 8332 23920 8372 23960
rect 8716 23920 8756 23960
rect 8908 23920 8948 23960
rect 12364 23920 12404 23960
rect 18796 23920 18836 23960
rect 20236 23920 20276 23960
rect 1612 23836 1652 23876
rect 6412 23836 6452 23876
rect 10924 23836 10964 23876
rect 19756 23836 19796 23876
rect 1900 23752 1940 23792
rect 2476 23752 2516 23792
rect 2572 23752 2612 23792
rect 2956 23752 2996 23792
rect 3052 23752 3092 23792
rect 3532 23752 3572 23792
rect 4012 23766 4052 23806
rect 4492 23752 4532 23792
rect 4588 23752 4628 23792
rect 4972 23752 5012 23792
rect 5068 23752 5108 23792
rect 5548 23752 5588 23792
rect 6076 23761 6116 23801
rect 6508 23752 6548 23792
rect 6892 23752 6932 23792
rect 8140 23752 8180 23792
rect 8524 23752 8564 23792
rect 8716 23752 8756 23792
rect 9196 23752 9236 23792
rect 9292 23752 9332 23792
rect 9580 23752 9620 23792
rect 9868 23752 9908 23792
rect 9964 23752 10004 23792
rect 10156 23752 10196 23792
rect 10444 23752 10484 23792
rect 10540 23752 10580 23792
rect 11020 23752 11060 23792
rect 11500 23752 11540 23792
rect 11980 23766 12020 23806
rect 12556 23752 12596 23792
rect 13804 23752 13844 23792
rect 14476 23752 14516 23792
rect 14572 23752 14612 23792
rect 14956 23752 14996 23792
rect 16060 23794 16100 23834
rect 15052 23752 15092 23792
rect 15532 23752 15572 23792
rect 16588 23752 16628 23792
rect 17836 23752 17876 23792
rect 18124 23752 18164 23792
rect 18412 23752 18452 23792
rect 19022 23767 19062 23807
rect 19180 23752 19220 23792
rect 19276 23752 19316 23792
rect 19468 23752 19508 23792
rect 19564 23752 19604 23792
rect 20140 23765 20180 23805
rect 4204 23668 4244 23708
rect 18508 23668 18548 23708
rect 1420 23584 1460 23624
rect 2188 23584 2228 23624
rect 6220 23584 6260 23624
rect 10156 23584 10196 23624
rect 12172 23584 12212 23624
rect 16204 23584 16244 23624
rect 16396 23584 16436 23624
rect 19372 23584 19412 23624
rect 19948 23584 19988 23624
rect 4928 23416 4968 23456
rect 5010 23416 5050 23456
rect 5092 23416 5132 23456
rect 5174 23416 5214 23456
rect 5256 23416 5296 23456
rect 20048 23416 20088 23456
rect 20130 23416 20170 23456
rect 20212 23416 20252 23456
rect 20294 23416 20334 23456
rect 20376 23416 20416 23456
rect 1324 23248 1364 23288
rect 3340 23248 3380 23288
rect 3628 23248 3668 23288
rect 4300 23248 4340 23288
rect 6316 23248 6356 23288
rect 10540 23248 10580 23288
rect 10924 23248 10964 23288
rect 18028 23248 18068 23288
rect 11596 23164 11636 23204
rect 12364 23164 12404 23204
rect 14284 23164 14324 23204
rect 16300 23164 16340 23204
rect 1900 23080 1940 23120
rect 3148 23080 3188 23120
rect 3820 23080 3860 23120
rect 4012 23080 4052 23120
rect 4108 23080 4148 23120
rect 4396 23080 4436 23120
rect 4492 23080 4532 23120
rect 4588 23080 4628 23120
rect 4876 23080 4916 23120
rect 6124 23080 6164 23120
rect 6700 23080 6740 23120
rect 7948 23080 7988 23120
rect 8524 23080 8564 23120
rect 8908 23080 8948 23120
rect 9100 23080 9140 23120
rect 10348 23080 10388 23120
rect 10732 23080 10772 23120
rect 10876 23070 10916 23110
rect 11020 23080 11060 23120
rect 11116 23080 11156 23120
rect 11273 23065 11313 23105
rect 11500 23080 11540 23120
rect 11980 23080 12020 23120
rect 12268 23080 12308 23120
rect 12844 23080 12884 23120
rect 14092 23080 14132 23120
rect 14572 23080 14612 23120
rect 14668 23080 14708 23120
rect 15628 23080 15668 23120
rect 16156 23070 16196 23110
rect 16588 23080 16628 23120
rect 17836 23080 17876 23120
rect 18412 23080 18452 23120
rect 19660 23080 19700 23120
rect 20044 23080 20084 23120
rect 20236 23080 20276 23120
rect 1708 22996 1748 23036
rect 8620 22996 8660 23036
rect 8812 22996 8852 23036
rect 15052 22996 15092 23036
rect 15148 22996 15188 23036
rect 20140 22996 20180 23036
rect 3628 22912 3668 22952
rect 8716 22912 8756 22952
rect 19852 22912 19892 22952
rect 1516 22828 1556 22868
rect 3820 22828 3860 22868
rect 8140 22828 8180 22868
rect 12652 22828 12692 22868
rect 18028 22828 18068 22868
rect 3688 22660 3728 22700
rect 3770 22660 3810 22700
rect 3852 22660 3892 22700
rect 3934 22660 3974 22700
rect 4016 22660 4056 22700
rect 18808 22660 18848 22700
rect 18890 22660 18930 22700
rect 18972 22660 19012 22700
rect 19054 22660 19094 22700
rect 19136 22660 19176 22700
rect 10732 22492 10772 22532
rect 11692 22492 11732 22532
rect 20236 22492 20276 22532
rect 3148 22408 3188 22448
rect 4492 22408 4532 22448
rect 4876 22408 4916 22448
rect 8908 22408 8948 22448
rect 18316 22408 18356 22448
rect 3052 22324 3092 22364
rect 3244 22324 3284 22364
rect 4396 22324 4436 22364
rect 4588 22324 4628 22364
rect 5452 22324 5492 22364
rect 6988 22324 7028 22364
rect 7084 22324 7124 22364
rect 8812 22324 8852 22364
rect 9004 22324 9044 22364
rect 11980 22324 12020 22364
rect 1228 22240 1268 22280
rect 2476 22240 2516 22280
rect 2956 22240 2996 22280
rect 3340 22240 3380 22280
rect 3532 22240 3572 22280
rect 3628 22240 3668 22280
rect 3820 22240 3860 22280
rect 3916 22240 3956 22280
rect 4071 22240 4111 22280
rect 4300 22240 4340 22280
rect 4684 22240 4724 22280
rect 6508 22240 6548 22280
rect 6604 22240 6644 22280
rect 7564 22240 7604 22280
rect 8044 22254 8084 22294
rect 8716 22240 8756 22280
rect 9100 22240 9140 22280
rect 9292 22240 9332 22280
rect 10540 22240 10580 22280
rect 11020 22240 11060 22280
rect 11308 22240 11348 22280
rect 11884 22240 11924 22280
rect 13516 22282 13556 22322
rect 12076 22240 12116 22280
rect 12268 22240 12308 22280
rect 14860 22240 14900 22280
rect 16108 22240 16148 22280
rect 16684 22240 16724 22280
rect 16876 22240 16916 22280
rect 17068 22240 17108 22280
rect 17164 22240 17204 22280
rect 17644 22240 17684 22280
rect 17932 22240 17972 22280
rect 18028 22240 18068 22280
rect 18508 22240 18548 22280
rect 19756 22240 19796 22280
rect 20127 22229 20167 22269
rect 5740 22156 5780 22196
rect 11404 22156 11444 22196
rect 19948 22156 19988 22196
rect 2668 22072 2708 22112
rect 3724 22072 3764 22112
rect 5260 22072 5300 22112
rect 6124 22072 6164 22112
rect 8236 22072 8276 22112
rect 8428 22072 8468 22112
rect 10732 22072 10772 22112
rect 13708 22072 13748 22112
rect 16300 22072 16340 22112
rect 16780 22072 16820 22112
rect 17356 22072 17396 22112
rect 20236 22072 20276 22112
rect 4928 21904 4968 21944
rect 5010 21904 5050 21944
rect 5092 21904 5132 21944
rect 5174 21904 5214 21944
rect 5256 21904 5296 21944
rect 20048 21904 20088 21944
rect 20130 21904 20170 21944
rect 20212 21904 20252 21944
rect 20294 21904 20334 21944
rect 20376 21904 20416 21944
rect 3052 21736 3092 21776
rect 3628 21736 3668 21776
rect 6028 21736 6068 21776
rect 9676 21736 9716 21776
rect 16396 21736 16436 21776
rect 18508 21736 18548 21776
rect 8044 21652 8084 21692
rect 11980 21652 12020 21692
rect 13996 21652 14036 21692
rect 1612 21568 1652 21608
rect 2860 21568 2900 21608
rect 4204 21568 4244 21608
rect 4396 21568 4436 21608
rect 4588 21568 4628 21608
rect 5836 21568 5876 21608
rect 6316 21568 6356 21608
rect 6412 21568 6452 21608
rect 6796 21568 6836 21608
rect 6892 21568 6932 21608
rect 7372 21568 7412 21608
rect 7852 21554 7892 21594
rect 8236 21568 8276 21608
rect 9484 21568 9524 21608
rect 9964 21568 10004 21608
rect 10348 21568 10388 21608
rect 10540 21568 10580 21608
rect 11788 21568 11828 21608
rect 12268 21568 12308 21608
rect 12364 21568 12404 21608
rect 12748 21568 12788 21608
rect 12844 21568 12884 21608
rect 13324 21568 13364 21608
rect 13804 21563 13844 21603
rect 14668 21568 14708 21608
rect 14764 21568 14804 21608
rect 15724 21568 15764 21608
rect 16252 21558 16292 21598
rect 16588 21568 16628 21608
rect 17836 21568 17876 21608
rect 18220 21568 18260 21608
rect 18316 21568 18356 21608
rect 18412 21568 18452 21608
rect 18700 21568 18740 21608
rect 19084 21568 19124 21608
rect 19276 21568 19316 21608
rect 19660 21568 19700 21608
rect 19852 21568 19892 21608
rect 19948 21568 19988 21608
rect 20140 21582 20180 21622
rect 1420 21484 1460 21524
rect 3340 21484 3380 21524
rect 3916 21484 3956 21524
rect 10060 21484 10100 21524
rect 10252 21484 10292 21524
rect 15148 21484 15188 21524
rect 15244 21484 15284 21524
rect 18796 21484 18836 21524
rect 18988 21484 19028 21524
rect 19372 21484 19412 21524
rect 19564 21484 19604 21524
rect 3532 21400 3572 21440
rect 4396 21400 4436 21440
rect 10156 21400 10196 21440
rect 18892 21400 18932 21440
rect 19468 21400 19508 21440
rect 19948 21400 19988 21440
rect 1228 21316 1268 21356
rect 18028 21316 18068 21356
rect 3688 21148 3728 21188
rect 3770 21148 3810 21188
rect 3852 21148 3892 21188
rect 3934 21148 3974 21188
rect 4016 21148 4056 21188
rect 18808 21148 18848 21188
rect 18890 21148 18930 21188
rect 18972 21148 19012 21188
rect 19054 21148 19094 21188
rect 19136 21148 19176 21188
rect 6124 20980 6164 21020
rect 7756 20980 7796 21020
rect 14860 20980 14900 21020
rect 15628 20980 15668 21020
rect 17260 20980 17300 21020
rect 2860 20896 2900 20936
rect 3148 20896 3188 20936
rect 3532 20896 3572 20936
rect 4012 20896 4052 20936
rect 3916 20812 3956 20852
rect 4108 20812 4148 20852
rect 15436 20812 15476 20852
rect 1228 20728 1268 20768
rect 2476 20728 2516 20768
rect 3820 20728 3860 20768
rect 4204 20728 4244 20768
rect 4396 20728 4436 20768
rect 4684 20728 4724 20768
rect 5932 20728 5972 20768
rect 6316 20728 6356 20768
rect 7564 20728 7604 20768
rect 9388 20728 9428 20768
rect 10636 20728 10676 20768
rect 11020 20728 11060 20768
rect 12268 20728 12308 20768
rect 13420 20728 13460 20768
rect 14668 20728 14708 20768
rect 15820 20728 15860 20768
rect 17068 20728 17108 20768
rect 17452 20728 17492 20768
rect 17548 20728 17588 20768
rect 17644 20728 17684 20768
rect 17740 20728 17780 20768
rect 17932 20728 17972 20768
rect 18124 20728 18164 20768
rect 18316 20728 18356 20768
rect 19564 20728 19604 20768
rect 19948 20728 19988 20768
rect 20140 20770 20180 20810
rect 20044 20728 20084 20768
rect 2668 20644 2708 20684
rect 19756 20644 19796 20684
rect 4492 20560 4532 20600
rect 10828 20560 10868 20600
rect 12460 20560 12500 20600
rect 18028 20560 18068 20600
rect 20236 20560 20276 20600
rect 4928 20392 4968 20432
rect 5010 20392 5050 20432
rect 5092 20392 5132 20432
rect 5174 20392 5214 20432
rect 5256 20392 5296 20432
rect 20048 20392 20088 20432
rect 20130 20392 20170 20432
rect 20212 20392 20252 20432
rect 20294 20392 20334 20432
rect 20376 20392 20416 20432
rect 19948 20224 19988 20264
rect 3724 20140 3764 20180
rect 8044 20140 8084 20180
rect 11020 20140 11060 20180
rect 13996 20140 14036 20180
rect 1228 20056 1268 20096
rect 2476 20056 2516 20096
rect 2860 20056 2900 20096
rect 3340 20056 3380 20096
rect 3628 20056 3668 20096
rect 4588 20056 4628 20096
rect 5836 20056 5876 20096
rect 6316 20056 6356 20096
rect 6412 20056 6452 20096
rect 7372 20056 7412 20096
rect 4396 19972 4436 20012
rect 6796 19972 6836 20012
rect 6892 19972 6932 20012
rect 7900 20014 7940 20054
rect 9292 20056 9332 20096
rect 9388 20056 9428 20096
rect 10348 20056 10388 20096
rect 10828 20051 10868 20091
rect 12268 20056 12308 20096
rect 12364 20056 12404 20096
rect 13324 20056 13364 20096
rect 13804 20042 13844 20082
rect 14380 20056 14420 20096
rect 15628 20056 15668 20096
rect 15820 20056 15860 20096
rect 17068 20035 17108 20075
rect 17644 20056 17684 20096
rect 18892 20056 18932 20096
rect 19276 20056 19316 20096
rect 19372 20056 19412 20096
rect 19468 20056 19508 20096
rect 19564 20056 19604 20096
rect 19756 20071 19796 20111
rect 19852 20056 19892 20096
rect 20044 20056 20084 20096
rect 9772 19972 9812 20012
rect 9868 19972 9908 20012
rect 12748 19972 12788 20012
rect 12844 19972 12884 20012
rect 4012 19888 4052 19928
rect 2668 19804 2708 19844
rect 2956 19804 2996 19844
rect 4204 19804 4244 19844
rect 6028 19804 6068 19844
rect 14188 19804 14228 19844
rect 17260 19804 17300 19844
rect 19084 19804 19124 19844
rect 3688 19636 3728 19676
rect 3770 19636 3810 19676
rect 3852 19636 3892 19676
rect 3934 19636 3974 19676
rect 4016 19636 4056 19676
rect 18808 19636 18848 19676
rect 18890 19636 18930 19676
rect 18972 19636 19012 19676
rect 19054 19636 19094 19676
rect 19136 19636 19176 19676
rect 5260 19468 5300 19508
rect 19660 19468 19700 19508
rect 3628 19384 3668 19424
rect 7660 19384 7700 19424
rect 16684 19384 16724 19424
rect 17452 19384 17492 19424
rect 1516 19300 1556 19340
rect 7564 19300 7604 19340
rect 7756 19300 7796 19340
rect 13900 19300 13940 19340
rect 1708 19216 1748 19256
rect 2956 19216 2996 19256
rect 3340 19216 3380 19256
rect 3436 19216 3476 19256
rect 3628 19216 3668 19256
rect 3820 19216 3860 19256
rect 5068 19216 5108 19256
rect 5548 19216 5588 19256
rect 5644 19216 5684 19256
rect 6028 19216 6068 19256
rect 6124 19216 6164 19256
rect 6604 19216 6644 19256
rect 7084 19230 7124 19270
rect 7468 19216 7508 19256
rect 7852 19216 7892 19256
rect 9100 19216 9140 19256
rect 9196 19216 9236 19256
rect 9580 19216 9620 19256
rect 9676 19216 9716 19256
rect 10156 19216 10196 19256
rect 10684 19225 10724 19265
rect 11596 19216 11636 19256
rect 12844 19216 12884 19256
rect 13324 19216 13364 19256
rect 13420 19216 13460 19256
rect 13804 19216 13844 19256
rect 14380 19216 14420 19256
rect 14860 19230 14900 19270
rect 15244 19216 15284 19256
rect 16492 19216 16532 19256
rect 17068 19216 17108 19256
rect 17164 19224 17204 19264
rect 17260 19216 17300 19256
rect 17452 19216 17492 19256
rect 17644 19216 17684 19256
rect 17740 19216 17780 19256
rect 18220 19216 18260 19256
rect 19468 19216 19508 19256
rect 19852 19216 19892 19256
rect 19948 19216 19988 19256
rect 20140 19227 20180 19267
rect 3148 19132 3188 19172
rect 10828 19132 10868 19172
rect 13036 19132 13076 19172
rect 1324 19048 1364 19088
rect 7276 19048 7316 19088
rect 15052 19048 15092 19088
rect 16972 19048 17012 19088
rect 20044 19048 20084 19088
rect 4928 18880 4968 18920
rect 5010 18880 5050 18920
rect 5092 18880 5132 18920
rect 5174 18880 5214 18920
rect 5256 18880 5296 18920
rect 20048 18880 20088 18920
rect 20130 18880 20170 18920
rect 20212 18880 20252 18920
rect 20294 18880 20334 18920
rect 20376 18880 20416 18920
rect 3916 18712 3956 18752
rect 5644 18712 5684 18752
rect 7564 18712 7604 18752
rect 9196 18712 9236 18752
rect 10828 18712 10868 18752
rect 14092 18712 14132 18752
rect 14956 18712 14996 18752
rect 20044 18712 20084 18752
rect 3340 18628 3380 18668
rect 15532 18628 15572 18668
rect 1228 18544 1268 18584
rect 2476 18544 2516 18584
rect 2956 18544 2996 18584
rect 3244 18544 3284 18584
rect 3820 18544 3860 18584
rect 4012 18544 4052 18584
rect 4204 18544 4244 18584
rect 5452 18544 5492 18584
rect 6124 18544 6164 18584
rect 7372 18544 7412 18584
rect 7756 18544 7796 18584
rect 9004 18544 9044 18584
rect 9388 18544 9428 18584
rect 10636 18544 10676 18584
rect 11020 18544 11060 18584
rect 12268 18544 12308 18584
rect 12652 18544 12692 18584
rect 15148 18544 15188 18584
rect 13900 18502 13940 18542
rect 15340 18544 15380 18584
rect 15724 18539 15764 18579
rect 16204 18544 16244 18584
rect 17164 18544 17204 18584
rect 17260 18544 17300 18584
rect 17548 18544 17588 18584
rect 17644 18544 17684 18584
rect 17740 18544 17780 18584
rect 17836 18544 17876 18584
rect 18316 18544 18356 18584
rect 18412 18544 18452 18584
rect 19372 18544 19412 18584
rect 19852 18539 19892 18579
rect 14764 18460 14804 18500
rect 16684 18460 16724 18500
rect 16780 18460 16820 18500
rect 18796 18460 18836 18500
rect 18892 18460 18932 18500
rect 3628 18376 3668 18416
rect 2668 18292 2708 18332
rect 12460 18292 12500 18332
rect 15340 18292 15380 18332
rect 3688 18124 3728 18164
rect 3770 18124 3810 18164
rect 3852 18124 3892 18164
rect 3934 18124 3974 18164
rect 4016 18124 4056 18164
rect 18808 18124 18848 18164
rect 18890 18124 18930 18164
rect 18972 18124 19012 18164
rect 19054 18124 19094 18164
rect 19136 18124 19176 18164
rect 14956 17956 14996 17996
rect 15628 17956 15668 17996
rect 20236 17956 20276 17996
rect 3916 17872 3956 17912
rect 7756 17872 7796 17912
rect 1228 17788 1268 17828
rect 6316 17788 6356 17828
rect 6412 17788 6452 17828
rect 7948 17788 7988 17828
rect 11308 17788 11348 17828
rect 11404 17788 11444 17828
rect 1516 17704 1556 17744
rect 2764 17704 2804 17744
rect 3244 17704 3284 17744
rect 3532 17704 3572 17744
rect 3628 17704 3668 17744
rect 4108 17704 4148 17744
rect 5356 17704 5396 17744
rect 5836 17704 5876 17744
rect 5932 17704 5972 17744
rect 6892 17704 6932 17744
rect 7372 17709 7412 17749
rect 8332 17704 8372 17744
rect 8428 17704 8468 17744
rect 8812 17704 8852 17744
rect 8908 17704 8948 17744
rect 9388 17704 9428 17744
rect 9868 17709 9908 17749
rect 10828 17704 10868 17744
rect 12412 17746 12452 17786
rect 13612 17788 13652 17828
rect 15148 17788 15188 17828
rect 18124 17788 18164 17828
rect 10924 17704 10964 17744
rect 11884 17704 11924 17744
rect 13036 17704 13076 17744
rect 13132 17704 13172 17744
rect 13516 17704 13556 17744
rect 14092 17704 14132 17744
rect 14620 17713 14660 17753
rect 15820 17704 15860 17744
rect 17068 17704 17108 17744
rect 17260 17704 17300 17744
rect 17356 17704 17396 17744
rect 17548 17704 17588 17744
rect 17932 17704 17972 17744
rect 18220 17704 18260 17744
rect 18412 17704 18452 17744
rect 19660 17704 19700 17744
rect 20044 17704 20084 17744
rect 20236 17704 20276 17744
rect 5548 17620 5588 17660
rect 7564 17620 7604 17660
rect 10060 17620 10100 17660
rect 14764 17620 14804 17660
rect 2956 17536 2996 17576
rect 12556 17536 12596 17576
rect 17452 17536 17492 17576
rect 19852 17536 19892 17576
rect 4928 17368 4968 17408
rect 5010 17368 5050 17408
rect 5092 17368 5132 17408
rect 5174 17368 5214 17408
rect 5256 17368 5296 17408
rect 20048 17368 20088 17408
rect 20130 17368 20170 17408
rect 20212 17368 20252 17408
rect 20294 17368 20334 17408
rect 20376 17368 20416 17408
rect 5836 17200 5876 17240
rect 8044 17200 8084 17240
rect 9676 17200 9716 17240
rect 9964 17200 10004 17240
rect 13132 17200 13172 17240
rect 14764 17200 14804 17240
rect 3436 17116 3476 17156
rect 17356 17116 17396 17156
rect 1804 17032 1844 17072
rect 3052 17032 3092 17072
rect 3628 17018 3668 17058
rect 4108 17032 4148 17072
rect 4588 17032 4628 17072
rect 5068 17032 5108 17072
rect 5164 17032 5204 17072
rect 5489 17032 5529 17072
rect 5644 17032 5684 17072
rect 5740 17032 5780 17072
rect 5932 17032 5972 17072
rect 6028 17032 6068 17072
rect 6220 17032 6260 17072
rect 6412 17032 6452 17072
rect 6604 17032 6644 17072
rect 7852 17032 7892 17072
rect 8236 17032 8276 17072
rect 9484 17032 9524 17072
rect 11692 17032 11732 17072
rect 12940 17032 12980 17072
rect 13324 17032 13364 17072
rect 14572 17032 14612 17072
rect 14956 17032 14996 17072
rect 16204 17032 16244 17072
rect 16780 17032 16820 17072
rect 17068 17032 17108 17072
rect 17260 17032 17300 17072
rect 17452 17032 17492 17072
rect 17644 17032 17684 17072
rect 17836 17032 17876 17072
rect 18124 17032 18164 17072
rect 19372 17032 19412 17072
rect 19756 17032 19796 17072
rect 20044 17032 20084 17072
rect 1612 16948 1652 16988
rect 4684 16948 4724 16988
rect 9868 16864 9908 16904
rect 17068 16864 17108 16904
rect 1420 16780 1460 16820
rect 3244 16780 3284 16820
rect 6412 16780 6452 16820
rect 16396 16780 16436 16820
rect 17644 16780 17684 16820
rect 19564 16780 19604 16820
rect 19756 16780 19796 16820
rect 3688 16612 3728 16652
rect 3770 16612 3810 16652
rect 3852 16612 3892 16652
rect 3934 16612 3974 16652
rect 4016 16612 4056 16652
rect 18808 16612 18848 16652
rect 18890 16612 18930 16652
rect 18972 16612 19012 16652
rect 19054 16612 19094 16652
rect 19136 16612 19176 16652
rect 2380 16444 2420 16484
rect 1420 16276 1460 16316
rect 4780 16276 4820 16316
rect 8044 16276 8084 16316
rect 9100 16276 9140 16316
rect 9484 16276 9524 16316
rect 10540 16276 10580 16316
rect 1708 16192 1748 16232
rect 1996 16192 2036 16232
rect 2092 16192 2132 16232
rect 2764 16206 2804 16246
rect 3244 16192 3284 16232
rect 3724 16192 3764 16232
rect 3820 16192 3860 16232
rect 4204 16192 4244 16232
rect 4300 16192 4340 16232
rect 5068 16192 5108 16232
rect 5260 16192 5300 16232
rect 6508 16192 6548 16232
rect 7084 16197 7124 16237
rect 7564 16192 7604 16232
rect 8140 16192 8180 16232
rect 8524 16192 8564 16232
rect 8620 16192 8660 16232
rect 9964 16192 10004 16232
rect 10060 16192 10100 16232
rect 11548 16234 11588 16274
rect 13996 16276 14036 16316
rect 16684 16276 16724 16316
rect 10444 16192 10484 16232
rect 11020 16192 11060 16232
rect 13516 16192 13556 16232
rect 13612 16192 13652 16232
rect 14092 16192 14132 16232
rect 14572 16192 14612 16232
rect 15100 16201 15140 16241
rect 15676 16201 15716 16241
rect 16204 16192 16244 16232
rect 16780 16192 16820 16232
rect 17164 16192 17204 16232
rect 17260 16192 17300 16232
rect 17548 16192 17588 16232
rect 18796 16192 18836 16232
rect 19180 16192 19220 16232
rect 19276 16192 19316 16232
rect 19660 16192 19700 16232
rect 19852 16192 19892 16232
rect 19948 16192 19988 16232
rect 6700 16108 6740 16148
rect 1228 16024 1268 16064
rect 2572 16024 2612 16064
rect 4588 16024 4628 16064
rect 4972 16024 5012 16064
rect 6892 16024 6932 16064
rect 8908 16024 8948 16064
rect 9292 16024 9332 16064
rect 11692 16024 11732 16064
rect 15244 16024 15284 16064
rect 15532 16024 15572 16064
rect 18988 16024 19028 16064
rect 19468 16024 19508 16064
rect 19756 16024 19796 16064
rect 4928 15856 4968 15896
rect 5010 15856 5050 15896
rect 5092 15856 5132 15896
rect 5174 15856 5214 15896
rect 5256 15856 5296 15896
rect 20048 15856 20088 15896
rect 20130 15856 20170 15896
rect 20212 15856 20252 15896
rect 20294 15856 20334 15896
rect 20376 15856 20416 15896
rect 4204 15688 4244 15728
rect 5836 15688 5876 15728
rect 7468 15688 7508 15728
rect 9676 15688 9716 15728
rect 9868 15688 9908 15728
rect 11692 15688 11732 15728
rect 15148 15688 15188 15728
rect 15628 15688 15668 15728
rect 18796 15692 18836 15732
rect 2284 15520 2324 15560
rect 2380 15520 2420 15560
rect 2476 15520 2516 15560
rect 2572 15520 2612 15560
rect 2764 15520 2804 15560
rect 4012 15520 4052 15560
rect 4396 15520 4436 15560
rect 5644 15520 5684 15560
rect 6028 15520 6068 15560
rect 7276 15520 7316 15560
rect 7660 15520 7700 15560
rect 7948 15520 7988 15560
rect 8236 15520 8276 15560
rect 9484 15520 9524 15560
rect 10252 15520 10292 15560
rect 11500 15520 11540 15560
rect 11980 15520 12020 15560
rect 13228 15520 13268 15560
rect 13708 15520 13748 15560
rect 14956 15520 14996 15560
rect 15820 15520 15860 15560
rect 17068 15520 17108 15560
rect 17356 15520 17396 15560
rect 17452 15520 17492 15560
rect 17548 15520 17588 15560
rect 17644 15520 17684 15560
rect 17836 15520 17876 15560
rect 18124 15520 18164 15560
rect 18604 15520 18644 15560
rect 18700 15520 18740 15560
rect 19084 15520 19124 15560
rect 19372 15520 19412 15560
rect 19468 15520 19508 15560
rect 19948 15520 19988 15560
rect 20140 15562 20180 15602
rect 20236 15520 20276 15560
rect 1708 15436 1748 15476
rect 2092 15436 2132 15476
rect 1324 15352 1364 15392
rect 1516 15352 1556 15392
rect 13420 15352 13460 15392
rect 19756 15352 19796 15392
rect 1900 15268 1940 15308
rect 7660 15268 7700 15308
rect 18124 15268 18164 15308
rect 18316 15268 18356 15308
rect 19948 15268 19988 15308
rect 3688 15100 3728 15140
rect 3770 15100 3810 15140
rect 3852 15100 3892 15140
rect 3934 15100 3974 15140
rect 4016 15100 4056 15140
rect 18808 15100 18848 15140
rect 18890 15100 18930 15140
rect 18972 15100 19012 15140
rect 19054 15100 19094 15140
rect 19136 15100 19176 15140
rect 2668 14932 2708 14972
rect 6028 14932 6068 14972
rect 7660 14932 7700 14972
rect 9868 14848 9908 14888
rect 18892 14848 18932 14888
rect 19756 14848 19796 14888
rect 3052 14764 3092 14804
rect 3916 14764 3956 14804
rect 4012 14764 4052 14804
rect 12556 14764 12596 14804
rect 12652 14764 12692 14804
rect 18796 14764 18836 14804
rect 18988 14764 19028 14804
rect 1228 14680 1268 14720
rect 2476 14680 2516 14720
rect 3436 14680 3476 14720
rect 3532 14680 3572 14720
rect 4492 14680 4532 14720
rect 4972 14685 5012 14725
rect 5548 14680 5588 14720
rect 5644 14680 5684 14720
rect 5740 14680 5780 14720
rect 5932 14680 5972 14720
rect 6220 14680 6260 14720
rect 7468 14680 7508 14720
rect 7948 14680 7988 14720
rect 8044 14680 8084 14720
rect 8428 14680 8468 14720
rect 8524 14680 8564 14720
rect 9004 14680 9044 14720
rect 9484 14685 9524 14725
rect 10348 14680 10388 14720
rect 11596 14680 11636 14720
rect 12076 14680 12116 14720
rect 12172 14680 12212 14720
rect 13132 14680 13172 14720
rect 13612 14685 13652 14725
rect 15628 14685 15668 14725
rect 16108 14680 16148 14720
rect 16588 14680 16628 14720
rect 16684 14680 16724 14720
rect 17068 14680 17108 14720
rect 17164 14680 17204 14720
rect 17740 14680 17780 14720
rect 17836 14680 17876 14720
rect 17932 14680 17972 14720
rect 18220 14680 18260 14720
rect 18316 14680 18356 14720
rect 18412 14680 18452 14720
rect 18700 14680 18740 14720
rect 19084 14680 19124 14720
rect 19276 14680 19316 14720
rect 19372 14680 19412 14720
rect 19468 14680 19508 14720
rect 19564 14680 19604 14720
rect 5164 14596 5204 14636
rect 19756 14638 19796 14678
rect 19948 14680 19988 14720
rect 20044 14680 20084 14720
rect 2860 14512 2900 14552
rect 5452 14512 5492 14552
rect 9676 14512 9716 14552
rect 11788 14512 11828 14552
rect 13804 14512 13844 14552
rect 15436 14512 15476 14552
rect 18028 14512 18068 14552
rect 18508 14512 18548 14552
rect 4928 14344 4968 14384
rect 5010 14344 5050 14384
rect 5092 14344 5132 14384
rect 5174 14344 5214 14384
rect 5256 14344 5296 14384
rect 20048 14344 20088 14384
rect 20130 14344 20170 14384
rect 20212 14344 20252 14384
rect 20294 14344 20334 14384
rect 20376 14344 20416 14384
rect 1228 14176 1268 14216
rect 9196 14176 9236 14216
rect 11212 14176 11252 14216
rect 11404 14176 11444 14216
rect 16204 14176 16244 14216
rect 1708 14092 1748 14132
rect 2380 14092 2420 14132
rect 2572 14092 2612 14132
rect 7468 14092 7508 14132
rect 14380 14092 14420 14132
rect 16012 14092 16052 14132
rect 20140 14092 20180 14132
rect 1612 14008 1652 14048
rect 1804 14008 1844 14048
rect 1900 14008 1940 14048
rect 2092 14008 2132 14048
rect 2188 13966 2228 14006
rect 2284 14000 2324 14040
rect 2764 13994 2804 14034
rect 3244 14008 3284 14048
rect 3820 14008 3860 14048
rect 4204 14008 4244 14048
rect 4300 14008 4340 14048
rect 4684 14008 4724 14048
rect 4780 14008 4820 14048
rect 4972 14008 5012 14048
rect 5164 14008 5204 14048
rect 5260 14008 5300 14048
rect 5356 14008 5396 14048
rect 5452 14008 5492 14048
rect 5740 14008 5780 14048
rect 5836 14008 5876 14048
rect 6796 14008 6836 14048
rect 7276 14003 7316 14043
rect 7756 14008 7796 14048
rect 9004 14008 9044 14048
rect 9484 14008 9524 14048
rect 9580 14008 9620 14048
rect 9964 14008 10004 14048
rect 10060 14008 10100 14048
rect 10540 14008 10580 14048
rect 11068 13998 11108 14038
rect 12652 14008 12692 14048
rect 12748 14008 12788 14048
rect 13132 14008 13172 14048
rect 13708 14008 13748 14048
rect 14188 13994 14228 14034
rect 14572 14008 14612 14048
rect 15820 14008 15860 14048
rect 16396 14008 16436 14048
rect 17644 14008 17684 14048
rect 17836 14008 17876 14048
rect 19084 14008 19124 14048
rect 19468 14008 19508 14048
rect 19852 14008 19892 14048
rect 20044 14008 20084 14048
rect 20236 14008 20276 14048
rect 1420 13924 1460 13964
rect 3724 13924 3764 13964
rect 6220 13924 6260 13964
rect 6316 13924 6356 13964
rect 11596 13924 11636 13964
rect 11980 13924 12020 13964
rect 12364 13924 12404 13964
rect 13228 13924 13268 13964
rect 19564 13924 19604 13964
rect 19756 13924 19796 13964
rect 11788 13840 11828 13880
rect 12172 13840 12212 13880
rect 19276 13840 19316 13880
rect 19660 13840 19700 13880
rect 4972 13756 5012 13796
rect 3688 13588 3728 13628
rect 3770 13588 3810 13628
rect 3852 13588 3892 13628
rect 3934 13588 3974 13628
rect 4016 13588 4056 13628
rect 18808 13588 18848 13628
rect 18890 13588 18930 13628
rect 18972 13588 19012 13628
rect 19054 13588 19094 13628
rect 19136 13588 19176 13628
rect 1228 13420 1268 13460
rect 3148 13420 3188 13460
rect 5740 13420 5780 13460
rect 7372 13420 7412 13460
rect 9580 13420 9620 13460
rect 11308 13420 11348 13460
rect 13420 13420 13460 13460
rect 18604 13420 18644 13460
rect 19852 13336 19892 13376
rect 1420 13252 1460 13292
rect 3532 13263 3572 13303
rect 3916 13252 3956 13292
rect 11692 13252 11732 13292
rect 1708 13168 1748 13208
rect 2956 13168 2996 13208
rect 4300 13168 4340 13208
rect 5548 13168 5588 13208
rect 5932 13168 5972 13208
rect 7180 13168 7220 13208
rect 7564 13168 7604 13208
rect 13228 13210 13268 13250
rect 7756 13168 7796 13208
rect 7852 13168 7892 13208
rect 8140 13168 8180 13208
rect 9388 13168 9428 13208
rect 9868 13168 9908 13208
rect 11116 13168 11156 13208
rect 11980 13168 12020 13208
rect 13804 13168 13844 13208
rect 15052 13168 15092 13208
rect 15244 13168 15284 13208
rect 16492 13168 16532 13208
rect 17164 13168 17204 13208
rect 18412 13168 18452 13208
rect 19180 13168 19220 13208
rect 19468 13168 19508 13208
rect 19564 13168 19604 13208
rect 20044 13168 20084 13208
rect 20236 13168 20276 13208
rect 13612 13084 13652 13124
rect 20140 13084 20180 13124
rect 3340 13000 3380 13040
rect 3724 13000 3764 13040
rect 7660 13000 7700 13040
rect 11500 13000 11540 13040
rect 16684 13000 16724 13040
rect 4928 12832 4968 12872
rect 5010 12832 5050 12872
rect 5092 12832 5132 12872
rect 5174 12832 5214 12872
rect 5256 12832 5296 12872
rect 20048 12832 20088 12872
rect 20130 12832 20170 12872
rect 20212 12832 20252 12872
rect 20294 12832 20334 12872
rect 20376 12832 20416 12872
rect 18892 12722 18932 12762
rect 2668 12664 2708 12704
rect 19564 12664 19604 12704
rect 2860 12580 2900 12620
rect 5452 12580 5492 12620
rect 9772 12580 9812 12620
rect 12556 12580 12596 12620
rect 15244 12580 15284 12620
rect 17260 12580 17300 12620
rect 1228 12496 1268 12536
rect 2476 12496 2516 12536
rect 3052 12482 3092 12522
rect 3532 12496 3572 12536
rect 4012 12496 4052 12536
rect 4108 12496 4148 12536
rect 4492 12496 4532 12536
rect 4588 12496 4628 12536
rect 4876 12496 4916 12536
rect 5068 12507 5108 12547
rect 5260 12496 5300 12536
rect 5356 12496 5396 12536
rect 5548 12496 5588 12536
rect 6220 12496 6260 12536
rect 7468 12496 7508 12536
rect 8044 12496 8084 12536
rect 9292 12496 9332 12536
rect 9868 12496 9908 12536
rect 10156 12487 10196 12527
rect 10444 12496 10484 12536
rect 10636 12496 10676 12536
rect 10732 12496 10772 12536
rect 11116 12496 11156 12536
rect 12364 12496 12404 12536
rect 12748 12496 12788 12536
rect 13996 12496 14036 12536
rect 14860 12496 14900 12536
rect 15052 12496 15092 12536
rect 15436 12491 15476 12531
rect 15916 12496 15956 12536
rect 16876 12496 16916 12536
rect 16972 12496 17012 12536
rect 17452 12496 17492 12536
rect 18700 12496 18740 12536
rect 18988 12496 19028 12536
rect 19084 12496 19124 12536
rect 19756 12496 19796 12536
rect 19852 12496 19892 12536
rect 5932 12412 5972 12452
rect 14668 12412 14708 12452
rect 16396 12412 16436 12452
rect 16492 12412 16532 12452
rect 20236 12412 20276 12452
rect 7852 12328 7892 12368
rect 9484 12328 9524 12368
rect 19372 12328 19412 12368
rect 5068 12244 5108 12284
rect 5740 12244 5780 12284
rect 7660 12244 7700 12284
rect 10444 12244 10484 12284
rect 14188 12244 14228 12284
rect 14476 12244 14516 12284
rect 14860 12244 14900 12284
rect 20044 12244 20084 12284
rect 3688 12076 3728 12116
rect 3770 12076 3810 12116
rect 3852 12076 3892 12116
rect 3934 12076 3974 12116
rect 4016 12076 4056 12116
rect 18808 12076 18848 12116
rect 18890 12076 18930 12116
rect 18972 12076 19012 12116
rect 19054 12076 19094 12116
rect 19136 12076 19176 12116
rect 2668 11908 2708 11948
rect 7468 11908 7508 11948
rect 7660 11908 7700 11948
rect 4588 11824 4628 11864
rect 10252 11824 10292 11864
rect 19084 11824 19124 11864
rect 5836 11740 5876 11780
rect 5932 11740 5972 11780
rect 12652 11740 12692 11780
rect 12748 11740 12788 11780
rect 14284 11740 14324 11780
rect 14764 11740 14804 11780
rect 15628 11740 15668 11780
rect 17164 11740 17204 11780
rect 20236 11740 20276 11780
rect 1228 11656 1268 11696
rect 2476 11656 2516 11696
rect 2860 11656 2900 11696
rect 2956 11656 2996 11696
rect 3148 11656 3188 11696
rect 4396 11656 4436 11696
rect 4780 11656 4820 11696
rect 4972 11656 5012 11696
rect 5068 11656 5108 11696
rect 5356 11656 5396 11696
rect 5452 11656 5492 11696
rect 6412 11656 6452 11696
rect 6892 11661 6932 11701
rect 7276 11656 7316 11696
rect 7468 11656 7508 11696
rect 7852 11656 7892 11696
rect 9100 11656 9140 11696
rect 9580 11656 9620 11696
rect 9868 11656 9908 11696
rect 10444 11656 10484 11696
rect 11692 11656 11732 11696
rect 12172 11656 12212 11696
rect 12268 11656 12308 11696
rect 13228 11656 13268 11696
rect 13708 11670 13748 11710
rect 15052 11656 15092 11696
rect 15148 11656 15188 11696
rect 16636 11698 16676 11738
rect 15532 11656 15572 11696
rect 16108 11656 16148 11696
rect 17356 11656 17396 11696
rect 18604 11656 18644 11696
rect 19468 11656 19508 11696
rect 19756 11656 19796 11696
rect 9964 11572 10004 11612
rect 11884 11572 11924 11612
rect 18796 11572 18836 11612
rect 19372 11572 19412 11612
rect 4876 11488 4916 11528
rect 7084 11488 7124 11528
rect 7660 11488 7700 11528
rect 13900 11488 13940 11528
rect 14092 11488 14132 11528
rect 14572 11488 14612 11528
rect 16780 11488 16820 11528
rect 16972 11488 17012 11528
rect 20044 11488 20084 11528
rect 4928 11320 4968 11360
rect 5010 11320 5050 11360
rect 5092 11320 5132 11360
rect 5174 11320 5214 11360
rect 5256 11320 5296 11360
rect 20048 11320 20088 11360
rect 20130 11320 20170 11360
rect 20212 11320 20252 11360
rect 20294 11320 20334 11360
rect 20376 11320 20416 11360
rect 1516 11152 1556 11192
rect 5260 11152 5300 11192
rect 5740 11152 5780 11192
rect 16780 11152 16820 11192
rect 18412 11152 18452 11192
rect 9484 11068 9524 11108
rect 13132 11068 13172 11108
rect 13324 11068 13364 11108
rect 1324 10984 1364 11024
rect 1612 10984 1652 11024
rect 2188 10984 2228 11024
rect 3436 10984 3476 11024
rect 3820 10984 3860 11024
rect 5068 10984 5108 11024
rect 5548 10984 5588 11024
rect 5932 10984 5972 11024
rect 7180 10984 7220 11024
rect 7372 10984 7412 11024
rect 8620 10984 8660 11024
rect 9100 10984 9140 11024
rect 9388 10984 9428 11024
rect 10252 10984 10292 11024
rect 11500 10984 11540 11024
rect 11692 10984 11732 11024
rect 12940 10984 12980 11024
rect 13516 10970 13556 11010
rect 13996 10984 14036 11024
rect 14476 10984 14516 11024
rect 14572 10984 14612 11024
rect 14956 10984 14996 11024
rect 15052 10984 15092 11024
rect 15340 10984 15380 11024
rect 16588 10984 16628 11024
rect 18220 10984 18260 11024
rect 18700 10984 18740 11024
rect 18988 10984 19028 11024
rect 16972 10942 17012 10982
rect 19084 10984 19124 11024
rect 19564 10984 19604 11024
rect 19948 10984 19988 11024
rect 20236 10984 20276 11024
rect 1996 10900 2036 10940
rect 19660 10900 19700 10940
rect 19852 10900 19892 10940
rect 5452 10816 5492 10856
rect 9772 10816 9812 10856
rect 19756 10816 19796 10856
rect 1804 10732 1844 10772
rect 3628 10732 3668 10772
rect 8812 10732 8852 10772
rect 10060 10732 10100 10772
rect 19372 10732 19412 10772
rect 20140 10732 20180 10772
rect 3688 10564 3728 10604
rect 3770 10564 3810 10604
rect 3852 10564 3892 10604
rect 3934 10564 3974 10604
rect 4016 10564 4056 10604
rect 18808 10564 18848 10604
rect 18890 10564 18930 10604
rect 18972 10564 19012 10604
rect 19054 10564 19094 10604
rect 19136 10564 19176 10604
rect 2860 10396 2900 10436
rect 3052 10396 3092 10436
rect 5068 10396 5108 10436
rect 6892 10396 6932 10436
rect 11788 10396 11828 10436
rect 14860 10396 14900 10436
rect 18892 10396 18932 10436
rect 4684 10312 4724 10352
rect 9964 10312 10004 10352
rect 12748 10312 12788 10352
rect 19084 10312 19124 10352
rect 20044 10312 20084 10352
rect 5260 10228 5300 10268
rect 9868 10228 9908 10268
rect 10060 10228 10100 10268
rect 20236 10228 20276 10268
rect 1420 10144 1460 10184
rect 2668 10144 2708 10184
rect 3244 10144 3284 10184
rect 4492 10144 4532 10184
rect 4684 10144 4724 10184
rect 4876 10144 4916 10184
rect 5452 10144 5492 10184
rect 6700 10144 6740 10184
rect 7180 10144 7220 10184
rect 7276 10144 7316 10184
rect 7372 10144 7412 10184
rect 7468 10144 7508 10184
rect 7660 10144 7700 10184
rect 7756 10144 7796 10184
rect 8140 10144 8180 10184
rect 9388 10144 9428 10184
rect 9772 10144 9812 10184
rect 10156 10144 10196 10184
rect 10348 10144 10388 10184
rect 11596 10144 11636 10184
rect 12076 10144 12116 10184
rect 12364 10144 12404 10184
rect 12460 10144 12500 10184
rect 12940 10144 12980 10184
rect 13132 10144 13172 10184
rect 13228 10144 13268 10184
rect 13420 10144 13460 10184
rect 14668 10144 14708 10184
rect 15052 10144 15092 10184
rect 15148 10144 15188 10184
rect 15340 10144 15380 10184
rect 16588 10144 16628 10184
rect 16972 10144 17012 10184
rect 17068 10144 17108 10184
rect 17260 10144 17300 10184
rect 17452 10144 17492 10184
rect 18700 10144 18740 10184
rect 19372 10144 19412 10184
rect 19468 10144 19508 10184
rect 19756 10144 19796 10184
rect 7948 9976 7988 10016
rect 9580 9976 9620 10016
rect 13036 9976 13076 10016
rect 16780 9976 16820 10016
rect 17164 9976 17204 10016
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 3052 9640 3092 9680
rect 13324 9640 13364 9680
rect 16780 9640 16820 9680
rect 17932 9640 17972 9680
rect 3244 9556 3284 9596
rect 7660 9556 7700 9596
rect 1228 9472 1268 9512
rect 1420 9472 1460 9512
rect 1612 9472 1652 9512
rect 2860 9451 2900 9491
rect 3436 9467 3476 9507
rect 3916 9472 3956 9512
rect 4492 9472 4532 9512
rect 4876 9472 4916 9512
rect 4972 9472 5012 9512
rect 5356 9472 5396 9512
rect 5548 9472 5588 9512
rect 5644 9470 5684 9510
rect 5932 9472 5972 9512
rect 6028 9472 6068 9512
rect 6988 9472 7028 9512
rect 7468 9458 7508 9498
rect 7852 9472 7892 9512
rect 8044 9472 8084 9512
rect 8524 9472 8564 9512
rect 8620 9472 8660 9512
rect 8908 9472 8948 9512
rect 9196 9472 9236 9512
rect 10444 9472 10484 9512
rect 10924 9472 10964 9512
rect 11308 9472 11348 9512
rect 11500 9472 11540 9512
rect 12748 9472 12788 9512
rect 13516 9472 13556 9512
rect 14764 9472 14804 9512
rect 15052 9472 15092 9512
rect 15148 9472 15188 9512
rect 16108 9472 16148 9512
rect 16588 9458 16628 9498
rect 16972 9472 17012 9512
rect 17068 9472 17108 9512
rect 17164 9472 17204 9512
rect 17260 9472 17300 9512
rect 17452 9472 17492 9512
rect 17644 9472 17684 9512
rect 17836 9472 17876 9512
rect 18028 9472 18068 9512
rect 18124 9472 18164 9512
rect 18316 9472 18356 9512
rect 19564 9472 19604 9512
rect 19948 9472 19988 9512
rect 20044 9472 20084 9512
rect 20236 9472 20276 9512
rect 4396 9388 4436 9428
rect 6412 9388 6452 9428
rect 6508 9388 6548 9428
rect 11020 9388 11060 9428
rect 8236 9304 8276 9344
rect 11116 9304 11156 9344
rect 11212 9346 11252 9386
rect 15532 9388 15572 9428
rect 15628 9388 15668 9428
rect 1420 9220 1460 9260
rect 5356 9220 5396 9260
rect 7852 9220 7892 9260
rect 10636 9220 10676 9260
rect 12940 9220 12980 9260
rect 17452 9220 17492 9260
rect 19756 9220 19796 9260
rect 20236 9220 20276 9260
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 6796 8884 6836 8924
rect 6988 8884 7028 8924
rect 11596 8884 11636 8924
rect 15052 8884 15092 8924
rect 16684 8884 16724 8924
rect 1228 8800 1268 8840
rect 1612 8800 1652 8840
rect 1996 8800 2036 8840
rect 4396 8800 4436 8840
rect 12556 8800 12596 8840
rect 13036 8800 13076 8840
rect 18220 8800 18260 8840
rect 1420 8716 1460 8756
rect 1804 8716 1844 8756
rect 2188 8703 2228 8743
rect 2956 8716 2996 8756
rect 4577 8727 4617 8767
rect 13420 8716 13460 8756
rect 2476 8632 2516 8672
rect 2572 8632 2612 8672
rect 3052 8632 3092 8672
rect 3532 8632 3572 8672
rect 4012 8637 4052 8677
rect 4972 8632 5012 8672
rect 5164 8632 5204 8672
rect 5356 8632 5396 8672
rect 6604 8632 6644 8672
rect 7180 8632 7220 8672
rect 8428 8632 8468 8672
rect 8716 8632 8756 8672
rect 8812 8611 8852 8651
rect 8908 8632 8948 8672
rect 9004 8632 9044 8672
rect 9292 8632 9332 8672
rect 9388 8632 9428 8672
rect 9772 8632 9812 8672
rect 9868 8632 9908 8672
rect 10348 8632 10388 8672
rect 10828 8646 10868 8686
rect 11308 8617 11348 8657
rect 11404 8632 11444 8672
rect 11596 8632 11636 8672
rect 11884 8632 11924 8672
rect 12172 8632 12212 8672
rect 12748 8632 12788 8672
rect 12844 8632 12884 8672
rect 13036 8632 13076 8672
rect 13612 8632 13652 8672
rect 14860 8632 14900 8672
rect 15244 8632 15284 8672
rect 16492 8632 16532 8672
rect 16876 8632 16916 8672
rect 16972 8611 17012 8651
rect 17068 8632 17108 8672
rect 17356 8632 17396 8672
rect 17644 8632 17684 8672
rect 17836 8632 17876 8672
rect 18028 8632 18068 8672
rect 18604 8632 18644 8672
rect 18892 8632 18932 8672
rect 19180 8632 19220 8672
rect 19372 8632 19412 8672
rect 19468 8632 19508 8672
rect 19660 8632 19700 8672
rect 19756 8611 19796 8651
rect 19852 8632 19892 8672
rect 19948 8632 19988 8672
rect 20127 8621 20167 8661
rect 4204 8548 4244 8588
rect 12268 8548 12308 8588
rect 17164 8548 17204 8588
rect 18508 8548 18548 8588
rect 5068 8464 5108 8504
rect 6796 8464 6836 8504
rect 6988 8464 7028 8504
rect 11020 8464 11060 8504
rect 13228 8464 13268 8504
rect 17452 8464 17492 8504
rect 17932 8464 17972 8504
rect 19276 8464 19316 8504
rect 20236 8464 20276 8504
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 1228 8128 1268 8168
rect 3052 8128 3092 8168
rect 5260 8128 5300 8168
rect 7276 8128 7316 8168
rect 12556 8128 12596 8168
rect 13132 8128 13172 8168
rect 14956 8128 14996 8168
rect 17164 8128 17204 8168
rect 17548 8128 17588 8168
rect 20140 8128 20180 8168
rect 14764 8044 14804 8084
rect 1612 7960 1652 8000
rect 2860 7939 2900 7979
rect 3436 7960 3476 8000
rect 3628 7960 3668 8000
rect 3820 7960 3860 8000
rect 5068 7960 5108 8000
rect 5452 7960 5492 8000
rect 6700 7960 6740 8000
rect 7084 7960 7124 8000
rect 7180 7960 7220 8000
rect 7372 7960 7412 8000
rect 7564 7960 7604 8000
rect 8812 7960 8852 8000
rect 9196 7960 9236 8000
rect 10444 7960 10484 8000
rect 10924 7960 10964 8000
rect 12172 7960 12212 8000
rect 12748 7960 12788 8000
rect 12844 7960 12884 8000
rect 13036 7960 13076 8000
rect 13324 7960 13364 8000
rect 14572 7960 14612 8000
rect 15148 7946 15188 7986
rect 15628 7960 15668 8000
rect 16108 7960 16148 8000
rect 16204 7960 16244 8000
rect 16588 7960 16628 8000
rect 16684 7960 16724 8000
rect 16972 7960 17012 8000
rect 17068 7960 17108 8000
rect 17260 7960 17300 8000
rect 17452 7960 17492 8000
rect 17644 7960 17684 8000
rect 17740 7960 17780 8000
rect 17932 7960 17972 8000
rect 18220 7960 18260 8000
rect 19468 7960 19508 8000
rect 19852 7960 19892 8000
rect 19948 7960 19988 8000
rect 1420 7876 1460 7916
rect 3532 7876 3572 7916
rect 6892 7708 6932 7748
rect 9004 7708 9044 7748
rect 10636 7708 10676 7748
rect 12364 7708 12404 7748
rect 18028 7708 18068 7748
rect 19660 7708 19700 7748
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 2764 7372 2804 7412
rect 5164 7372 5204 7412
rect 14764 7372 14804 7412
rect 20140 7372 20180 7412
rect 18604 7288 18644 7328
rect 19756 7288 19796 7328
rect 3532 7204 3572 7244
rect 10636 7204 10676 7244
rect 10732 7204 10772 7244
rect 12748 7204 12788 7244
rect 17068 7204 17108 7244
rect 19660 7204 19700 7244
rect 19852 7204 19892 7244
rect 1324 7120 1364 7160
rect 2572 7120 2612 7160
rect 3052 7120 3092 7160
rect 3148 7120 3188 7160
rect 3628 7120 3668 7160
rect 4108 7120 4148 7160
rect 4588 7125 4628 7165
rect 4972 7120 5012 7160
rect 5164 7120 5204 7160
rect 5452 7120 5492 7160
rect 5548 7120 5588 7160
rect 5932 7120 5972 7160
rect 6028 7120 6068 7160
rect 6508 7120 6548 7160
rect 6988 7134 7028 7174
rect 7564 7120 7604 7160
rect 8812 7120 8852 7160
rect 9004 7120 9044 7160
rect 9100 7120 9140 7160
rect 9292 7120 9332 7160
rect 9484 7120 9524 7160
rect 9580 7120 9620 7160
rect 9772 7120 9812 7160
rect 10156 7120 10196 7160
rect 10252 7120 10292 7160
rect 11212 7120 11252 7160
rect 11740 7129 11780 7169
rect 12268 7120 12308 7160
rect 12364 7120 12404 7160
rect 12844 7120 12884 7160
rect 13324 7120 13364 7160
rect 13852 7129 13892 7169
rect 14285 7122 14325 7162
rect 14380 7120 14420 7160
rect 14572 7120 14612 7160
rect 14956 7120 14996 7160
rect 16204 7120 16244 7160
rect 16492 7120 16532 7160
rect 16588 7120 16628 7160
rect 16972 7120 17012 7160
rect 17548 7120 17588 7160
rect 18028 7125 18068 7165
rect 18892 7120 18932 7160
rect 18988 7120 19028 7160
rect 19276 7120 19316 7160
rect 19564 7120 19604 7160
rect 19948 7120 19988 7160
rect 20236 7120 20276 7160
rect 7180 7036 7220 7076
rect 9676 7036 9716 7076
rect 11884 7036 11924 7076
rect 13996 7036 14036 7076
rect 4780 6952 4820 6992
rect 7372 6952 7412 6992
rect 9196 6952 9236 6992
rect 14476 6952 14516 6992
rect 18220 6952 18260 6992
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 8428 6674 8468 6714
rect 1228 6616 1268 6656
rect 1612 6616 1652 6656
rect 2092 6616 2132 6656
rect 9388 6658 9428 6698
rect 4204 6616 4244 6656
rect 6508 6616 6548 6656
rect 11884 6616 11924 6656
rect 12076 6616 12116 6656
rect 13900 6616 13940 6656
rect 15820 6616 15860 6656
rect 18508 6616 18548 6656
rect 4396 6532 4436 6572
rect 6892 6532 6932 6572
rect 9100 6532 9140 6572
rect 1996 6448 2036 6488
rect 2188 6448 2228 6488
rect 2380 6448 2420 6488
rect 2572 6448 2612 6488
rect 2764 6448 2804 6488
rect 4012 6448 4052 6488
rect 4588 6434 4628 6474
rect 5068 6448 5108 6488
rect 5548 6448 5588 6488
rect 5644 6448 5684 6488
rect 6028 6448 6068 6488
rect 6124 6448 6164 6488
rect 6412 6448 6452 6488
rect 6604 6448 6644 6488
rect 6700 6448 6740 6488
rect 6988 6448 7028 6488
rect 7084 6448 7124 6488
rect 7180 6448 7220 6488
rect 7372 6448 7412 6488
rect 7756 6448 7796 6488
rect 8236 6448 8276 6488
rect 8332 6448 8372 6488
rect 8716 6448 8756 6488
rect 9004 6448 9044 6488
rect 9580 6448 9620 6488
rect 9868 6448 9908 6488
rect 10060 6448 10100 6488
rect 10252 6447 10292 6487
rect 10444 6448 10484 6488
rect 11692 6448 11732 6488
rect 12460 6448 12500 6488
rect 13708 6448 13748 6488
rect 14092 6448 14132 6488
rect 15340 6448 15380 6488
rect 15724 6448 15764 6488
rect 15916 6448 15956 6488
rect 16108 6448 16148 6488
rect 16300 6448 16340 6488
rect 16396 6448 16436 6488
rect 16972 6448 17012 6488
rect 17260 6448 17300 6488
rect 17356 6448 17396 6488
rect 17836 6448 17876 6488
rect 18028 6448 18068 6488
rect 18124 6448 18164 6488
rect 18316 6448 18356 6488
rect 18412 6448 18452 6488
rect 18604 6437 18644 6477
rect 19188 6448 19228 6488
rect 19468 6448 19508 6488
rect 19564 6448 19604 6488
rect 20044 6448 20084 6488
rect 20236 6448 20276 6488
rect 1420 6364 1460 6404
rect 1804 6364 1844 6404
rect 7468 6364 7508 6404
rect 7660 6364 7700 6404
rect 12268 6364 12308 6404
rect 2380 6280 2420 6320
rect 7564 6280 7604 6320
rect 7948 6280 7988 6320
rect 9580 6280 9620 6320
rect 16588 6280 16628 6320
rect 17644 6280 17684 6320
rect 19852 6280 19892 6320
rect 10060 6196 10100 6236
rect 15532 6196 15572 6236
rect 16108 6196 16148 6236
rect 17836 6196 17876 6236
rect 20044 6196 20084 6236
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 3148 5860 3188 5900
rect 5260 5860 5300 5900
rect 6220 5860 6260 5900
rect 9292 5860 9332 5900
rect 20140 5860 20180 5900
rect 2668 5776 2708 5816
rect 9676 5776 9716 5816
rect 15436 5776 15476 5816
rect 13996 5692 14036 5732
rect 1228 5608 1268 5648
rect 2476 5608 2516 5648
rect 2860 5608 2900 5648
rect 3148 5608 3188 5648
rect 3436 5608 3476 5648
rect 3532 5608 3572 5648
rect 3628 5608 3668 5648
rect 3820 5608 3860 5648
rect 5068 5608 5108 5648
rect 5452 5608 5492 5648
rect 5644 5608 5684 5648
rect 5740 5608 5780 5648
rect 5932 5608 5972 5648
rect 6220 5608 6260 5648
rect 6412 5608 6452 5648
rect 6508 5608 6548 5648
rect 6604 5608 6644 5648
rect 6700 5608 6740 5648
rect 6892 5608 6932 5648
rect 8140 5608 8180 5648
rect 8620 5608 8660 5648
rect 8908 5608 8948 5648
rect 9484 5608 9524 5648
rect 9676 5608 9716 5648
rect 9772 5608 9812 5648
rect 10156 5608 10196 5648
rect 11404 5608 11444 5648
rect 11788 5608 11828 5648
rect 13036 5608 13076 5648
rect 13516 5608 13556 5648
rect 13612 5608 13652 5648
rect 14092 5608 14132 5648
rect 14572 5608 14612 5648
rect 15052 5622 15092 5662
rect 15820 5608 15860 5648
rect 16108 5608 16148 5648
rect 16396 5608 16436 5648
rect 17644 5608 17684 5648
rect 18028 5608 18068 5648
rect 18124 5608 18164 5648
rect 18220 5608 18260 5648
rect 18316 5608 18356 5648
rect 18508 5608 18548 5648
rect 19756 5608 19796 5648
rect 20236 5608 20276 5648
rect 9004 5524 9044 5564
rect 13228 5524 13268 5564
rect 15244 5524 15284 5564
rect 15724 5524 15764 5564
rect 19948 5524 19988 5564
rect 3340 5440 3380 5480
rect 5548 5440 5588 5480
rect 8332 5440 8372 5480
rect 11596 5440 11636 5480
rect 17836 5440 17876 5480
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 4492 5104 4532 5144
rect 15628 5104 15668 5144
rect 4300 5020 4340 5060
rect 6124 5020 6164 5060
rect 11308 5020 11348 5060
rect 11500 5020 11540 5060
rect 13612 5020 13652 5060
rect 17548 5020 17588 5060
rect 2572 4936 2612 4976
rect 2668 4936 2708 4976
rect 3628 4936 3668 4976
rect 4108 4922 4148 4962
rect 4684 4936 4724 4976
rect 5932 4936 5972 4976
rect 6316 4936 6356 4976
rect 7564 4936 7604 4976
rect 7948 4936 7988 4976
rect 9196 4936 9236 4976
rect 9580 4936 9620 4976
rect 9676 4936 9716 4976
rect 10156 4936 10196 4976
rect 10636 4936 10676 4976
rect 11116 4931 11156 4971
rect 11596 4936 11636 4976
rect 11884 4936 11924 4976
rect 11980 4936 12020 4976
rect 12364 4936 12404 4976
rect 12940 4936 12980 4976
rect 13420 4922 13460 4962
rect 13900 4936 13940 4976
rect 13996 4936 14036 4976
rect 14956 4936 14996 4976
rect 15436 4931 15476 4971
rect 16108 4936 16148 4976
rect 17356 4936 17396 4976
rect 17740 4936 17780 4976
rect 18028 4936 18068 4976
rect 18124 4936 18164 4976
rect 18316 4936 18356 4976
rect 18508 4936 18548 4976
rect 19756 4936 19796 4976
rect 1420 4852 1460 4892
rect 1900 4852 1940 4892
rect 2092 4852 2132 4892
rect 3052 4852 3092 4892
rect 3148 4852 3188 4892
rect 10060 4852 10100 4892
rect 12460 4852 12500 4892
rect 14380 4852 14420 4892
rect 14476 4852 14516 4892
rect 1228 4768 1268 4808
rect 1708 4768 1748 4808
rect 15820 4768 15860 4808
rect 18316 4768 18356 4808
rect 2284 4684 2324 4724
rect 7756 4684 7796 4724
rect 19948 4684 19988 4724
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 2764 4348 2804 4388
rect 4396 4348 4436 4388
rect 10252 4348 10292 4388
rect 13324 4348 13364 4388
rect 15532 4348 15572 4388
rect 17836 4348 17876 4388
rect 11116 4264 11156 4304
rect 7276 4180 7316 4220
rect 7372 4180 7412 4220
rect 11884 4180 11924 4220
rect 13516 4180 13556 4220
rect 13900 4180 13940 4220
rect 1324 4096 1364 4136
rect 2572 4096 2612 4136
rect 2956 4096 2996 4136
rect 4204 4096 4244 4136
rect 4588 4096 4628 4136
rect 5836 4096 5876 4136
rect 6220 4096 6260 4136
rect 6316 4096 6356 4136
rect 6412 4096 6452 4136
rect 6508 4096 6548 4136
rect 6796 4096 6836 4136
rect 6892 4096 6932 4136
rect 7852 4096 7892 4136
rect 8380 4105 8420 4145
rect 8812 4096 8852 4136
rect 10060 4096 10100 4136
rect 10444 4096 10484 4136
rect 10540 4096 10580 4136
rect 10636 4096 10676 4136
rect 10732 4096 10772 4136
rect 10924 4096 10964 4136
rect 11116 4096 11156 4136
rect 11404 4096 11444 4136
rect 11500 4096 11540 4136
rect 11980 4096 12020 4136
rect 12460 4096 12500 4136
rect 12988 4105 13028 4145
rect 14092 4096 14132 4136
rect 15340 4096 15380 4136
rect 15916 4096 15956 4136
rect 16012 4096 16052 4136
rect 16396 4096 16436 4136
rect 17644 4096 17684 4136
rect 18028 4096 18068 4136
rect 18124 4096 18164 4136
rect 18316 4096 18356 4136
rect 18508 4096 18548 4136
rect 19756 4096 19796 4136
rect 8524 4012 8564 4052
rect 18220 4012 18260 4052
rect 6028 3928 6068 3968
rect 13132 3928 13172 3968
rect 13708 3928 13748 3968
rect 16204 3928 16244 3968
rect 17836 3928 17876 3968
rect 19948 3928 19988 3968
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 1324 3592 1364 3632
rect 1996 3592 2036 3632
rect 4300 3592 4340 3632
rect 6412 3592 6452 3632
rect 8620 3592 8660 3632
rect 8812 3592 8852 3632
rect 10444 3592 10484 3632
rect 11212 3592 11252 3632
rect 13228 3592 13268 3632
rect 16972 3592 17012 3632
rect 17356 3592 17396 3632
rect 19948 3592 19988 3632
rect 4012 3508 4052 3548
rect 4588 3508 4628 3548
rect 13900 3508 13940 3548
rect 19468 3508 19508 3548
rect 2188 3419 2228 3459
rect 2668 3424 2708 3464
rect 3244 3424 3284 3464
rect 3628 3424 3668 3464
rect 3724 3424 3764 3464
rect 4396 3424 4436 3464
rect 4780 3424 4820 3464
rect 6028 3424 6068 3464
rect 6316 3424 6356 3464
rect 6508 3424 6548 3464
rect 6604 3424 6644 3464
rect 6892 3424 6932 3464
rect 6988 3424 7028 3464
rect 7468 3424 7508 3464
rect 7948 3424 7988 3464
rect 8428 3410 8468 3450
rect 9004 3424 9044 3464
rect 10252 3424 10292 3464
rect 11020 3424 11060 3464
rect 11116 3424 11156 3464
rect 11308 3424 11348 3464
rect 11404 3424 11444 3464
rect 11505 3424 11545 3464
rect 11788 3424 11828 3464
rect 13036 3424 13076 3464
rect 13516 3424 13556 3464
rect 13804 3424 13844 3464
rect 15244 3424 15284 3464
rect 15340 3424 15380 3464
rect 15724 3424 15764 3464
rect 15820 3424 15860 3464
rect 16300 3424 16340 3464
rect 16780 3410 16820 3450
rect 17164 3424 17204 3464
rect 17452 3424 17492 3464
rect 17740 3424 17780 3464
rect 17836 3424 17876 3464
rect 18220 3424 18260 3464
rect 18316 3424 18356 3464
rect 18796 3424 18836 3464
rect 19324 3414 19364 3454
rect 19660 3424 19700 3464
rect 19756 3424 19796 3464
rect 19852 3424 19892 3464
rect 1516 3340 1556 3380
rect 3148 3340 3188 3380
rect 7372 3340 7412 3380
rect 10636 3340 10676 3380
rect 14380 3340 14420 3380
rect 14956 3340 14996 3380
rect 20140 3340 20180 3380
rect 1804 3256 1844 3296
rect 14188 3256 14228 3296
rect 14572 3172 14612 3212
rect 14764 3172 14804 3212
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 2860 2836 2900 2876
rect 9196 2836 9236 2876
rect 9964 2836 10004 2876
rect 14188 2836 14228 2876
rect 14380 2836 14420 2876
rect 3820 2752 3860 2792
rect 4396 2752 4436 2792
rect 9676 2752 9716 2792
rect 17644 2752 17684 2792
rect 3148 2668 3188 2708
rect 3628 2668 3668 2708
rect 4204 2668 4244 2708
rect 5644 2668 5684 2708
rect 6988 2668 7028 2708
rect 7372 2668 7412 2708
rect 10156 2668 10196 2708
rect 10540 2668 10580 2708
rect 11404 2668 11444 2708
rect 14572 2668 14612 2708
rect 15436 2668 15476 2708
rect 15532 2668 15572 2708
rect 17068 2668 17108 2708
rect 17452 2668 17492 2708
rect 18508 2668 18548 2708
rect 1420 2584 1460 2624
rect 2668 2584 2708 2624
rect 3052 2584 3092 2624
rect 3244 2584 3284 2624
rect 4684 2584 4724 2624
rect 5068 2584 5108 2624
rect 5164 2584 5204 2624
rect 5548 2584 5588 2624
rect 6124 2584 6164 2624
rect 6604 2589 6644 2629
rect 7756 2584 7796 2624
rect 9004 2584 9044 2624
rect 9388 2584 9428 2624
rect 9580 2584 9620 2624
rect 9676 2584 9716 2624
rect 10828 2584 10868 2624
rect 10924 2584 10964 2624
rect 11308 2584 11348 2624
rect 11884 2584 11924 2624
rect 12364 2589 12404 2629
rect 12748 2584 12788 2624
rect 13996 2584 14036 2624
rect 14956 2564 14996 2604
rect 15052 2603 15092 2643
rect 16540 2626 16580 2666
rect 16012 2584 16052 2624
rect 18028 2584 18068 2624
rect 18124 2584 18164 2624
rect 18604 2584 18644 2624
rect 19084 2584 19124 2624
rect 19564 2598 19604 2638
rect 19948 2584 19988 2624
rect 20044 2584 20084 2624
rect 20140 2584 20180 2624
rect 20236 2584 20276 2624
rect 6796 2500 6836 2540
rect 12556 2500 12596 2540
rect 16684 2500 16724 2540
rect 4012 2416 4052 2456
rect 7180 2416 7220 2456
rect 7564 2416 7604 2456
rect 10348 2416 10388 2456
rect 16876 2416 16916 2456
rect 17260 2416 17300 2456
rect 19756 2416 19796 2456
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 4300 2080 4340 2120
rect 5452 2080 5492 2120
rect 9004 2080 9044 2120
rect 9292 2080 9332 2120
rect 11692 2080 11732 2120
rect 11980 2080 12020 2120
rect 15244 2080 15284 2120
rect 15436 2080 15476 2120
rect 17164 2080 17204 2120
rect 19660 2080 19700 2120
rect 3820 1996 3860 2036
rect 2380 1912 2420 1952
rect 3628 1912 3668 1952
rect 4012 1912 4052 1952
rect 4108 1912 4148 1952
rect 5548 1912 5588 1952
rect 5644 1912 5684 1952
rect 5740 1912 5780 1952
rect 5932 1912 5972 1952
rect 7180 1912 7220 1952
rect 7564 1912 7604 1952
rect 8812 1912 8852 1952
rect 9964 1912 10004 1952
rect 10060 1912 10100 1952
rect 10540 1912 10580 1952
rect 11020 1912 11060 1952
rect 11500 1898 11540 1938
rect 12172 1912 12212 1952
rect 13420 1912 13460 1952
rect 13804 1912 13844 1952
rect 15052 1912 15092 1952
rect 15724 1912 15764 1952
rect 16972 1912 17012 1952
rect 17932 1912 17972 1952
rect 19180 1912 19220 1952
rect 19564 1912 19604 1952
rect 19756 1912 19796 1952
rect 19948 1912 19988 1952
rect 20044 1912 20084 1952
rect 20236 1912 20276 1952
rect 1228 1828 1268 1868
rect 1612 1828 1652 1868
rect 1996 1828 2036 1868
rect 4684 1828 4724 1868
rect 5068 1828 5108 1868
rect 9484 1828 9524 1868
rect 10444 1828 10484 1868
rect 17548 1828 17588 1868
rect 4876 1744 4916 1784
rect 7372 1744 7412 1784
rect 20236 1744 20276 1784
rect 1420 1660 1460 1700
rect 1804 1660 1844 1700
rect 2188 1660 2228 1700
rect 5260 1660 5300 1700
rect 9676 1660 9716 1700
rect 17356 1660 17396 1700
rect 19372 1660 19412 1700
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 20044 1324 20084 1364
rect 2860 1240 2900 1280
rect 4492 1240 4532 1280
rect 5836 1240 5876 1280
rect 7564 1240 7604 1280
rect 11020 1240 11060 1280
rect 12844 1240 12884 1280
rect 14572 1240 14612 1280
rect 16684 1240 16724 1280
rect 17452 1240 17492 1280
rect 17644 1240 17684 1280
rect 5068 1156 5108 1196
rect 5644 1156 5684 1196
rect 14956 1156 14996 1196
rect 17068 1156 17108 1196
rect 1420 1072 1460 1112
rect 2668 1072 2708 1112
rect 3052 1072 3092 1112
rect 4300 1072 4340 1112
rect 6124 1072 6164 1112
rect 7372 1072 7412 1112
rect 7756 1072 7796 1112
rect 9004 1072 9044 1112
rect 9580 1072 9620 1112
rect 10828 1072 10868 1112
rect 11212 1072 11252 1112
rect 12460 1072 12500 1112
rect 13036 1072 13076 1112
rect 14284 1072 14324 1112
rect 15244 1072 15284 1112
rect 16492 1072 16532 1112
rect 17836 1072 17876 1112
rect 19084 1072 19124 1112
rect 19372 1072 19412 1112
rect 19660 1072 19700 1112
rect 19756 1072 19796 1112
rect 4876 988 4916 1028
rect 9196 988 9236 1028
rect 5260 904 5300 944
rect 5452 904 5492 944
rect 9388 904 9428 944
rect 14764 904 14804 944
rect 16876 904 16916 944
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
<< metal2 >>
rect 1784 42928 1864 43008
rect 1976 42928 2056 43008
rect 2168 42944 2248 43008
rect 2168 42928 2188 42944
rect 75 42776 117 42785
rect 75 42736 76 42776
rect 116 42736 117 42776
rect 75 42727 117 42736
rect 76 28841 116 42727
rect 1611 42608 1653 42617
rect 1611 42568 1612 42608
rect 1652 42568 1653 42608
rect 1611 42559 1653 42568
rect 747 42440 789 42449
rect 747 42400 748 42440
rect 788 42400 789 42440
rect 747 42391 789 42400
rect 267 42104 309 42113
rect 267 42064 268 42104
rect 308 42064 309 42104
rect 267 42055 309 42064
rect 171 39668 213 39677
rect 171 39628 172 39668
rect 212 39628 213 39668
rect 171 39619 213 39628
rect 172 29009 212 39619
rect 268 33629 308 42055
rect 363 40424 405 40433
rect 363 40384 364 40424
rect 404 40384 405 40424
rect 363 40375 405 40384
rect 267 33620 309 33629
rect 267 33580 268 33620
rect 308 33580 309 33620
rect 267 33571 309 33580
rect 364 31949 404 40375
rect 363 31940 405 31949
rect 363 31900 364 31940
rect 404 31900 405 31940
rect 363 31891 405 31900
rect 748 29933 788 42391
rect 1419 41768 1461 41777
rect 1419 41728 1420 41768
rect 1460 41728 1461 41768
rect 1419 41719 1461 41728
rect 1323 41180 1365 41189
rect 1323 41140 1324 41180
rect 1364 41140 1365 41180
rect 1323 41131 1365 41140
rect 1324 41046 1364 41131
rect 1420 40928 1460 41719
rect 1515 41600 1557 41609
rect 1515 41560 1516 41600
rect 1556 41560 1557 41600
rect 1515 41551 1557 41560
rect 1516 41432 1556 41551
rect 1516 41383 1556 41392
rect 1515 41180 1557 41189
rect 1515 41140 1516 41180
rect 1556 41140 1557 41180
rect 1515 41131 1557 41140
rect 1324 40888 1460 40928
rect 1324 39920 1364 40888
rect 1419 40508 1461 40517
rect 1419 40468 1420 40508
rect 1460 40468 1461 40508
rect 1419 40459 1461 40468
rect 1420 40374 1460 40459
rect 1228 39880 1364 39920
rect 1228 39509 1268 39880
rect 1420 39836 1460 39845
rect 1324 39796 1420 39836
rect 1227 39500 1269 39509
rect 1227 39460 1228 39500
rect 1268 39460 1269 39500
rect 1227 39451 1269 39460
rect 1228 38996 1268 39005
rect 1228 37829 1268 38956
rect 1324 38240 1364 39796
rect 1420 39787 1460 39796
rect 1420 39080 1460 39089
rect 1516 39080 1556 41131
rect 1612 40676 1652 42559
rect 1804 42281 1844 42928
rect 1899 42440 1941 42449
rect 1899 42400 1900 42440
rect 1940 42400 1941 42440
rect 1899 42391 1941 42400
rect 1803 42272 1845 42281
rect 1803 42232 1804 42272
rect 1844 42232 1845 42272
rect 1803 42223 1845 42232
rect 1612 40627 1652 40636
rect 1708 41264 1748 41273
rect 1612 39738 1652 39747
rect 1612 39425 1652 39698
rect 1611 39416 1653 39425
rect 1611 39376 1612 39416
rect 1652 39376 1653 39416
rect 1611 39367 1653 39376
rect 1708 39257 1748 41224
rect 1900 40676 1940 42391
rect 1804 40636 1940 40676
rect 1707 39248 1749 39257
rect 1707 39208 1708 39248
rect 1748 39208 1749 39248
rect 1707 39199 1749 39208
rect 1804 39080 1844 40636
rect 1900 40508 1940 40517
rect 1900 40349 1940 40468
rect 1899 40340 1941 40349
rect 1899 40300 1900 40340
rect 1940 40300 1941 40340
rect 1899 40291 1941 40300
rect 1996 40181 2036 42928
rect 2187 42904 2188 42928
rect 2228 42928 2248 42944
rect 2360 42928 2440 43008
rect 2552 42928 2632 43008
rect 2744 42928 2824 43008
rect 2936 42928 3016 43008
rect 3128 42928 3208 43008
rect 3320 42928 3400 43008
rect 3512 42928 3592 43008
rect 3704 42928 3784 43008
rect 3896 42928 3976 43008
rect 4088 42928 4168 43008
rect 4280 42928 4360 43008
rect 4472 42928 4552 43008
rect 4664 42928 4744 43008
rect 4856 42928 4936 43008
rect 5048 42928 5128 43008
rect 5240 42928 5320 43008
rect 5432 42928 5512 43008
rect 5624 42928 5704 43008
rect 5816 42928 5896 43008
rect 6008 42928 6088 43008
rect 6200 42928 6280 43008
rect 6392 42928 6472 43008
rect 6584 42928 6664 43008
rect 6776 42928 6856 43008
rect 6968 42928 7048 43008
rect 7160 42928 7240 43008
rect 7352 42928 7432 43008
rect 7544 42928 7624 43008
rect 7736 42928 7816 43008
rect 7928 42928 8008 43008
rect 8120 42928 8200 43008
rect 8312 42928 8392 43008
rect 8504 42928 8584 43008
rect 8696 42928 8776 43008
rect 8888 42928 8968 43008
rect 9080 42928 9160 43008
rect 9272 42928 9352 43008
rect 9464 42928 9544 43008
rect 9656 42928 9736 43008
rect 9848 42928 9928 43008
rect 10040 42928 10120 43008
rect 10232 42928 10312 43008
rect 10424 42928 10504 43008
rect 10616 42928 10696 43008
rect 10808 42928 10888 43008
rect 11000 42928 11080 43008
rect 11192 42928 11272 43008
rect 11384 42928 11464 43008
rect 11576 42928 11656 43008
rect 11768 42928 11848 43008
rect 11960 42928 12040 43008
rect 12152 42928 12232 43008
rect 12344 42928 12424 43008
rect 12536 42928 12616 43008
rect 12728 42928 12808 43008
rect 12920 42928 13000 43008
rect 13112 42928 13192 43008
rect 13304 42928 13384 43008
rect 13496 42928 13576 43008
rect 13688 42928 13768 43008
rect 13880 42928 13960 43008
rect 14072 42928 14152 43008
rect 14264 42928 14344 43008
rect 14456 42928 14536 43008
rect 14648 42928 14728 43008
rect 14840 42928 14920 43008
rect 15032 42928 15112 43008
rect 15224 42928 15304 43008
rect 15416 42928 15496 43008
rect 15608 42928 15688 43008
rect 15800 42928 15880 43008
rect 15992 42928 16072 43008
rect 16184 42928 16264 43008
rect 16376 42928 16456 43008
rect 16568 42928 16648 43008
rect 16760 42928 16840 43008
rect 16952 42928 17032 43008
rect 17144 42928 17224 43008
rect 17336 42928 17416 43008
rect 17528 42928 17608 43008
rect 17720 42928 17800 43008
rect 17912 42928 17992 43008
rect 18104 42928 18184 43008
rect 18296 42928 18376 43008
rect 18488 42928 18568 43008
rect 18680 42928 18760 43008
rect 18872 42928 18952 43008
rect 19064 42928 19144 43008
rect 19256 42928 19336 43008
rect 19448 42928 19528 43008
rect 2228 42904 2229 42928
rect 2187 42895 2229 42904
rect 2187 42020 2229 42029
rect 2187 41980 2188 42020
rect 2228 41980 2229 42020
rect 2187 41971 2229 41980
rect 2091 40592 2133 40601
rect 2091 40552 2092 40592
rect 2132 40552 2133 40592
rect 2091 40543 2133 40552
rect 2092 40458 2132 40543
rect 2091 40340 2133 40349
rect 2091 40300 2092 40340
rect 2132 40300 2133 40340
rect 2091 40291 2133 40300
rect 1995 40172 2037 40181
rect 1995 40132 1996 40172
rect 2036 40132 2037 40172
rect 1995 40123 2037 40132
rect 2092 39920 2132 40291
rect 1460 39040 1556 39080
rect 1708 39040 1844 39080
rect 1900 39880 2132 39920
rect 1420 39031 1460 39040
rect 1612 38996 1652 39005
rect 1515 38912 1557 38921
rect 1515 38872 1516 38912
rect 1556 38872 1557 38912
rect 1515 38863 1557 38872
rect 1516 38324 1556 38863
rect 1612 38501 1652 38956
rect 1708 38921 1748 39040
rect 1707 38912 1749 38921
rect 1707 38872 1708 38912
rect 1748 38872 1749 38912
rect 1707 38863 1749 38872
rect 1804 38744 1844 38753
rect 1707 38660 1749 38669
rect 1707 38620 1708 38660
rect 1748 38620 1749 38660
rect 1707 38611 1749 38620
rect 1611 38492 1653 38501
rect 1611 38452 1612 38492
rect 1652 38452 1653 38492
rect 1611 38443 1653 38452
rect 1708 38408 1748 38611
rect 1804 38585 1844 38704
rect 1900 38660 1940 39880
rect 2091 39752 2133 39761
rect 2091 39712 2092 39752
rect 2132 39712 2133 39752
rect 2091 39703 2133 39712
rect 2092 39618 2132 39703
rect 2091 39500 2133 39509
rect 2091 39460 2092 39500
rect 2132 39460 2133 39500
rect 2091 39451 2133 39460
rect 1995 38996 2037 39005
rect 1995 38956 1996 38996
rect 2036 38956 2037 38996
rect 1995 38947 2037 38956
rect 1996 38862 2036 38947
rect 1900 38620 2036 38660
rect 1803 38576 1845 38585
rect 1803 38536 1804 38576
rect 1844 38536 1845 38576
rect 1803 38527 1845 38536
rect 1708 38359 1748 38368
rect 1803 38408 1845 38417
rect 1803 38368 1804 38408
rect 1844 38368 1845 38408
rect 1803 38359 1845 38368
rect 1516 38284 1652 38324
rect 1324 38200 1460 38240
rect 1324 38072 1364 38081
rect 1227 37820 1269 37829
rect 1227 37780 1228 37820
rect 1268 37780 1269 37820
rect 1227 37771 1269 37780
rect 1227 37652 1269 37661
rect 1227 37612 1228 37652
rect 1268 37612 1269 37652
rect 1324 37652 1364 38032
rect 1420 37820 1460 38200
rect 1515 38156 1557 38165
rect 1515 38116 1516 38156
rect 1556 38116 1557 38156
rect 1515 38107 1557 38116
rect 1516 38022 1556 38107
rect 1420 37780 1556 37820
rect 1324 37612 1460 37652
rect 1227 37603 1269 37612
rect 1228 36644 1268 37603
rect 1323 37484 1365 37493
rect 1323 37444 1324 37484
rect 1364 37444 1365 37484
rect 1323 37435 1365 37444
rect 1324 37350 1364 37435
rect 1323 37232 1365 37241
rect 1323 37192 1324 37232
rect 1364 37192 1365 37232
rect 1323 37183 1365 37192
rect 1228 36595 1268 36604
rect 1324 36392 1364 37183
rect 1420 37073 1460 37612
rect 1516 37484 1556 37780
rect 1516 37435 1556 37444
rect 1419 37064 1461 37073
rect 1419 37024 1420 37064
rect 1460 37024 1461 37064
rect 1419 37015 1461 37024
rect 1420 36896 1460 36905
rect 1612 36896 1652 38284
rect 1708 37652 1748 37661
rect 1804 37652 1844 38359
rect 1899 37736 1941 37745
rect 1899 37696 1900 37736
rect 1940 37696 1941 37736
rect 1899 37687 1941 37696
rect 1748 37612 1844 37652
rect 1708 37603 1748 37612
rect 1900 37316 1940 37687
rect 1900 37267 1940 37276
rect 1707 37232 1749 37241
rect 1707 37192 1708 37232
rect 1748 37192 1749 37232
rect 1707 37183 1749 37192
rect 1460 36856 1652 36896
rect 1708 36896 1748 37183
rect 1899 37064 1941 37073
rect 1899 37024 1900 37064
rect 1940 37024 1941 37064
rect 1899 37015 1941 37024
rect 1420 36847 1460 36856
rect 1708 36847 1748 36856
rect 1612 36569 1652 36654
rect 1900 36569 1940 37015
rect 1611 36560 1653 36569
rect 1611 36520 1612 36560
rect 1652 36520 1653 36560
rect 1611 36511 1653 36520
rect 1899 36560 1941 36569
rect 1899 36520 1900 36560
rect 1940 36520 1941 36560
rect 1899 36511 1941 36520
rect 1324 36352 1652 36392
rect 939 35972 981 35981
rect 939 35932 940 35972
rect 980 35932 981 35972
rect 939 35923 981 35932
rect 1516 35972 1556 35981
rect 1612 35972 1652 36352
rect 1708 36149 1748 36234
rect 1707 36140 1749 36149
rect 1707 36100 1708 36140
rect 1748 36100 1749 36140
rect 1707 36091 1749 36100
rect 1612 35932 1748 35972
rect 843 31016 885 31025
rect 843 30976 844 31016
rect 884 30976 885 31016
rect 843 30967 885 30976
rect 747 29924 789 29933
rect 747 29884 748 29924
rect 788 29884 789 29924
rect 747 29875 789 29884
rect 459 29588 501 29597
rect 459 29548 460 29588
rect 500 29548 501 29588
rect 459 29539 501 29548
rect 171 29000 213 29009
rect 171 28960 172 29000
rect 212 28960 213 29000
rect 171 28951 213 28960
rect 75 28832 117 28841
rect 75 28792 76 28832
rect 116 28792 117 28832
rect 75 28783 117 28792
rect 460 23633 500 29539
rect 651 26732 693 26741
rect 651 26692 652 26732
rect 692 26692 693 26732
rect 651 26683 693 26692
rect 652 23969 692 26683
rect 844 24053 884 30967
rect 940 29093 980 35923
rect 1324 35720 1364 35731
rect 1324 35645 1364 35680
rect 1323 35636 1365 35645
rect 1323 35596 1324 35636
rect 1364 35596 1365 35636
rect 1323 35587 1365 35596
rect 1324 35216 1364 35225
rect 1324 34805 1364 35176
rect 1420 35216 1460 35225
rect 1323 34796 1365 34805
rect 1323 34756 1324 34796
rect 1364 34756 1365 34796
rect 1323 34747 1365 34756
rect 1420 34628 1460 35176
rect 1324 34588 1460 34628
rect 1035 34460 1077 34469
rect 1035 34420 1036 34460
rect 1076 34420 1077 34460
rect 1035 34411 1077 34420
rect 939 29084 981 29093
rect 939 29044 940 29084
rect 980 29044 981 29084
rect 939 29035 981 29044
rect 1036 28253 1076 34411
rect 1131 33620 1173 33629
rect 1131 33580 1132 33620
rect 1172 33580 1173 33620
rect 1131 33571 1173 33580
rect 1228 33620 1268 33629
rect 1132 32864 1172 33571
rect 1228 33209 1268 33580
rect 1227 33200 1269 33209
rect 1227 33160 1228 33200
rect 1268 33160 1269 33200
rect 1227 33151 1269 33160
rect 1324 33032 1364 34588
rect 1419 34460 1461 34469
rect 1419 34420 1420 34460
rect 1460 34420 1461 34460
rect 1419 34411 1461 34420
rect 1420 34326 1460 34411
rect 1516 34301 1556 35932
rect 1611 34628 1653 34637
rect 1611 34588 1612 34628
rect 1652 34588 1653 34628
rect 1611 34579 1653 34588
rect 1612 34494 1652 34579
rect 1611 34376 1653 34385
rect 1611 34336 1612 34376
rect 1652 34336 1653 34376
rect 1611 34327 1653 34336
rect 1515 34292 1557 34301
rect 1515 34252 1516 34292
rect 1556 34252 1557 34292
rect 1515 34243 1557 34252
rect 1419 33872 1461 33881
rect 1419 33832 1420 33872
rect 1460 33832 1461 33872
rect 1419 33823 1461 33832
rect 1420 33738 1460 33823
rect 1612 33704 1652 34327
rect 1612 33655 1652 33664
rect 1708 33536 1748 35932
rect 1900 35720 1940 36511
rect 1996 36149 2036 38620
rect 2092 38492 2132 39451
rect 2188 39080 2228 41971
rect 2283 40424 2325 40433
rect 2283 40384 2284 40424
rect 2324 40384 2325 40424
rect 2283 40375 2325 40384
rect 2284 40290 2324 40375
rect 2380 39164 2420 42928
rect 2475 42524 2517 42533
rect 2475 42484 2476 42524
rect 2516 42484 2517 42524
rect 2475 42475 2517 42484
rect 2188 39031 2228 39040
rect 2284 39124 2420 39164
rect 2284 38669 2324 39124
rect 2379 38996 2421 39005
rect 2379 38956 2380 38996
rect 2420 38956 2421 38996
rect 2379 38947 2421 38956
rect 2380 38862 2420 38947
rect 2283 38660 2325 38669
rect 2283 38620 2284 38660
rect 2324 38620 2325 38660
rect 2283 38611 2325 38620
rect 2092 38452 2324 38492
rect 2187 38156 2229 38165
rect 2187 38116 2188 38156
rect 2228 38116 2229 38156
rect 2187 38107 2229 38116
rect 2188 38022 2228 38107
rect 2284 37820 2324 38452
rect 2379 38156 2421 38165
rect 2379 38116 2380 38156
rect 2420 38116 2421 38156
rect 2379 38107 2421 38116
rect 2380 38022 2420 38107
rect 2284 37780 2420 37820
rect 2091 37568 2133 37577
rect 2091 37528 2092 37568
rect 2132 37528 2133 37568
rect 2091 37519 2133 37528
rect 2092 37414 2132 37519
rect 2092 37365 2132 37374
rect 2188 36728 2228 36737
rect 2228 36688 2324 36728
rect 2188 36679 2228 36688
rect 2091 36644 2133 36653
rect 2091 36604 2092 36644
rect 2132 36604 2133 36644
rect 2091 36595 2133 36604
rect 1995 36140 2037 36149
rect 1995 36100 1996 36140
rect 2036 36100 2037 36140
rect 1995 36091 2037 36100
rect 2092 35972 2132 36595
rect 1804 35680 1900 35720
rect 1804 35309 1844 35680
rect 1900 35671 1940 35680
rect 1996 35932 2132 35972
rect 1899 35552 1941 35561
rect 1899 35512 1900 35552
rect 1940 35512 1941 35552
rect 1899 35503 1941 35512
rect 1803 35300 1845 35309
rect 1803 35260 1804 35300
rect 1844 35260 1845 35300
rect 1803 35251 1845 35260
rect 1900 35216 1940 35503
rect 1900 35167 1940 35176
rect 1804 35132 1844 35141
rect 1804 34889 1844 35092
rect 1803 34880 1845 34889
rect 1803 34840 1804 34880
rect 1844 34840 1845 34880
rect 1803 34831 1845 34840
rect 1996 34628 2036 35932
rect 2188 35720 2228 35729
rect 1996 34579 2036 34588
rect 2092 35680 2188 35720
rect 1804 34460 1844 34469
rect 1804 34133 1844 34420
rect 1803 34124 1845 34133
rect 1803 34084 1804 34124
rect 1844 34084 1845 34124
rect 1803 34075 1845 34084
rect 2092 33956 2132 35680
rect 2188 35671 2228 35680
rect 2284 35552 2324 36688
rect 2380 36476 2420 37780
rect 2476 36653 2516 42475
rect 2572 40424 2612 42928
rect 2764 42533 2804 42928
rect 2763 42524 2805 42533
rect 2763 42484 2764 42524
rect 2804 42484 2805 42524
rect 2763 42475 2805 42484
rect 2956 41432 2996 42928
rect 2956 41392 3092 41432
rect 2956 41264 2996 41273
rect 2860 41224 2956 41264
rect 2572 40384 2804 40424
rect 2667 40004 2709 40013
rect 2667 39964 2668 40004
rect 2708 39964 2709 40004
rect 2667 39955 2709 39964
rect 2668 39752 2708 39955
rect 2668 39677 2708 39712
rect 2572 39668 2612 39677
rect 2572 39416 2612 39628
rect 2667 39668 2709 39677
rect 2667 39628 2668 39668
rect 2708 39628 2709 39668
rect 2667 39619 2709 39628
rect 2668 39617 2708 39619
rect 2667 39416 2709 39425
rect 2572 39376 2668 39416
rect 2708 39376 2709 39416
rect 2667 39367 2709 39376
rect 2764 39173 2804 40384
rect 2763 39164 2805 39173
rect 2763 39124 2764 39164
rect 2804 39124 2805 39164
rect 2763 39115 2805 39124
rect 2764 38996 2804 39005
rect 2668 38956 2764 38996
rect 2572 38744 2612 38753
rect 2572 38333 2612 38704
rect 2571 38324 2613 38333
rect 2571 38284 2572 38324
rect 2612 38284 2613 38324
rect 2571 38275 2613 38284
rect 2571 38156 2613 38165
rect 2571 38116 2572 38156
rect 2612 38116 2613 38156
rect 2571 38107 2613 38116
rect 2572 38072 2612 38107
rect 2572 38021 2612 38032
rect 2572 37400 2612 37411
rect 2572 37325 2612 37360
rect 2571 37316 2613 37325
rect 2571 37276 2572 37316
rect 2612 37276 2613 37316
rect 2571 37267 2613 37276
rect 2475 36644 2517 36653
rect 2475 36604 2476 36644
rect 2516 36604 2517 36644
rect 2475 36595 2517 36604
rect 2380 36436 2516 36476
rect 2379 36140 2421 36149
rect 2379 36100 2380 36140
rect 2420 36100 2421 36140
rect 2379 36091 2421 36100
rect 2380 35888 2420 36091
rect 2380 35839 2420 35848
rect 2188 35512 2324 35552
rect 2188 35225 2228 35512
rect 2379 35300 2421 35309
rect 2476 35300 2516 36436
rect 2571 35636 2613 35645
rect 2571 35596 2572 35636
rect 2612 35596 2613 35636
rect 2571 35587 2613 35596
rect 2379 35260 2380 35300
rect 2420 35260 2516 35300
rect 2379 35251 2421 35260
rect 2187 35216 2229 35225
rect 2187 35176 2188 35216
rect 2228 35176 2229 35216
rect 2187 35167 2229 35176
rect 2367 35189 2407 35198
rect 2188 34721 2228 35167
rect 2367 34880 2407 35149
rect 2572 34880 2612 35587
rect 2668 35057 2708 38956
rect 2764 38947 2804 38956
rect 2860 38240 2900 41224
rect 2956 41215 2996 41224
rect 3052 40508 3092 41392
rect 3148 41180 3188 42928
rect 3340 41684 3380 42928
rect 3340 41644 3476 41684
rect 3339 41264 3381 41273
rect 3339 41224 3340 41264
rect 3380 41224 3381 41264
rect 3339 41215 3381 41224
rect 3148 41140 3284 41180
rect 3147 41012 3189 41021
rect 3147 40972 3148 41012
rect 3188 40972 3189 41012
rect 3147 40963 3189 40972
rect 3148 40878 3188 40963
rect 3147 40760 3189 40769
rect 3147 40720 3148 40760
rect 3188 40720 3189 40760
rect 3147 40711 3189 40720
rect 2956 40468 3092 40508
rect 2956 39173 2996 40468
rect 3052 39752 3092 39761
rect 2955 39164 2997 39173
rect 2955 39124 2956 39164
rect 2996 39124 2997 39164
rect 2955 39115 2997 39124
rect 2956 38753 2996 38838
rect 2955 38744 2997 38753
rect 2955 38704 2956 38744
rect 2996 38704 2997 38744
rect 2955 38695 2997 38704
rect 2955 38576 2997 38585
rect 2955 38536 2956 38576
rect 2996 38536 2997 38576
rect 2955 38527 2997 38536
rect 2956 38408 2996 38527
rect 2956 38359 2996 38368
rect 2860 38200 2996 38240
rect 2763 38156 2805 38165
rect 2763 38116 2764 38156
rect 2804 38116 2805 38156
rect 2763 38107 2805 38116
rect 2764 38022 2804 38107
rect 2956 37913 2996 38200
rect 2955 37904 2997 37913
rect 2955 37864 2956 37904
rect 2996 37864 2997 37904
rect 2955 37855 2997 37864
rect 2763 37820 2805 37829
rect 2763 37780 2764 37820
rect 2804 37780 2805 37820
rect 2763 37771 2805 37780
rect 2667 35048 2709 35057
rect 2667 35008 2668 35048
rect 2708 35008 2709 35048
rect 2667 34999 2709 35008
rect 2367 34840 2612 34880
rect 2187 34712 2229 34721
rect 2187 34672 2188 34712
rect 2228 34672 2229 34712
rect 2187 34663 2229 34672
rect 2380 34385 2420 34390
rect 2379 34381 2421 34385
rect 2379 34336 2380 34381
rect 2420 34336 2421 34381
rect 2379 34327 2421 34336
rect 2187 34292 2229 34301
rect 2187 34252 2188 34292
rect 2228 34252 2229 34292
rect 2187 34243 2229 34252
rect 2380 34246 2420 34327
rect 2188 34158 2228 34243
rect 2283 34124 2325 34133
rect 2283 34084 2284 34124
rect 2324 34084 2325 34124
rect 2283 34075 2325 34084
rect 1612 33496 1748 33536
rect 1996 33916 2132 33956
rect 2187 33956 2229 33965
rect 2187 33916 2188 33956
rect 2228 33916 2229 33956
rect 1324 32992 1460 33032
rect 1324 32864 1364 32873
rect 1132 32824 1324 32864
rect 1324 32815 1364 32824
rect 1323 32612 1365 32621
rect 1323 32572 1324 32612
rect 1364 32572 1365 32612
rect 1323 32563 1365 32572
rect 1324 32360 1364 32563
rect 1324 32311 1364 32320
rect 1228 32192 1268 32201
rect 1228 31781 1268 32152
rect 1420 32033 1460 32992
rect 1515 32108 1557 32117
rect 1515 32068 1516 32108
rect 1556 32068 1557 32108
rect 1515 32059 1557 32068
rect 1419 32024 1461 32033
rect 1419 31984 1420 32024
rect 1460 31984 1461 32024
rect 1419 31975 1461 31984
rect 1516 31974 1556 32059
rect 1612 31856 1652 33496
rect 1707 32444 1749 32453
rect 1707 32404 1708 32444
rect 1748 32404 1749 32444
rect 1707 32395 1749 32404
rect 1708 32360 1748 32395
rect 1708 32309 1748 32320
rect 1996 32192 2036 33916
rect 2187 33907 2229 33916
rect 1996 32143 2036 32152
rect 2091 32192 2133 32201
rect 2091 32152 2092 32192
rect 2132 32152 2133 32192
rect 2091 32143 2133 32152
rect 2092 32058 2132 32143
rect 1707 32024 1749 32033
rect 1707 31984 1708 32024
rect 1748 31984 1749 32024
rect 1707 31975 1749 31984
rect 1516 31816 1652 31856
rect 1227 31772 1269 31781
rect 1227 31732 1228 31772
rect 1268 31732 1269 31772
rect 1227 31723 1269 31732
rect 1419 31520 1461 31529
rect 1419 31480 1420 31520
rect 1460 31480 1461 31520
rect 1419 31471 1461 31480
rect 1131 31436 1173 31445
rect 1131 31396 1132 31436
rect 1172 31396 1173 31436
rect 1131 31387 1173 31396
rect 1132 30353 1172 31387
rect 1323 31184 1365 31193
rect 1323 31144 1324 31184
rect 1364 31144 1365 31184
rect 1323 31135 1365 31144
rect 1324 31050 1364 31135
rect 1323 30932 1365 30941
rect 1228 30892 1324 30932
rect 1364 30892 1365 30932
rect 1228 30680 1268 30892
rect 1323 30883 1365 30892
rect 1228 30631 1268 30640
rect 1323 30428 1365 30437
rect 1323 30388 1324 30428
rect 1364 30388 1365 30428
rect 1323 30379 1365 30388
rect 1131 30344 1173 30353
rect 1131 30304 1132 30344
rect 1172 30304 1173 30344
rect 1131 30295 1173 30304
rect 1227 29924 1269 29933
rect 1227 29884 1228 29924
rect 1268 29884 1269 29924
rect 1227 29875 1269 29884
rect 1228 29840 1268 29875
rect 1228 29681 1268 29800
rect 1227 29672 1269 29681
rect 1227 29632 1228 29672
rect 1268 29632 1269 29672
rect 1227 29623 1269 29632
rect 1131 29000 1173 29009
rect 1131 28960 1132 29000
rect 1172 28960 1173 29000
rect 1324 29000 1364 30379
rect 1420 29168 1460 31471
rect 1516 30437 1556 31816
rect 1611 31268 1653 31277
rect 1611 31228 1612 31268
rect 1652 31228 1653 31268
rect 1611 31219 1653 31228
rect 1612 31134 1652 31219
rect 1515 30428 1557 30437
rect 1515 30388 1516 30428
rect 1556 30388 1557 30428
rect 1515 30379 1557 30388
rect 1708 30269 1748 31975
rect 2188 31940 2228 33907
rect 2284 33881 2324 34075
rect 2572 33965 2612 34840
rect 2764 34637 2804 37771
rect 3052 37652 3092 39712
rect 3148 39752 3188 40711
rect 3148 39703 3188 39712
rect 3147 39080 3189 39089
rect 3147 39040 3148 39080
rect 3188 39040 3189 39080
rect 3147 39031 3189 39040
rect 3148 38996 3188 39031
rect 3148 38945 3188 38956
rect 3147 38828 3189 38837
rect 3147 38788 3148 38828
rect 3188 38788 3189 38828
rect 3147 38779 3189 38788
rect 3148 38417 3188 38779
rect 3147 38408 3189 38417
rect 3147 38368 3148 38408
rect 3188 38368 3189 38408
rect 3147 38359 3189 38368
rect 3148 38240 3188 38249
rect 3148 37997 3188 38200
rect 3147 37988 3189 37997
rect 3147 37948 3148 37988
rect 3188 37948 3189 37988
rect 3147 37939 3189 37948
rect 2956 37612 3092 37652
rect 2859 36896 2901 36905
rect 2859 36856 2860 36896
rect 2900 36856 2901 36896
rect 2859 36847 2901 36856
rect 2860 35981 2900 36847
rect 2859 35972 2901 35981
rect 2859 35932 2860 35972
rect 2900 35932 2901 35972
rect 2859 35923 2901 35932
rect 2956 35477 2996 37612
rect 3052 37484 3092 37493
rect 3052 36569 3092 37444
rect 3147 37400 3189 37409
rect 3147 37360 3148 37400
rect 3188 37360 3189 37400
rect 3147 37351 3189 37360
rect 3148 37266 3188 37351
rect 3051 36560 3093 36569
rect 3051 36520 3052 36560
rect 3092 36520 3093 36560
rect 3051 36511 3093 36520
rect 3147 36224 3189 36233
rect 3147 36184 3148 36224
rect 3188 36184 3189 36224
rect 3147 36175 3189 36184
rect 3148 35561 3188 36175
rect 3147 35552 3189 35561
rect 3147 35512 3148 35552
rect 3188 35512 3189 35552
rect 3147 35503 3189 35512
rect 2955 35468 2997 35477
rect 2955 35428 2956 35468
rect 2996 35428 2997 35468
rect 2955 35419 2997 35428
rect 3052 35300 3092 35309
rect 2908 35174 2948 35183
rect 3052 35141 3092 35260
rect 3147 35216 3189 35225
rect 3147 35176 3148 35216
rect 3188 35176 3189 35216
rect 3244 35216 3284 41140
rect 3340 41130 3380 41215
rect 3339 40676 3381 40685
rect 3339 40636 3340 40676
rect 3380 40636 3381 40676
rect 3339 40627 3381 40636
rect 3340 38921 3380 40627
rect 3436 40433 3476 41644
rect 3532 40685 3572 42928
rect 3724 42365 3764 42928
rect 3723 42356 3765 42365
rect 3723 42316 3724 42356
rect 3764 42316 3765 42356
rect 3723 42307 3765 42316
rect 3916 41189 3956 42928
rect 4108 42449 4148 42928
rect 4107 42440 4149 42449
rect 4107 42400 4108 42440
rect 4148 42400 4149 42440
rect 4107 42391 4149 42400
rect 3915 41180 3957 41189
rect 3915 41140 3916 41180
rect 3956 41140 3957 41180
rect 3915 41131 3957 41140
rect 3688 40844 4056 40853
rect 3728 40804 3770 40844
rect 3810 40804 3852 40844
rect 3892 40804 3934 40844
rect 3974 40804 4016 40844
rect 3688 40795 4056 40804
rect 3531 40676 3573 40685
rect 3531 40636 3532 40676
rect 3572 40636 3573 40676
rect 3531 40627 3573 40636
rect 4107 40676 4149 40685
rect 4107 40636 4108 40676
rect 4148 40636 4149 40676
rect 4107 40627 4149 40636
rect 3531 40508 3573 40517
rect 3531 40468 3532 40508
rect 3572 40468 3573 40508
rect 3531 40459 3573 40468
rect 3435 40424 3477 40433
rect 3435 40384 3436 40424
rect 3476 40384 3477 40424
rect 3435 40375 3477 40384
rect 3532 40424 3572 40459
rect 3532 40373 3572 40384
rect 3916 40424 3956 40435
rect 3916 40349 3956 40384
rect 3915 40340 3957 40349
rect 3915 40300 3916 40340
rect 3956 40300 3957 40340
rect 3915 40291 3957 40300
rect 3724 40256 3764 40265
rect 3436 40216 3724 40256
rect 3339 38912 3381 38921
rect 3339 38872 3340 38912
rect 3380 38872 3381 38912
rect 3339 38863 3381 38872
rect 3339 38744 3381 38753
rect 3339 38704 3340 38744
rect 3380 38704 3381 38744
rect 3339 38695 3381 38704
rect 3340 38610 3380 38695
rect 3436 36896 3476 40216
rect 3724 40207 3764 40216
rect 3915 40172 3957 40181
rect 3915 40132 3916 40172
rect 3956 40132 3957 40172
rect 3915 40123 3957 40132
rect 3916 39920 3956 40123
rect 3916 39871 3956 39880
rect 3531 39836 3573 39845
rect 3531 39796 3532 39836
rect 3572 39796 3573 39836
rect 3531 39787 3573 39796
rect 3532 39702 3572 39787
rect 3723 39668 3765 39677
rect 3723 39628 3724 39668
rect 3764 39628 3765 39668
rect 3723 39619 3765 39628
rect 4108 39668 4148 40627
rect 4300 40424 4340 42928
rect 4395 41768 4437 41777
rect 4395 41728 4396 41768
rect 4436 41728 4437 41768
rect 4395 41719 4437 41728
rect 3724 39534 3764 39619
rect 3688 39332 4056 39341
rect 3728 39292 3770 39332
rect 3810 39292 3852 39332
rect 3892 39292 3934 39332
rect 3974 39292 4016 39332
rect 3688 39283 4056 39292
rect 4011 39164 4053 39173
rect 4011 39124 4012 39164
rect 4052 39124 4053 39164
rect 4011 39115 4053 39124
rect 3627 39080 3669 39089
rect 3627 39040 3628 39080
rect 3668 39040 3669 39080
rect 3627 39031 3669 39040
rect 3531 38996 3573 39005
rect 3531 38956 3532 38996
rect 3572 38956 3573 38996
rect 3531 38947 3573 38956
rect 3532 38862 3572 38947
rect 3628 38501 3668 39031
rect 4012 38931 4052 39115
rect 4108 39089 4148 39628
rect 4204 40384 4340 40424
rect 4204 39332 4244 40384
rect 4299 40088 4341 40097
rect 4299 40048 4300 40088
rect 4340 40048 4341 40088
rect 4299 40039 4341 40048
rect 4300 39920 4340 40039
rect 4300 39871 4340 39880
rect 4204 39292 4340 39332
rect 4203 39164 4245 39173
rect 4203 39124 4204 39164
rect 4244 39124 4245 39164
rect 4203 39115 4245 39124
rect 4107 39080 4149 39089
rect 4107 39040 4108 39080
rect 4148 39040 4149 39080
rect 4107 39031 4149 39040
rect 4012 38882 4052 38891
rect 4107 38912 4149 38921
rect 4107 38872 4108 38912
rect 4148 38872 4149 38912
rect 4107 38863 4149 38872
rect 3819 38828 3861 38837
rect 3819 38788 3820 38828
rect 3860 38788 3861 38828
rect 3819 38779 3861 38788
rect 3724 38744 3764 38753
rect 3627 38492 3669 38501
rect 3627 38452 3628 38492
rect 3668 38452 3669 38492
rect 3627 38443 3669 38452
rect 3628 38081 3668 38443
rect 3724 38165 3764 38704
rect 3723 38156 3765 38165
rect 3723 38116 3724 38156
rect 3764 38116 3765 38156
rect 3723 38107 3765 38116
rect 3627 38072 3669 38081
rect 3627 38032 3628 38072
rect 3668 38032 3669 38072
rect 3627 38023 3669 38032
rect 3820 37997 3860 38779
rect 4108 38778 4148 38863
rect 4011 38660 4053 38669
rect 4011 38620 4012 38660
rect 4052 38620 4053 38660
rect 4011 38611 4053 38620
rect 3819 37988 3861 37997
rect 3819 37948 3820 37988
rect 3860 37948 3861 37988
rect 4012 37988 4052 38611
rect 4012 37948 4148 37988
rect 3819 37939 3861 37948
rect 3688 37820 4056 37829
rect 3728 37780 3770 37820
rect 3810 37780 3852 37820
rect 3892 37780 3934 37820
rect 3974 37780 4016 37820
rect 3688 37771 4056 37780
rect 4108 37652 4148 37948
rect 4012 37612 4148 37652
rect 3532 37400 3572 37409
rect 3532 37157 3572 37360
rect 3628 37400 3668 37409
rect 3531 37148 3573 37157
rect 3531 37108 3532 37148
rect 3572 37108 3573 37148
rect 3531 37099 3573 37108
rect 3340 36856 3476 36896
rect 3531 36896 3573 36905
rect 3531 36856 3532 36896
rect 3572 36856 3573 36896
rect 3340 36569 3380 36856
rect 3531 36847 3573 36856
rect 3436 36728 3476 36737
rect 3532 36728 3572 36847
rect 3476 36688 3572 36728
rect 3436 36679 3476 36688
rect 3628 36644 3668 37360
rect 3819 37400 3861 37409
rect 3819 37360 3820 37400
rect 3860 37360 3861 37400
rect 3819 37351 3861 37360
rect 3820 37241 3860 37351
rect 3819 37232 3861 37241
rect 3819 37192 3820 37232
rect 3860 37192 3861 37232
rect 3819 37183 3861 37192
rect 3532 36604 3668 36644
rect 3820 36644 3860 37183
rect 4012 36896 4052 37612
rect 4107 37484 4149 37493
rect 4107 37444 4108 37484
rect 4148 37444 4149 37484
rect 4107 37435 4149 37444
rect 4108 37350 4148 37435
rect 4012 36847 4052 36856
rect 4204 36812 4244 39115
rect 4300 37820 4340 39292
rect 4396 38669 4436 41719
rect 4492 41609 4532 42928
rect 4491 41600 4533 41609
rect 4491 41560 4492 41600
rect 4532 41560 4533 41600
rect 4491 41551 4533 41560
rect 4587 41516 4629 41525
rect 4587 41476 4588 41516
rect 4628 41476 4629 41516
rect 4587 41467 4629 41476
rect 4588 41264 4628 41467
rect 4588 41215 4628 41224
rect 4491 40760 4533 40769
rect 4491 40720 4492 40760
rect 4532 40720 4533 40760
rect 4491 40711 4533 40720
rect 4492 40265 4532 40711
rect 4684 40424 4724 42928
rect 4876 41777 4916 42928
rect 5068 42617 5108 42928
rect 5067 42608 5109 42617
rect 5067 42568 5068 42608
rect 5108 42568 5109 42608
rect 5067 42559 5109 42568
rect 5260 41852 5300 42928
rect 5452 42869 5492 42928
rect 5451 42860 5493 42869
rect 5451 42820 5452 42860
rect 5492 42820 5493 42860
rect 5451 42811 5493 42820
rect 5260 41812 5588 41852
rect 4875 41768 4917 41777
rect 4875 41728 4876 41768
rect 4916 41728 4917 41768
rect 4875 41719 4917 41728
rect 5451 41684 5493 41693
rect 5451 41644 5452 41684
rect 5492 41644 5493 41684
rect 5451 41635 5493 41644
rect 4928 41600 5296 41609
rect 4968 41560 5010 41600
rect 5050 41560 5092 41600
rect 5132 41560 5174 41600
rect 5214 41560 5256 41600
rect 4928 41551 5296 41560
rect 5355 41516 5397 41525
rect 5355 41476 5356 41516
rect 5396 41476 5397 41516
rect 5355 41467 5397 41476
rect 4972 41264 5012 41273
rect 4588 40384 4724 40424
rect 4780 41012 4820 41021
rect 4491 40256 4533 40265
rect 4491 40216 4492 40256
rect 4532 40216 4533 40256
rect 4491 40207 4533 40216
rect 4491 39668 4533 39677
rect 4491 39628 4492 39668
rect 4532 39628 4533 39668
rect 4491 39619 4533 39628
rect 4492 39534 4532 39619
rect 4588 39173 4628 40384
rect 4683 40256 4725 40265
rect 4683 40216 4684 40256
rect 4724 40216 4725 40256
rect 4683 40207 4725 40216
rect 4684 39920 4724 40207
rect 4684 39871 4724 39880
rect 4683 39668 4725 39677
rect 4683 39628 4684 39668
rect 4724 39628 4725 39668
rect 4683 39619 4725 39628
rect 4587 39164 4629 39173
rect 4587 39124 4588 39164
rect 4628 39124 4629 39164
rect 4587 39115 4629 39124
rect 4588 38996 4628 39005
rect 4684 38996 4724 39619
rect 4628 38956 4724 38996
rect 4491 38912 4533 38921
rect 4491 38872 4492 38912
rect 4532 38872 4533 38912
rect 4491 38863 4533 38872
rect 4492 38778 4532 38863
rect 4395 38660 4437 38669
rect 4588 38660 4628 38956
rect 4395 38620 4396 38660
rect 4436 38620 4437 38660
rect 4395 38611 4437 38620
rect 4492 38620 4628 38660
rect 4395 38492 4437 38501
rect 4395 38452 4396 38492
rect 4436 38452 4437 38492
rect 4395 38443 4437 38452
rect 4396 38240 4436 38443
rect 4396 38191 4436 38200
rect 4300 37780 4436 37820
rect 4299 37652 4341 37661
rect 4299 37612 4300 37652
rect 4340 37612 4341 37652
rect 4299 37603 4341 37612
rect 4300 37518 4340 37603
rect 4396 36896 4436 37780
rect 4492 37493 4532 38620
rect 4588 37997 4628 38082
rect 4587 37988 4629 37997
rect 4587 37948 4588 37988
rect 4628 37948 4629 37988
rect 4587 37939 4629 37948
rect 4587 37736 4629 37745
rect 4587 37696 4588 37736
rect 4628 37696 4629 37736
rect 4587 37687 4629 37696
rect 4491 37484 4533 37493
rect 4491 37444 4492 37484
rect 4532 37444 4533 37484
rect 4491 37435 4533 37444
rect 4492 37232 4532 37243
rect 4492 37157 4532 37192
rect 4491 37148 4533 37157
rect 4491 37108 4492 37148
rect 4532 37108 4533 37148
rect 4491 37099 4533 37108
rect 4396 36847 4436 36856
rect 4588 36896 4628 37687
rect 4780 37414 4820 40972
rect 4972 40769 5012 41224
rect 4971 40760 5013 40769
rect 4971 40720 4972 40760
rect 5012 40720 5013 40760
rect 4971 40711 5013 40720
rect 5067 40592 5109 40601
rect 5067 40552 5068 40592
rect 5108 40552 5109 40592
rect 5067 40543 5109 40552
rect 5068 40424 5108 40543
rect 5356 40438 5396 41467
rect 5164 40424 5204 40433
rect 5068 40384 5164 40424
rect 5164 40340 5204 40384
rect 5260 40398 5396 40438
rect 5260 40340 5300 40398
rect 5164 40300 5300 40340
rect 5355 40340 5397 40349
rect 5355 40300 5356 40340
rect 5396 40300 5397 40340
rect 5355 40291 5397 40300
rect 5356 40206 5396 40291
rect 4928 40088 5296 40097
rect 4968 40048 5010 40088
rect 5050 40048 5092 40088
rect 5132 40048 5174 40088
rect 5214 40048 5256 40088
rect 4928 40039 5296 40048
rect 5068 39920 5108 39929
rect 5452 39920 5492 41635
rect 5548 41180 5588 41812
rect 5644 41777 5684 42928
rect 5643 41768 5685 41777
rect 5836 41768 5876 42928
rect 6028 41861 6068 42928
rect 6027 41852 6069 41861
rect 6027 41812 6028 41852
rect 6068 41812 6069 41852
rect 6027 41803 6069 41812
rect 5643 41728 5644 41768
rect 5684 41728 5685 41768
rect 5643 41719 5685 41728
rect 5740 41728 5876 41768
rect 5931 41768 5973 41777
rect 5931 41728 5932 41768
rect 5972 41728 5973 41768
rect 5740 41441 5780 41728
rect 5931 41719 5973 41728
rect 5835 41600 5877 41609
rect 5835 41560 5836 41600
rect 5876 41560 5877 41600
rect 5835 41551 5877 41560
rect 5739 41432 5781 41441
rect 5739 41392 5740 41432
rect 5780 41392 5781 41432
rect 5739 41383 5781 41392
rect 5548 41140 5780 41180
rect 5547 40844 5589 40853
rect 5547 40804 5548 40844
rect 5588 40804 5589 40844
rect 5547 40795 5589 40804
rect 5108 39880 5492 39920
rect 5068 39871 5108 39880
rect 5067 39752 5109 39761
rect 5067 39712 5068 39752
rect 5108 39712 5109 39752
rect 5067 39703 5109 39712
rect 5356 39752 5396 39761
rect 4875 39668 4917 39677
rect 4875 39628 4876 39668
rect 4916 39628 4917 39668
rect 4875 39619 4917 39628
rect 4876 39534 4916 39619
rect 5068 38912 5108 39703
rect 5259 39500 5301 39509
rect 5259 39460 5260 39500
rect 5300 39460 5301 39500
rect 5259 39451 5301 39460
rect 5260 39366 5300 39451
rect 5356 39173 5396 39712
rect 5355 39164 5397 39173
rect 5355 39124 5356 39164
rect 5396 39124 5397 39164
rect 5355 39115 5397 39124
rect 5548 38926 5588 40795
rect 5643 40508 5685 40517
rect 5643 40468 5644 40508
rect 5684 40468 5685 40508
rect 5740 40508 5780 41140
rect 5836 40676 5876 41551
rect 5836 40627 5876 40636
rect 5740 40468 5876 40508
rect 5643 40459 5685 40468
rect 5644 40374 5684 40459
rect 5548 38877 5588 38886
rect 5644 39752 5684 39761
rect 5068 38863 5108 38872
rect 4928 38576 5296 38585
rect 4968 38536 5010 38576
rect 5050 38536 5092 38576
rect 5132 38536 5174 38576
rect 5214 38536 5256 38576
rect 4928 38527 5296 38536
rect 5067 38240 5109 38249
rect 5067 38200 5068 38240
rect 5108 38200 5109 38240
rect 5067 38191 5109 38200
rect 5068 38106 5108 38191
rect 4875 38072 4917 38081
rect 4875 38032 4876 38072
rect 4916 38032 4917 38072
rect 4875 38023 4917 38032
rect 4876 37938 4916 38023
rect 5644 37820 5684 39712
rect 5739 39752 5781 39761
rect 5739 39712 5740 39752
rect 5780 39712 5781 39752
rect 5739 39703 5781 39712
rect 5740 39618 5780 39703
rect 5836 39257 5876 40468
rect 5932 39416 5972 41719
rect 6220 41600 6260 42928
rect 6315 41768 6357 41777
rect 6315 41728 6316 41768
rect 6356 41728 6357 41768
rect 6315 41719 6357 41728
rect 6124 41560 6260 41600
rect 6027 41348 6069 41357
rect 6027 41308 6028 41348
rect 6068 41308 6069 41348
rect 6027 41299 6069 41308
rect 6028 40424 6068 41299
rect 6028 40375 6068 40384
rect 6124 40256 6164 41560
rect 6219 41432 6261 41441
rect 6219 41392 6220 41432
rect 6260 41392 6261 41432
rect 6219 41383 6261 41392
rect 6220 41264 6260 41383
rect 6220 41215 6260 41224
rect 6316 41096 6356 41719
rect 6412 41180 6452 42928
rect 6604 41441 6644 42928
rect 6699 42524 6741 42533
rect 6699 42484 6700 42524
rect 6740 42484 6741 42524
rect 6699 42475 6741 42484
rect 6603 41432 6645 41441
rect 6603 41392 6604 41432
rect 6644 41392 6645 41432
rect 6603 41383 6645 41392
rect 6603 41264 6645 41273
rect 6603 41224 6604 41264
rect 6644 41224 6645 41264
rect 6603 41215 6645 41224
rect 6412 41140 6548 41180
rect 6028 40216 6164 40256
rect 6220 41056 6356 41096
rect 6028 39500 6068 40216
rect 6220 39845 6260 41056
rect 6412 41012 6452 41021
rect 6412 40433 6452 40972
rect 6508 40844 6548 41140
rect 6604 41130 6644 41215
rect 6508 40804 6644 40844
rect 6411 40424 6453 40433
rect 6411 40384 6412 40424
rect 6452 40384 6453 40424
rect 6411 40375 6453 40384
rect 6219 39836 6261 39845
rect 6219 39796 6220 39836
rect 6260 39796 6261 39836
rect 6219 39787 6261 39796
rect 6124 39677 6164 39762
rect 6123 39668 6165 39677
rect 6123 39628 6124 39668
rect 6164 39628 6165 39668
rect 6123 39619 6165 39628
rect 6220 39668 6260 39677
rect 6028 39460 6164 39500
rect 5932 39376 6068 39416
rect 5835 39248 5877 39257
rect 5835 39208 5836 39248
rect 5876 39208 5877 39248
rect 5835 39199 5877 39208
rect 5932 38912 5972 38921
rect 5740 38744 5780 38753
rect 5780 38704 5876 38744
rect 5740 38695 5780 38704
rect 5739 37988 5781 37997
rect 5739 37948 5740 37988
rect 5780 37948 5781 37988
rect 5739 37939 5781 37948
rect 5548 37780 5684 37820
rect 5259 37736 5301 37745
rect 5259 37696 5260 37736
rect 5300 37696 5301 37736
rect 5259 37687 5301 37696
rect 5260 37577 5300 37687
rect 5259 37568 5301 37577
rect 5259 37528 5260 37568
rect 5300 37528 5301 37568
rect 5259 37519 5301 37528
rect 5451 37568 5493 37577
rect 5451 37528 5452 37568
rect 5492 37528 5493 37568
rect 5451 37519 5493 37528
rect 4924 37414 4964 37418
rect 4780 37409 4964 37414
rect 4780 37374 4924 37409
rect 4924 37360 4964 37369
rect 5452 37400 5492 37519
rect 5452 37351 5492 37360
rect 4780 37232 4820 37241
rect 4588 36847 4628 36856
rect 4684 37192 4780 37232
rect 3339 36560 3381 36569
rect 3532 36560 3572 36604
rect 3820 36595 3860 36604
rect 4108 36772 4244 36812
rect 3339 36520 3340 36560
rect 3380 36520 3381 36560
rect 3339 36511 3381 36520
rect 3436 36520 3572 36560
rect 3244 35176 3380 35216
rect 3147 35167 3189 35176
rect 2908 35132 2948 35134
rect 3051 35132 3093 35141
rect 2908 35092 2996 35132
rect 2763 34628 2805 34637
rect 2763 34588 2764 34628
rect 2804 34588 2805 34628
rect 2763 34579 2805 34588
rect 2667 34376 2709 34385
rect 2667 34336 2668 34376
rect 2708 34336 2709 34376
rect 2667 34327 2709 34336
rect 2860 34376 2900 34387
rect 2571 33956 2613 33965
rect 2571 33916 2572 33956
rect 2612 33916 2613 33956
rect 2571 33907 2613 33916
rect 2283 33872 2325 33881
rect 2283 33832 2284 33872
rect 2324 33832 2325 33872
rect 2283 33823 2325 33832
rect 2668 33788 2708 34327
rect 2860 34301 2900 34336
rect 2859 34292 2901 34301
rect 2859 34252 2860 34292
rect 2900 34252 2901 34292
rect 2859 34243 2901 34252
rect 2956 33797 2996 35092
rect 3051 35092 3052 35132
rect 3092 35092 3093 35132
rect 3051 35083 3093 35092
rect 3148 34469 3188 35167
rect 3244 35048 3284 35057
rect 3244 34637 3284 35008
rect 3340 34973 3380 35176
rect 3339 34964 3381 34973
rect 3339 34924 3340 34964
rect 3380 34924 3381 34964
rect 3339 34915 3381 34924
rect 3243 34628 3285 34637
rect 3243 34588 3244 34628
rect 3284 34588 3285 34628
rect 3243 34579 3285 34588
rect 3436 34544 3476 36520
rect 3628 36476 3668 36485
rect 3532 36436 3628 36476
rect 3532 35477 3572 36436
rect 3628 36427 3668 36436
rect 3688 36308 4056 36317
rect 3728 36268 3770 36308
rect 3810 36268 3852 36308
rect 3892 36268 3934 36308
rect 3974 36268 4016 36308
rect 3688 36259 4056 36268
rect 4012 36140 4052 36149
rect 4108 36140 4148 36772
rect 4684 36728 4724 37192
rect 4780 37183 4820 37192
rect 4928 37064 5296 37073
rect 4968 37024 5010 37064
rect 5050 37024 5092 37064
rect 5132 37024 5174 37064
rect 5214 37024 5256 37064
rect 4928 37015 5296 37024
rect 4492 36688 4724 36728
rect 4052 36100 4148 36140
rect 4204 36644 4244 36653
rect 4012 36091 4052 36100
rect 3819 36056 3861 36065
rect 3819 36016 3820 36056
rect 3860 36016 3861 36056
rect 3819 36007 3861 36016
rect 3820 35972 3860 36007
rect 3628 35888 3668 35897
rect 3628 35561 3668 35848
rect 3820 35813 3860 35932
rect 4204 35897 4244 36604
rect 4299 36560 4341 36569
rect 4299 36520 4300 36560
rect 4340 36520 4341 36560
rect 4299 36511 4341 36520
rect 4203 35888 4245 35897
rect 4203 35848 4204 35888
rect 4244 35848 4245 35888
rect 4203 35839 4245 35848
rect 4300 35888 4340 36511
rect 4300 35839 4340 35848
rect 4395 35888 4437 35897
rect 4395 35848 4396 35888
rect 4436 35848 4437 35888
rect 4395 35839 4437 35848
rect 3819 35804 3861 35813
rect 3819 35764 3820 35804
rect 3860 35764 3861 35804
rect 3819 35755 3861 35764
rect 4396 35754 4436 35839
rect 4299 35636 4341 35645
rect 4299 35596 4300 35636
rect 4340 35596 4341 35636
rect 4299 35587 4341 35596
rect 3627 35552 3669 35561
rect 3627 35512 3628 35552
rect 3668 35512 3669 35552
rect 3627 35503 3669 35512
rect 3531 35468 3573 35477
rect 3531 35428 3532 35468
rect 3572 35428 3573 35468
rect 3531 35419 3573 35428
rect 3819 35384 3861 35393
rect 3819 35344 3820 35384
rect 3860 35344 3861 35384
rect 3819 35335 3861 35344
rect 3820 35141 3860 35335
rect 4012 35216 4052 35225
rect 3916 35176 4012 35216
rect 3723 35132 3765 35141
rect 3723 35092 3724 35132
rect 3764 35092 3765 35132
rect 3820 35132 3868 35141
rect 3820 35092 3827 35132
rect 3867 35092 3868 35132
rect 3723 35083 3765 35092
rect 3826 35083 3868 35092
rect 3724 34998 3764 35083
rect 3916 34973 3956 35176
rect 4012 35167 4052 35176
rect 4203 35216 4245 35225
rect 4203 35176 4204 35216
rect 4244 35176 4245 35216
rect 4203 35167 4245 35176
rect 4204 35082 4244 35167
rect 4059 35048 4101 35057
rect 4022 35008 4060 35048
rect 4100 35008 4101 35048
rect 4022 34999 4101 35008
rect 4022 34973 4062 34999
rect 3531 34964 3573 34973
rect 3531 34924 3532 34964
rect 3572 34924 3573 34964
rect 3531 34915 3573 34924
rect 3915 34964 3957 34973
rect 3915 34924 3916 34964
rect 3956 34924 3957 34964
rect 3915 34915 3957 34924
rect 4012 34964 4062 34973
rect 4052 34924 4062 34964
rect 4012 34915 4052 34924
rect 3532 34830 3572 34915
rect 3688 34796 4056 34805
rect 3728 34756 3770 34796
rect 3810 34756 3852 34796
rect 3892 34756 3934 34796
rect 3974 34756 4016 34796
rect 3688 34747 4056 34756
rect 3436 34504 3572 34544
rect 3147 34460 3189 34469
rect 3147 34420 3148 34460
rect 3188 34420 3189 34460
rect 3147 34411 3189 34420
rect 3340 34376 3380 34385
rect 3340 34208 3380 34336
rect 3435 34376 3477 34385
rect 3435 34336 3436 34376
rect 3476 34336 3477 34376
rect 3435 34327 3477 34336
rect 3436 34242 3476 34327
rect 3052 34168 3380 34208
rect 2572 33748 2708 33788
rect 2955 33788 2997 33797
rect 2955 33748 2956 33788
rect 2996 33748 2997 33788
rect 2572 33116 2612 33748
rect 2955 33739 2997 33748
rect 2860 33704 2900 33713
rect 2561 33076 2612 33116
rect 2668 33664 2860 33704
rect 2561 33032 2601 33076
rect 2476 32992 2601 33032
rect 2283 32696 2325 32705
rect 2283 32656 2284 32696
rect 2324 32656 2325 32696
rect 2283 32647 2325 32656
rect 2092 31900 2228 31940
rect 2092 31394 2132 31900
rect 2188 31529 2228 31614
rect 2187 31520 2229 31529
rect 2187 31480 2188 31520
rect 2228 31480 2229 31520
rect 2187 31471 2229 31480
rect 1900 31352 2036 31361
rect 1940 31321 2036 31352
rect 2092 31345 2132 31354
rect 2188 31352 2228 31361
rect 2284 31352 2324 32647
rect 2476 32528 2516 32992
rect 2572 32864 2612 32873
rect 2668 32864 2708 33664
rect 2860 33655 2900 33664
rect 3052 33620 3092 34168
rect 3147 34040 3189 34049
rect 3147 34000 3148 34040
rect 3188 34000 3189 34040
rect 3147 33991 3189 34000
rect 2956 33580 3092 33620
rect 2859 33284 2901 33293
rect 2859 33244 2860 33284
rect 2900 33244 2901 33284
rect 2859 33235 2901 33244
rect 2612 32824 2708 32864
rect 2572 32815 2612 32824
rect 2476 32488 2612 32528
rect 2572 32369 2612 32488
rect 2571 32360 2613 32369
rect 2571 32320 2572 32360
rect 2612 32320 2613 32360
rect 2571 32311 2613 32320
rect 2476 32108 2516 32117
rect 1900 31303 1940 31312
rect 1996 31268 2036 31321
rect 2228 31312 2324 31352
rect 2380 31352 2420 31361
rect 2188 31268 2228 31312
rect 1996 31228 2228 31268
rect 1804 31184 1844 31193
rect 2380 31184 2420 31312
rect 1804 30773 1844 31144
rect 2284 31144 2420 31184
rect 2187 31100 2229 31109
rect 2187 31060 2188 31100
rect 2228 31060 2229 31100
rect 2187 31051 2229 31060
rect 2091 30848 2133 30857
rect 2091 30808 2092 30848
rect 2132 30808 2133 30848
rect 2091 30799 2133 30808
rect 1803 30764 1845 30773
rect 1803 30724 1804 30764
rect 1844 30724 1845 30764
rect 1803 30715 1845 30724
rect 1707 30260 1749 30269
rect 1707 30220 1708 30260
rect 1748 30220 1749 30260
rect 1707 30211 1749 30220
rect 1803 30176 1845 30185
rect 1803 30136 1804 30176
rect 1844 30136 1845 30176
rect 1803 30127 1845 30136
rect 1707 30092 1749 30101
rect 1707 30052 1708 30092
rect 1748 30052 1749 30092
rect 1707 30043 1749 30052
rect 1420 29119 1460 29128
rect 1516 29093 1556 29178
rect 1611 29168 1653 29177
rect 1611 29128 1612 29168
rect 1652 29128 1653 29168
rect 1611 29119 1653 29128
rect 1515 29084 1557 29093
rect 1515 29044 1516 29084
rect 1556 29044 1557 29084
rect 1515 29035 1557 29044
rect 1612 29000 1652 29119
rect 1708 29084 1748 30043
rect 1804 29168 1844 30127
rect 2092 30017 2132 30799
rect 2091 30008 2133 30017
rect 2091 29968 2092 30008
rect 2132 29968 2133 30008
rect 2091 29959 2133 29968
rect 1804 29119 1844 29128
rect 1996 29168 2036 29177
rect 2036 29128 2132 29168
rect 1996 29119 2036 29128
rect 1708 29035 1748 29044
rect 1324 28960 1460 29000
rect 1131 28951 1173 28960
rect 1035 28244 1077 28253
rect 1035 28204 1036 28244
rect 1076 28204 1077 28244
rect 1035 28195 1077 28204
rect 939 25640 981 25649
rect 939 25600 940 25640
rect 980 25600 981 25640
rect 939 25591 981 25600
rect 843 24044 885 24053
rect 843 24004 844 24044
rect 884 24004 885 24044
rect 843 23995 885 24004
rect 651 23960 693 23969
rect 651 23920 652 23960
rect 692 23920 693 23960
rect 651 23911 693 23920
rect 459 23624 501 23633
rect 459 23584 460 23624
rect 500 23584 501 23624
rect 459 23575 501 23584
rect 555 22868 597 22877
rect 555 22828 556 22868
rect 596 22828 597 22868
rect 555 22819 597 22828
rect 171 21356 213 21365
rect 171 21316 172 21356
rect 212 21316 213 21356
rect 171 21307 213 21316
rect 172 12545 212 21307
rect 267 14132 309 14141
rect 267 14092 268 14132
rect 308 14092 309 14132
rect 267 14083 309 14092
rect 171 12536 213 12545
rect 171 12496 172 12536
rect 212 12496 213 12536
rect 171 12487 213 12496
rect 171 10184 213 10193
rect 171 10144 172 10184
rect 212 10144 213 10184
rect 171 10135 213 10144
rect 172 944 212 10135
rect 268 5825 308 14083
rect 459 13880 501 13889
rect 459 13840 460 13880
rect 500 13840 501 13880
rect 459 13831 501 13840
rect 363 12620 405 12629
rect 363 12580 364 12620
rect 404 12580 405 12620
rect 363 12571 405 12580
rect 364 10361 404 12571
rect 363 10352 405 10361
rect 363 10312 364 10352
rect 404 10312 405 10352
rect 363 10303 405 10312
rect 460 8849 500 13831
rect 556 11873 596 22819
rect 940 18677 980 25591
rect 1035 23036 1077 23045
rect 1035 22996 1036 23036
rect 1076 22996 1077 23036
rect 1035 22987 1077 22996
rect 939 18668 981 18677
rect 939 18628 940 18668
rect 980 18628 981 18668
rect 939 18619 981 18628
rect 939 13208 981 13217
rect 939 13168 940 13208
rect 980 13168 981 13208
rect 939 13159 981 13168
rect 747 13040 789 13049
rect 747 13000 748 13040
rect 788 13000 789 13040
rect 747 12991 789 13000
rect 651 12788 693 12797
rect 651 12748 652 12788
rect 692 12748 693 12788
rect 651 12739 693 12748
rect 555 11864 597 11873
rect 555 11824 556 11864
rect 596 11824 597 11864
rect 555 11815 597 11824
rect 459 8840 501 8849
rect 459 8800 460 8840
rect 500 8800 501 8840
rect 459 8791 501 8800
rect 555 7580 597 7589
rect 555 7540 556 7580
rect 596 7540 597 7580
rect 555 7531 597 7540
rect 267 5816 309 5825
rect 267 5776 268 5816
rect 308 5776 309 5816
rect 267 5767 309 5776
rect 556 2549 596 7531
rect 652 6497 692 12739
rect 748 7505 788 12991
rect 940 11360 980 13159
rect 1036 11621 1076 22987
rect 1035 11612 1077 11621
rect 1035 11572 1036 11612
rect 1076 11572 1077 11612
rect 1035 11563 1077 11572
rect 940 11320 1076 11360
rect 939 11192 981 11201
rect 939 11152 940 11192
rect 980 11152 981 11192
rect 939 11143 981 11152
rect 843 9512 885 9521
rect 843 9472 844 9512
rect 884 9472 885 9512
rect 843 9463 885 9472
rect 747 7496 789 7505
rect 747 7456 748 7496
rect 788 7456 789 7496
rect 747 7447 789 7456
rect 844 7160 884 9463
rect 940 8000 980 11143
rect 1036 8168 1076 11320
rect 1132 10865 1172 28951
rect 1323 28160 1365 28169
rect 1323 28120 1324 28160
rect 1364 28120 1365 28160
rect 1323 28111 1365 28120
rect 1324 28026 1364 28111
rect 1323 27740 1365 27749
rect 1228 27700 1324 27740
rect 1364 27700 1365 27740
rect 1228 27656 1268 27700
rect 1323 27691 1365 27700
rect 1228 27607 1268 27616
rect 1323 27404 1365 27413
rect 1323 27364 1324 27404
rect 1364 27364 1365 27404
rect 1323 27355 1365 27364
rect 1227 26816 1269 26825
rect 1227 26776 1228 26816
rect 1268 26776 1269 26816
rect 1227 26767 1269 26776
rect 1228 26682 1268 26767
rect 1324 26144 1364 27355
rect 1420 26648 1460 28960
rect 1612 28951 1652 28960
rect 1995 29000 2037 29009
rect 1995 28960 1996 29000
rect 2036 28960 2037 29000
rect 1995 28951 2037 28960
rect 1707 28916 1749 28925
rect 1707 28876 1708 28916
rect 1748 28876 1749 28916
rect 1707 28867 1749 28876
rect 1708 28337 1748 28867
rect 1899 28496 1941 28505
rect 1899 28456 1900 28496
rect 1940 28456 1941 28496
rect 1899 28447 1941 28456
rect 1707 28328 1749 28337
rect 1707 28288 1708 28328
rect 1748 28288 1749 28328
rect 1707 28279 1749 28288
rect 1611 28160 1653 28169
rect 1611 28120 1612 28160
rect 1652 28120 1653 28160
rect 1611 28111 1653 28120
rect 1420 26608 1556 26648
rect 1419 26480 1461 26489
rect 1419 26440 1420 26480
rect 1460 26440 1461 26480
rect 1419 26431 1461 26440
rect 1324 26095 1364 26104
rect 1227 26060 1269 26069
rect 1227 26020 1228 26060
rect 1268 26020 1269 26060
rect 1227 26011 1269 26020
rect 1228 25926 1268 26011
rect 1323 25388 1365 25397
rect 1228 25348 1324 25388
rect 1364 25348 1365 25388
rect 1228 25304 1268 25348
rect 1323 25339 1365 25348
rect 1228 25255 1268 25264
rect 1420 24800 1460 26431
rect 1324 24760 1460 24800
rect 1516 26144 1556 26608
rect 1324 23288 1364 24760
rect 1419 24632 1461 24641
rect 1419 24592 1420 24632
rect 1460 24592 1461 24632
rect 1419 24583 1461 24592
rect 1420 24498 1460 24583
rect 1324 22541 1364 23248
rect 1420 23624 1460 23633
rect 1420 22709 1460 23584
rect 1516 23213 1556 26104
rect 1612 24968 1652 28111
rect 1708 25145 1748 28279
rect 1803 27824 1845 27833
rect 1803 27784 1804 27824
rect 1844 27784 1845 27824
rect 1803 27775 1845 27784
rect 1804 26909 1844 27775
rect 1803 26900 1845 26909
rect 1803 26860 1804 26900
rect 1844 26860 1845 26900
rect 1803 26851 1845 26860
rect 1707 25136 1749 25145
rect 1707 25096 1708 25136
rect 1748 25096 1749 25136
rect 1707 25087 1749 25096
rect 1612 24928 1748 24968
rect 1611 23876 1653 23885
rect 1611 23836 1612 23876
rect 1652 23836 1653 23876
rect 1611 23827 1653 23836
rect 1612 23742 1652 23827
rect 1708 23381 1748 24928
rect 1707 23372 1749 23381
rect 1707 23332 1708 23372
rect 1748 23332 1749 23372
rect 1707 23323 1749 23332
rect 1515 23204 1557 23213
rect 1515 23164 1516 23204
rect 1556 23164 1557 23204
rect 1515 23155 1557 23164
rect 1516 23036 1556 23155
rect 1707 23036 1749 23045
rect 1516 22996 1652 23036
rect 1515 22868 1557 22877
rect 1515 22828 1516 22868
rect 1556 22828 1557 22868
rect 1515 22819 1557 22828
rect 1516 22734 1556 22819
rect 1419 22700 1461 22709
rect 1419 22660 1420 22700
rect 1460 22660 1461 22700
rect 1419 22651 1461 22660
rect 1323 22532 1365 22541
rect 1323 22492 1324 22532
rect 1364 22492 1365 22532
rect 1323 22483 1365 22492
rect 1612 22364 1652 22996
rect 1707 22996 1708 23036
rect 1748 22996 1749 23036
rect 1707 22987 1749 22996
rect 1708 22902 1748 22987
rect 1804 22625 1844 26851
rect 1900 24800 1940 28447
rect 1996 28328 2036 28951
rect 2092 28841 2132 29128
rect 2091 28832 2133 28841
rect 2091 28792 2092 28832
rect 2132 28792 2133 28832
rect 2091 28783 2133 28792
rect 1996 28279 2036 28288
rect 2092 28328 2132 28337
rect 2092 26405 2132 28288
rect 2188 26825 2228 31051
rect 2284 30521 2324 31144
rect 2476 30857 2516 32068
rect 2572 32108 2612 32117
rect 2572 31865 2612 32068
rect 2571 31856 2613 31865
rect 2571 31816 2572 31856
rect 2612 31816 2613 31856
rect 2571 31807 2613 31816
rect 2572 31613 2612 31807
rect 2571 31604 2613 31613
rect 2571 31564 2572 31604
rect 2612 31564 2613 31604
rect 2571 31555 2613 31564
rect 2572 31352 2612 31361
rect 2572 31193 2612 31312
rect 2571 31184 2613 31193
rect 2571 31144 2572 31184
rect 2612 31144 2613 31184
rect 2571 31135 2613 31144
rect 2668 31016 2708 32824
rect 2763 32696 2805 32705
rect 2763 32656 2764 32696
rect 2804 32656 2805 32696
rect 2763 32647 2805 32656
rect 2764 32562 2804 32647
rect 2763 32192 2805 32201
rect 2860 32192 2900 33235
rect 2956 33041 2996 33580
rect 3052 33452 3092 33461
rect 3052 33293 3092 33412
rect 3051 33284 3093 33293
rect 3051 33244 3052 33284
rect 3092 33244 3093 33284
rect 3051 33235 3093 33244
rect 2955 33032 2997 33041
rect 2955 32992 2956 33032
rect 2996 32992 2997 33032
rect 2955 32983 2997 32992
rect 3052 32864 3092 32873
rect 2955 32696 2997 32705
rect 2955 32656 2956 32696
rect 2996 32656 2997 32696
rect 2955 32647 2997 32656
rect 2956 32562 2996 32647
rect 3052 32453 3092 32824
rect 3051 32444 3093 32453
rect 3051 32404 3052 32444
rect 3092 32404 3093 32444
rect 3051 32395 3093 32404
rect 3148 32369 3188 33991
rect 3532 33704 3572 34504
rect 3820 34376 3860 34385
rect 3820 33965 3860 34336
rect 3915 34376 3957 34385
rect 3915 34336 3916 34376
rect 3956 34336 3957 34376
rect 3915 34327 3957 34336
rect 4204 34376 4244 34385
rect 4300 34376 4340 35587
rect 4395 35468 4437 35477
rect 4395 35428 4396 35468
rect 4436 35428 4437 35468
rect 4395 35419 4437 35428
rect 4396 35216 4436 35419
rect 4492 35393 4532 36688
rect 4780 36644 4820 36653
rect 4684 36604 4780 36644
rect 4587 35888 4629 35897
rect 4587 35848 4588 35888
rect 4628 35848 4629 35888
rect 4587 35839 4629 35848
rect 4491 35384 4533 35393
rect 4491 35344 4492 35384
rect 4532 35344 4533 35384
rect 4491 35335 4533 35344
rect 4588 35300 4628 35839
rect 4684 35384 4724 36604
rect 4780 36595 4820 36604
rect 5068 36644 5108 36653
rect 5068 36485 5108 36604
rect 5451 36644 5493 36653
rect 5451 36604 5452 36644
rect 5492 36604 5493 36644
rect 5451 36595 5493 36604
rect 5259 36560 5301 36569
rect 5259 36520 5260 36560
rect 5300 36520 5301 36560
rect 5259 36511 5301 36520
rect 5067 36476 5109 36485
rect 5067 36436 5068 36476
rect 5108 36436 5109 36476
rect 5067 36427 5109 36436
rect 5260 36426 5300 36511
rect 5452 36510 5492 36595
rect 5355 36476 5397 36485
rect 5355 36436 5356 36476
rect 5396 36436 5397 36476
rect 5355 36427 5397 36436
rect 4875 36140 4917 36149
rect 4875 36100 4876 36140
rect 4916 36100 4917 36140
rect 4875 36091 4917 36100
rect 4876 35972 4916 36091
rect 4876 35923 4916 35932
rect 4780 35888 4820 35897
rect 4780 35729 4820 35848
rect 5356 35888 5396 36427
rect 5356 35839 5396 35848
rect 4779 35720 4821 35729
rect 4779 35680 4780 35720
rect 4820 35680 4821 35720
rect 4779 35671 4821 35680
rect 4928 35552 5296 35561
rect 4968 35512 5010 35552
rect 5050 35512 5092 35552
rect 5132 35512 5174 35552
rect 5214 35512 5256 35552
rect 4928 35503 5296 35512
rect 4684 35344 4820 35384
rect 4588 35251 4628 35260
rect 4396 35167 4436 35176
rect 4492 35216 4532 35225
rect 4492 35141 4532 35176
rect 4684 35216 4724 35225
rect 4491 35132 4533 35141
rect 4491 35092 4492 35132
rect 4532 35092 4533 35132
rect 4491 35083 4533 35092
rect 4395 34964 4437 34973
rect 4395 34924 4396 34964
rect 4436 34924 4437 34964
rect 4395 34915 4437 34924
rect 4244 34336 4340 34376
rect 4204 34327 4244 34336
rect 3916 34242 3956 34327
rect 4203 34208 4245 34217
rect 4203 34168 4204 34208
rect 4244 34168 4245 34208
rect 4203 34159 4245 34168
rect 3627 33956 3669 33965
rect 3627 33916 3628 33956
rect 3668 33916 3669 33956
rect 3627 33907 3669 33916
rect 3819 33956 3861 33965
rect 3819 33916 3820 33956
rect 3860 33916 3861 33956
rect 3819 33907 3861 33916
rect 3628 33872 3668 33907
rect 3628 33821 3668 33832
rect 4107 33872 4149 33881
rect 4107 33832 4108 33872
rect 4148 33832 4149 33872
rect 4107 33823 4149 33832
rect 4108 33738 4148 33823
rect 3532 33664 3671 33704
rect 3244 33620 3284 33629
rect 3244 33041 3284 33580
rect 3531 33536 3573 33545
rect 3436 33496 3532 33536
rect 3572 33496 3573 33536
rect 3436 33452 3476 33496
rect 3531 33487 3573 33496
rect 3631 33452 3671 33664
rect 3819 33620 3861 33629
rect 3819 33580 3820 33620
rect 3860 33580 3861 33620
rect 3819 33571 3861 33580
rect 3820 33486 3860 33571
rect 3436 33403 3476 33412
rect 3623 33412 3671 33452
rect 3623 33368 3663 33412
rect 3532 33328 3663 33368
rect 3435 33284 3477 33293
rect 3435 33244 3436 33284
rect 3476 33244 3477 33284
rect 3435 33235 3477 33244
rect 3436 33116 3476 33235
rect 3436 33067 3476 33076
rect 3243 33032 3285 33041
rect 3243 32992 3244 33032
rect 3284 32992 3285 33032
rect 3243 32983 3285 32992
rect 3244 32864 3284 32873
rect 3244 32453 3284 32824
rect 3435 32864 3477 32873
rect 3435 32824 3436 32864
rect 3476 32824 3477 32864
rect 3435 32815 3477 32824
rect 3436 32730 3476 32815
rect 3243 32444 3285 32453
rect 3243 32404 3244 32444
rect 3284 32404 3285 32444
rect 3243 32395 3285 32404
rect 2955 32360 2997 32369
rect 2955 32320 2956 32360
rect 2996 32320 2997 32360
rect 2955 32311 2997 32320
rect 3147 32360 3189 32369
rect 3147 32320 3148 32360
rect 3188 32320 3189 32360
rect 3147 32311 3189 32320
rect 2763 32152 2764 32192
rect 2804 32152 2900 32192
rect 2763 32143 2805 32152
rect 2572 30976 2708 31016
rect 2475 30848 2517 30857
rect 2475 30808 2476 30848
rect 2516 30808 2517 30848
rect 2475 30799 2517 30808
rect 2476 30680 2516 30691
rect 2476 30605 2516 30640
rect 2572 30605 2612 30976
rect 2667 30764 2709 30773
rect 2667 30724 2668 30764
rect 2708 30724 2709 30764
rect 2667 30715 2709 30724
rect 2475 30596 2517 30605
rect 2475 30556 2476 30596
rect 2516 30556 2517 30596
rect 2475 30547 2517 30556
rect 2571 30596 2613 30605
rect 2571 30556 2572 30596
rect 2612 30556 2613 30596
rect 2571 30547 2613 30556
rect 2668 30521 2708 30715
rect 2283 30512 2325 30521
rect 2283 30472 2284 30512
rect 2324 30472 2325 30512
rect 2283 30463 2325 30472
rect 2667 30512 2709 30521
rect 2667 30472 2668 30512
rect 2708 30472 2709 30512
rect 2667 30463 2709 30472
rect 2571 30428 2613 30437
rect 2571 30388 2572 30428
rect 2612 30388 2613 30428
rect 2571 30379 2613 30388
rect 2379 30260 2421 30269
rect 2379 30220 2380 30260
rect 2420 30220 2421 30260
rect 2379 30211 2421 30220
rect 2283 29756 2325 29765
rect 2283 29716 2284 29756
rect 2324 29716 2325 29756
rect 2283 29707 2325 29716
rect 2187 26816 2229 26825
rect 2187 26776 2188 26816
rect 2228 26776 2229 26816
rect 2187 26767 2229 26776
rect 2091 26396 2133 26405
rect 2091 26356 2092 26396
rect 2132 26356 2133 26396
rect 2091 26347 2133 26356
rect 1900 24760 2132 24800
rect 1995 24632 2037 24641
rect 1995 24592 1996 24632
rect 2036 24592 2037 24632
rect 1995 24583 2037 24592
rect 1899 23792 1941 23801
rect 1899 23752 1900 23792
rect 1940 23752 1941 23792
rect 1899 23743 1941 23752
rect 1900 23658 1940 23743
rect 1900 23120 1940 23129
rect 1803 22616 1845 22625
rect 1803 22576 1804 22616
rect 1844 22576 1845 22616
rect 1803 22567 1845 22576
rect 1516 22324 1652 22364
rect 1228 22280 1268 22289
rect 1516 22280 1556 22324
rect 1268 22240 1556 22280
rect 1707 22280 1749 22289
rect 1707 22240 1708 22280
rect 1748 22240 1749 22280
rect 1228 22231 1268 22240
rect 1707 22231 1749 22240
rect 1419 21692 1461 21701
rect 1419 21652 1420 21692
rect 1460 21652 1461 21692
rect 1419 21643 1461 21652
rect 1420 21524 1460 21643
rect 1611 21608 1653 21617
rect 1611 21568 1612 21608
rect 1652 21568 1653 21608
rect 1611 21559 1653 21568
rect 1420 21475 1460 21484
rect 1612 21474 1652 21559
rect 1227 21356 1269 21365
rect 1227 21316 1228 21356
rect 1268 21316 1269 21356
rect 1227 21307 1269 21316
rect 1228 21222 1268 21307
rect 1228 20768 1268 20777
rect 1323 20768 1365 20777
rect 1268 20728 1324 20768
rect 1364 20728 1365 20768
rect 1228 20719 1268 20728
rect 1323 20719 1365 20728
rect 1515 20348 1557 20357
rect 1515 20308 1516 20348
rect 1556 20308 1557 20348
rect 1515 20299 1557 20308
rect 1228 20096 1268 20105
rect 1268 20056 1364 20096
rect 1228 20047 1268 20056
rect 1324 19769 1364 20056
rect 1323 19760 1365 19769
rect 1323 19720 1324 19760
rect 1364 19720 1365 19760
rect 1323 19711 1365 19720
rect 1516 19340 1556 20299
rect 1708 20180 1748 22231
rect 1900 20693 1940 23080
rect 1899 20684 1941 20693
rect 1899 20644 1900 20684
rect 1940 20644 1941 20684
rect 1899 20635 1941 20644
rect 1516 19291 1556 19300
rect 1612 20140 1748 20180
rect 1324 19088 1364 19097
rect 1228 18584 1268 18595
rect 1228 18509 1268 18544
rect 1227 18500 1269 18509
rect 1227 18460 1228 18500
rect 1268 18460 1269 18500
rect 1227 18451 1269 18460
rect 1227 18248 1269 18257
rect 1227 18208 1228 18248
rect 1268 18208 1269 18248
rect 1227 18199 1269 18208
rect 1228 17837 1268 18199
rect 1227 17828 1269 17837
rect 1227 17788 1228 17828
rect 1268 17788 1269 17828
rect 1227 17779 1269 17788
rect 1228 17694 1268 17779
rect 1324 17333 1364 19048
rect 1515 18500 1557 18509
rect 1515 18460 1516 18500
rect 1556 18460 1557 18500
rect 1515 18451 1557 18460
rect 1516 17753 1556 18451
rect 1515 17744 1557 17753
rect 1515 17704 1516 17744
rect 1556 17704 1557 17744
rect 1515 17695 1557 17704
rect 1516 17610 1556 17695
rect 1323 17324 1365 17333
rect 1323 17284 1324 17324
rect 1364 17284 1365 17324
rect 1323 17275 1365 17284
rect 1612 17165 1652 20140
rect 1708 19256 1748 19267
rect 1708 19181 1748 19216
rect 1707 19172 1749 19181
rect 1707 19132 1708 19172
rect 1748 19132 1749 19172
rect 1707 19123 1749 19132
rect 1996 17912 2036 24583
rect 2092 22037 2132 24760
rect 2284 24221 2324 29707
rect 2380 28505 2420 30211
rect 2476 29840 2516 29849
rect 2476 29177 2516 29800
rect 2475 29168 2517 29177
rect 2475 29128 2476 29168
rect 2516 29128 2517 29168
rect 2475 29119 2517 29128
rect 2379 28496 2421 28505
rect 2379 28456 2380 28496
rect 2420 28456 2421 28496
rect 2379 28447 2421 28456
rect 2572 28412 2612 30379
rect 2764 30344 2804 32143
rect 2956 31781 2996 32311
rect 3532 32276 3572 33328
rect 3688 33284 4056 33293
rect 3728 33244 3770 33284
rect 3810 33244 3852 33284
rect 3892 33244 3934 33284
rect 3974 33244 4016 33284
rect 3688 33235 4056 33244
rect 3819 33116 3861 33125
rect 4204 33116 4244 34159
rect 4300 33690 4340 33699
rect 4300 33125 4340 33650
rect 4396 33377 4436 34915
rect 4492 34217 4532 35083
rect 4684 35057 4724 35176
rect 4683 35048 4725 35057
rect 4683 35008 4684 35048
rect 4724 35008 4725 35048
rect 4683 34999 4725 35008
rect 4683 34796 4725 34805
rect 4683 34756 4684 34796
rect 4724 34756 4725 34796
rect 4683 34747 4725 34756
rect 4587 34376 4629 34385
rect 4587 34336 4588 34376
rect 4628 34336 4629 34376
rect 4587 34327 4629 34336
rect 4491 34208 4533 34217
rect 4491 34168 4492 34208
rect 4532 34168 4533 34208
rect 4491 34159 4533 34168
rect 4395 33368 4437 33377
rect 4395 33328 4396 33368
rect 4436 33328 4437 33368
rect 4395 33319 4437 33328
rect 4588 33200 4628 34327
rect 4684 34133 4724 34747
rect 4683 34124 4725 34133
rect 4683 34084 4684 34124
rect 4724 34084 4725 34124
rect 4683 34075 4725 34084
rect 4780 34049 4820 35344
rect 4876 35216 4916 35225
rect 4876 34805 4916 35176
rect 4971 35216 5013 35225
rect 4971 35176 4972 35216
rect 5012 35176 5013 35216
rect 4971 35167 5013 35176
rect 4875 34796 4917 34805
rect 4875 34756 4876 34796
rect 4916 34756 4917 34796
rect 4875 34747 4917 34756
rect 4972 34217 5012 35167
rect 5355 34712 5397 34721
rect 5355 34672 5356 34712
rect 5396 34672 5397 34712
rect 5355 34663 5397 34672
rect 4971 34208 5013 34217
rect 4971 34168 4972 34208
rect 5012 34168 5013 34208
rect 4971 34159 5013 34168
rect 4779 34040 4821 34049
rect 4779 34000 4780 34040
rect 4820 34000 4821 34040
rect 4779 33991 4821 34000
rect 4928 34040 5296 34049
rect 4968 34000 5010 34040
rect 5050 34000 5092 34040
rect 5132 34000 5174 34040
rect 5214 34000 5256 34040
rect 4928 33991 5296 34000
rect 4683 33956 4725 33965
rect 4683 33916 4684 33956
rect 4724 33916 4725 33956
rect 4683 33907 4725 33916
rect 4396 33160 4628 33200
rect 3819 33076 3820 33116
rect 3860 33076 3861 33116
rect 3819 33067 3861 33076
rect 4012 33076 4244 33116
rect 4299 33116 4341 33125
rect 4299 33076 4300 33116
rect 4340 33076 4341 33116
rect 3820 32982 3860 33067
rect 3628 32864 3668 32873
rect 3628 32705 3668 32824
rect 3820 32864 3860 32873
rect 4012 32864 4052 33076
rect 4299 33067 4341 33076
rect 4107 32948 4149 32957
rect 4107 32908 4108 32948
rect 4148 32908 4149 32948
rect 4107 32899 4149 32908
rect 4299 32948 4341 32957
rect 4299 32908 4300 32948
rect 4340 32908 4341 32948
rect 4299 32899 4341 32908
rect 3860 32824 4012 32864
rect 3820 32815 3860 32824
rect 4012 32815 4052 32824
rect 4108 32864 4148 32899
rect 4108 32813 4148 32824
rect 4204 32864 4244 32873
rect 4204 32705 4244 32824
rect 4300 32864 4340 32899
rect 4300 32813 4340 32824
rect 4396 32705 4436 33160
rect 4492 32864 4532 32875
rect 4492 32789 4532 32824
rect 4587 32864 4629 32873
rect 4587 32824 4588 32864
rect 4628 32824 4629 32864
rect 4587 32815 4629 32824
rect 4491 32780 4533 32789
rect 4491 32740 4492 32780
rect 4532 32740 4533 32780
rect 4491 32731 4533 32740
rect 3627 32696 3669 32705
rect 3627 32656 3628 32696
rect 3668 32656 3669 32696
rect 3627 32647 3669 32656
rect 4203 32696 4245 32705
rect 4203 32656 4204 32696
rect 4244 32656 4245 32696
rect 4203 32647 4245 32656
rect 4395 32696 4437 32705
rect 4395 32656 4396 32696
rect 4436 32656 4437 32696
rect 4395 32647 4437 32656
rect 3723 32360 3765 32369
rect 3723 32320 3724 32360
rect 3764 32320 3765 32360
rect 3723 32311 3765 32320
rect 4011 32360 4053 32369
rect 4011 32320 4012 32360
rect 4052 32320 4053 32360
rect 4011 32311 4053 32320
rect 4396 32360 4436 32369
rect 4436 32320 4532 32360
rect 4396 32311 4436 32320
rect 3436 32236 3572 32276
rect 3052 32192 3092 32201
rect 3052 31865 3092 32152
rect 3051 31856 3093 31865
rect 3051 31816 3052 31856
rect 3092 31816 3093 31856
rect 3051 31807 3093 31816
rect 2955 31772 2997 31781
rect 2955 31732 2956 31772
rect 2996 31732 2997 31772
rect 2955 31723 2997 31732
rect 2859 30764 2901 30773
rect 2859 30724 2860 30764
rect 2900 30724 2901 30764
rect 2859 30715 2901 30724
rect 2860 30680 2900 30715
rect 2860 30629 2900 30640
rect 2668 30304 2804 30344
rect 2668 30185 2708 30304
rect 2859 30260 2901 30269
rect 2859 30220 2860 30260
rect 2900 30220 2901 30260
rect 2859 30211 2901 30220
rect 2667 30176 2709 30185
rect 2667 30136 2668 30176
rect 2708 30136 2709 30176
rect 2667 30127 2709 30136
rect 2763 30092 2805 30101
rect 2763 30052 2764 30092
rect 2804 30052 2805 30092
rect 2763 30043 2805 30052
rect 2860 30092 2900 30211
rect 2860 30043 2900 30052
rect 2668 29672 2708 29681
rect 2668 29009 2708 29632
rect 2667 29000 2709 29009
rect 2667 28960 2668 29000
rect 2708 28960 2709 29000
rect 2667 28951 2709 28960
rect 2572 28363 2612 28372
rect 2476 28328 2516 28337
rect 2476 27833 2516 28288
rect 2764 27917 2804 30043
rect 2956 29924 2996 31723
rect 3147 31268 3189 31277
rect 3147 31228 3148 31268
rect 3188 31228 3189 31268
rect 3147 31219 3189 31228
rect 3051 30848 3093 30857
rect 3051 30808 3052 30848
rect 3092 30808 3093 30848
rect 3051 30799 3093 30808
rect 3052 30680 3092 30799
rect 3052 30631 3092 30640
rect 3052 30428 3092 30439
rect 3052 30353 3092 30388
rect 3051 30344 3093 30353
rect 3051 30304 3052 30344
rect 3092 30304 3093 30344
rect 3051 30295 3093 30304
rect 2860 29884 2996 29924
rect 2860 29261 2900 29884
rect 3052 29840 3092 29849
rect 3148 29840 3188 31219
rect 3339 30764 3381 30773
rect 3339 30724 3340 30764
rect 3380 30724 3381 30764
rect 3339 30715 3381 30724
rect 3340 30680 3380 30715
rect 3340 30629 3380 30640
rect 3339 30512 3381 30521
rect 3339 30472 3340 30512
rect 3380 30472 3381 30512
rect 3339 30463 3381 30472
rect 3092 29800 3188 29840
rect 2955 29420 2997 29429
rect 2955 29380 2956 29420
rect 2996 29380 2997 29420
rect 2955 29371 2997 29380
rect 2859 29252 2901 29261
rect 2859 29212 2860 29252
rect 2900 29212 2901 29252
rect 2859 29203 2901 29212
rect 2763 27908 2805 27917
rect 2763 27868 2764 27908
rect 2804 27868 2805 27908
rect 2763 27859 2805 27868
rect 2860 27833 2900 29203
rect 2475 27824 2517 27833
rect 2475 27784 2476 27824
rect 2516 27784 2517 27824
rect 2475 27775 2517 27784
rect 2859 27824 2901 27833
rect 2859 27784 2860 27824
rect 2900 27784 2901 27824
rect 2859 27775 2901 27784
rect 2571 27740 2613 27749
rect 2571 27700 2572 27740
rect 2612 27700 2613 27740
rect 2571 27691 2613 27700
rect 2476 27656 2516 27665
rect 2476 26816 2516 27616
rect 2476 26153 2516 26776
rect 2572 26657 2612 27691
rect 2763 27656 2805 27665
rect 2763 27616 2764 27656
rect 2804 27616 2805 27656
rect 2763 27607 2805 27616
rect 2667 27488 2709 27497
rect 2667 27448 2668 27488
rect 2708 27448 2709 27488
rect 2667 27439 2709 27448
rect 2668 27354 2708 27439
rect 2764 27413 2804 27607
rect 2865 27413 2905 27494
rect 2763 27404 2805 27413
rect 2763 27364 2764 27404
rect 2804 27364 2805 27404
rect 2763 27355 2805 27364
rect 2860 27404 2906 27413
rect 2905 27364 2906 27404
rect 2860 27355 2906 27364
rect 2668 27068 2708 27077
rect 2764 27068 2804 27355
rect 2859 27236 2901 27245
rect 2859 27196 2860 27236
rect 2900 27196 2901 27236
rect 2859 27187 2901 27196
rect 2708 27028 2804 27068
rect 2668 27019 2708 27028
rect 2571 26648 2613 26657
rect 2571 26608 2572 26648
rect 2612 26608 2613 26648
rect 2571 26599 2613 26608
rect 2764 26153 2804 26238
rect 2475 26144 2517 26153
rect 2475 26104 2476 26144
rect 2516 26104 2517 26144
rect 2475 26095 2517 26104
rect 2763 26144 2805 26153
rect 2763 26104 2764 26144
rect 2804 26104 2805 26144
rect 2763 26095 2805 26104
rect 2860 25976 2900 27187
rect 2956 26312 2996 29371
rect 3052 29009 3092 29800
rect 3243 29756 3285 29765
rect 3243 29716 3244 29756
rect 3284 29716 3285 29756
rect 3243 29707 3285 29716
rect 3147 29504 3189 29513
rect 3147 29464 3148 29504
rect 3188 29464 3189 29504
rect 3147 29455 3189 29464
rect 3051 29000 3093 29009
rect 3051 28960 3052 29000
rect 3092 28960 3093 29000
rect 3051 28951 3093 28960
rect 3148 28421 3188 29455
rect 3244 29345 3284 29707
rect 3243 29336 3285 29345
rect 3243 29296 3244 29336
rect 3284 29296 3285 29336
rect 3243 29287 3285 29296
rect 3244 29168 3284 29287
rect 3147 28412 3189 28421
rect 3147 28372 3148 28412
rect 3188 28372 3189 28412
rect 3147 28363 3189 28372
rect 3052 28328 3092 28337
rect 3052 28169 3092 28288
rect 3051 28160 3093 28169
rect 3051 28120 3052 28160
rect 3092 28120 3093 28160
rect 3051 28111 3093 28120
rect 3244 28001 3284 29128
rect 3243 27992 3285 28001
rect 3243 27952 3244 27992
rect 3284 27952 3285 27992
rect 3243 27943 3285 27952
rect 3243 27824 3285 27833
rect 3243 27784 3244 27824
rect 3284 27784 3285 27824
rect 3243 27775 3285 27784
rect 3147 27740 3189 27749
rect 3147 27700 3148 27740
rect 3188 27700 3189 27740
rect 3147 27691 3189 27700
rect 3148 27606 3188 27691
rect 3244 27656 3284 27775
rect 3147 27488 3189 27497
rect 3147 27448 3148 27488
rect 3188 27448 3189 27488
rect 3147 27439 3189 27448
rect 3051 27404 3093 27413
rect 3051 27364 3052 27404
rect 3092 27364 3093 27404
rect 3051 27355 3093 27364
rect 3052 26480 3092 27355
rect 3148 26816 3188 27439
rect 3244 27245 3284 27616
rect 3243 27236 3285 27245
rect 3243 27196 3244 27236
rect 3284 27196 3285 27236
rect 3243 27187 3285 27196
rect 3243 26984 3285 26993
rect 3243 26944 3244 26984
rect 3284 26944 3285 26984
rect 3243 26935 3285 26944
rect 3148 26767 3188 26776
rect 3244 26480 3284 26935
rect 3340 26816 3380 30463
rect 3436 30092 3476 32236
rect 3724 32226 3764 32311
rect 3915 32192 3957 32201
rect 3532 32178 3572 32187
rect 3915 32152 3916 32192
rect 3956 32152 3957 32192
rect 3915 32143 3957 32152
rect 4012 32192 4052 32311
rect 4204 32192 4244 32201
rect 4012 32143 4052 32152
rect 4108 32152 4204 32192
rect 3532 30269 3572 32138
rect 3916 32058 3956 32143
rect 3688 31772 4056 31781
rect 3728 31732 3770 31772
rect 3810 31732 3852 31772
rect 3892 31732 3934 31772
rect 3974 31732 4016 31772
rect 3688 31723 4056 31732
rect 3627 31520 3669 31529
rect 3627 31480 3628 31520
rect 3668 31480 3669 31520
rect 3627 31471 3669 31480
rect 3628 30680 3668 31471
rect 3820 31352 3860 31363
rect 3820 31277 3860 31312
rect 3819 31268 3861 31277
rect 3819 31228 3820 31268
rect 3860 31228 3861 31268
rect 3819 31219 3861 31228
rect 3628 30521 3668 30640
rect 3723 30680 3765 30689
rect 3723 30640 3724 30680
rect 3764 30640 3765 30680
rect 3723 30631 3765 30640
rect 3724 30546 3764 30631
rect 3820 30521 3860 31219
rect 4011 31184 4053 31193
rect 4011 31144 4012 31184
rect 4052 31144 4053 31184
rect 4011 31135 4053 31144
rect 4012 31050 4052 31135
rect 3627 30512 3669 30521
rect 3627 30472 3628 30512
rect 3668 30472 3669 30512
rect 3627 30463 3669 30472
rect 3819 30512 3861 30521
rect 3819 30472 3820 30512
rect 3860 30472 3861 30512
rect 3819 30463 3861 30472
rect 4012 30437 4052 30522
rect 4011 30428 4053 30437
rect 4011 30388 4012 30428
rect 4052 30388 4053 30428
rect 4011 30379 4053 30388
rect 4108 30344 4148 32152
rect 4204 32143 4244 32152
rect 4300 32192 4340 32201
rect 4401 32192 4441 32201
rect 4204 31352 4244 31363
rect 4204 31277 4244 31312
rect 4203 31268 4245 31277
rect 4203 31228 4204 31268
rect 4244 31228 4245 31268
rect 4203 31219 4245 31228
rect 4203 30932 4245 30941
rect 4203 30892 4204 30932
rect 4244 30892 4245 30932
rect 4203 30883 4245 30892
rect 4204 30680 4244 30883
rect 4300 30857 4340 32152
rect 4396 32152 4401 32192
rect 4396 32143 4441 32152
rect 4299 30848 4341 30857
rect 4299 30808 4300 30848
rect 4340 30808 4341 30848
rect 4299 30799 4341 30808
rect 4204 30631 4244 30640
rect 4396 30437 4436 32143
rect 4395 30428 4437 30437
rect 4395 30388 4396 30428
rect 4436 30388 4437 30428
rect 4395 30379 4437 30388
rect 4203 30344 4245 30353
rect 4108 30304 4204 30344
rect 4244 30304 4245 30344
rect 4203 30295 4245 30304
rect 3531 30260 3573 30269
rect 3531 30220 3532 30260
rect 3572 30220 3573 30260
rect 3531 30211 3573 30220
rect 3688 30260 4056 30269
rect 3728 30220 3770 30260
rect 3810 30220 3852 30260
rect 3892 30220 3934 30260
rect 3974 30220 4016 30260
rect 3688 30211 4056 30220
rect 3436 30052 3668 30092
rect 3628 29336 3668 30052
rect 3628 29287 3668 29296
rect 3820 29168 3860 29177
rect 3820 29009 3860 29128
rect 4107 29084 4149 29093
rect 4107 29044 4108 29084
rect 4148 29044 4149 29084
rect 4107 29035 4149 29044
rect 3819 29000 3861 29009
rect 3819 28960 3820 29000
rect 3860 28960 3861 29000
rect 3819 28951 3861 28960
rect 3436 28916 3476 28925
rect 3476 28876 3572 28916
rect 3436 28867 3476 28876
rect 3435 28748 3477 28757
rect 3435 28708 3436 28748
rect 3476 28708 3477 28748
rect 3435 28699 3477 28708
rect 3436 27077 3476 28699
rect 3532 28342 3572 28876
rect 3688 28748 4056 28757
rect 3728 28708 3770 28748
rect 3810 28708 3852 28748
rect 3892 28708 3934 28748
rect 3974 28708 4016 28748
rect 3688 28699 4056 28708
rect 3915 28580 3957 28589
rect 3915 28540 3916 28580
rect 3956 28540 3957 28580
rect 3915 28531 3957 28540
rect 3532 28293 3572 28302
rect 3916 28328 3956 28531
rect 4108 28496 4148 29035
rect 4204 28589 4244 30295
rect 4492 30185 4532 32320
rect 4491 30176 4533 30185
rect 4491 30136 4492 30176
rect 4532 30136 4533 30176
rect 4491 30127 4533 30136
rect 4299 29924 4341 29933
rect 4299 29884 4300 29924
rect 4340 29884 4341 29924
rect 4299 29875 4341 29884
rect 4300 29840 4340 29875
rect 4300 29789 4340 29800
rect 4588 29756 4628 32815
rect 4684 31529 4724 33907
rect 5356 33788 5396 34663
rect 5548 34628 5588 37780
rect 5643 36896 5685 36905
rect 5643 36856 5644 36896
rect 5684 36856 5685 36896
rect 5643 36847 5685 36856
rect 5644 36762 5684 36847
rect 5740 36560 5780 37939
rect 5836 36980 5876 38704
rect 5932 37745 5972 38872
rect 5931 37736 5973 37745
rect 5931 37696 5932 37736
rect 5972 37696 5973 37736
rect 5931 37687 5973 37696
rect 6028 37661 6068 39376
rect 6027 37652 6069 37661
rect 6027 37612 6028 37652
rect 6068 37612 6069 37652
rect 6027 37603 6069 37612
rect 5932 37400 5972 37411
rect 5932 37325 5972 37360
rect 6028 37400 6068 37409
rect 5931 37316 5973 37325
rect 5931 37276 5932 37316
rect 5972 37276 5973 37316
rect 5931 37267 5973 37276
rect 6028 37157 6068 37360
rect 6027 37148 6069 37157
rect 6027 37108 6028 37148
rect 6068 37108 6069 37148
rect 6027 37099 6069 37108
rect 5836 36940 6068 36980
rect 5836 36737 5876 36822
rect 5931 36812 5973 36821
rect 5931 36772 5932 36812
rect 5972 36772 5973 36812
rect 5931 36763 5973 36772
rect 5835 36728 5877 36737
rect 5835 36688 5836 36728
rect 5876 36688 5877 36728
rect 5835 36679 5877 36688
rect 5932 36678 5972 36763
rect 5740 36520 5876 36560
rect 5836 35902 5876 36520
rect 6028 35888 6068 36940
rect 6124 36896 6164 39460
rect 6220 39257 6260 39628
rect 6219 39248 6261 39257
rect 6219 39208 6220 39248
rect 6260 39208 6261 39248
rect 6219 39199 6261 39208
rect 6316 38240 6356 38249
rect 6316 37997 6356 38200
rect 6315 37988 6357 37997
rect 6315 37948 6316 37988
rect 6356 37948 6357 37988
rect 6315 37939 6357 37948
rect 6508 37988 6548 37997
rect 6508 37820 6548 37948
rect 6316 37780 6548 37820
rect 6604 37820 6644 40804
rect 6700 39752 6740 42475
rect 6796 41693 6836 42928
rect 6795 41684 6837 41693
rect 6795 41644 6796 41684
rect 6836 41644 6837 41684
rect 6795 41635 6837 41644
rect 6988 40517 7028 42928
rect 6987 40508 7029 40517
rect 6987 40468 6988 40508
rect 7028 40468 7029 40508
rect 6987 40459 7029 40468
rect 6987 40340 7029 40349
rect 7180 40340 7220 42928
rect 7275 41516 7317 41525
rect 7275 41476 7276 41516
rect 7316 41476 7317 41516
rect 7275 41467 7317 41476
rect 7276 41273 7316 41467
rect 7275 41264 7317 41273
rect 7275 41224 7276 41264
rect 7316 41224 7317 41264
rect 7275 41215 7317 41224
rect 7276 40424 7316 41215
rect 7372 41021 7412 42928
rect 7371 41012 7413 41021
rect 7371 40972 7372 41012
rect 7412 40972 7413 41012
rect 7371 40963 7413 40972
rect 7564 40685 7604 42928
rect 7756 42029 7796 42928
rect 7755 42020 7797 42029
rect 7755 41980 7756 42020
rect 7796 41980 7797 42020
rect 7755 41971 7797 41980
rect 7659 41432 7701 41441
rect 7659 41392 7660 41432
rect 7700 41392 7701 41432
rect 7659 41383 7701 41392
rect 7563 40676 7605 40685
rect 7563 40636 7564 40676
rect 7604 40636 7605 40676
rect 7563 40627 7605 40636
rect 7660 40676 7700 41383
rect 7851 41264 7893 41273
rect 7851 41224 7852 41264
rect 7892 41224 7893 41264
rect 7851 41215 7893 41224
rect 7852 41130 7892 41215
rect 7660 40627 7700 40636
rect 7755 40508 7797 40517
rect 7755 40468 7756 40508
rect 7796 40468 7797 40508
rect 7755 40459 7797 40468
rect 7852 40508 7892 40517
rect 7276 40349 7316 40384
rect 6987 40300 6988 40340
rect 7028 40300 7029 40340
rect 6987 40291 7029 40300
rect 7084 40300 7220 40340
rect 7275 40340 7317 40349
rect 7275 40300 7276 40340
rect 7316 40300 7317 40340
rect 6988 39761 7028 40291
rect 6700 39703 6740 39712
rect 6987 39752 7029 39761
rect 6987 39712 6988 39752
rect 7028 39712 7029 39752
rect 6987 39703 7029 39712
rect 6795 39164 6837 39173
rect 6795 39124 6796 39164
rect 6836 39124 6837 39164
rect 6795 39115 6837 39124
rect 6604 37780 6740 37820
rect 6219 37736 6261 37745
rect 6219 37696 6220 37736
rect 6260 37696 6261 37736
rect 6219 37687 6261 37696
rect 6124 36847 6164 36856
rect 6220 36821 6260 37687
rect 6219 36812 6261 36821
rect 6219 36772 6220 36812
rect 6260 36772 6261 36812
rect 6316 36812 6356 37780
rect 6411 37400 6453 37409
rect 6411 37360 6412 37400
rect 6452 37360 6453 37400
rect 6411 37351 6453 37360
rect 6508 37400 6548 37409
rect 6548 37360 6644 37400
rect 6508 37351 6548 37360
rect 6412 37266 6452 37351
rect 6507 37064 6549 37073
rect 6507 37024 6508 37064
rect 6548 37024 6549 37064
rect 6507 37015 6549 37024
rect 6316 36772 6452 36812
rect 6219 36763 6261 36772
rect 6315 36644 6357 36653
rect 6315 36604 6316 36644
rect 6356 36604 6357 36644
rect 6315 36595 6357 36604
rect 6316 36510 6356 36595
rect 6412 36392 6452 36772
rect 6508 36728 6548 37015
rect 6508 36679 6548 36688
rect 6507 36560 6549 36569
rect 6507 36520 6508 36560
rect 6548 36520 6549 36560
rect 6507 36511 6549 36520
rect 6316 36352 6452 36392
rect 5836 35853 5876 35862
rect 5932 35848 6068 35888
rect 6220 35888 6260 35897
rect 6316 35888 6356 36352
rect 6260 35848 6356 35888
rect 6412 35888 6452 35897
rect 5932 35384 5972 35848
rect 6028 35720 6068 35729
rect 6028 35468 6068 35680
rect 6220 35645 6260 35848
rect 6412 35729 6452 35848
rect 6508 35888 6548 36511
rect 6508 35839 6548 35848
rect 6316 35720 6356 35729
rect 6219 35636 6261 35645
rect 6219 35596 6220 35636
rect 6260 35596 6261 35636
rect 6219 35587 6261 35596
rect 6028 35428 6260 35468
rect 5740 35344 5972 35384
rect 5644 34628 5684 34637
rect 5548 34588 5644 34628
rect 5644 34579 5684 34588
rect 5452 34376 5492 34385
rect 5452 34049 5492 34336
rect 5451 34040 5493 34049
rect 5451 34000 5452 34040
rect 5492 34000 5493 34040
rect 5451 33991 5493 34000
rect 5740 33872 5780 35344
rect 6027 35300 6069 35309
rect 6027 35260 6028 35300
rect 6068 35260 6069 35300
rect 6027 35251 6069 35260
rect 6028 34292 6068 35251
rect 6123 35216 6165 35225
rect 6123 35176 6124 35216
rect 6164 35176 6165 35216
rect 6123 35167 6165 35176
rect 6124 35082 6164 35167
rect 6220 34964 6260 35428
rect 6316 35393 6356 35680
rect 6411 35720 6453 35729
rect 6411 35680 6412 35720
rect 6452 35680 6453 35720
rect 6411 35671 6453 35680
rect 6411 35552 6453 35561
rect 6411 35512 6412 35552
rect 6452 35512 6453 35552
rect 6411 35503 6453 35512
rect 6315 35384 6357 35393
rect 6315 35344 6316 35384
rect 6356 35344 6357 35384
rect 6315 35335 6357 35344
rect 6028 34243 6068 34252
rect 6124 34924 6260 34964
rect 6316 34964 6356 34973
rect 5548 33832 5780 33872
rect 5356 33748 5492 33788
rect 4780 33704 4820 33713
rect 4780 33377 4820 33664
rect 5259 33704 5301 33713
rect 5259 33664 5260 33704
rect 5300 33664 5301 33704
rect 5259 33655 5301 33664
rect 4875 33620 4917 33629
rect 4875 33580 4876 33620
rect 4916 33580 4917 33620
rect 4875 33571 4917 33580
rect 4779 33368 4821 33377
rect 4779 33328 4780 33368
rect 4820 33328 4821 33368
rect 4779 33319 4821 33328
rect 4779 32780 4821 32789
rect 4779 32740 4780 32780
rect 4820 32740 4821 32780
rect 4779 32731 4821 32740
rect 4780 32369 4820 32731
rect 4876 32705 4916 33571
rect 5260 33570 5300 33655
rect 5355 33620 5397 33629
rect 5355 33580 5356 33620
rect 5396 33580 5397 33620
rect 5355 33571 5397 33580
rect 5356 33486 5396 33571
rect 4875 32696 4917 32705
rect 4875 32656 4876 32696
rect 4916 32656 4917 32696
rect 4875 32647 4917 32656
rect 4928 32528 5296 32537
rect 4968 32488 5010 32528
rect 5050 32488 5092 32528
rect 5132 32488 5174 32528
rect 5214 32488 5256 32528
rect 4928 32479 5296 32488
rect 4779 32360 4821 32369
rect 4779 32320 4780 32360
rect 4820 32320 4821 32360
rect 4779 32311 4821 32320
rect 5355 32276 5397 32285
rect 5355 32236 5356 32276
rect 5396 32236 5397 32276
rect 5355 32227 5397 32236
rect 4780 32192 4820 32201
rect 4780 31949 4820 32152
rect 4779 31940 4821 31949
rect 4779 31900 4780 31940
rect 4820 31900 4821 31940
rect 4779 31891 4821 31900
rect 4683 31520 4725 31529
rect 4683 31480 4684 31520
rect 4724 31480 4725 31520
rect 4683 31471 4725 31480
rect 4928 31016 5296 31025
rect 4968 30976 5010 31016
rect 5050 30976 5092 31016
rect 5132 30976 5174 31016
rect 5214 30976 5256 31016
rect 4928 30967 5296 30976
rect 5067 30848 5109 30857
rect 5067 30808 5068 30848
rect 5108 30808 5109 30848
rect 5067 30799 5109 30808
rect 4779 30260 4821 30269
rect 4779 30220 4780 30260
rect 4820 30220 4821 30260
rect 4779 30211 4821 30220
rect 4780 29854 4820 30211
rect 4780 29805 4820 29814
rect 5068 29765 5108 30799
rect 5356 30269 5396 32227
rect 5452 31529 5492 33748
rect 5451 31520 5493 31529
rect 5451 31480 5452 31520
rect 5492 31480 5493 31520
rect 5451 31471 5493 31480
rect 5452 31352 5492 31361
rect 5452 31025 5492 31312
rect 5451 31016 5493 31025
rect 5451 30976 5452 31016
rect 5492 30976 5493 31016
rect 5451 30967 5493 30976
rect 5452 30857 5492 30967
rect 5451 30848 5493 30857
rect 5451 30808 5452 30848
rect 5492 30808 5493 30848
rect 5451 30799 5493 30808
rect 5452 30680 5492 30689
rect 5452 30521 5492 30640
rect 5451 30512 5493 30521
rect 5451 30472 5452 30512
rect 5492 30472 5493 30512
rect 5451 30463 5493 30472
rect 5355 30260 5397 30269
rect 5355 30220 5356 30260
rect 5396 30220 5397 30260
rect 5355 30211 5397 30220
rect 5260 29840 5300 29849
rect 5300 29800 5396 29840
rect 5260 29791 5300 29800
rect 4588 29707 4628 29716
rect 5067 29756 5109 29765
rect 5067 29716 5068 29756
rect 5108 29716 5109 29756
rect 5067 29707 5109 29716
rect 4928 29504 5296 29513
rect 4968 29464 5010 29504
rect 5050 29464 5092 29504
rect 5132 29464 5174 29504
rect 5214 29464 5256 29504
rect 4928 29455 5296 29464
rect 5356 29429 5396 29800
rect 5451 29756 5493 29765
rect 5451 29716 5452 29756
rect 5492 29716 5493 29756
rect 5451 29707 5493 29716
rect 5355 29420 5397 29429
rect 5355 29380 5356 29420
rect 5396 29380 5397 29420
rect 5355 29371 5397 29380
rect 5067 29336 5109 29345
rect 5067 29296 5068 29336
rect 5108 29296 5109 29336
rect 5067 29287 5109 29296
rect 5068 29168 5108 29287
rect 5068 29119 5108 29128
rect 4683 29000 4725 29009
rect 4683 28960 4684 29000
rect 4724 28960 4725 29000
rect 4683 28951 4725 28960
rect 4491 28832 4533 28841
rect 4491 28792 4492 28832
rect 4532 28792 4533 28832
rect 4491 28783 4533 28792
rect 4203 28580 4245 28589
rect 4203 28540 4204 28580
rect 4244 28540 4245 28580
rect 4203 28531 4245 28540
rect 4108 28447 4148 28456
rect 4011 28412 4053 28421
rect 4011 28372 4012 28412
rect 4052 28372 4053 28412
rect 4011 28363 4053 28372
rect 4203 28412 4245 28421
rect 4203 28372 4204 28412
rect 4244 28372 4245 28412
rect 4203 28363 4245 28372
rect 3916 28279 3956 28288
rect 4012 28278 4052 28363
rect 4204 28278 4244 28363
rect 4300 28337 4340 28422
rect 4299 28328 4341 28337
rect 4299 28288 4300 28328
rect 4340 28288 4341 28328
rect 4299 28279 4341 28288
rect 4492 28328 4532 28783
rect 4492 28279 4532 28288
rect 3723 28244 3765 28253
rect 3723 28204 3724 28244
rect 3764 28204 3765 28244
rect 3723 28195 3765 28204
rect 3724 28110 3764 28195
rect 4491 28160 4533 28169
rect 4491 28120 4492 28160
rect 4532 28120 4533 28160
rect 4491 28111 4533 28120
rect 4299 27824 4341 27833
rect 4299 27784 4300 27824
rect 4340 27784 4341 27824
rect 4299 27775 4341 27784
rect 3532 27656 3572 27667
rect 3532 27581 3572 27616
rect 3820 27656 3860 27665
rect 3531 27572 3573 27581
rect 3531 27532 3532 27572
rect 3572 27532 3573 27572
rect 3531 27523 3573 27532
rect 3820 27497 3860 27616
rect 3915 27656 3957 27665
rect 3915 27616 3916 27656
rect 3956 27616 3957 27656
rect 3915 27607 3957 27616
rect 4107 27656 4149 27665
rect 4107 27616 4108 27656
rect 4148 27616 4149 27656
rect 4107 27607 4149 27616
rect 4300 27656 4340 27775
rect 4300 27607 4340 27616
rect 3916 27522 3956 27607
rect 4108 27522 4148 27607
rect 3819 27488 3861 27497
rect 3819 27448 3820 27488
rect 3860 27448 3861 27488
rect 3819 27439 3861 27448
rect 4108 27404 4148 27413
rect 4148 27364 4340 27404
rect 4108 27355 4148 27364
rect 3688 27236 4056 27245
rect 3728 27196 3770 27236
rect 3810 27196 3852 27236
rect 3892 27196 3934 27236
rect 3974 27196 4016 27236
rect 3688 27187 4056 27196
rect 3435 27068 3477 27077
rect 3435 27028 3436 27068
rect 3476 27028 3477 27068
rect 3435 27019 3477 27028
rect 4204 26993 4244 27078
rect 3820 26984 3860 26993
rect 3436 26816 3476 26825
rect 3340 26776 3436 26816
rect 3436 26489 3476 26776
rect 3531 26732 3573 26741
rect 3531 26692 3532 26732
rect 3572 26692 3573 26732
rect 3531 26683 3573 26692
rect 3532 26598 3572 26683
rect 3435 26480 3477 26489
rect 3820 26480 3860 26944
rect 4203 26984 4245 26993
rect 4203 26944 4204 26984
rect 4244 26944 4245 26984
rect 4203 26935 4245 26944
rect 4012 26816 4052 26827
rect 4012 26741 4052 26776
rect 4204 26816 4244 26825
rect 4011 26732 4053 26741
rect 4011 26692 4012 26732
rect 4052 26692 4053 26732
rect 4011 26683 4053 26692
rect 4204 26573 4244 26776
rect 4300 26648 4340 27364
rect 4395 26900 4437 26909
rect 4395 26860 4396 26900
rect 4436 26860 4437 26900
rect 4395 26851 4437 26860
rect 4396 26816 4436 26851
rect 4396 26765 4436 26776
rect 4300 26608 4436 26648
rect 4203 26564 4245 26573
rect 4203 26524 4204 26564
rect 4244 26524 4245 26564
rect 4203 26515 4245 26524
rect 3052 26440 3188 26480
rect 3244 26440 3362 26480
rect 2956 26272 3092 26312
rect 3052 26228 3092 26272
rect 3047 26188 3092 26228
rect 3148 26228 3188 26440
rect 3322 26396 3362 26440
rect 3435 26440 3436 26480
rect 3476 26440 3477 26480
rect 3435 26431 3477 26440
rect 3780 26440 3860 26480
rect 3322 26356 3388 26396
rect 3348 26312 3388 26356
rect 3628 26321 3668 26406
rect 3340 26272 3388 26312
rect 3627 26312 3669 26321
rect 3627 26272 3628 26312
rect 3668 26272 3669 26312
rect 3241 26237 3281 26243
rect 3240 26228 3282 26237
rect 3148 26188 3198 26228
rect 2955 26144 2997 26153
rect 2955 26104 2956 26144
rect 2996 26104 2997 26144
rect 2955 26095 2997 26104
rect 2764 25936 2900 25976
rect 2956 25976 2996 26095
rect 3047 25976 3087 26188
rect 3047 25936 3092 25976
rect 2476 25304 2516 25313
rect 2476 25220 2516 25264
rect 2476 25180 2612 25220
rect 2475 25052 2517 25061
rect 2475 25012 2476 25052
rect 2516 25012 2517 25052
rect 2475 25003 2517 25012
rect 2476 24641 2516 25003
rect 2572 24800 2612 25180
rect 2667 25136 2709 25145
rect 2667 25096 2668 25136
rect 2708 25096 2709 25136
rect 2667 25087 2709 25096
rect 2668 25002 2708 25087
rect 2667 24800 2709 24809
rect 2572 24760 2668 24800
rect 2708 24760 2709 24800
rect 2667 24751 2709 24760
rect 2475 24632 2517 24641
rect 2475 24592 2476 24632
rect 2516 24592 2517 24632
rect 2475 24583 2517 24592
rect 2668 24632 2708 24751
rect 2668 24583 2708 24592
rect 2283 24212 2325 24221
rect 2283 24172 2284 24212
rect 2324 24172 2325 24212
rect 2283 24163 2325 24172
rect 2476 23792 2516 24583
rect 2667 24464 2709 24473
rect 2667 24424 2668 24464
rect 2708 24424 2709 24464
rect 2667 24415 2709 24424
rect 2476 23743 2516 23752
rect 2571 23792 2613 23801
rect 2571 23752 2572 23792
rect 2612 23752 2613 23792
rect 2571 23743 2613 23752
rect 2572 23658 2612 23743
rect 2187 23624 2229 23633
rect 2187 23584 2188 23624
rect 2228 23584 2229 23624
rect 2187 23575 2229 23584
rect 2188 23490 2228 23575
rect 2187 23372 2229 23381
rect 2187 23332 2188 23372
rect 2228 23332 2229 23372
rect 2187 23323 2229 23332
rect 2188 22289 2228 23323
rect 2475 22616 2517 22625
rect 2475 22576 2476 22616
rect 2516 22576 2517 22616
rect 2475 22567 2517 22576
rect 2379 22364 2421 22373
rect 2379 22324 2380 22364
rect 2420 22324 2421 22364
rect 2379 22315 2421 22324
rect 2187 22280 2229 22289
rect 2187 22240 2188 22280
rect 2228 22240 2229 22280
rect 2187 22231 2229 22240
rect 2091 22028 2133 22037
rect 2091 21988 2092 22028
rect 2132 21988 2133 22028
rect 2091 21979 2133 21988
rect 2092 18929 2132 21979
rect 2283 21524 2325 21533
rect 2283 21484 2284 21524
rect 2324 21484 2325 21524
rect 2283 21475 2325 21484
rect 2284 19853 2324 21475
rect 2283 19844 2325 19853
rect 2283 19804 2284 19844
rect 2324 19804 2325 19844
rect 2283 19795 2325 19804
rect 2283 19676 2325 19685
rect 2283 19636 2284 19676
rect 2324 19636 2325 19676
rect 2283 19627 2325 19636
rect 2091 18920 2133 18929
rect 2091 18880 2092 18920
rect 2132 18880 2133 18920
rect 2091 18871 2133 18880
rect 2091 18668 2133 18677
rect 2091 18628 2092 18668
rect 2132 18628 2133 18668
rect 2091 18619 2133 18628
rect 1804 17872 2036 17912
rect 1323 17156 1365 17165
rect 1323 17116 1324 17156
rect 1364 17116 1365 17156
rect 1323 17107 1365 17116
rect 1611 17156 1653 17165
rect 1611 17116 1612 17156
rect 1652 17116 1653 17156
rect 1611 17107 1653 17116
rect 1228 16064 1268 16073
rect 1228 14981 1268 16024
rect 1324 15392 1364 17107
rect 1804 17081 1844 17872
rect 1899 17744 1941 17753
rect 1899 17704 1900 17744
rect 1940 17704 1941 17744
rect 1899 17695 1941 17704
rect 1803 17072 1845 17081
rect 1803 17032 1804 17072
rect 1844 17032 1845 17072
rect 1803 17023 1845 17032
rect 1612 16988 1652 16997
rect 1652 16948 1748 16988
rect 1612 16939 1652 16948
rect 1420 16820 1460 16829
rect 1460 16780 1556 16820
rect 1420 16771 1460 16780
rect 1419 16484 1461 16493
rect 1419 16444 1420 16484
rect 1460 16444 1461 16484
rect 1419 16435 1461 16444
rect 1420 16316 1460 16435
rect 1420 16267 1460 16276
rect 1516 15905 1556 16780
rect 1708 16400 1748 16948
rect 1804 16938 1844 17023
rect 1708 16360 1844 16400
rect 1708 16232 1748 16241
rect 1708 15980 1748 16192
rect 1804 16157 1844 16360
rect 1803 16148 1845 16157
rect 1803 16108 1804 16148
rect 1844 16108 1845 16148
rect 1803 16099 1845 16108
rect 1900 15980 1940 17695
rect 1996 16232 2036 16241
rect 1996 15989 2036 16192
rect 2092 16232 2132 18619
rect 2284 17837 2324 19627
rect 2283 17828 2325 17837
rect 2283 17788 2284 17828
rect 2324 17788 2325 17828
rect 2283 17779 2325 17788
rect 2284 17333 2324 17779
rect 2283 17324 2325 17333
rect 2283 17284 2284 17324
rect 2324 17284 2325 17324
rect 2283 17275 2325 17284
rect 2187 16484 2229 16493
rect 2187 16444 2188 16484
rect 2228 16444 2229 16484
rect 2187 16435 2229 16444
rect 2380 16484 2420 22315
rect 2476 22280 2516 22567
rect 2668 22280 2708 24415
rect 2764 24212 2804 25936
rect 2956 25927 2996 25936
rect 3052 25304 3092 25936
rect 3158 25892 3198 26188
rect 3240 26188 3241 26228
rect 3281 26188 3282 26228
rect 3240 26179 3282 26188
rect 3241 26148 3281 26179
rect 3241 26099 3281 26108
rect 3340 26144 3380 26272
rect 3627 26263 3669 26272
rect 3780 26153 3820 26440
rect 4011 26312 4053 26321
rect 4011 26272 4012 26312
rect 4052 26272 4053 26312
rect 4011 26263 4053 26272
rect 3506 26144 3546 26153
rect 3772 26144 3820 26153
rect 3380 26129 3388 26144
rect 3380 26104 3428 26129
rect 3340 26095 3428 26104
rect 3546 26129 3547 26144
rect 3546 26104 3569 26129
rect 3506 26095 3569 26104
rect 3348 26089 3428 26095
rect 3507 26089 3569 26095
rect 3388 26060 3428 26089
rect 3388 26020 3476 26060
rect 3148 25852 3198 25892
rect 3339 25892 3381 25901
rect 3339 25852 3340 25892
rect 3380 25852 3381 25892
rect 3148 25388 3188 25852
rect 3339 25843 3381 25852
rect 3243 25472 3285 25481
rect 3243 25432 3244 25472
rect 3284 25432 3285 25472
rect 3243 25423 3285 25432
rect 3148 25339 3188 25348
rect 3244 25338 3284 25423
rect 3340 25388 3380 25843
rect 3436 25817 3476 26020
rect 3529 25976 3569 26089
rect 3628 26115 3668 26124
rect 3812 26104 3820 26144
rect 4012 26144 4052 26263
rect 3772 26095 3812 26104
rect 4012 26095 4052 26104
rect 4107 26144 4149 26153
rect 4107 26104 4108 26144
rect 4148 26104 4149 26144
rect 4107 26095 4149 26104
rect 4396 26144 4436 26608
rect 4396 26095 4436 26104
rect 3628 26069 3668 26075
rect 3627 26060 3669 26069
rect 3627 26020 3628 26060
rect 3668 26020 3669 26060
rect 3627 26011 3669 26020
rect 4108 26060 4148 26095
rect 3628 25980 3668 26011
rect 4108 26009 4148 26020
rect 4300 26060 4340 26069
rect 4203 25976 4245 25985
rect 3529 25936 3575 25976
rect 3535 25892 3575 25936
rect 4203 25936 4204 25976
rect 4244 25936 4245 25976
rect 4203 25927 4245 25936
rect 3627 25892 3669 25901
rect 3535 25852 3628 25892
rect 3668 25852 3669 25892
rect 3435 25808 3477 25817
rect 3535 25808 3575 25852
rect 3627 25843 3669 25852
rect 4204 25842 4244 25927
rect 3435 25768 3436 25808
rect 3476 25768 3477 25808
rect 3435 25759 3477 25768
rect 3532 25768 3575 25808
rect 3340 25339 3380 25348
rect 3052 25255 3092 25264
rect 3436 25304 3476 25313
rect 3532 25304 3572 25768
rect 3688 25724 4056 25733
rect 3728 25684 3770 25724
rect 3810 25684 3852 25724
rect 3892 25684 3934 25724
rect 3974 25684 4016 25724
rect 3688 25675 4056 25684
rect 3627 25556 3669 25565
rect 3627 25516 3628 25556
rect 3668 25516 3669 25556
rect 3627 25507 3669 25516
rect 3476 25264 3572 25304
rect 3628 25304 3668 25507
rect 4300 25481 4340 26020
rect 4492 25640 4532 28111
rect 4684 26237 4724 28951
rect 5260 28916 5300 28925
rect 5260 28421 5300 28876
rect 5259 28412 5301 28421
rect 5259 28372 5260 28412
rect 5300 28372 5301 28412
rect 5259 28363 5301 28372
rect 5452 28337 5492 29707
rect 5548 29672 5588 33832
rect 5643 33704 5685 33713
rect 5643 33664 5644 33704
rect 5684 33664 5685 33704
rect 5643 33655 5685 33664
rect 5740 33704 5780 33713
rect 5644 31445 5684 33655
rect 5740 33545 5780 33664
rect 5836 33704 5876 33713
rect 5739 33536 5781 33545
rect 5739 33496 5740 33536
rect 5780 33496 5781 33536
rect 5739 33487 5781 33496
rect 5836 33284 5876 33664
rect 6124 33368 6164 34924
rect 6220 34390 6260 34471
rect 6316 34390 6356 34924
rect 6220 34385 6356 34390
rect 6219 34381 6356 34385
rect 6219 34336 6220 34381
rect 6260 34350 6356 34381
rect 6260 34336 6261 34350
rect 6219 34327 6261 34336
rect 6412 34133 6452 35503
rect 6507 35216 6549 35225
rect 6507 35176 6508 35216
rect 6548 35176 6549 35216
rect 6507 35167 6549 35176
rect 6508 35082 6548 35167
rect 6507 34376 6549 34385
rect 6507 34336 6508 34376
rect 6548 34336 6549 34376
rect 6507 34327 6549 34336
rect 6219 34124 6261 34133
rect 6219 34084 6220 34124
rect 6260 34084 6261 34124
rect 6219 34075 6261 34084
rect 6411 34124 6453 34133
rect 6411 34084 6412 34124
rect 6452 34084 6453 34124
rect 6411 34075 6453 34084
rect 6220 33704 6260 34075
rect 6315 33956 6357 33965
rect 6315 33916 6316 33956
rect 6356 33916 6357 33956
rect 6315 33907 6357 33916
rect 6220 33655 6260 33664
rect 6316 33704 6356 33907
rect 6508 33881 6548 34327
rect 6507 33872 6549 33881
rect 6507 33832 6508 33872
rect 6548 33832 6549 33872
rect 6507 33823 6549 33832
rect 6316 33655 6356 33664
rect 6411 33620 6453 33629
rect 6411 33580 6412 33620
rect 6452 33580 6453 33620
rect 6411 33571 6453 33580
rect 6219 33368 6261 33377
rect 6124 33328 6220 33368
rect 6260 33328 6261 33368
rect 6219 33319 6261 33328
rect 5836 33244 6164 33284
rect 5932 33041 5972 33126
rect 6124 33116 6164 33244
rect 6315 33200 6357 33209
rect 6315 33160 6316 33200
rect 6356 33160 6357 33200
rect 6315 33151 6357 33160
rect 6124 33067 6164 33076
rect 5931 33032 5973 33041
rect 5931 32992 5932 33032
rect 5972 32992 5973 33032
rect 5931 32983 5973 32992
rect 6316 32873 6356 33151
rect 5739 32864 5781 32873
rect 5739 32824 5740 32864
rect 5780 32824 5781 32864
rect 5739 32815 5781 32824
rect 6315 32864 6357 32873
rect 6315 32824 6316 32864
rect 6356 32824 6357 32864
rect 6315 32815 6357 32824
rect 5740 32192 5780 32815
rect 6316 32730 6356 32815
rect 6219 32444 6261 32453
rect 6219 32404 6220 32444
rect 6260 32404 6261 32444
rect 6219 32395 6261 32404
rect 6220 32360 6260 32395
rect 6220 32309 6260 32320
rect 6412 32285 6452 33571
rect 6604 33125 6644 37360
rect 6700 36905 6740 37780
rect 6796 37073 6836 39115
rect 7084 38408 7124 40300
rect 7275 40291 7317 40300
rect 7371 40256 7413 40265
rect 7371 40216 7372 40256
rect 7412 40216 7413 40256
rect 7371 40207 7413 40216
rect 7468 40256 7508 40265
rect 7275 40088 7317 40097
rect 7372 40088 7412 40207
rect 7275 40048 7276 40088
rect 7316 40048 7412 40088
rect 7275 40039 7317 40048
rect 7372 39836 7412 39845
rect 7276 39796 7372 39836
rect 7179 39752 7221 39761
rect 7179 39707 7180 39752
rect 7220 39707 7221 39752
rect 7179 39703 7221 39707
rect 7180 39617 7220 39703
rect 7179 39080 7221 39089
rect 7179 39040 7180 39080
rect 7220 39040 7221 39080
rect 7179 39031 7221 39040
rect 7180 38912 7220 39031
rect 7180 38585 7220 38872
rect 7179 38576 7221 38585
rect 7179 38536 7180 38576
rect 7220 38536 7221 38576
rect 7179 38527 7221 38536
rect 7084 38359 7124 38368
rect 7276 38240 7316 39796
rect 7372 39787 7412 39796
rect 7468 38921 7508 40216
rect 7659 39836 7701 39845
rect 7659 39796 7660 39836
rect 7700 39796 7701 39836
rect 7659 39787 7701 39796
rect 7564 39752 7604 39761
rect 7467 38912 7509 38921
rect 7467 38872 7468 38912
rect 7508 38872 7509 38912
rect 7564 38912 7604 39712
rect 7660 39752 7700 39787
rect 7660 39701 7700 39712
rect 7756 39164 7796 40459
rect 7852 40097 7892 40468
rect 7851 40088 7893 40097
rect 7851 40048 7852 40088
rect 7892 40048 7893 40088
rect 7851 40039 7893 40048
rect 7851 39920 7893 39929
rect 7851 39880 7852 39920
rect 7892 39880 7893 39920
rect 7851 39871 7893 39880
rect 7852 39786 7892 39871
rect 7756 39124 7892 39164
rect 7756 38996 7796 39005
rect 7564 38872 7700 38912
rect 7467 38863 7509 38872
rect 7084 38200 7316 38240
rect 7372 38744 7412 38753
rect 6892 38156 6932 38165
rect 6892 37568 6932 38116
rect 6892 37519 6932 37528
rect 7084 37493 7124 38200
rect 7372 37820 7412 38704
rect 7563 38744 7605 38753
rect 7563 38704 7564 38744
rect 7604 38704 7605 38744
rect 7563 38695 7605 38704
rect 7564 38610 7604 38695
rect 7563 38072 7605 38081
rect 7563 38032 7564 38072
rect 7604 38032 7605 38072
rect 7563 38023 7605 38032
rect 7564 37938 7604 38023
rect 7276 37780 7412 37820
rect 7563 37820 7605 37829
rect 7563 37780 7564 37820
rect 7604 37780 7605 37820
rect 7083 37484 7125 37493
rect 7083 37444 7084 37484
rect 7124 37444 7125 37484
rect 7083 37435 7125 37444
rect 7180 37400 7220 37409
rect 6891 37232 6933 37241
rect 6891 37192 6892 37232
rect 6932 37192 6933 37232
rect 6891 37183 6933 37192
rect 6988 37232 7028 37241
rect 7028 37192 7124 37232
rect 6988 37183 7028 37192
rect 6795 37064 6837 37073
rect 6795 37024 6796 37064
rect 6836 37024 6837 37064
rect 6795 37015 6837 37024
rect 6699 36896 6741 36905
rect 6699 36856 6700 36896
rect 6740 36856 6741 36896
rect 6699 36847 6741 36856
rect 6892 36569 6932 37183
rect 6891 36560 6933 36569
rect 6891 36520 6892 36560
rect 6932 36520 6933 36560
rect 6891 36511 6933 36520
rect 6700 35888 6740 35897
rect 6700 35141 6740 35848
rect 6796 35888 6836 35897
rect 6796 35309 6836 35848
rect 6891 35888 6933 35897
rect 6891 35848 6892 35888
rect 6932 35848 6933 35888
rect 6891 35839 6933 35848
rect 6892 35754 6932 35839
rect 6988 35720 7028 35729
rect 6891 35636 6933 35645
rect 6891 35596 6892 35636
rect 6932 35596 6933 35636
rect 6891 35587 6933 35596
rect 6795 35300 6837 35309
rect 6795 35260 6796 35300
rect 6836 35260 6837 35300
rect 6795 35251 6837 35260
rect 6699 35132 6741 35141
rect 6699 35092 6700 35132
rect 6740 35092 6741 35132
rect 6699 35083 6741 35092
rect 6892 34721 6932 35587
rect 6988 35309 7028 35680
rect 6987 35300 7029 35309
rect 6987 35260 6988 35300
rect 7028 35260 7029 35300
rect 6987 35251 7029 35260
rect 6891 34712 6933 34721
rect 6891 34672 6892 34712
rect 6932 34672 6933 34712
rect 6891 34663 6933 34672
rect 6987 34544 7029 34553
rect 6987 34504 6988 34544
rect 7028 34504 7029 34544
rect 6987 34495 7029 34504
rect 6699 34460 6741 34469
rect 6699 34420 6700 34460
rect 6740 34420 6741 34460
rect 6699 34411 6741 34420
rect 6700 34376 6740 34411
rect 6700 34325 6740 34336
rect 6891 34292 6933 34301
rect 6891 34252 6892 34292
rect 6932 34252 6933 34292
rect 6891 34243 6933 34252
rect 6700 33620 6740 33629
rect 6700 33545 6740 33580
rect 6795 33620 6837 33629
rect 6795 33580 6796 33620
rect 6836 33580 6837 33620
rect 6795 33571 6837 33580
rect 6699 33536 6741 33545
rect 6699 33496 6700 33536
rect 6740 33496 6741 33536
rect 6699 33487 6741 33496
rect 6603 33116 6645 33125
rect 6603 33076 6604 33116
rect 6644 33076 6645 33116
rect 6603 33067 6645 33076
rect 6700 32369 6740 33487
rect 6796 33486 6836 33571
rect 6699 32360 6741 32369
rect 6699 32320 6700 32360
rect 6740 32320 6741 32360
rect 6699 32311 6741 32320
rect 6411 32276 6453 32285
rect 6411 32236 6412 32276
rect 6452 32236 6453 32276
rect 6411 32227 6453 32236
rect 6028 32192 6068 32201
rect 5740 32152 6028 32192
rect 5739 31688 5781 31697
rect 5739 31648 5740 31688
rect 5780 31648 5781 31688
rect 5739 31639 5781 31648
rect 5643 31436 5685 31445
rect 5643 31396 5644 31436
rect 5684 31396 5685 31436
rect 5643 31387 5685 31396
rect 5644 31268 5684 31277
rect 5740 31268 5780 31639
rect 5835 31520 5877 31529
rect 5835 31480 5836 31520
rect 5876 31480 5877 31520
rect 5835 31471 5877 31480
rect 5684 31228 5780 31268
rect 5644 31219 5684 31228
rect 5836 30848 5876 31471
rect 5932 31100 5972 32152
rect 6028 32143 6068 32152
rect 6412 32192 6452 32227
rect 6123 31688 6165 31697
rect 6123 31648 6124 31688
rect 6164 31648 6165 31688
rect 6123 31639 6165 31648
rect 6124 31352 6164 31639
rect 6412 31529 6452 32152
rect 6892 31604 6932 34243
rect 6988 33461 7028 34495
rect 6987 33452 7029 33461
rect 6987 33412 6988 33452
rect 7028 33412 7029 33452
rect 6987 33403 7029 33412
rect 6700 31564 6932 31604
rect 6411 31520 6453 31529
rect 6411 31480 6412 31520
rect 6452 31480 6453 31520
rect 6411 31471 6453 31480
rect 6700 31436 6740 31564
rect 6700 31387 6740 31396
rect 6795 31436 6837 31445
rect 6795 31396 6796 31436
rect 6836 31396 6837 31436
rect 6795 31387 6837 31396
rect 6124 31303 6164 31312
rect 6220 31352 6260 31361
rect 5932 31060 6068 31100
rect 5836 30799 5876 30808
rect 5931 30764 5973 30773
rect 5931 30724 5932 30764
rect 5972 30724 5973 30764
rect 5931 30715 5973 30724
rect 5644 30428 5684 30437
rect 5644 30269 5684 30388
rect 5643 30260 5685 30269
rect 5643 30220 5644 30260
rect 5684 30220 5685 30260
rect 5643 30211 5685 30220
rect 5739 29924 5781 29933
rect 5739 29884 5740 29924
rect 5780 29884 5781 29924
rect 5739 29875 5781 29884
rect 5740 29790 5780 29875
rect 5835 29840 5877 29849
rect 5835 29800 5836 29840
rect 5876 29800 5877 29840
rect 5835 29791 5877 29800
rect 5836 29706 5876 29791
rect 5548 29632 5780 29672
rect 5548 29168 5588 29177
rect 5451 28328 5493 28337
rect 5451 28288 5452 28328
rect 5492 28288 5493 28328
rect 5451 28279 5493 28288
rect 4928 27992 5296 28001
rect 4968 27952 5010 27992
rect 5050 27952 5092 27992
rect 5132 27952 5174 27992
rect 5214 27952 5256 27992
rect 4928 27943 5296 27952
rect 5355 27992 5397 28001
rect 5355 27952 5356 27992
rect 5396 27952 5397 27992
rect 5355 27943 5397 27952
rect 4779 27656 4821 27665
rect 4779 27616 4780 27656
rect 4820 27616 4821 27656
rect 4779 27607 4821 27616
rect 4683 26228 4725 26237
rect 4683 26188 4684 26228
rect 4724 26188 4725 26228
rect 4683 26179 4725 26188
rect 4588 26144 4628 26155
rect 4588 26069 4628 26104
rect 4780 26144 4820 27607
rect 5356 26732 5396 27943
rect 5452 27833 5492 28279
rect 5548 27917 5588 29128
rect 5643 29168 5685 29177
rect 5643 29128 5644 29168
rect 5684 29128 5685 29168
rect 5643 29119 5685 29128
rect 5644 29034 5684 29119
rect 5740 28496 5780 29632
rect 5835 29420 5877 29429
rect 5835 29380 5836 29420
rect 5876 29380 5877 29420
rect 5835 29371 5877 29380
rect 5644 28456 5780 28496
rect 5644 28169 5684 28456
rect 5740 28328 5780 28337
rect 5643 28160 5685 28169
rect 5643 28120 5644 28160
rect 5684 28120 5685 28160
rect 5643 28111 5685 28120
rect 5547 27908 5589 27917
rect 5547 27868 5548 27908
rect 5588 27868 5589 27908
rect 5547 27859 5589 27868
rect 5451 27824 5493 27833
rect 5451 27784 5452 27824
rect 5492 27784 5493 27824
rect 5451 27775 5493 27784
rect 5740 27749 5780 28288
rect 5836 27917 5876 29371
rect 5932 29168 5972 30715
rect 6028 30680 6068 31060
rect 6028 30521 6068 30640
rect 6027 30512 6069 30521
rect 6027 30472 6028 30512
rect 6068 30472 6069 30512
rect 6027 30463 6069 30472
rect 5932 29119 5972 29128
rect 6220 29840 6260 31312
rect 6604 31352 6644 31361
rect 6315 31184 6357 31193
rect 6315 31144 6316 31184
rect 6356 31144 6357 31184
rect 6315 31135 6357 31144
rect 6316 30689 6356 31135
rect 6604 31109 6644 31312
rect 6603 31100 6645 31109
rect 6603 31060 6604 31100
rect 6644 31060 6645 31100
rect 6603 31051 6645 31060
rect 6315 30680 6357 30689
rect 6315 30640 6316 30680
rect 6356 30640 6357 30680
rect 6315 30631 6357 30640
rect 6220 29168 6260 29800
rect 6316 29840 6356 30631
rect 6316 29791 6356 29800
rect 6604 29168 6644 31051
rect 6699 30092 6741 30101
rect 6699 30052 6700 30092
rect 6740 30052 6741 30092
rect 6699 30043 6741 30052
rect 6700 29840 6740 30043
rect 6700 29791 6740 29800
rect 6699 29336 6741 29345
rect 6699 29296 6700 29336
rect 6740 29296 6741 29336
rect 6699 29287 6741 29296
rect 5932 28496 5972 28507
rect 6220 28496 6260 29128
rect 6508 29128 6604 29168
rect 6316 28916 6356 28925
rect 6316 28589 6356 28876
rect 6508 28664 6548 29128
rect 6604 29119 6644 29128
rect 6604 29000 6644 29009
rect 6700 29000 6740 29287
rect 6796 29168 6836 31387
rect 6892 29513 6932 31564
rect 6988 30101 7028 33403
rect 7084 31184 7124 37192
rect 7180 36989 7220 37360
rect 7179 36980 7221 36989
rect 7179 36940 7180 36980
rect 7220 36940 7221 36980
rect 7179 36931 7221 36940
rect 7179 36560 7221 36569
rect 7179 36520 7180 36560
rect 7220 36520 7221 36560
rect 7179 36511 7221 36520
rect 7180 34637 7220 36511
rect 7276 35888 7316 37780
rect 7563 37771 7605 37780
rect 7371 37652 7413 37661
rect 7371 37612 7372 37652
rect 7412 37612 7413 37652
rect 7371 37603 7413 37612
rect 7372 37325 7412 37603
rect 7564 37484 7604 37771
rect 7660 37661 7700 38872
rect 7756 38081 7796 38956
rect 7852 38753 7892 39124
rect 7851 38744 7893 38753
rect 7851 38704 7852 38744
rect 7892 38704 7893 38744
rect 7851 38695 7893 38704
rect 7851 38492 7893 38501
rect 7851 38452 7852 38492
rect 7892 38452 7893 38492
rect 7851 38443 7893 38452
rect 7852 38408 7892 38443
rect 7852 38357 7892 38368
rect 7755 38072 7797 38081
rect 7755 38032 7756 38072
rect 7796 38032 7797 38072
rect 7755 38023 7797 38032
rect 7851 37904 7893 37913
rect 7851 37864 7852 37904
rect 7892 37864 7893 37904
rect 7851 37855 7893 37864
rect 7852 37736 7892 37855
rect 7756 37696 7892 37736
rect 7659 37652 7701 37661
rect 7659 37612 7660 37652
rect 7700 37612 7701 37652
rect 7659 37603 7701 37612
rect 7564 37444 7700 37484
rect 7371 37316 7413 37325
rect 7371 37276 7372 37316
rect 7412 37276 7413 37316
rect 7371 37267 7413 37276
rect 7563 37064 7605 37073
rect 7563 37024 7564 37064
rect 7604 37024 7605 37064
rect 7563 37015 7605 37024
rect 7371 36056 7413 36065
rect 7371 36016 7372 36056
rect 7412 36016 7413 36056
rect 7371 36007 7413 36016
rect 7276 35839 7316 35848
rect 7372 35888 7412 36007
rect 7372 35839 7412 35848
rect 7371 34796 7413 34805
rect 7371 34756 7372 34796
rect 7412 34756 7413 34796
rect 7371 34747 7413 34756
rect 7179 34628 7221 34637
rect 7179 34588 7180 34628
rect 7220 34588 7221 34628
rect 7179 34579 7221 34588
rect 7179 34376 7221 34385
rect 7179 34336 7180 34376
rect 7220 34336 7221 34376
rect 7179 34327 7221 34336
rect 7276 34376 7316 34385
rect 7180 34242 7220 34327
rect 7276 34049 7316 34336
rect 7275 34040 7317 34049
rect 7275 34000 7276 34040
rect 7316 34000 7317 34040
rect 7275 33991 7317 34000
rect 7276 33704 7316 33713
rect 7276 33545 7316 33664
rect 7275 33536 7317 33545
rect 7275 33496 7276 33536
rect 7316 33496 7317 33536
rect 7275 33487 7317 33496
rect 7372 32957 7412 34747
rect 7564 33881 7604 37015
rect 7660 35216 7700 37444
rect 7756 36728 7796 37696
rect 7948 36728 7988 42928
rect 8140 41609 8180 42928
rect 8332 42785 8372 42928
rect 8331 42776 8373 42785
rect 8331 42736 8332 42776
rect 8372 42736 8373 42776
rect 8331 42727 8373 42736
rect 8524 41945 8564 42928
rect 8523 41936 8565 41945
rect 8523 41896 8524 41936
rect 8564 41896 8565 41936
rect 8523 41887 8565 41896
rect 8716 41861 8756 42928
rect 8715 41852 8757 41861
rect 8715 41812 8716 41852
rect 8756 41812 8757 41852
rect 8715 41803 8757 41812
rect 8139 41600 8181 41609
rect 8139 41560 8140 41600
rect 8180 41560 8181 41600
rect 8139 41551 8181 41560
rect 8235 41264 8277 41273
rect 8235 41224 8236 41264
rect 8276 41224 8277 41264
rect 8235 41215 8277 41224
rect 8044 41012 8084 41021
rect 8044 40601 8084 40972
rect 8139 40676 8181 40685
rect 8139 40636 8140 40676
rect 8180 40636 8181 40676
rect 8139 40627 8181 40636
rect 8043 40592 8085 40601
rect 8043 40552 8044 40592
rect 8084 40552 8085 40592
rect 8043 40543 8085 40552
rect 8044 40424 8084 40433
rect 8140 40424 8180 40627
rect 8084 40384 8180 40424
rect 8044 40375 8084 40384
rect 8236 40340 8276 41215
rect 8331 40508 8373 40517
rect 8331 40468 8332 40508
rect 8372 40468 8373 40508
rect 8331 40459 8373 40468
rect 8140 40300 8276 40340
rect 8140 39341 8180 40300
rect 8236 39752 8276 39761
rect 8236 39593 8276 39712
rect 8235 39584 8277 39593
rect 8235 39544 8236 39584
rect 8276 39544 8277 39584
rect 8235 39535 8277 39544
rect 8139 39332 8181 39341
rect 8139 39292 8140 39332
rect 8180 39292 8181 39332
rect 8139 39283 8181 39292
rect 8043 39080 8085 39089
rect 8043 39040 8044 39080
rect 8084 39040 8085 39080
rect 8043 39031 8085 39040
rect 8044 38501 8084 39031
rect 8235 38996 8277 39005
rect 8235 38956 8236 38996
rect 8276 38956 8277 38996
rect 8235 38947 8277 38956
rect 8139 38912 8181 38921
rect 8139 38872 8140 38912
rect 8180 38872 8181 38912
rect 8139 38863 8181 38872
rect 8236 38912 8276 38947
rect 8140 38778 8180 38863
rect 8236 38861 8276 38872
rect 8332 38744 8372 40459
rect 8523 39920 8565 39929
rect 8523 39880 8524 39920
rect 8564 39880 8565 39920
rect 8523 39871 8565 39880
rect 8427 39416 8469 39425
rect 8427 39376 8428 39416
rect 8468 39376 8469 39416
rect 8427 39367 8469 39376
rect 8236 38704 8372 38744
rect 8043 38492 8085 38501
rect 8043 38452 8044 38492
rect 8084 38452 8085 38492
rect 8043 38443 8085 38452
rect 8139 38408 8181 38417
rect 8139 38368 8140 38408
rect 8180 38368 8181 38408
rect 8139 38359 8181 38368
rect 8043 38324 8085 38333
rect 8043 38284 8044 38324
rect 8084 38284 8085 38324
rect 8043 38275 8085 38284
rect 8044 38190 8084 38275
rect 8140 37820 8180 38359
rect 7756 36317 7796 36688
rect 7852 36688 7988 36728
rect 8044 37780 8180 37820
rect 7755 36308 7797 36317
rect 7755 36268 7756 36308
rect 7796 36268 7797 36308
rect 7755 36259 7797 36268
rect 7852 36065 7892 36688
rect 7947 36560 7989 36569
rect 7947 36520 7948 36560
rect 7988 36520 7989 36560
rect 7947 36511 7989 36520
rect 7948 36426 7988 36511
rect 7851 36056 7893 36065
rect 7851 36016 7852 36056
rect 7892 36016 7893 36056
rect 7851 36007 7893 36016
rect 7755 35972 7797 35981
rect 7755 35932 7756 35972
rect 7796 35932 7797 35972
rect 7755 35923 7797 35932
rect 7756 35838 7796 35923
rect 7851 35888 7893 35897
rect 7851 35848 7852 35888
rect 7892 35848 7893 35888
rect 7851 35839 7893 35848
rect 7852 35754 7892 35839
rect 7755 35216 7797 35225
rect 7660 35176 7756 35216
rect 7796 35176 7797 35216
rect 7755 35167 7797 35176
rect 7756 34889 7796 35167
rect 7947 35132 7989 35141
rect 7947 35092 7948 35132
rect 7988 35092 7989 35132
rect 7947 35083 7989 35092
rect 7851 35048 7893 35057
rect 7851 35008 7852 35048
rect 7892 35008 7893 35048
rect 7851 34999 7893 35008
rect 7948 35048 7988 35083
rect 7755 34880 7797 34889
rect 7755 34840 7756 34880
rect 7796 34840 7797 34880
rect 7755 34831 7797 34840
rect 7659 34376 7701 34385
rect 7659 34336 7660 34376
rect 7700 34336 7701 34376
rect 7659 34327 7701 34336
rect 7756 34376 7796 34385
rect 7660 34242 7700 34327
rect 7756 34133 7796 34336
rect 7755 34124 7797 34133
rect 7755 34084 7756 34124
rect 7796 34084 7797 34124
rect 7755 34075 7797 34084
rect 7563 33872 7605 33881
rect 7563 33832 7564 33872
rect 7604 33832 7605 33872
rect 7563 33823 7605 33832
rect 7755 33872 7797 33881
rect 7755 33832 7756 33872
rect 7796 33832 7797 33872
rect 7755 33823 7797 33832
rect 7756 33699 7796 33823
rect 7756 33650 7796 33659
rect 7755 33116 7797 33125
rect 7755 33076 7756 33116
rect 7796 33076 7797 33116
rect 7755 33067 7797 33076
rect 7756 32982 7796 33067
rect 7371 32948 7413 32957
rect 7371 32908 7372 32948
rect 7412 32908 7413 32948
rect 7371 32899 7413 32908
rect 7180 31352 7220 31361
rect 7220 31312 7316 31352
rect 7180 31303 7220 31312
rect 7084 31144 7220 31184
rect 6987 30092 7029 30101
rect 6987 30052 6988 30092
rect 7028 30052 7029 30092
rect 6987 30043 7029 30052
rect 6987 29840 7029 29849
rect 6987 29800 6988 29840
rect 7028 29800 7029 29840
rect 6987 29791 7029 29800
rect 6988 29706 7028 29791
rect 7084 29765 7124 29850
rect 7083 29756 7125 29765
rect 7083 29716 7084 29756
rect 7124 29716 7125 29756
rect 7083 29707 7125 29716
rect 7180 29588 7220 31144
rect 7276 30857 7316 31312
rect 7275 30848 7317 30857
rect 7275 30808 7276 30848
rect 7316 30808 7317 30848
rect 7275 30799 7317 30808
rect 7276 30680 7316 30689
rect 7372 30680 7412 32899
rect 7563 32864 7605 32873
rect 7563 32824 7564 32864
rect 7604 32824 7605 32864
rect 7563 32815 7605 32824
rect 7564 32730 7604 32815
rect 7563 32444 7605 32453
rect 7563 32404 7564 32444
rect 7604 32404 7605 32444
rect 7563 32395 7605 32404
rect 7467 31520 7509 31529
rect 7467 31480 7468 31520
rect 7508 31480 7509 31520
rect 7467 31471 7509 31480
rect 7468 31025 7508 31471
rect 7467 31016 7509 31025
rect 7467 30976 7468 31016
rect 7508 30976 7509 31016
rect 7467 30967 7509 30976
rect 7316 30640 7412 30680
rect 7468 30680 7508 30689
rect 7276 30631 7316 30640
rect 7084 29548 7220 29588
rect 7372 30008 7412 30017
rect 7468 30008 7508 30640
rect 7564 30680 7604 32395
rect 7660 32192 7700 32201
rect 7660 31697 7700 32152
rect 7852 32117 7892 34999
rect 7948 34997 7988 35008
rect 7947 34880 7989 34889
rect 7947 34840 7948 34880
rect 7988 34840 7989 34880
rect 7947 34831 7989 34840
rect 7948 34049 7988 34831
rect 7947 34040 7989 34049
rect 7947 34000 7948 34040
rect 7988 34000 7989 34040
rect 7947 33991 7989 34000
rect 7948 33872 7988 33881
rect 8044 33872 8084 37780
rect 8139 37652 8181 37661
rect 8139 37612 8140 37652
rect 8180 37612 8181 37652
rect 8139 37603 8181 37612
rect 8140 37073 8180 37603
rect 8139 37064 8181 37073
rect 8139 37024 8140 37064
rect 8180 37024 8181 37064
rect 8139 37015 8181 37024
rect 8139 36896 8181 36905
rect 8139 36856 8140 36896
rect 8180 36856 8181 36896
rect 8139 36847 8181 36856
rect 8140 36762 8180 36847
rect 8139 36308 8181 36317
rect 8139 36268 8140 36308
rect 8180 36268 8181 36308
rect 8139 36259 8181 36268
rect 8140 35300 8180 36259
rect 8236 35477 8276 38704
rect 8428 38660 8468 39367
rect 8524 38744 8564 39871
rect 8715 39080 8757 39089
rect 8715 39040 8716 39080
rect 8756 39040 8757 39080
rect 8715 39031 8757 39040
rect 8620 38921 8660 39006
rect 8716 38996 8756 39031
rect 8716 38945 8756 38956
rect 8619 38912 8661 38921
rect 8619 38872 8620 38912
rect 8660 38872 8661 38912
rect 8619 38863 8661 38872
rect 8524 38704 8756 38744
rect 8428 38620 8564 38660
rect 8427 38492 8469 38501
rect 8427 38452 8428 38492
rect 8468 38452 8469 38492
rect 8427 38443 8469 38452
rect 8331 38324 8373 38333
rect 8331 38284 8332 38324
rect 8372 38284 8373 38324
rect 8331 38275 8373 38284
rect 8332 38240 8372 38275
rect 8332 36401 8372 38200
rect 8428 37913 8468 38443
rect 8427 37904 8469 37913
rect 8427 37864 8428 37904
rect 8468 37864 8469 37904
rect 8427 37855 8469 37864
rect 8428 37442 8468 37855
rect 8428 37393 8468 37402
rect 8524 37316 8564 38620
rect 8428 37276 8564 37316
rect 8331 36392 8373 36401
rect 8331 36352 8332 36392
rect 8372 36352 8373 36392
rect 8331 36343 8373 36352
rect 8331 35888 8373 35897
rect 8331 35848 8332 35888
rect 8372 35848 8373 35888
rect 8331 35839 8373 35848
rect 8332 35754 8372 35839
rect 8235 35468 8277 35477
rect 8235 35428 8236 35468
rect 8276 35428 8277 35468
rect 8235 35419 8277 35428
rect 8140 35260 8276 35300
rect 8139 35048 8181 35057
rect 8139 35008 8140 35048
rect 8180 35008 8181 35048
rect 8139 34999 8181 35008
rect 8140 34914 8180 34999
rect 8236 34889 8276 35260
rect 8331 35216 8373 35225
rect 8331 35176 8332 35216
rect 8372 35176 8373 35216
rect 8331 35167 8373 35176
rect 8332 35082 8372 35167
rect 8235 34880 8277 34889
rect 8235 34840 8236 34880
rect 8276 34840 8277 34880
rect 8235 34831 8277 34840
rect 8428 34721 8468 37276
rect 8620 37232 8660 37241
rect 8524 37192 8620 37232
rect 8524 36728 8564 37192
rect 8620 37183 8660 37192
rect 8524 36679 8564 36688
rect 8619 36728 8661 36737
rect 8619 36688 8620 36728
rect 8660 36688 8661 36728
rect 8619 36679 8661 36688
rect 8620 36594 8660 36679
rect 8427 34712 8469 34721
rect 8427 34672 8428 34712
rect 8468 34672 8469 34712
rect 8427 34663 8469 34672
rect 8139 34544 8181 34553
rect 8139 34504 8140 34544
rect 8180 34504 8181 34544
rect 8139 34495 8181 34504
rect 8331 34544 8373 34553
rect 8331 34504 8332 34544
rect 8372 34504 8373 34544
rect 8331 34495 8373 34504
rect 8140 34376 8180 34495
rect 8236 34385 8276 34470
rect 8140 34327 8180 34336
rect 8235 34376 8277 34385
rect 8235 34336 8236 34376
rect 8276 34336 8277 34376
rect 8235 34327 8277 34336
rect 8332 34376 8372 34495
rect 8716 34460 8756 38704
rect 8908 37820 8948 42928
rect 9100 42281 9140 42928
rect 9099 42272 9141 42281
rect 9099 42232 9100 42272
rect 9140 42232 9141 42272
rect 9099 42223 9141 42232
rect 9195 42104 9237 42113
rect 9195 42064 9196 42104
rect 9236 42064 9237 42104
rect 9195 42055 9237 42064
rect 9099 41096 9141 41105
rect 9099 41056 9100 41096
rect 9140 41056 9141 41096
rect 9099 41047 9141 41056
rect 9100 40349 9140 41047
rect 9099 40340 9141 40349
rect 9099 40300 9100 40340
rect 9140 40300 9141 40340
rect 9099 40291 9141 40300
rect 9099 39752 9141 39761
rect 9099 39712 9100 39752
rect 9140 39712 9141 39752
rect 9099 39703 9141 39712
rect 9100 39341 9140 39703
rect 9099 39332 9141 39341
rect 9099 39292 9100 39332
rect 9140 39292 9141 39332
rect 9099 39283 9141 39292
rect 9003 38912 9045 38921
rect 9003 38872 9004 38912
rect 9044 38872 9045 38912
rect 9003 38863 9045 38872
rect 9004 37997 9044 38863
rect 9003 37988 9045 37997
rect 9003 37948 9004 37988
rect 9044 37948 9045 37988
rect 9003 37939 9045 37948
rect 8812 37780 8948 37820
rect 9100 37820 9140 39283
rect 9196 38912 9236 42055
rect 9292 40592 9332 42928
rect 9484 42197 9524 42928
rect 9676 42701 9716 42928
rect 9675 42692 9717 42701
rect 9675 42652 9676 42692
rect 9716 42652 9717 42692
rect 9675 42643 9717 42652
rect 9483 42188 9525 42197
rect 9483 42148 9484 42188
rect 9524 42148 9525 42188
rect 9483 42139 9525 42148
rect 9484 41264 9524 41275
rect 9868 41264 9908 42928
rect 10060 42197 10100 42928
rect 10059 42188 10101 42197
rect 10059 42148 10060 42188
rect 10100 42148 10101 42188
rect 10059 42139 10101 42148
rect 10252 41441 10292 42928
rect 10444 41525 10484 42928
rect 10443 41516 10485 41525
rect 10636 41516 10676 42928
rect 10828 41684 10868 42928
rect 11020 41777 11060 42928
rect 11019 41768 11061 41777
rect 11019 41728 11020 41768
rect 11060 41728 11061 41768
rect 11019 41719 11061 41728
rect 10443 41476 10444 41516
rect 10484 41476 10485 41516
rect 10443 41467 10485 41476
rect 10540 41476 10676 41516
rect 10732 41644 10868 41684
rect 10251 41432 10293 41441
rect 10251 41392 10252 41432
rect 10292 41392 10293 41432
rect 10251 41383 10293 41392
rect 9484 41189 9524 41224
rect 9772 41224 9908 41264
rect 10252 41264 10292 41273
rect 9483 41180 9525 41189
rect 9483 41140 9484 41180
rect 9524 41140 9525 41180
rect 9483 41131 9525 41140
rect 9675 41012 9717 41021
rect 9675 40972 9676 41012
rect 9716 40972 9717 41012
rect 9675 40963 9717 40972
rect 9676 40878 9716 40963
rect 9579 40592 9621 40601
rect 9292 40552 9428 40592
rect 9292 40424 9332 40435
rect 9292 40349 9332 40384
rect 9291 40340 9333 40349
rect 9291 40300 9292 40340
rect 9332 40300 9333 40340
rect 9291 40291 9333 40300
rect 9292 39929 9332 40291
rect 9291 39920 9333 39929
rect 9291 39880 9292 39920
rect 9332 39880 9333 39920
rect 9291 39871 9333 39880
rect 9291 39668 9333 39677
rect 9291 39628 9292 39668
rect 9332 39628 9333 39668
rect 9291 39619 9333 39628
rect 9196 38863 9236 38872
rect 9292 38249 9332 39619
rect 9291 38240 9333 38249
rect 9291 38200 9292 38240
rect 9332 38200 9333 38240
rect 9291 38191 9333 38200
rect 9100 37780 9236 37820
rect 8812 36989 8852 37780
rect 9196 37661 9236 37780
rect 9003 37652 9045 37661
rect 9195 37652 9237 37661
rect 9388 37652 9428 40552
rect 9579 40552 9580 40592
rect 9620 40552 9621 40592
rect 9579 40543 9621 40552
rect 9483 40340 9525 40349
rect 9483 40300 9484 40340
rect 9524 40300 9525 40340
rect 9483 40291 9525 40300
rect 9484 40206 9524 40291
rect 9483 39920 9525 39929
rect 9483 39880 9484 39920
rect 9524 39880 9525 39920
rect 9483 39871 9525 39880
rect 9484 39752 9524 39871
rect 9484 39005 9524 39712
rect 9580 39332 9620 40543
rect 9675 40172 9717 40181
rect 9675 40132 9676 40172
rect 9716 40132 9717 40172
rect 9675 40123 9717 40132
rect 9676 39929 9716 40123
rect 9675 39920 9717 39929
rect 9675 39880 9676 39920
rect 9716 39880 9717 39920
rect 9675 39871 9717 39880
rect 9676 39509 9716 39594
rect 9675 39500 9717 39509
rect 9675 39460 9676 39500
rect 9716 39460 9717 39500
rect 9675 39451 9717 39460
rect 9580 39292 9716 39332
rect 9483 38996 9525 39005
rect 9483 38956 9484 38996
rect 9524 38956 9525 38996
rect 9483 38947 9525 38956
rect 9676 38926 9716 39292
rect 9676 38877 9716 38886
rect 9772 38828 9812 41224
rect 10155 41180 10197 41189
rect 10060 41140 10156 41180
rect 10196 41140 10197 41180
rect 9868 41096 9908 41105
rect 10060 41096 10100 41140
rect 10155 41131 10197 41140
rect 9908 41056 10100 41096
rect 9868 39584 9908 41056
rect 10156 41012 10196 41021
rect 10156 40769 10196 40972
rect 10155 40760 10197 40769
rect 10155 40720 10156 40760
rect 10196 40720 10197 40760
rect 10155 40711 10197 40720
rect 9963 40424 10005 40433
rect 9963 40384 9964 40424
rect 10004 40384 10005 40424
rect 9963 40375 10005 40384
rect 10060 40424 10100 40433
rect 9964 40290 10004 40375
rect 10060 40181 10100 40384
rect 10059 40172 10101 40181
rect 10059 40132 10060 40172
rect 10100 40132 10101 40172
rect 10059 40123 10101 40132
rect 10155 39920 10197 39929
rect 10155 39880 10156 39920
rect 10196 39880 10197 39920
rect 10155 39871 10197 39880
rect 9963 39836 10005 39845
rect 9963 39796 9964 39836
rect 10004 39796 10005 39836
rect 9963 39787 10005 39796
rect 9868 39509 9908 39544
rect 9867 39500 9909 39509
rect 9867 39460 9868 39500
rect 9908 39460 9909 39500
rect 9867 39451 9909 39460
rect 9867 39332 9909 39341
rect 9867 39292 9868 39332
rect 9908 39292 9909 39332
rect 9867 39283 9909 39292
rect 9484 38788 9812 38828
rect 9868 38828 9908 39283
rect 9484 37829 9524 38788
rect 9868 38779 9908 38788
rect 9964 38576 10004 39787
rect 10060 39761 10100 39780
rect 10059 39752 10101 39761
rect 10156 39752 10196 39871
rect 10059 39712 10060 39752
rect 10100 39712 10196 39752
rect 10059 39703 10101 39712
rect 10156 39665 10196 39712
rect 10156 39616 10196 39625
rect 10252 39080 10292 41224
rect 10540 41189 10580 41476
rect 10636 41273 10676 41358
rect 10635 41264 10677 41273
rect 10635 41224 10636 41264
rect 10676 41224 10677 41264
rect 10635 41215 10677 41224
rect 10539 41180 10581 41189
rect 10539 41140 10540 41180
rect 10580 41140 10581 41180
rect 10539 41131 10581 41140
rect 10444 40508 10484 40532
rect 10444 40447 10484 40468
rect 10540 40508 10580 41131
rect 10732 40517 10772 41644
rect 10827 41516 10869 41525
rect 10827 41476 10828 41516
rect 10868 41476 10869 41516
rect 10827 41467 10869 41476
rect 10540 40459 10580 40468
rect 10731 40508 10773 40517
rect 10731 40468 10732 40508
rect 10772 40468 10773 40508
rect 10731 40459 10773 40468
rect 10442 40438 10484 40447
rect 10442 40398 10443 40438
rect 10483 40398 10484 40438
rect 10442 40389 10484 40398
rect 10731 40340 10773 40349
rect 10731 40300 10732 40340
rect 10772 40300 10773 40340
rect 10731 40291 10773 40300
rect 10347 40088 10389 40097
rect 10347 40048 10348 40088
rect 10388 40048 10389 40088
rect 10347 40039 10389 40048
rect 10348 39929 10388 40039
rect 10347 39920 10389 39929
rect 10347 39880 10348 39920
rect 10388 39880 10389 39920
rect 10347 39871 10389 39880
rect 10539 39920 10581 39929
rect 10539 39880 10540 39920
rect 10580 39880 10581 39920
rect 10539 39871 10581 39880
rect 10540 39786 10580 39871
rect 10347 39500 10389 39509
rect 10347 39460 10348 39500
rect 10388 39460 10389 39500
rect 10347 39451 10389 39460
rect 10348 39366 10388 39451
rect 10732 39416 10772 40291
rect 10828 39920 10868 41467
rect 11019 41180 11061 41189
rect 11019 41140 11020 41180
rect 11060 41140 11061 41180
rect 11019 41131 11061 41140
rect 11020 40424 11060 41131
rect 11020 40375 11060 40384
rect 11019 40172 11061 40181
rect 11019 40132 11020 40172
rect 11060 40132 11061 40172
rect 11019 40123 11061 40132
rect 10828 39871 10868 39880
rect 10924 39584 10964 39593
rect 10732 39376 10868 39416
rect 10156 39040 10292 39080
rect 10059 38744 10101 38753
rect 10059 38704 10060 38744
rect 10100 38704 10101 38744
rect 10059 38695 10101 38704
rect 10060 38610 10100 38695
rect 9676 38536 10004 38576
rect 9579 38492 9621 38501
rect 9579 38452 9580 38492
rect 9620 38452 9621 38492
rect 9579 38443 9621 38452
rect 9580 38240 9620 38443
rect 9580 38191 9620 38200
rect 9579 38072 9621 38081
rect 9579 38032 9580 38072
rect 9620 38032 9621 38072
rect 9579 38023 9621 38032
rect 9483 37820 9525 37829
rect 9483 37780 9484 37820
rect 9524 37780 9525 37820
rect 9483 37771 9525 37780
rect 9003 37612 9004 37652
rect 9044 37612 9140 37652
rect 9003 37603 9045 37612
rect 9003 37400 9045 37409
rect 9003 37360 9004 37400
rect 9044 37360 9045 37400
rect 9003 37351 9045 37360
rect 9100 37400 9140 37612
rect 9195 37612 9196 37652
rect 9236 37612 9237 37652
rect 9195 37603 9237 37612
rect 9292 37612 9428 37652
rect 9483 37652 9525 37661
rect 9483 37612 9484 37652
rect 9524 37612 9525 37652
rect 9100 37351 9140 37360
rect 9196 37400 9236 37409
rect 8908 37232 8948 37241
rect 8811 36980 8853 36989
rect 8811 36940 8812 36980
rect 8852 36940 8853 36980
rect 8811 36931 8853 36940
rect 8908 36653 8948 37192
rect 9004 36905 9044 37351
rect 9003 36896 9045 36905
rect 9003 36856 9004 36896
rect 9044 36856 9045 36896
rect 9003 36847 9045 36856
rect 9004 36728 9044 36847
rect 9004 36679 9044 36688
rect 9099 36728 9141 36737
rect 9099 36688 9100 36728
rect 9140 36688 9141 36728
rect 9099 36679 9141 36688
rect 8907 36644 8949 36653
rect 8907 36604 8908 36644
rect 8948 36604 8949 36644
rect 8907 36595 8949 36604
rect 9100 36594 9140 36679
rect 9196 36569 9236 37360
rect 8811 36560 8853 36569
rect 8811 36520 8812 36560
rect 8852 36520 8853 36560
rect 8811 36511 8853 36520
rect 9195 36560 9237 36569
rect 9195 36520 9196 36560
rect 9236 36520 9237 36560
rect 9195 36511 9237 36520
rect 8812 35902 8852 36511
rect 9292 36140 9332 37612
rect 9483 37603 9525 37612
rect 9580 37652 9620 38023
rect 9580 37603 9620 37612
rect 9387 37484 9429 37493
rect 9387 37444 9388 37484
rect 9428 37444 9429 37484
rect 9387 37435 9429 37444
rect 9388 37350 9428 37435
rect 9484 36560 9524 37603
rect 9580 36728 9620 36737
rect 9676 36728 9716 38536
rect 9867 38240 9909 38249
rect 9867 38200 9868 38240
rect 9908 38200 9909 38240
rect 9867 38191 9909 38200
rect 10059 38240 10101 38249
rect 10059 38200 10060 38240
rect 10100 38200 10101 38240
rect 10059 38191 10101 38200
rect 9771 37988 9813 37997
rect 9771 37948 9772 37988
rect 9812 37948 9813 37988
rect 9771 37939 9813 37948
rect 9772 37854 9812 37939
rect 9771 37652 9813 37661
rect 9771 37612 9772 37652
rect 9812 37612 9813 37652
rect 9771 37603 9813 37612
rect 9772 37400 9812 37603
rect 9772 37351 9812 37360
rect 9771 36980 9813 36989
rect 9771 36940 9772 36980
rect 9812 36940 9813 36980
rect 9771 36931 9813 36940
rect 9620 36688 9716 36728
rect 9580 36679 9620 36688
rect 9484 36520 9716 36560
rect 8812 35853 8852 35862
rect 9100 36100 9332 36140
rect 9003 35804 9045 35813
rect 9003 35764 9004 35804
rect 9044 35764 9045 35804
rect 9003 35755 9045 35764
rect 8811 35720 8853 35729
rect 8811 35680 8812 35720
rect 8852 35680 8853 35720
rect 8811 35671 8853 35680
rect 8812 34544 8852 35671
rect 9004 35670 9044 35755
rect 8907 35132 8949 35141
rect 8907 35092 8908 35132
rect 8948 35092 8949 35132
rect 8907 35083 8949 35092
rect 8812 34495 8852 34504
rect 8716 34411 8756 34420
rect 8908 34460 8948 35083
rect 8908 34411 8948 34420
rect 8620 34376 8660 34385
rect 8332 34327 8372 34336
rect 8524 34336 8620 34376
rect 8428 34208 8468 34217
rect 7988 33832 8084 33872
rect 8140 34168 8428 34208
rect 7948 33823 7988 33832
rect 8140 33690 8180 34168
rect 8428 34159 8468 34168
rect 8331 33956 8373 33965
rect 8331 33916 8332 33956
rect 8372 33916 8373 33956
rect 8331 33907 8373 33916
rect 8044 33650 8180 33690
rect 7947 33116 7989 33125
rect 7947 33076 7948 33116
rect 7988 33076 7989 33116
rect 7947 33067 7989 33076
rect 7948 32864 7988 33067
rect 7948 32815 7988 32824
rect 8044 32276 8084 33650
rect 8140 33536 8180 33545
rect 8140 32360 8180 33496
rect 8235 33452 8277 33461
rect 8235 33412 8236 33452
rect 8276 33412 8277 33452
rect 8235 33403 8277 33412
rect 8140 32311 8180 32320
rect 7948 32236 8084 32276
rect 7851 32108 7893 32117
rect 7851 32068 7852 32108
rect 7892 32068 7893 32108
rect 7851 32059 7893 32068
rect 7852 31940 7892 31949
rect 7756 31900 7852 31940
rect 7659 31688 7701 31697
rect 7659 31648 7660 31688
rect 7700 31648 7701 31688
rect 7659 31639 7701 31648
rect 7660 31529 7700 31639
rect 7659 31520 7701 31529
rect 7659 31480 7660 31520
rect 7700 31480 7701 31520
rect 7659 31471 7701 31480
rect 7756 31394 7796 31900
rect 7852 31891 7892 31900
rect 7660 31366 7796 31394
rect 7700 31354 7796 31366
rect 7660 31317 7700 31326
rect 7851 31268 7893 31277
rect 7851 31228 7852 31268
rect 7892 31228 7893 31268
rect 7851 31219 7893 31228
rect 7852 31134 7892 31219
rect 7948 31016 7988 32236
rect 8044 32033 8084 32118
rect 8139 32108 8181 32117
rect 8139 32068 8140 32108
rect 8180 32068 8181 32108
rect 8139 32059 8181 32068
rect 8043 32024 8085 32033
rect 8043 31984 8044 32024
rect 8084 31984 8085 32024
rect 8043 31975 8085 31984
rect 8140 31856 8180 32059
rect 8044 31816 8180 31856
rect 8044 31352 8084 31816
rect 8139 31436 8181 31445
rect 8139 31396 8140 31436
rect 8180 31396 8181 31436
rect 8139 31387 8181 31396
rect 8044 31303 8084 31312
rect 8140 31302 8180 31387
rect 8236 31352 8276 33403
rect 8332 33125 8372 33907
rect 8427 33788 8469 33797
rect 8427 33748 8428 33788
rect 8468 33748 8469 33788
rect 8427 33739 8469 33748
rect 8428 33654 8468 33739
rect 8331 33116 8373 33125
rect 8331 33076 8332 33116
rect 8372 33076 8373 33116
rect 8331 33067 8373 33076
rect 8427 32696 8469 32705
rect 8427 32656 8428 32696
rect 8468 32656 8469 32696
rect 8427 32647 8469 32656
rect 8331 32192 8373 32201
rect 8331 32152 8332 32192
rect 8372 32152 8373 32192
rect 8331 32143 8373 32152
rect 8332 32058 8372 32143
rect 8428 31520 8468 32647
rect 8524 32621 8564 34336
rect 8620 34327 8660 34336
rect 9004 34376 9044 34385
rect 8811 34292 8853 34301
rect 8811 34252 8812 34292
rect 8852 34252 8853 34292
rect 8811 34243 8853 34252
rect 8715 34208 8757 34217
rect 8715 34168 8716 34208
rect 8756 34168 8757 34208
rect 8715 34159 8757 34168
rect 8619 33956 8661 33965
rect 8619 33916 8620 33956
rect 8660 33916 8661 33956
rect 8619 33907 8661 33916
rect 8620 33704 8660 33907
rect 8620 33209 8660 33664
rect 8619 33200 8661 33209
rect 8619 33160 8620 33200
rect 8660 33160 8661 33200
rect 8619 33151 8661 33160
rect 8523 32612 8565 32621
rect 8523 32572 8524 32612
rect 8564 32572 8565 32612
rect 8523 32563 8565 32572
rect 8619 32528 8661 32537
rect 8619 32488 8620 32528
rect 8660 32488 8661 32528
rect 8619 32479 8661 32488
rect 8523 32192 8565 32201
rect 8523 32152 8524 32192
rect 8564 32152 8565 32192
rect 8523 32143 8565 32152
rect 8620 32192 8660 32479
rect 8620 32143 8660 32152
rect 8524 32058 8564 32143
rect 8619 32024 8661 32033
rect 8619 31984 8620 32024
rect 8660 31984 8661 32024
rect 8619 31975 8661 31984
rect 8620 31890 8660 31975
rect 8236 31303 8276 31312
rect 8332 31480 8468 31520
rect 7564 30631 7604 30640
rect 7660 30976 7988 31016
rect 7660 30680 7700 30976
rect 7660 30631 7700 30640
rect 7755 30680 7797 30689
rect 7948 30680 7988 30689
rect 7755 30640 7756 30680
rect 7796 30640 7892 30680
rect 7755 30631 7797 30640
rect 7756 30546 7796 30631
rect 7468 29968 7796 30008
rect 6891 29504 6933 29513
rect 6891 29464 6892 29504
rect 6932 29464 6933 29504
rect 6891 29455 6933 29464
rect 6988 29168 7028 29177
rect 6796 29128 6988 29168
rect 6988 29119 7028 29128
rect 6644 28960 6740 29000
rect 6604 28951 6644 28960
rect 6796 28916 6836 28925
rect 6508 28624 6644 28664
rect 6315 28580 6357 28589
rect 6315 28540 6316 28580
rect 6356 28540 6357 28580
rect 6315 28531 6357 28540
rect 6604 28505 6644 28624
rect 5932 28421 5972 28456
rect 6124 28456 6260 28496
rect 6412 28496 6452 28505
rect 5931 28412 5973 28421
rect 5931 28372 5932 28412
rect 5972 28372 5973 28412
rect 5931 28363 5973 28372
rect 6027 28328 6069 28337
rect 6027 28288 6028 28328
rect 6068 28288 6069 28328
rect 6027 28279 6069 28288
rect 5835 27908 5877 27917
rect 5835 27868 5836 27908
rect 5876 27868 5877 27908
rect 5835 27859 5877 27868
rect 5739 27740 5781 27749
rect 5739 27700 5740 27740
rect 5780 27700 5781 27740
rect 5739 27691 5781 27700
rect 5548 27656 5588 27665
rect 5588 27616 5684 27656
rect 5548 27607 5588 27616
rect 5644 27077 5684 27616
rect 5740 27404 5780 27413
rect 5780 27364 5972 27404
rect 5740 27355 5780 27364
rect 5739 27152 5781 27161
rect 5739 27112 5740 27152
rect 5780 27112 5781 27152
rect 5739 27103 5781 27112
rect 5643 27068 5685 27077
rect 5643 27028 5644 27068
rect 5684 27028 5685 27068
rect 5643 27019 5685 27028
rect 5644 26816 5684 27019
rect 5644 26767 5684 26776
rect 5356 26692 5588 26732
rect 5451 26564 5493 26573
rect 5451 26524 5452 26564
rect 5492 26524 5493 26564
rect 5451 26515 5493 26524
rect 4928 26480 5296 26489
rect 4968 26440 5010 26480
rect 5050 26440 5092 26480
rect 5132 26440 5174 26480
rect 5214 26440 5256 26480
rect 4928 26431 5296 26440
rect 4875 26228 4917 26237
rect 4875 26188 4876 26228
rect 4916 26188 4917 26228
rect 4875 26179 4917 26188
rect 4780 26095 4820 26104
rect 4587 26060 4629 26069
rect 4587 26020 4588 26060
rect 4628 26020 4629 26060
rect 4587 26011 4629 26020
rect 4587 25892 4629 25901
rect 4587 25852 4588 25892
rect 4628 25852 4629 25892
rect 4587 25843 4629 25852
rect 4588 25758 4628 25843
rect 4492 25600 4724 25640
rect 4299 25472 4341 25481
rect 4299 25432 4300 25472
rect 4340 25432 4341 25472
rect 4299 25423 4341 25432
rect 3436 25255 3476 25264
rect 3243 25136 3285 25145
rect 3243 25096 3244 25136
rect 3284 25096 3285 25136
rect 3243 25087 3285 25096
rect 3531 25136 3573 25145
rect 3531 25096 3532 25136
rect 3572 25096 3573 25136
rect 3531 25087 3573 25096
rect 3147 24716 3189 24725
rect 3147 24676 3148 24716
rect 3188 24676 3189 24716
rect 3147 24667 3189 24676
rect 3052 24632 3092 24641
rect 3052 24473 3092 24592
rect 3148 24582 3188 24667
rect 2859 24464 2901 24473
rect 2859 24424 2860 24464
rect 2900 24424 2901 24464
rect 2859 24415 2901 24424
rect 3051 24464 3093 24473
rect 3051 24424 3052 24464
rect 3092 24424 3093 24464
rect 3051 24415 3093 24424
rect 2860 24330 2900 24415
rect 2764 24172 2900 24212
rect 2860 23129 2900 24172
rect 2956 23792 2996 23801
rect 2859 23120 2901 23129
rect 2859 23080 2860 23120
rect 2900 23080 2901 23120
rect 2859 23071 2901 23080
rect 2956 23045 2996 23752
rect 3051 23792 3093 23801
rect 3051 23752 3052 23792
rect 3092 23752 3093 23792
rect 3051 23743 3093 23752
rect 3052 23658 3092 23743
rect 3244 23129 3284 25087
rect 3436 24632 3476 24641
rect 3340 24592 3436 24632
rect 3340 23969 3380 24592
rect 3436 24583 3476 24592
rect 3435 24464 3477 24473
rect 3435 24424 3436 24464
rect 3476 24424 3477 24464
rect 3435 24415 3477 24424
rect 3436 24053 3476 24415
rect 3435 24044 3477 24053
rect 3435 24004 3436 24044
rect 3476 24004 3477 24044
rect 3435 23995 3477 24004
rect 3339 23960 3381 23969
rect 3339 23920 3340 23960
rect 3380 23920 3381 23960
rect 3532 23960 3572 25087
rect 3628 24893 3668 25264
rect 4011 25220 4053 25229
rect 4011 25180 4012 25220
rect 4052 25180 4053 25220
rect 4011 25171 4053 25180
rect 3627 24884 3669 24893
rect 3627 24844 3628 24884
rect 3668 24844 3669 24884
rect 3627 24835 3669 24844
rect 3819 24632 3861 24641
rect 3819 24592 3820 24632
rect 3860 24592 3861 24632
rect 3819 24583 3861 24592
rect 3916 24632 3956 24641
rect 3820 24498 3860 24583
rect 3628 24389 3668 24474
rect 3627 24380 3669 24389
rect 3627 24340 3628 24380
rect 3668 24340 3669 24380
rect 3916 24380 3956 24592
rect 4012 24632 4052 25171
rect 4395 24716 4437 24725
rect 4378 24676 4396 24716
rect 4436 24676 4628 24716
rect 4378 24667 4437 24676
rect 4378 24647 4418 24667
rect 4012 24583 4052 24592
rect 4107 24632 4149 24641
rect 4107 24592 4108 24632
rect 4148 24592 4149 24632
rect 4378 24598 4418 24607
rect 4107 24583 4149 24592
rect 4108 24498 4148 24583
rect 4395 24380 4437 24389
rect 3916 24340 4340 24380
rect 3627 24331 3669 24340
rect 3688 24212 4056 24221
rect 3728 24172 3770 24212
rect 3810 24172 3852 24212
rect 3892 24172 3934 24212
rect 3974 24172 4016 24212
rect 3688 24163 4056 24172
rect 4011 24044 4053 24053
rect 4011 24004 4012 24044
rect 4052 24004 4053 24044
rect 4011 23995 4053 24004
rect 3532 23920 3668 23960
rect 3339 23911 3381 23920
rect 3339 23792 3381 23801
rect 3532 23792 3572 23801
rect 3339 23752 3340 23792
rect 3380 23752 3381 23792
rect 3339 23743 3381 23752
rect 3436 23752 3532 23792
rect 3340 23288 3380 23743
rect 3340 23239 3380 23248
rect 3148 23120 3188 23129
rect 3243 23120 3285 23129
rect 3436 23120 3476 23752
rect 3532 23743 3572 23752
rect 3628 23288 3668 23920
rect 4012 23806 4052 23995
rect 4203 23960 4245 23969
rect 4203 23920 4204 23960
rect 4244 23920 4245 23960
rect 4203 23911 4245 23920
rect 4012 23757 4052 23766
rect 4204 23708 4244 23911
rect 4204 23659 4244 23668
rect 3628 23239 3668 23248
rect 4300 23288 4340 24340
rect 4395 24340 4396 24380
rect 4436 24340 4437 24380
rect 4395 24331 4437 24340
rect 4300 23239 4340 23248
rect 3820 23120 3860 23129
rect 3188 23080 3244 23120
rect 3284 23080 3285 23120
rect 3148 23071 3188 23080
rect 3243 23071 3285 23080
rect 3340 23080 3476 23120
rect 3532 23080 3820 23120
rect 2955 23036 2997 23045
rect 2955 22996 2956 23036
rect 2996 22996 2997 23036
rect 2955 22987 2997 22996
rect 3244 22986 3284 23071
rect 2955 22868 2997 22877
rect 2955 22828 2956 22868
rect 2996 22828 2997 22868
rect 2955 22819 2997 22828
rect 2859 22700 2901 22709
rect 2859 22660 2860 22700
rect 2900 22660 2901 22700
rect 2859 22651 2901 22660
rect 2476 21533 2516 22240
rect 2572 22240 2708 22280
rect 2572 21953 2612 22240
rect 2860 22121 2900 22651
rect 2956 22280 2996 22819
rect 3340 22625 3380 23080
rect 3532 23036 3572 23080
rect 3820 23071 3860 23080
rect 4012 23120 4052 23129
rect 3436 22996 3572 23036
rect 3436 22709 3476 22996
rect 3628 22952 3668 22961
rect 3532 22912 3628 22952
rect 3435 22700 3477 22709
rect 3435 22660 3436 22700
rect 3476 22660 3477 22700
rect 3435 22651 3477 22660
rect 3339 22616 3381 22625
rect 3339 22576 3340 22616
rect 3380 22576 3381 22616
rect 3339 22567 3381 22576
rect 3532 22532 3572 22912
rect 3628 22903 3668 22912
rect 3820 22877 3860 22962
rect 3819 22868 3861 22877
rect 3819 22828 3820 22868
rect 3860 22828 3861 22868
rect 4012 22868 4052 23080
rect 4108 23120 4148 23131
rect 4108 23045 4148 23080
rect 4396 23120 4436 24331
rect 4588 23960 4628 24676
rect 4684 24632 4724 25600
rect 4876 25397 4916 26179
rect 5068 26144 5108 26155
rect 5356 26153 5396 26238
rect 5068 26069 5108 26104
rect 5355 26144 5397 26153
rect 5355 26104 5356 26144
rect 5396 26104 5397 26144
rect 5355 26095 5397 26104
rect 5452 26144 5492 26515
rect 5067 26060 5109 26069
rect 5067 26020 5068 26060
rect 5108 26020 5109 26060
rect 5067 26011 5109 26020
rect 5452 25976 5492 26104
rect 5164 25936 5492 25976
rect 4875 25388 4917 25397
rect 4875 25348 4876 25388
rect 4916 25348 4917 25388
rect 4875 25339 4917 25348
rect 4876 25304 4916 25339
rect 5164 25313 5204 25936
rect 4876 25253 4916 25264
rect 5163 25304 5205 25313
rect 5163 25264 5164 25304
rect 5204 25264 5205 25304
rect 5163 25255 5205 25264
rect 5260 25304 5300 25315
rect 5548 25313 5588 26692
rect 5643 26480 5685 26489
rect 5643 26440 5644 26480
rect 5684 26440 5685 26480
rect 5643 26431 5685 26440
rect 5644 25556 5684 26431
rect 5740 25976 5780 27103
rect 5932 26741 5972 27364
rect 5931 26732 5973 26741
rect 5931 26692 5932 26732
rect 5972 26692 5973 26732
rect 5931 26683 5973 26692
rect 5740 25927 5780 25936
rect 5836 26648 5876 26657
rect 5644 25507 5684 25516
rect 5836 25472 5876 26608
rect 5932 26228 5972 26683
rect 6028 26648 6068 28279
rect 6124 27833 6164 28456
rect 6316 28412 6356 28421
rect 6219 28328 6261 28337
rect 6219 28288 6220 28328
rect 6260 28288 6261 28328
rect 6219 28279 6261 28288
rect 6220 28194 6260 28279
rect 6123 27824 6165 27833
rect 6123 27784 6124 27824
rect 6164 27784 6165 27824
rect 6123 27775 6165 27784
rect 6124 27656 6164 27665
rect 6124 27413 6164 27616
rect 6123 27404 6165 27413
rect 6123 27364 6124 27404
rect 6164 27364 6165 27404
rect 6123 27355 6165 27364
rect 6219 27152 6261 27161
rect 6219 27112 6220 27152
rect 6260 27112 6261 27152
rect 6219 27103 6261 27112
rect 6220 27026 6260 27103
rect 6220 26986 6270 27026
rect 6124 26825 6164 26910
rect 6230 26900 6270 26986
rect 6316 26984 6356 28372
rect 6412 28085 6452 28456
rect 6603 28496 6645 28505
rect 6603 28456 6604 28496
rect 6644 28456 6645 28496
rect 6603 28447 6645 28456
rect 6507 28412 6549 28421
rect 6507 28372 6508 28412
rect 6548 28372 6549 28412
rect 6507 28363 6549 28372
rect 6508 28278 6548 28363
rect 6796 28337 6836 28876
rect 6604 28328 6644 28337
rect 6795 28328 6837 28337
rect 6644 28288 6740 28328
rect 6604 28279 6644 28288
rect 6411 28076 6453 28085
rect 6411 28036 6412 28076
rect 6452 28036 6453 28076
rect 6411 28027 6453 28036
rect 6603 27824 6645 27833
rect 6603 27784 6604 27824
rect 6644 27784 6645 27824
rect 6603 27775 6645 27784
rect 6411 27152 6453 27161
rect 6411 27112 6412 27152
rect 6452 27112 6453 27152
rect 6411 27103 6453 27112
rect 6316 26935 6356 26944
rect 6230 26851 6270 26860
rect 6412 26900 6452 27103
rect 6507 26984 6549 26993
rect 6507 26944 6508 26984
rect 6548 26944 6549 26984
rect 6507 26935 6549 26944
rect 6123 26816 6165 26825
rect 6123 26776 6124 26816
rect 6164 26776 6165 26816
rect 6123 26767 6165 26776
rect 6412 26741 6452 26860
rect 6508 26816 6548 26935
rect 6508 26741 6548 26776
rect 6411 26732 6453 26741
rect 6411 26692 6412 26732
rect 6452 26692 6453 26732
rect 6508 26732 6554 26741
rect 6508 26692 6513 26732
rect 6553 26692 6554 26732
rect 6411 26683 6453 26692
rect 6512 26683 6554 26692
rect 6513 26657 6553 26683
rect 6028 26608 6260 26648
rect 5932 26188 6164 26228
rect 5932 26069 5972 26188
rect 6028 26144 6068 26188
rect 6028 26095 6068 26104
rect 5931 26060 5973 26069
rect 5931 26020 5932 26060
rect 5972 26020 5973 26060
rect 5931 26011 5973 26020
rect 5836 25432 6068 25472
rect 5260 25229 5300 25264
rect 5452 25304 5492 25313
rect 5067 25220 5109 25229
rect 5067 25180 5068 25220
rect 5108 25180 5109 25220
rect 5067 25171 5109 25180
rect 5259 25220 5301 25229
rect 5259 25180 5260 25220
rect 5300 25180 5301 25220
rect 5259 25171 5301 25180
rect 5068 25086 5108 25171
rect 5356 25145 5396 25230
rect 5355 25136 5397 25145
rect 5355 25096 5356 25136
rect 5396 25096 5397 25136
rect 5355 25087 5397 25096
rect 4928 24968 5296 24977
rect 5452 24968 5492 25264
rect 5547 25304 5589 25313
rect 5547 25264 5548 25304
rect 5588 25264 5589 25304
rect 5547 25255 5589 25264
rect 5740 25304 5780 25313
rect 5836 25304 5876 25432
rect 5780 25264 5876 25304
rect 5931 25304 5973 25313
rect 5931 25264 5932 25304
rect 5972 25264 5973 25304
rect 5740 25255 5780 25264
rect 5931 25255 5973 25264
rect 6028 25304 6068 25432
rect 6124 25304 6164 26188
rect 6220 25556 6260 26608
rect 6507 26480 6549 26489
rect 6507 26440 6508 26480
rect 6548 26440 6549 26480
rect 6507 26431 6549 26440
rect 6315 26396 6357 26405
rect 6315 26356 6316 26396
rect 6356 26356 6357 26396
rect 6315 26347 6357 26356
rect 6220 25507 6260 25516
rect 6316 26144 6356 26347
rect 6411 26312 6453 26321
rect 6411 26272 6412 26312
rect 6452 26272 6453 26312
rect 6411 26263 6453 26272
rect 6220 25304 6260 25313
rect 6124 25264 6220 25304
rect 6028 25255 6068 25264
rect 6220 25255 6260 25264
rect 5643 25136 5685 25145
rect 5643 25096 5644 25136
rect 5684 25096 5685 25136
rect 5643 25087 5685 25096
rect 5835 25136 5877 25145
rect 5835 25096 5836 25136
rect 5876 25096 5877 25136
rect 5835 25087 5877 25096
rect 4968 24928 5010 24968
rect 5050 24928 5092 24968
rect 5132 24928 5174 24968
rect 5214 24928 5256 24968
rect 4928 24919 5296 24928
rect 5356 24928 5492 24968
rect 5356 24800 5396 24928
rect 5164 24760 5396 24800
rect 4779 24716 4821 24725
rect 4779 24676 4780 24716
rect 4820 24676 4821 24716
rect 4779 24667 4821 24676
rect 4684 24464 4724 24592
rect 4780 24582 4820 24667
rect 5164 24632 5204 24760
rect 4972 24592 5204 24632
rect 5260 24632 5300 24641
rect 4684 24424 4820 24464
rect 4588 23920 4724 23960
rect 4491 23792 4533 23801
rect 4491 23752 4492 23792
rect 4532 23752 4533 23792
rect 4491 23743 4533 23752
rect 4588 23792 4628 23803
rect 4492 23658 4532 23743
rect 4588 23717 4628 23752
rect 4587 23708 4629 23717
rect 4587 23668 4588 23708
rect 4628 23668 4629 23708
rect 4587 23659 4629 23668
rect 4396 23071 4436 23080
rect 4492 23120 4532 23131
rect 4492 23045 4532 23080
rect 4588 23120 4628 23129
rect 4684 23120 4724 23920
rect 4780 23885 4820 24424
rect 4875 24128 4917 24137
rect 4875 24088 4876 24128
rect 4916 24088 4917 24128
rect 4875 24079 4917 24088
rect 4779 23876 4821 23885
rect 4779 23836 4780 23876
rect 4820 23836 4821 23876
rect 4779 23827 4821 23836
rect 4876 23792 4916 24079
rect 4972 23969 5012 24592
rect 5068 24464 5108 24473
rect 5260 24464 5300 24592
rect 5356 24632 5396 24643
rect 5356 24557 5396 24592
rect 5547 24632 5589 24641
rect 5547 24592 5548 24632
rect 5588 24592 5589 24632
rect 5644 24632 5684 25087
rect 5740 24632 5780 24641
rect 5644 24592 5740 24632
rect 5547 24583 5589 24592
rect 5740 24583 5780 24592
rect 5355 24548 5397 24557
rect 5355 24508 5356 24548
rect 5396 24508 5397 24548
rect 5355 24499 5397 24508
rect 5548 24498 5588 24583
rect 5836 24548 5876 25087
rect 5932 24800 5972 25255
rect 6219 25136 6261 25145
rect 6219 25096 6220 25136
rect 6260 25096 6261 25136
rect 6219 25087 6261 25096
rect 5932 24760 6068 24800
rect 5836 24499 5876 24508
rect 5932 24632 5972 24641
rect 5108 24424 5300 24464
rect 5068 24415 5108 24424
rect 5548 24380 5588 24389
rect 5932 24380 5972 24592
rect 5588 24340 5972 24380
rect 5548 24331 5588 24340
rect 5643 24044 5685 24053
rect 5643 24004 5644 24044
rect 5684 24004 5685 24044
rect 5643 23995 5685 24004
rect 4971 23960 5013 23969
rect 4971 23920 4972 23960
rect 5012 23920 5013 23960
rect 4971 23911 5013 23920
rect 4972 23792 5012 23801
rect 4876 23752 4972 23792
rect 4972 23743 5012 23752
rect 5068 23792 5108 23801
rect 5548 23792 5588 23801
rect 5108 23752 5396 23792
rect 5068 23743 5108 23752
rect 4779 23456 4821 23465
rect 4779 23416 4780 23456
rect 4820 23416 4821 23456
rect 4779 23407 4821 23416
rect 4928 23456 5296 23465
rect 4968 23416 5010 23456
rect 5050 23416 5092 23456
rect 5132 23416 5174 23456
rect 5214 23416 5256 23456
rect 4928 23407 5296 23416
rect 4628 23080 4724 23120
rect 4780 23120 4820 23407
rect 4876 23120 4916 23129
rect 4780 23080 4876 23120
rect 4588 23071 4628 23080
rect 4107 23036 4149 23045
rect 4107 22996 4108 23036
rect 4148 22996 4149 23036
rect 4107 22987 4149 22996
rect 4491 23036 4533 23045
rect 4491 22996 4492 23036
rect 4532 22996 4533 23036
rect 4491 22987 4533 22996
rect 4876 22877 4916 23080
rect 5356 23045 5396 23752
rect 5355 23036 5397 23045
rect 5355 22996 5356 23036
rect 5396 22996 5397 23036
rect 5355 22987 5397 22996
rect 4875 22868 4917 22877
rect 4012 22828 4820 22868
rect 3819 22819 3861 22828
rect 3688 22700 4056 22709
rect 3728 22660 3770 22700
rect 3810 22660 3852 22700
rect 3892 22660 3934 22700
rect 3974 22660 4016 22700
rect 3688 22651 4056 22660
rect 4299 22616 4341 22625
rect 4299 22576 4300 22616
rect 4340 22576 4341 22616
rect 4299 22567 4341 22576
rect 3532 22492 3668 22532
rect 3147 22448 3189 22457
rect 3147 22408 3148 22448
rect 3188 22408 3189 22448
rect 3147 22399 3189 22408
rect 3244 22408 3572 22448
rect 2956 22231 2996 22240
rect 3052 22364 3092 22373
rect 2667 22112 2709 22121
rect 2667 22072 2668 22112
rect 2708 22072 2709 22112
rect 2667 22063 2709 22072
rect 2859 22112 2901 22121
rect 2859 22072 2860 22112
rect 2900 22072 2901 22112
rect 2859 22063 2901 22072
rect 2571 21944 2613 21953
rect 2571 21904 2572 21944
rect 2612 21904 2613 21944
rect 2571 21895 2613 21904
rect 2668 21617 2708 22063
rect 3052 21944 3092 22324
rect 3148 22314 3188 22399
rect 3244 22364 3284 22408
rect 2956 21904 3092 21944
rect 2667 21608 2709 21617
rect 2667 21568 2668 21608
rect 2708 21568 2709 21608
rect 2667 21559 2709 21568
rect 2860 21608 2900 21619
rect 2860 21533 2900 21568
rect 2475 21524 2517 21533
rect 2475 21484 2476 21524
rect 2516 21484 2517 21524
rect 2475 21475 2517 21484
rect 2859 21524 2901 21533
rect 2859 21484 2860 21524
rect 2900 21484 2901 21524
rect 2859 21475 2901 21484
rect 2476 20768 2516 21475
rect 2571 21188 2613 21197
rect 2571 21148 2572 21188
rect 2612 21148 2613 21188
rect 2571 21139 2613 21148
rect 2476 20719 2516 20728
rect 2572 20441 2612 21139
rect 2956 21029 2996 21904
rect 3052 21776 3092 21785
rect 3244 21776 3284 22324
rect 3340 22280 3380 22289
rect 3340 21869 3380 22240
rect 3532 22280 3572 22408
rect 3532 22231 3572 22240
rect 3628 22280 3668 22492
rect 3435 21944 3477 21953
rect 3435 21904 3436 21944
rect 3476 21904 3477 21944
rect 3435 21895 3477 21904
rect 3339 21860 3381 21869
rect 3339 21820 3340 21860
rect 3380 21820 3381 21860
rect 3339 21811 3381 21820
rect 3092 21736 3284 21776
rect 3052 21727 3092 21736
rect 3051 21608 3093 21617
rect 3051 21568 3052 21608
rect 3092 21568 3093 21608
rect 3051 21559 3093 21568
rect 2955 21020 2997 21029
rect 2955 20980 2956 21020
rect 2996 20980 2997 21020
rect 2955 20971 2997 20980
rect 2859 20936 2901 20945
rect 2859 20896 2860 20936
rect 2900 20896 2901 20936
rect 2859 20887 2901 20896
rect 2860 20802 2900 20887
rect 2667 20684 2709 20693
rect 2667 20644 2668 20684
rect 2708 20644 2709 20684
rect 2667 20635 2709 20644
rect 2668 20550 2708 20635
rect 3052 20441 3092 21559
rect 3339 21524 3381 21533
rect 3339 21484 3340 21524
rect 3380 21484 3381 21524
rect 3339 21475 3381 21484
rect 3147 21440 3189 21449
rect 3147 21400 3148 21440
rect 3188 21400 3189 21440
rect 3147 21391 3189 21400
rect 3148 20936 3188 21391
rect 3340 21390 3380 21475
rect 2571 20432 2613 20441
rect 2571 20392 2572 20432
rect 2612 20392 2613 20432
rect 2571 20383 2613 20392
rect 3051 20432 3093 20441
rect 3051 20392 3052 20432
rect 3092 20392 3093 20432
rect 3051 20383 3093 20392
rect 2955 20264 2997 20273
rect 2955 20224 2956 20264
rect 2996 20224 2997 20264
rect 2955 20215 2997 20224
rect 2956 20105 2996 20215
rect 2475 20096 2517 20105
rect 2475 20056 2476 20096
rect 2516 20056 2517 20096
rect 2475 20047 2517 20056
rect 2860 20096 2900 20105
rect 2476 19265 2516 20047
rect 2668 19844 2708 19853
rect 2860 19844 2900 20056
rect 2955 20096 2997 20105
rect 2955 20056 2956 20096
rect 2996 20056 2997 20096
rect 2955 20047 2997 20056
rect 2708 19804 2900 19844
rect 2668 19795 2708 19804
rect 2667 19508 2709 19517
rect 2667 19468 2668 19508
rect 2708 19468 2709 19508
rect 2667 19459 2709 19468
rect 2475 19256 2517 19265
rect 2475 19216 2476 19256
rect 2516 19216 2517 19256
rect 2475 19207 2517 19216
rect 2476 18584 2516 19207
rect 2668 18752 2708 19459
rect 2763 19424 2805 19433
rect 2763 19384 2764 19424
rect 2804 19384 2805 19424
rect 2763 19375 2805 19384
rect 2476 18535 2516 18544
rect 2572 18712 2708 18752
rect 2475 17828 2517 17837
rect 2475 17788 2476 17828
rect 2516 17788 2517 17828
rect 2475 17779 2517 17788
rect 2476 17669 2516 17779
rect 2475 17660 2517 17669
rect 2475 17620 2476 17660
rect 2516 17620 2517 17660
rect 2475 17611 2517 17620
rect 2380 16435 2420 16444
rect 2092 16183 2132 16192
rect 1708 15940 1940 15980
rect 1995 15980 2037 15989
rect 1995 15940 1996 15980
rect 2036 15940 2037 15980
rect 1995 15931 2037 15940
rect 1515 15896 1557 15905
rect 1515 15856 1516 15896
rect 1556 15856 1557 15896
rect 1515 15847 1557 15856
rect 1515 15560 1557 15569
rect 1515 15520 1516 15560
rect 1556 15520 1557 15560
rect 1515 15511 1557 15520
rect 1227 14972 1269 14981
rect 1227 14932 1228 14972
rect 1268 14932 1269 14972
rect 1227 14923 1269 14932
rect 1228 14729 1268 14814
rect 1227 14720 1269 14729
rect 1227 14680 1228 14720
rect 1268 14680 1269 14720
rect 1227 14671 1269 14680
rect 1227 14552 1269 14561
rect 1227 14512 1228 14552
rect 1268 14512 1269 14552
rect 1227 14503 1269 14512
rect 1228 14216 1268 14503
rect 1228 14167 1268 14176
rect 1227 14048 1269 14057
rect 1227 14008 1228 14048
rect 1268 14008 1269 14048
rect 1227 13999 1269 14008
rect 1228 13460 1268 13999
rect 1228 13411 1268 13420
rect 1324 13124 1364 15352
rect 1516 15392 1556 15511
rect 1707 15476 1749 15485
rect 1707 15436 1708 15476
rect 1748 15436 1749 15476
rect 1707 15427 1749 15436
rect 2092 15476 2132 15485
rect 2188 15476 2228 16435
rect 2572 16274 2612 18712
rect 2667 18584 2709 18593
rect 2667 18544 2668 18584
rect 2708 18544 2709 18584
rect 2667 18535 2709 18544
rect 2668 18332 2708 18535
rect 2668 17753 2708 18292
rect 2667 17744 2709 17753
rect 2667 17704 2668 17744
rect 2708 17704 2709 17744
rect 2667 17695 2709 17704
rect 2764 17744 2804 19375
rect 2860 19181 2900 19804
rect 2956 19844 2996 19853
rect 2956 19517 2996 19804
rect 2955 19508 2997 19517
rect 2955 19468 2956 19508
rect 2996 19468 2997 19508
rect 2955 19459 2997 19468
rect 2955 19256 2997 19265
rect 2955 19216 2956 19256
rect 2996 19216 2997 19256
rect 2955 19207 2997 19216
rect 2859 19172 2901 19181
rect 2859 19132 2860 19172
rect 2900 19132 2901 19172
rect 2859 19123 2901 19132
rect 2956 19122 2996 19207
rect 2956 18584 2996 18593
rect 3052 18584 3092 20383
rect 3148 19685 3188 20896
rect 3243 20852 3285 20861
rect 3243 20812 3244 20852
rect 3284 20812 3285 20852
rect 3243 20803 3285 20812
rect 3147 19676 3189 19685
rect 3147 19636 3148 19676
rect 3188 19636 3189 19676
rect 3147 19627 3189 19636
rect 3147 19172 3189 19181
rect 3147 19132 3148 19172
rect 3188 19132 3189 19172
rect 3147 19123 3189 19132
rect 3148 19038 3188 19123
rect 3244 18752 3284 20803
rect 3339 20432 3381 20441
rect 3339 20392 3340 20432
rect 3380 20392 3381 20432
rect 3339 20383 3381 20392
rect 3340 20096 3380 20383
rect 3436 20273 3476 21895
rect 3628 21776 3668 22240
rect 3820 22280 3860 22289
rect 3724 22112 3764 22121
rect 3724 21869 3764 22072
rect 3723 21860 3765 21869
rect 3723 21820 3724 21860
rect 3764 21820 3765 21860
rect 3723 21811 3765 21820
rect 3628 21727 3668 21736
rect 3820 21449 3860 22240
rect 3916 22280 3956 22289
rect 3916 21785 3956 22240
rect 4071 22280 4111 22289
rect 4300 22280 4340 22567
rect 4491 22448 4533 22457
rect 4491 22408 4492 22448
rect 4532 22408 4533 22448
rect 4491 22399 4533 22408
rect 4395 22364 4437 22373
rect 4395 22324 4396 22364
rect 4436 22324 4437 22364
rect 4395 22315 4437 22324
rect 4111 22240 4148 22280
rect 4071 22231 4148 22240
rect 3915 21776 3957 21785
rect 3915 21736 3916 21776
rect 3956 21736 3957 21776
rect 3915 21727 3957 21736
rect 3915 21524 3957 21533
rect 3915 21484 3916 21524
rect 3956 21484 3957 21524
rect 3915 21475 3957 21484
rect 3532 21440 3572 21449
rect 3532 20936 3572 21400
rect 3819 21440 3861 21449
rect 3819 21400 3820 21440
rect 3860 21400 3861 21440
rect 3819 21391 3861 21400
rect 3916 21390 3956 21475
rect 4108 21356 4148 22231
rect 4300 21869 4340 22240
rect 4396 22230 4436 22315
rect 4492 22314 4532 22399
rect 4588 22364 4628 22373
rect 4299 21860 4341 21869
rect 4299 21820 4300 21860
rect 4340 21820 4341 21860
rect 4299 21811 4341 21820
rect 4395 21776 4437 21785
rect 4395 21736 4396 21776
rect 4436 21736 4437 21776
rect 4588 21776 4628 22324
rect 4683 22280 4725 22289
rect 4683 22240 4684 22280
rect 4724 22240 4725 22280
rect 4683 22231 4725 22240
rect 4684 22146 4724 22231
rect 4588 21736 4724 21776
rect 4395 21727 4437 21736
rect 4203 21608 4245 21617
rect 4203 21568 4204 21608
rect 4244 21568 4245 21608
rect 4203 21559 4245 21568
rect 4396 21608 4436 21727
rect 4396 21559 4436 21568
rect 4587 21608 4629 21617
rect 4587 21568 4588 21608
rect 4628 21568 4629 21608
rect 4587 21559 4629 21568
rect 4204 21474 4244 21559
rect 4588 21474 4628 21559
rect 4395 21440 4437 21449
rect 4395 21400 4396 21440
rect 4436 21400 4437 21440
rect 4395 21391 4437 21400
rect 4108 21316 4340 21356
rect 3688 21188 4056 21197
rect 3728 21148 3770 21188
rect 3810 21148 3852 21188
rect 3892 21148 3934 21188
rect 3974 21148 4016 21188
rect 3688 21139 4056 21148
rect 3532 20861 3572 20896
rect 4011 20936 4053 20945
rect 4011 20896 4012 20936
rect 4052 20896 4053 20936
rect 4011 20887 4053 20896
rect 3531 20852 3573 20861
rect 3531 20812 3532 20852
rect 3572 20812 3573 20852
rect 3531 20803 3573 20812
rect 3916 20852 3956 20861
rect 3532 20772 3572 20803
rect 3820 20768 3860 20777
rect 3820 20609 3860 20728
rect 3819 20600 3861 20609
rect 3819 20560 3820 20600
rect 3860 20560 3861 20600
rect 3819 20551 3861 20560
rect 3435 20264 3477 20273
rect 3435 20224 3436 20264
rect 3476 20224 3477 20264
rect 3435 20215 3477 20224
rect 3627 20264 3669 20273
rect 3627 20224 3628 20264
rect 3668 20224 3764 20264
rect 3627 20215 3669 20224
rect 3724 20180 3764 20224
rect 3724 20131 3764 20140
rect 3340 20045 3380 20056
rect 3531 20096 3573 20105
rect 3531 20056 3532 20096
rect 3572 20056 3573 20096
rect 3531 20047 3573 20056
rect 3628 20096 3668 20105
rect 3435 19760 3477 19769
rect 3435 19720 3436 19760
rect 3476 19720 3477 19760
rect 3435 19711 3477 19720
rect 3436 19433 3476 19711
rect 3435 19424 3477 19433
rect 3435 19384 3436 19424
rect 3476 19384 3477 19424
rect 3435 19375 3477 19384
rect 3340 19256 3380 19265
rect 3340 19097 3380 19216
rect 3435 19256 3477 19265
rect 3435 19216 3436 19256
rect 3476 19216 3477 19256
rect 3435 19207 3477 19216
rect 3436 19122 3476 19207
rect 3339 19088 3381 19097
rect 3339 19048 3340 19088
rect 3380 19048 3381 19088
rect 3339 19039 3381 19048
rect 2996 18544 3092 18584
rect 3148 18712 3284 18752
rect 2956 18535 2996 18544
rect 3148 18164 3188 18712
rect 3339 18668 3381 18677
rect 3339 18628 3340 18668
rect 3380 18628 3381 18668
rect 3339 18619 3381 18628
rect 3244 18584 3284 18593
rect 3244 18341 3284 18544
rect 3340 18534 3380 18619
rect 3243 18332 3285 18341
rect 3243 18292 3244 18332
rect 3284 18292 3285 18332
rect 3243 18283 3285 18292
rect 3148 18124 3380 18164
rect 3243 17744 3285 17753
rect 2804 17704 3092 17744
rect 2764 17695 2804 17704
rect 2956 17576 2996 17585
rect 2956 17081 2996 17536
rect 2955 17072 2997 17081
rect 2955 17032 2956 17072
rect 2996 17032 2997 17072
rect 2955 17023 2997 17032
rect 3052 17072 3092 17704
rect 3243 17704 3244 17744
rect 3284 17704 3285 17744
rect 3243 17695 3285 17704
rect 3244 17610 3284 17695
rect 2763 16820 2805 16829
rect 2763 16780 2764 16820
rect 2804 16780 2805 16820
rect 2763 16771 2805 16780
rect 2572 16234 2708 16274
rect 2571 16064 2613 16073
rect 2571 16024 2572 16064
rect 2612 16024 2613 16064
rect 2571 16015 2613 16024
rect 2572 15930 2612 16015
rect 2132 15436 2228 15476
rect 2284 15560 2324 15569
rect 2092 15427 2132 15436
rect 1516 15343 1556 15352
rect 1708 15342 1748 15427
rect 1900 15308 1940 15317
rect 1900 14561 1940 15268
rect 1995 14888 2037 14897
rect 1995 14848 1996 14888
rect 2036 14848 2037 14888
rect 1995 14839 2037 14848
rect 1899 14552 1941 14561
rect 1899 14512 1900 14552
rect 1940 14512 1941 14552
rect 1899 14503 1941 14512
rect 1707 14300 1749 14309
rect 1707 14260 1708 14300
rect 1748 14260 1749 14300
rect 1707 14251 1749 14260
rect 1708 14132 1748 14251
rect 1708 14083 1748 14092
rect 1612 14048 1652 14057
rect 1516 14008 1612 14048
rect 1419 13964 1461 13973
rect 1419 13924 1420 13964
rect 1460 13924 1461 13964
rect 1419 13915 1461 13924
rect 1420 13830 1460 13915
rect 1419 13712 1461 13721
rect 1419 13672 1420 13712
rect 1460 13672 1461 13712
rect 1419 13663 1461 13672
rect 1420 13292 1460 13663
rect 1420 13243 1460 13252
rect 1324 13084 1460 13124
rect 1228 12536 1268 12545
rect 1268 12496 1364 12536
rect 1228 12487 1268 12496
rect 1324 12041 1364 12496
rect 1323 12032 1365 12041
rect 1323 11992 1324 12032
rect 1364 11992 1365 12032
rect 1323 11983 1365 11992
rect 1228 11696 1268 11705
rect 1323 11696 1365 11705
rect 1268 11656 1324 11696
rect 1364 11656 1365 11696
rect 1228 11647 1268 11656
rect 1323 11647 1365 11656
rect 1323 11024 1365 11033
rect 1323 10984 1324 11024
rect 1364 10984 1365 11024
rect 1323 10975 1365 10984
rect 1324 10890 1364 10975
rect 1131 10856 1173 10865
rect 1131 10816 1132 10856
rect 1172 10816 1173 10856
rect 1131 10807 1173 10816
rect 1420 10772 1460 13084
rect 1516 11192 1556 14008
rect 1612 13999 1652 14008
rect 1803 14048 1845 14057
rect 1803 14008 1804 14048
rect 1844 14008 1845 14048
rect 1803 13999 1845 14008
rect 1900 14048 1940 14057
rect 1996 14048 2036 14839
rect 2284 14225 2324 15520
rect 2380 15560 2420 15569
rect 2380 14393 2420 15520
rect 2476 15560 2516 15569
rect 2476 14981 2516 15520
rect 2572 15560 2612 15569
rect 2475 14972 2517 14981
rect 2475 14932 2476 14972
rect 2516 14932 2517 14972
rect 2475 14923 2517 14932
rect 2475 14720 2517 14729
rect 2475 14680 2476 14720
rect 2516 14680 2517 14720
rect 2475 14671 2517 14680
rect 2476 14586 2516 14671
rect 2379 14384 2421 14393
rect 2379 14344 2380 14384
rect 2420 14344 2421 14384
rect 2379 14335 2421 14344
rect 2572 14300 2612 15520
rect 2668 15401 2708 16234
rect 2764 16246 2804 16771
rect 2764 16197 2804 16206
rect 3052 15569 3092 17032
rect 3243 16820 3285 16829
rect 3243 16780 3244 16820
rect 3284 16780 3285 16820
rect 3243 16771 3285 16780
rect 3244 16686 3284 16771
rect 3244 16232 3284 16241
rect 3244 15653 3284 16192
rect 3243 15644 3285 15653
rect 3243 15604 3244 15644
rect 3284 15604 3285 15644
rect 3243 15595 3285 15604
rect 2763 15560 2805 15569
rect 2763 15520 2764 15560
rect 2804 15520 2805 15560
rect 2763 15511 2805 15520
rect 3051 15560 3093 15569
rect 3051 15520 3052 15560
rect 3092 15520 3093 15560
rect 3051 15511 3093 15520
rect 2764 15426 2804 15511
rect 2667 15392 2709 15401
rect 2667 15352 2668 15392
rect 2708 15352 2709 15392
rect 2667 15343 2709 15352
rect 2667 14972 2709 14981
rect 3052 14972 3092 15511
rect 2667 14932 2668 14972
rect 2708 14932 2709 14972
rect 2667 14923 2709 14932
rect 2956 14932 3092 14972
rect 2668 14838 2708 14923
rect 2956 14729 2996 14932
rect 3051 14804 3093 14813
rect 3051 14764 3052 14804
rect 3092 14764 3093 14804
rect 3051 14755 3093 14764
rect 2955 14720 2997 14729
rect 2955 14680 2956 14720
rect 2996 14680 2997 14720
rect 2955 14671 2997 14680
rect 2476 14260 2612 14300
rect 2860 14552 2900 14561
rect 2283 14216 2325 14225
rect 2283 14176 2284 14216
rect 2324 14176 2325 14216
rect 2283 14167 2325 14176
rect 2092 14057 2132 14142
rect 1940 14008 2036 14048
rect 2091 14048 2133 14057
rect 2091 14008 2092 14048
rect 2132 14008 2133 14048
rect 2284 14040 2324 14167
rect 2380 14132 2420 14141
rect 1900 13999 1940 14008
rect 2091 13999 2133 14008
rect 2188 14006 2228 14015
rect 1707 13208 1749 13217
rect 1707 13168 1708 13208
rect 1748 13168 1749 13208
rect 1707 13159 1749 13168
rect 1708 13074 1748 13159
rect 1707 12620 1749 12629
rect 1707 12580 1708 12620
rect 1748 12580 1749 12620
rect 1707 12571 1749 12580
rect 1516 11143 1556 11152
rect 1611 11108 1653 11117
rect 1611 11068 1612 11108
rect 1652 11068 1653 11108
rect 1611 11059 1653 11068
rect 1612 11024 1652 11059
rect 1612 10973 1652 10984
rect 1708 10856 1748 12571
rect 1804 11117 1844 13999
rect 2177 13966 2188 14006
rect 2284 13991 2324 14000
rect 2373 14092 2380 14132
rect 2373 14083 2420 14092
rect 2373 14037 2413 14083
rect 2373 13997 2420 14037
rect 2177 13957 2228 13966
rect 2380 13964 2420 13997
rect 2177 13889 2217 13957
rect 2380 13924 2421 13964
rect 2177 13880 2229 13889
rect 2381 13880 2421 13924
rect 2177 13840 2188 13880
rect 2228 13840 2229 13880
rect 2187 13831 2229 13840
rect 2380 13840 2421 13880
rect 2380 13796 2420 13840
rect 2284 13756 2420 13796
rect 2476 13796 2516 14260
rect 2860 14141 2900 14512
rect 2572 14132 2612 14141
rect 2572 13973 2612 14092
rect 2859 14132 2901 14141
rect 2859 14092 2860 14132
rect 2900 14092 2901 14132
rect 2859 14083 2901 14092
rect 2764 14034 2804 14043
rect 2804 13994 2900 14006
rect 2571 13964 2613 13973
rect 2764 13966 2900 13994
rect 2571 13924 2572 13964
rect 2612 13924 2613 13964
rect 2571 13915 2613 13924
rect 2763 13880 2805 13889
rect 2763 13840 2764 13880
rect 2804 13840 2805 13880
rect 2763 13831 2805 13840
rect 2476 13756 2612 13796
rect 2284 12293 2324 13756
rect 2379 13628 2421 13637
rect 2379 13588 2380 13628
rect 2420 13588 2421 13628
rect 2379 13579 2421 13588
rect 2283 12284 2325 12293
rect 2283 12244 2284 12284
rect 2324 12244 2325 12284
rect 2283 12235 2325 12244
rect 2091 12200 2133 12209
rect 2091 12160 2092 12200
rect 2132 12160 2133 12200
rect 2091 12151 2133 12160
rect 1899 11528 1941 11537
rect 1899 11488 1900 11528
rect 1940 11488 1941 11528
rect 1899 11479 1941 11488
rect 1803 11108 1845 11117
rect 1803 11068 1804 11108
rect 1844 11068 1845 11108
rect 1803 11059 1845 11068
rect 1324 10732 1460 10772
rect 1516 10816 1748 10856
rect 1227 9512 1269 9521
rect 1227 9472 1228 9512
rect 1268 9472 1269 9512
rect 1227 9463 1269 9472
rect 1228 9378 1268 9463
rect 1324 9008 1364 10732
rect 1419 10184 1461 10193
rect 1419 10144 1420 10184
rect 1460 10144 1461 10184
rect 1419 10135 1461 10144
rect 1420 10050 1460 10135
rect 1420 9512 1460 9521
rect 1516 9512 1556 10816
rect 1804 10772 1844 10781
rect 1611 9764 1653 9773
rect 1611 9724 1612 9764
rect 1652 9724 1653 9764
rect 1611 9715 1653 9724
rect 1460 9472 1556 9512
rect 1612 9512 1652 9715
rect 1420 9463 1460 9472
rect 1612 9463 1652 9472
rect 1611 9344 1653 9353
rect 1611 9304 1612 9344
rect 1652 9304 1653 9344
rect 1611 9295 1653 9304
rect 1419 9260 1461 9269
rect 1419 9220 1420 9260
rect 1460 9220 1461 9260
rect 1419 9211 1461 9220
rect 1420 9126 1460 9211
rect 1324 8968 1556 9008
rect 1227 8840 1269 8849
rect 1330 8840 1372 8849
rect 1227 8800 1228 8840
rect 1268 8800 1269 8840
rect 1227 8791 1269 8800
rect 1324 8800 1331 8840
rect 1371 8800 1372 8840
rect 1324 8791 1372 8800
rect 1228 8706 1268 8791
rect 1228 8168 1268 8177
rect 1036 8128 1228 8168
rect 1228 8119 1268 8128
rect 940 7960 1268 8000
rect 844 7120 1172 7160
rect 843 6992 885 7001
rect 843 6952 844 6992
rect 884 6952 885 6992
rect 843 6943 885 6952
rect 651 6488 693 6497
rect 651 6448 652 6488
rect 692 6448 693 6488
rect 651 6439 693 6448
rect 651 6236 693 6245
rect 651 6196 652 6236
rect 692 6196 693 6236
rect 651 6187 693 6196
rect 555 2540 597 2549
rect 555 2500 556 2540
rect 596 2500 597 2540
rect 555 2491 597 2500
rect 267 944 309 953
rect 172 904 268 944
rect 308 904 309 944
rect 267 895 309 904
rect 652 449 692 6187
rect 747 2540 789 2549
rect 747 2500 748 2540
rect 788 2500 789 2540
rect 747 2491 789 2500
rect 748 2129 788 2491
rect 747 2120 789 2129
rect 747 2080 748 2120
rect 788 2080 789 2120
rect 747 2071 789 2080
rect 844 1877 884 6943
rect 1035 5396 1077 5405
rect 1035 5356 1036 5396
rect 1076 5356 1077 5396
rect 1035 5347 1077 5356
rect 843 1868 885 1877
rect 843 1828 844 1868
rect 884 1828 885 1868
rect 843 1819 885 1828
rect 651 440 693 449
rect 651 400 652 440
rect 692 400 693 440
rect 651 391 693 400
rect 1036 365 1076 5347
rect 1132 4808 1172 7120
rect 1228 6656 1268 7960
rect 1324 7916 1364 8791
rect 1419 8756 1461 8765
rect 1419 8716 1420 8756
rect 1460 8716 1461 8756
rect 1419 8707 1461 8716
rect 1420 8622 1460 8707
rect 1516 8672 1556 8968
rect 1612 8840 1652 9295
rect 1804 9101 1844 10732
rect 1900 9353 1940 11479
rect 1995 10940 2037 10949
rect 1995 10900 1996 10940
rect 2036 10900 2037 10940
rect 1995 10891 2037 10900
rect 1996 10806 2036 10891
rect 1995 9848 2037 9857
rect 1995 9808 1996 9848
rect 2036 9808 2037 9848
rect 1995 9799 2037 9808
rect 1899 9344 1941 9353
rect 1899 9304 1900 9344
rect 1940 9304 1941 9344
rect 1899 9295 1941 9304
rect 1803 9092 1845 9101
rect 1803 9052 1804 9092
rect 1844 9052 1845 9092
rect 1803 9043 1845 9052
rect 1996 9008 2036 9799
rect 2092 9008 2132 12151
rect 2188 11024 2228 11033
rect 2188 10445 2228 10984
rect 2187 10436 2229 10445
rect 2187 10396 2188 10436
rect 2228 10396 2229 10436
rect 2187 10387 2229 10396
rect 2187 10268 2229 10277
rect 2187 10228 2188 10268
rect 2228 10228 2229 10268
rect 2187 10219 2229 10228
rect 1612 8791 1652 8800
rect 1900 8968 2036 9008
rect 2082 8968 2132 9008
rect 1803 8756 1845 8765
rect 1803 8716 1804 8756
rect 1844 8716 1845 8756
rect 1803 8707 1845 8716
rect 1516 8632 1748 8672
rect 1515 8504 1557 8513
rect 1515 8464 1516 8504
rect 1556 8464 1557 8504
rect 1515 8455 1557 8464
rect 1420 7916 1460 7925
rect 1324 7876 1420 7916
rect 1420 7867 1460 7876
rect 1419 7496 1461 7505
rect 1419 7456 1420 7496
rect 1460 7456 1461 7496
rect 1419 7447 1461 7456
rect 1324 7169 1364 7254
rect 1323 7160 1365 7169
rect 1323 7120 1324 7160
rect 1364 7120 1365 7160
rect 1323 7111 1365 7120
rect 1323 6992 1365 7001
rect 1323 6952 1324 6992
rect 1364 6952 1365 6992
rect 1323 6943 1365 6952
rect 1228 6607 1268 6616
rect 1227 5648 1269 5657
rect 1227 5608 1228 5648
rect 1268 5608 1269 5648
rect 1227 5599 1269 5608
rect 1228 5514 1268 5599
rect 1228 4808 1268 4817
rect 1132 4768 1228 4808
rect 1228 4759 1268 4768
rect 1324 4304 1364 6943
rect 1420 6404 1460 7447
rect 1516 6656 1556 8455
rect 1611 8000 1653 8009
rect 1611 7960 1612 8000
rect 1652 7960 1653 8000
rect 1611 7951 1653 7960
rect 1612 7866 1652 7951
rect 1612 6656 1652 6665
rect 1516 6616 1612 6656
rect 1612 6607 1652 6616
rect 1515 6488 1557 6497
rect 1708 6488 1748 8632
rect 1804 8622 1844 8707
rect 1900 7001 1940 8968
rect 2082 8924 2122 8968
rect 1996 8884 2122 8924
rect 1996 8840 2036 8884
rect 2188 8840 2228 10219
rect 2283 9932 2325 9941
rect 2283 9892 2284 9932
rect 2324 9892 2325 9932
rect 2283 9883 2325 9892
rect 2284 8849 2324 9883
rect 2380 9857 2420 13579
rect 2476 12536 2516 12576
rect 2476 12461 2516 12496
rect 2475 12452 2517 12461
rect 2475 12412 2476 12452
rect 2516 12412 2517 12452
rect 2475 12403 2517 12412
rect 2476 11696 2516 12403
rect 2476 11453 2516 11656
rect 2475 11444 2517 11453
rect 2475 11404 2476 11444
rect 2516 11404 2517 11444
rect 2475 11395 2517 11404
rect 2475 11024 2517 11033
rect 2475 10984 2476 11024
rect 2516 10984 2517 11024
rect 2475 10975 2517 10984
rect 2379 9848 2421 9857
rect 2379 9808 2380 9848
rect 2420 9808 2421 9848
rect 2379 9799 2421 9808
rect 2380 9521 2420 9799
rect 2379 9512 2421 9521
rect 2379 9472 2380 9512
rect 2420 9472 2421 9512
rect 2379 9463 2421 9472
rect 1996 8791 2036 8800
rect 2103 8800 2228 8840
rect 2283 8840 2325 8849
rect 2476 8840 2516 10975
rect 2572 10193 2612 13756
rect 2667 13376 2709 13385
rect 2667 13336 2668 13376
rect 2708 13336 2709 13376
rect 2667 13327 2709 13336
rect 2668 12704 2708 13327
rect 2668 12655 2708 12664
rect 2668 11948 2708 11957
rect 2764 11948 2804 13831
rect 2860 13385 2900 13966
rect 2859 13376 2901 13385
rect 2859 13336 2860 13376
rect 2900 13336 2901 13376
rect 2859 13327 2901 13336
rect 2956 13208 2996 14671
rect 3052 14670 3092 14755
rect 3147 14552 3189 14561
rect 3147 14512 3148 14552
rect 3188 14512 3189 14552
rect 3147 14503 3189 14512
rect 3051 14216 3093 14225
rect 3051 14176 3052 14216
rect 3092 14176 3093 14216
rect 3051 14167 3093 14176
rect 2956 13133 2996 13168
rect 2955 13124 2997 13133
rect 2955 13084 2956 13124
rect 2996 13084 2997 13124
rect 2955 13075 2997 13084
rect 2956 13044 2996 13075
rect 2859 12620 2901 12629
rect 2859 12580 2860 12620
rect 2900 12580 2901 12620
rect 2859 12571 2901 12580
rect 2860 12486 2900 12571
rect 3052 12522 3092 14167
rect 3148 13460 3188 14503
rect 3244 14048 3284 14057
rect 3244 13805 3284 14008
rect 3243 13796 3285 13805
rect 3243 13756 3244 13796
rect 3284 13756 3285 13796
rect 3243 13747 3285 13756
rect 3243 13628 3285 13637
rect 3243 13588 3244 13628
rect 3284 13588 3285 13628
rect 3243 13579 3285 13588
rect 3148 13411 3188 13420
rect 3244 12788 3284 13579
rect 3340 13469 3380 18124
rect 3435 17996 3477 18005
rect 3435 17956 3436 17996
rect 3476 17956 3477 17996
rect 3532 17996 3572 20047
rect 3628 19853 3668 20056
rect 3916 19937 3956 20812
rect 4012 20802 4052 20887
rect 4108 20852 4148 20861
rect 4108 20441 4148 20812
rect 4203 20768 4245 20777
rect 4203 20728 4204 20768
rect 4244 20728 4245 20768
rect 4203 20719 4245 20728
rect 4204 20634 4244 20719
rect 4107 20432 4149 20441
rect 4107 20392 4108 20432
rect 4148 20392 4149 20432
rect 4107 20383 4149 20392
rect 4300 20264 4340 21316
rect 4396 20945 4436 21391
rect 4684 21356 4724 21736
rect 4588 21316 4724 21356
rect 4395 20936 4437 20945
rect 4395 20896 4396 20936
rect 4436 20896 4437 20936
rect 4395 20887 4437 20896
rect 4396 20768 4436 20779
rect 4396 20693 4436 20728
rect 4395 20684 4437 20693
rect 4395 20644 4396 20684
rect 4436 20644 4437 20684
rect 4395 20635 4437 20644
rect 4492 20600 4532 20609
rect 4405 20432 4447 20441
rect 4492 20432 4532 20560
rect 4405 20392 4406 20432
rect 4446 20392 4532 20432
rect 4588 20432 4628 21316
rect 4684 20777 4724 20862
rect 4683 20768 4725 20777
rect 4683 20728 4684 20768
rect 4724 20728 4725 20768
rect 4683 20719 4725 20728
rect 4780 20693 4820 22828
rect 4875 22828 4876 22868
rect 4916 22828 4917 22868
rect 4875 22819 4917 22828
rect 5356 22793 5396 22987
rect 5355 22784 5397 22793
rect 5355 22744 5356 22784
rect 5396 22744 5397 22784
rect 5355 22735 5397 22744
rect 4875 22616 4917 22625
rect 4875 22576 4876 22616
rect 4916 22576 4917 22616
rect 4875 22567 4917 22576
rect 4876 22448 4916 22567
rect 4876 22399 4916 22408
rect 5452 22373 5492 22458
rect 5451 22364 5493 22373
rect 5451 22324 5452 22364
rect 5492 22324 5493 22364
rect 5451 22315 5493 22324
rect 5260 22112 5300 22121
rect 5300 22072 5396 22112
rect 5260 22063 5300 22072
rect 4928 21944 5296 21953
rect 4968 21904 5010 21944
rect 5050 21904 5092 21944
rect 5132 21904 5174 21944
rect 5214 21904 5256 21944
rect 4928 21895 5296 21904
rect 5356 21449 5396 22072
rect 5355 21440 5397 21449
rect 5355 21400 5356 21440
rect 5396 21400 5397 21440
rect 5355 21391 5397 21400
rect 4875 21104 4917 21113
rect 4875 21064 4876 21104
rect 4916 21064 4917 21104
rect 4875 21055 4917 21064
rect 4779 20684 4821 20693
rect 4779 20644 4780 20684
rect 4820 20644 4821 20684
rect 4779 20635 4821 20644
rect 4876 20609 4916 21055
rect 5355 20768 5397 20777
rect 5355 20728 5356 20768
rect 5396 20728 5397 20768
rect 5355 20719 5397 20728
rect 4683 20600 4725 20609
rect 4683 20560 4684 20600
rect 4724 20560 4725 20600
rect 4683 20551 4725 20560
rect 4875 20600 4917 20609
rect 4875 20560 4876 20600
rect 4916 20560 4917 20600
rect 4875 20551 4917 20560
rect 4588 20392 4629 20432
rect 4405 20383 4447 20392
rect 4589 20348 4629 20392
rect 4588 20308 4629 20348
rect 4588 20264 4628 20308
rect 4012 20224 4340 20264
rect 4492 20224 4628 20264
rect 3915 19928 3957 19937
rect 3915 19888 3916 19928
rect 3956 19888 3957 19928
rect 3915 19879 3957 19888
rect 4012 19928 4052 20224
rect 4395 20012 4437 20021
rect 4395 19972 4396 20012
rect 4436 19972 4437 20012
rect 4395 19963 4437 19972
rect 4012 19879 4052 19888
rect 4107 19928 4149 19937
rect 4107 19888 4108 19928
rect 4148 19888 4149 19928
rect 4107 19879 4149 19888
rect 3627 19844 3669 19853
rect 3627 19804 3628 19844
rect 3668 19804 3669 19844
rect 3627 19795 3669 19804
rect 3688 19676 4056 19685
rect 3728 19636 3770 19676
rect 3810 19636 3852 19676
rect 3892 19636 3934 19676
rect 3974 19636 4016 19676
rect 3688 19627 4056 19636
rect 3628 19433 3668 19518
rect 4011 19508 4053 19517
rect 4011 19468 4012 19508
rect 4052 19468 4053 19508
rect 4011 19459 4053 19468
rect 3627 19424 3669 19433
rect 3627 19384 3628 19424
rect 3668 19384 3669 19424
rect 3627 19375 3669 19384
rect 3628 19256 3668 19265
rect 3628 18593 3668 19216
rect 3819 19256 3861 19265
rect 3819 19216 3820 19256
rect 3860 19216 3861 19256
rect 3819 19207 3861 19216
rect 3820 19122 3860 19207
rect 3915 18752 3957 18761
rect 3915 18712 3916 18752
rect 3956 18712 3957 18752
rect 3915 18703 3957 18712
rect 3916 18618 3956 18703
rect 3627 18584 3669 18593
rect 3627 18544 3628 18584
rect 3668 18544 3669 18584
rect 3627 18535 3669 18544
rect 3819 18584 3861 18593
rect 3819 18544 3820 18584
rect 3860 18544 3861 18584
rect 3819 18535 3861 18544
rect 4012 18584 4052 19459
rect 3820 18450 3860 18535
rect 3627 18416 3669 18425
rect 3627 18376 3628 18416
rect 3668 18376 3669 18416
rect 3627 18367 3669 18376
rect 3628 18282 3668 18367
rect 4012 18341 4052 18544
rect 4108 18425 4148 19879
rect 4396 19878 4436 19963
rect 4203 19844 4245 19853
rect 4203 19804 4204 19844
rect 4244 19804 4245 19844
rect 4203 19795 4245 19804
rect 4204 19710 4244 19795
rect 4492 19517 4532 20224
rect 4684 20180 4724 20551
rect 4928 20432 5296 20441
rect 4968 20392 5010 20432
rect 5050 20392 5092 20432
rect 5132 20392 5174 20432
rect 5214 20392 5256 20432
rect 4928 20383 5296 20392
rect 4588 20140 4724 20180
rect 4588 20096 4628 20140
rect 4588 20047 4628 20056
rect 4491 19508 4533 19517
rect 4491 19468 4492 19508
rect 4532 19468 4533 19508
rect 4491 19459 4533 19468
rect 5259 19508 5301 19517
rect 5259 19468 5260 19508
rect 5300 19468 5301 19508
rect 5259 19459 5301 19468
rect 5260 19374 5300 19459
rect 5068 19256 5108 19265
rect 5356 19256 5396 20719
rect 5548 20273 5588 23752
rect 5547 20264 5589 20273
rect 5547 20224 5548 20264
rect 5588 20224 5589 20264
rect 5547 20215 5589 20224
rect 5644 20180 5684 23995
rect 6028 23960 6068 24760
rect 5932 23920 6068 23960
rect 5739 22196 5781 22205
rect 5739 22156 5740 22196
rect 5780 22156 5781 22196
rect 5739 22147 5781 22156
rect 5740 22062 5780 22147
rect 5835 22112 5877 22121
rect 5835 22072 5836 22112
rect 5876 22072 5877 22112
rect 5835 22063 5877 22072
rect 5836 21608 5876 22063
rect 5836 20777 5876 21568
rect 5932 21524 5972 23920
rect 6076 23801 6116 23810
rect 6116 23761 6164 23792
rect 6076 23752 6164 23761
rect 6124 23288 6164 23752
rect 6220 23624 6260 25087
rect 6316 24800 6356 26104
rect 6412 26144 6452 26263
rect 6412 25052 6452 26104
rect 6508 25817 6548 26431
rect 6604 26405 6644 27775
rect 6700 27068 6740 28288
rect 6795 28288 6796 28328
rect 6836 28288 6837 28328
rect 6795 28279 6837 28288
rect 6892 28328 6932 28339
rect 6892 28253 6932 28288
rect 6891 28244 6933 28253
rect 6891 28204 6892 28244
rect 6932 28204 6933 28244
rect 6891 28195 6933 28204
rect 7084 27161 7124 29548
rect 7275 28412 7317 28421
rect 7275 28372 7276 28412
rect 7316 28372 7317 28412
rect 7275 28363 7317 28372
rect 7276 27488 7316 28363
rect 7372 28328 7412 29968
rect 7564 29840 7604 29849
rect 7564 28925 7604 29800
rect 7659 29840 7701 29849
rect 7659 29800 7660 29840
rect 7700 29800 7701 29840
rect 7659 29791 7701 29800
rect 7563 28916 7605 28925
rect 7563 28876 7564 28916
rect 7604 28876 7605 28916
rect 7563 28867 7605 28876
rect 7372 28288 7508 28328
rect 7371 27740 7413 27749
rect 7371 27700 7372 27740
rect 7412 27700 7413 27740
rect 7371 27691 7413 27700
rect 7372 27656 7412 27691
rect 7468 27665 7508 28288
rect 7563 27740 7605 27749
rect 7563 27700 7564 27740
rect 7604 27700 7605 27740
rect 7563 27691 7605 27700
rect 7372 27605 7412 27616
rect 7467 27656 7509 27665
rect 7467 27616 7468 27656
rect 7508 27616 7509 27656
rect 7467 27607 7509 27616
rect 7276 27448 7508 27488
rect 7083 27152 7125 27161
rect 7083 27112 7084 27152
rect 7124 27112 7125 27152
rect 7083 27103 7125 27112
rect 7179 27068 7221 27077
rect 6700 27028 7028 27068
rect 6795 26816 6837 26825
rect 6795 26776 6796 26816
rect 6836 26776 6837 26816
rect 6795 26767 6837 26776
rect 6892 26816 6932 26825
rect 6796 26682 6836 26767
rect 6603 26396 6645 26405
rect 6603 26356 6604 26396
rect 6644 26356 6645 26396
rect 6603 26347 6645 26356
rect 6892 26321 6932 26776
rect 6891 26312 6933 26321
rect 6891 26272 6892 26312
rect 6932 26272 6933 26312
rect 6891 26263 6933 26272
rect 6988 26312 7028 27028
rect 7179 27028 7180 27068
rect 7220 27028 7221 27068
rect 7179 27019 7221 27028
rect 7180 26830 7220 27019
rect 7276 26909 7316 26911
rect 7275 26900 7317 26909
rect 7275 26860 7276 26900
rect 7316 26860 7317 26900
rect 7275 26851 7317 26860
rect 6988 26263 7028 26272
rect 7084 26790 7220 26830
rect 7276 26816 7316 26851
rect 7372 26816 7412 26825
rect 6603 26144 6645 26153
rect 6603 26104 6604 26144
rect 6644 26104 6645 26144
rect 7084 26144 7124 26790
rect 7276 26767 7316 26776
rect 7371 26776 7372 26816
rect 7179 26732 7221 26741
rect 7371 26734 7412 26776
rect 7179 26692 7180 26732
rect 7220 26692 7221 26732
rect 7179 26683 7221 26692
rect 6603 26095 6645 26104
rect 6926 26129 6966 26138
rect 6507 25808 6549 25817
rect 6507 25768 6508 25808
rect 6548 25768 6549 25808
rect 6507 25759 6549 25768
rect 6604 25472 6644 26095
rect 7084 26095 7124 26104
rect 7180 26144 7220 26683
rect 7372 26573 7412 26734
rect 7371 26564 7413 26573
rect 7371 26524 7372 26564
rect 7412 26524 7413 26564
rect 7371 26515 7413 26524
rect 7275 26480 7317 26489
rect 7275 26440 7276 26480
rect 7316 26440 7317 26480
rect 7275 26431 7317 26440
rect 7180 26095 7220 26104
rect 6700 25976 6740 25985
rect 6926 25976 6966 26089
rect 6740 25936 6966 25976
rect 6700 25927 6740 25936
rect 6987 25808 7029 25817
rect 6987 25768 6988 25808
rect 7028 25768 7029 25808
rect 6987 25759 7029 25768
rect 7179 25808 7221 25817
rect 7179 25768 7180 25808
rect 7220 25768 7221 25808
rect 7179 25759 7221 25768
rect 6604 25432 6740 25472
rect 6603 25304 6645 25313
rect 6603 25264 6604 25304
rect 6644 25264 6645 25304
rect 6603 25255 6645 25264
rect 6604 25170 6644 25255
rect 6412 25012 6644 25052
rect 6507 24800 6549 24809
rect 6316 24760 6452 24800
rect 6315 24632 6357 24641
rect 6315 24592 6316 24632
rect 6356 24592 6357 24632
rect 6315 24583 6357 24592
rect 6316 24498 6356 24583
rect 6412 24380 6452 24760
rect 6507 24760 6508 24800
rect 6548 24760 6549 24800
rect 6507 24751 6549 24760
rect 6508 24632 6548 24751
rect 6604 24632 6644 25012
rect 6700 24800 6740 25432
rect 6700 24751 6740 24760
rect 6892 24632 6932 24643
rect 6604 24592 6836 24632
rect 6508 24583 6548 24592
rect 6507 24464 6549 24473
rect 6507 24424 6508 24464
rect 6548 24424 6549 24464
rect 6507 24415 6549 24424
rect 6220 23575 6260 23584
rect 6316 24340 6452 24380
rect 6316 23456 6356 24340
rect 6508 24330 6548 24415
rect 6700 24380 6740 24389
rect 6604 24340 6700 24380
rect 6412 23885 6452 23970
rect 6411 23876 6453 23885
rect 6411 23836 6412 23876
rect 6452 23836 6453 23876
rect 6411 23827 6453 23836
rect 6508 23792 6548 23801
rect 6604 23792 6644 24340
rect 6700 24331 6740 24340
rect 6548 23752 6644 23792
rect 6508 23743 6548 23752
rect 6316 23416 6452 23456
rect 6316 23288 6356 23297
rect 6124 23248 6316 23288
rect 6316 23239 6356 23248
rect 6123 23120 6165 23129
rect 6123 23080 6124 23120
rect 6164 23080 6165 23120
rect 6123 23071 6165 23080
rect 6124 22986 6164 23071
rect 6219 22784 6261 22793
rect 6219 22744 6220 22784
rect 6260 22744 6261 22784
rect 6219 22735 6261 22744
rect 6124 22112 6164 22121
rect 6124 21953 6164 22072
rect 6123 21944 6165 21953
rect 6123 21904 6124 21944
rect 6164 21904 6165 21944
rect 6123 21895 6165 21904
rect 6027 21776 6069 21785
rect 6027 21736 6028 21776
rect 6068 21736 6069 21776
rect 6027 21727 6069 21736
rect 6028 21642 6068 21727
rect 6123 21608 6165 21617
rect 6123 21568 6124 21608
rect 6164 21568 6165 21608
rect 6123 21559 6165 21568
rect 5932 21484 6068 21524
rect 5835 20768 5877 20777
rect 5932 20768 5972 20777
rect 5835 20728 5836 20768
rect 5876 20728 5932 20768
rect 5835 20719 5877 20728
rect 5932 20719 5972 20728
rect 5836 20634 5876 20719
rect 5835 20432 5877 20441
rect 5835 20392 5836 20432
rect 5876 20392 5877 20432
rect 5835 20383 5877 20392
rect 5644 20140 5780 20180
rect 5740 19937 5780 20140
rect 5836 20096 5876 20383
rect 5739 19928 5781 19937
rect 5739 19888 5740 19928
rect 5780 19888 5781 19928
rect 5739 19879 5781 19888
rect 5740 19265 5780 19879
rect 5108 19216 5396 19256
rect 5068 19207 5108 19216
rect 4395 19088 4437 19097
rect 4395 19048 4396 19088
rect 4436 19048 4437 19088
rect 4395 19039 4437 19048
rect 4203 18836 4245 18845
rect 4203 18796 4204 18836
rect 4244 18796 4245 18836
rect 4203 18787 4245 18796
rect 4204 18584 4244 18787
rect 4204 18535 4244 18544
rect 4107 18416 4149 18425
rect 4107 18376 4108 18416
rect 4148 18376 4149 18416
rect 4107 18367 4149 18376
rect 4011 18332 4053 18341
rect 4011 18292 4012 18332
rect 4052 18292 4053 18332
rect 4011 18283 4053 18292
rect 3688 18164 4056 18173
rect 3728 18124 3770 18164
rect 3810 18124 3852 18164
rect 3892 18124 3934 18164
rect 3974 18124 4016 18164
rect 4396 18164 4436 19039
rect 4928 18920 5296 18929
rect 4968 18880 5010 18920
rect 5050 18880 5092 18920
rect 5132 18880 5174 18920
rect 5214 18880 5256 18920
rect 4928 18871 5296 18880
rect 5259 18668 5301 18677
rect 5259 18628 5260 18668
rect 5300 18628 5301 18668
rect 5259 18619 5301 18628
rect 4396 18124 4532 18164
rect 3688 18115 4056 18124
rect 3532 17956 3668 17996
rect 3435 17947 3477 17956
rect 3436 17744 3476 17947
rect 3532 17744 3572 17753
rect 3436 17704 3532 17744
rect 3532 17585 3572 17704
rect 3628 17744 3668 17956
rect 3628 17695 3668 17704
rect 3916 17912 3956 17921
rect 3531 17576 3573 17585
rect 3531 17536 3532 17576
rect 3572 17536 3573 17576
rect 3531 17527 3573 17536
rect 3916 17165 3956 17872
rect 4108 17744 4148 17753
rect 4148 17704 4244 17744
rect 4108 17695 4148 17704
rect 3436 17156 3476 17165
rect 3436 16409 3476 17116
rect 3915 17156 3957 17165
rect 3915 17116 3916 17156
rect 3956 17116 3957 17156
rect 3915 17107 3957 17116
rect 4108 17072 4148 17083
rect 3628 17058 3668 17067
rect 3628 16829 3668 17018
rect 4108 16997 4148 17032
rect 4107 16988 4149 16997
rect 4107 16948 4108 16988
rect 4148 16948 4149 16988
rect 4107 16939 4149 16948
rect 3627 16820 3669 16829
rect 3627 16780 3628 16820
rect 3668 16780 3669 16820
rect 3627 16771 3669 16780
rect 4107 16820 4149 16829
rect 4107 16780 4108 16820
rect 4148 16780 4149 16820
rect 4107 16771 4149 16780
rect 3688 16652 4056 16661
rect 3728 16612 3770 16652
rect 3810 16612 3852 16652
rect 3892 16612 3934 16652
rect 3974 16612 4016 16652
rect 3688 16603 4056 16612
rect 3435 16400 3477 16409
rect 3435 16360 3436 16400
rect 3476 16360 3477 16400
rect 3435 16351 3477 16360
rect 3915 16400 3957 16409
rect 3915 16360 3916 16400
rect 3956 16360 3957 16400
rect 3820 16325 3860 16356
rect 3915 16351 3957 16360
rect 3819 16316 3861 16325
rect 3819 16276 3820 16316
rect 3860 16276 3861 16316
rect 3819 16267 3861 16276
rect 3723 16232 3765 16241
rect 3723 16192 3724 16232
rect 3764 16192 3765 16232
rect 3723 16183 3765 16192
rect 3820 16232 3860 16267
rect 3724 15821 3764 16183
rect 3723 15812 3765 15821
rect 3723 15772 3724 15812
rect 3764 15772 3765 15812
rect 3723 15763 3765 15772
rect 3820 15308 3860 16192
rect 3916 15392 3956 16351
rect 4108 15728 4148 16771
rect 4204 16409 4244 17704
rect 4203 16400 4245 16409
rect 4203 16360 4204 16400
rect 4244 16360 4245 16400
rect 4203 16351 4245 16360
rect 4203 16232 4245 16241
rect 4203 16192 4204 16232
rect 4244 16192 4245 16232
rect 4203 16183 4245 16192
rect 4300 16232 4340 16241
rect 4204 16098 4244 16183
rect 4204 15728 4244 15737
rect 4108 15688 4204 15728
rect 4204 15679 4244 15688
rect 4012 15569 4052 15654
rect 4011 15560 4053 15569
rect 4011 15520 4012 15560
rect 4052 15520 4053 15560
rect 4011 15511 4053 15520
rect 3916 15352 4148 15392
rect 3532 15268 3860 15308
rect 3532 14972 3572 15268
rect 3688 15140 4056 15149
rect 3728 15100 3770 15140
rect 3810 15100 3852 15140
rect 3892 15100 3934 15140
rect 3974 15100 4016 15140
rect 3688 15091 4056 15100
rect 3532 14932 3668 14972
rect 3436 14720 3476 14729
rect 3339 13460 3381 13469
rect 3339 13420 3340 13460
rect 3380 13420 3381 13460
rect 3339 13411 3381 13420
rect 3339 13040 3381 13049
rect 3339 13000 3340 13040
rect 3380 13000 3381 13040
rect 3339 12991 3381 13000
rect 3340 12906 3380 12991
rect 3244 12748 3380 12788
rect 2708 11908 2804 11948
rect 2668 11899 2708 11908
rect 2955 11780 2997 11789
rect 2955 11740 2956 11780
rect 2996 11740 2997 11780
rect 2955 11731 2997 11740
rect 2859 11696 2901 11705
rect 2859 11656 2860 11696
rect 2900 11656 2901 11696
rect 2859 11647 2901 11656
rect 2956 11696 2996 11731
rect 2763 11612 2805 11621
rect 2763 11572 2764 11612
rect 2804 11572 2805 11612
rect 2763 11563 2805 11572
rect 2667 11444 2709 11453
rect 2667 11404 2668 11444
rect 2708 11404 2709 11444
rect 2667 11395 2709 11404
rect 2571 10184 2613 10193
rect 2571 10144 2572 10184
rect 2612 10144 2613 10184
rect 2571 10135 2613 10144
rect 2668 10184 2708 11395
rect 2764 11117 2804 11563
rect 2860 11562 2900 11647
rect 2956 11645 2996 11656
rect 2859 11276 2901 11285
rect 2859 11236 2860 11276
rect 2900 11236 2901 11276
rect 2859 11227 2901 11236
rect 2763 11108 2805 11117
rect 2763 11068 2764 11108
rect 2804 11068 2805 11108
rect 2763 11059 2805 11068
rect 2668 10135 2708 10144
rect 2667 9512 2709 9521
rect 2667 9472 2668 9512
rect 2708 9472 2709 9512
rect 2667 9463 2709 9472
rect 2283 8800 2284 8840
rect 2324 8800 2325 8840
rect 2103 8672 2143 8800
rect 2283 8791 2325 8800
rect 2380 8800 2516 8840
rect 2380 8756 2420 8800
rect 2092 8632 2143 8672
rect 2188 8743 2228 8752
rect 1995 8168 2037 8177
rect 1995 8128 1996 8168
rect 2036 8128 2037 8168
rect 1995 8119 2037 8128
rect 1899 6992 1941 7001
rect 1899 6952 1900 6992
rect 1940 6952 1941 6992
rect 1899 6943 1941 6952
rect 1803 6908 1845 6917
rect 1803 6868 1804 6908
rect 1844 6868 1845 6908
rect 1803 6859 1845 6868
rect 1515 6448 1516 6488
rect 1556 6448 1557 6488
rect 1515 6439 1557 6448
rect 1612 6448 1748 6488
rect 1420 6355 1460 6364
rect 1420 4892 1460 4901
rect 1516 4892 1556 6439
rect 1460 4852 1556 4892
rect 1420 4843 1460 4852
rect 1324 4264 1460 4304
rect 1323 4136 1365 4145
rect 1323 4096 1324 4136
rect 1364 4096 1365 4136
rect 1323 4087 1365 4096
rect 1324 4002 1364 4087
rect 1324 3632 1364 3641
rect 1420 3632 1460 4264
rect 1515 4220 1557 4229
rect 1515 4180 1516 4220
rect 1556 4180 1557 4220
rect 1515 4171 1557 4180
rect 1364 3592 1460 3632
rect 1324 3583 1364 3592
rect 1516 3548 1556 4171
rect 1420 3508 1556 3548
rect 1420 2624 1460 3508
rect 1515 3380 1557 3389
rect 1515 3340 1516 3380
rect 1556 3340 1557 3380
rect 1515 3331 1557 3340
rect 1516 3246 1556 3331
rect 1420 2575 1460 2584
rect 1515 2036 1557 2045
rect 1515 1996 1516 2036
rect 1556 1996 1557 2036
rect 1515 1987 1557 1996
rect 1227 1868 1269 1877
rect 1227 1828 1228 1868
rect 1268 1828 1269 1868
rect 1227 1819 1269 1828
rect 1228 1734 1268 1819
rect 1419 1700 1461 1709
rect 1419 1660 1420 1700
rect 1460 1660 1461 1700
rect 1419 1651 1461 1660
rect 1420 1566 1460 1651
rect 1420 1112 1460 1121
rect 1516 1112 1556 1987
rect 1612 1868 1652 6448
rect 1804 6404 1844 6859
rect 1899 6824 1941 6833
rect 1899 6784 1900 6824
rect 1940 6784 1941 6824
rect 1899 6775 1941 6784
rect 1804 6355 1844 6364
rect 1707 6320 1749 6329
rect 1707 6280 1708 6320
rect 1748 6280 1749 6320
rect 1707 6271 1749 6280
rect 1708 4808 1748 6271
rect 1900 4892 1940 6775
rect 1996 6749 2036 8119
rect 2092 7169 2132 8632
rect 2188 7925 2228 8703
rect 2373 8716 2420 8756
rect 2373 8672 2413 8716
rect 2284 8632 2413 8672
rect 2476 8672 2516 8681
rect 2187 7916 2229 7925
rect 2187 7876 2188 7916
rect 2228 7876 2229 7916
rect 2187 7867 2229 7876
rect 2091 7160 2133 7169
rect 2091 7120 2092 7160
rect 2132 7120 2133 7160
rect 2091 7111 2133 7120
rect 1995 6740 2037 6749
rect 1995 6700 1996 6740
rect 2036 6700 2037 6740
rect 1995 6691 2037 6700
rect 2091 6656 2133 6665
rect 2091 6616 2092 6656
rect 2132 6616 2133 6656
rect 2091 6607 2133 6616
rect 2092 6522 2132 6607
rect 1900 4843 1940 4852
rect 1996 6488 2036 6497
rect 1708 4759 1748 4768
rect 1996 3800 2036 6448
rect 2188 6488 2228 6497
rect 2188 6329 2228 6448
rect 2187 6320 2229 6329
rect 2187 6280 2188 6320
rect 2228 6280 2229 6320
rect 2187 6271 2229 6280
rect 2091 4892 2133 4901
rect 2091 4852 2092 4892
rect 2132 4852 2133 4892
rect 2284 4892 2324 8632
rect 2380 6497 2420 6582
rect 2379 6488 2421 6497
rect 2379 6448 2380 6488
rect 2420 6448 2421 6488
rect 2379 6439 2421 6448
rect 2379 6320 2421 6329
rect 2379 6280 2380 6320
rect 2420 6280 2421 6320
rect 2379 6271 2421 6280
rect 2380 6186 2420 6271
rect 2476 5816 2516 8632
rect 2572 8672 2612 8683
rect 2572 8597 2612 8632
rect 2571 8588 2613 8597
rect 2571 8548 2572 8588
rect 2612 8548 2613 8588
rect 2571 8539 2613 8548
rect 2572 7160 2612 7169
rect 2572 7001 2612 7120
rect 2571 6992 2613 7001
rect 2571 6952 2572 6992
rect 2612 6952 2613 6992
rect 2571 6943 2613 6952
rect 2572 6488 2612 6497
rect 2572 6329 2612 6448
rect 2571 6320 2613 6329
rect 2571 6280 2572 6320
rect 2612 6280 2613 6320
rect 2668 6320 2708 9463
rect 2764 8177 2804 11059
rect 2860 10436 2900 11227
rect 2860 10387 2900 10396
rect 3052 10436 3092 12482
rect 3147 11948 3189 11957
rect 3147 11908 3148 11948
rect 3188 11908 3189 11948
rect 3147 11899 3189 11908
rect 3148 11696 3188 11899
rect 3148 11647 3188 11656
rect 3243 10856 3285 10865
rect 3243 10816 3244 10856
rect 3284 10816 3285 10856
rect 3243 10807 3285 10816
rect 3052 10387 3092 10396
rect 3244 10184 3284 10807
rect 3244 10100 3284 10144
rect 2860 10060 3284 10100
rect 2860 9491 2900 10060
rect 3051 9848 3093 9857
rect 3051 9808 3052 9848
rect 3092 9808 3093 9848
rect 3051 9799 3093 9808
rect 3052 9680 3092 9799
rect 3052 9631 3092 9640
rect 3340 9605 3380 12748
rect 3436 11453 3476 14680
rect 3531 14720 3573 14729
rect 3531 14680 3532 14720
rect 3572 14680 3573 14720
rect 3531 14671 3573 14680
rect 3532 14586 3572 14671
rect 3628 13964 3668 14932
rect 3915 14888 3957 14897
rect 3915 14848 3916 14888
rect 3956 14848 3957 14888
rect 3915 14839 3957 14848
rect 3916 14804 3956 14839
rect 3916 14753 3956 14764
rect 4011 14804 4053 14813
rect 4011 14764 4012 14804
rect 4052 14764 4053 14804
rect 4011 14755 4053 14764
rect 4012 14670 4052 14755
rect 4108 14645 4148 15352
rect 4300 14981 4340 16192
rect 4396 15560 4436 15569
rect 4396 15317 4436 15520
rect 4395 15308 4437 15317
rect 4395 15268 4396 15308
rect 4436 15268 4437 15308
rect 4395 15259 4437 15268
rect 4299 14972 4341 14981
rect 4299 14932 4300 14972
rect 4340 14932 4341 14972
rect 4299 14923 4341 14932
rect 4492 14720 4532 18124
rect 5260 17576 5300 18619
rect 5356 17744 5396 19216
rect 5548 19256 5588 19265
rect 5548 18752 5588 19216
rect 5644 19256 5684 19265
rect 5644 19013 5684 19216
rect 5739 19256 5781 19265
rect 5739 19216 5740 19256
rect 5780 19216 5781 19256
rect 5739 19207 5781 19216
rect 5643 19004 5685 19013
rect 5643 18964 5644 19004
rect 5684 18964 5685 19004
rect 5643 18955 5685 18964
rect 5644 18752 5684 18761
rect 5548 18712 5644 18752
rect 5644 18703 5684 18712
rect 5836 18593 5876 20056
rect 6028 20012 6068 21484
rect 6124 21020 6164 21559
rect 6124 20971 6164 20980
rect 6220 20180 6260 22735
rect 6315 21608 6357 21617
rect 6315 21568 6316 21608
rect 6356 21568 6357 21608
rect 6315 21559 6357 21568
rect 6412 21608 6452 23416
rect 6603 23372 6645 23381
rect 6603 23332 6604 23372
rect 6644 23332 6645 23372
rect 6603 23323 6645 23332
rect 6508 22280 6548 22289
rect 6508 21785 6548 22240
rect 6604 22280 6644 23323
rect 6699 23120 6741 23129
rect 6699 23080 6700 23120
rect 6740 23080 6741 23120
rect 6699 23071 6741 23080
rect 6700 22986 6740 23071
rect 6796 22868 6836 24592
rect 6892 24557 6932 24592
rect 6891 24548 6933 24557
rect 6891 24508 6892 24548
rect 6932 24508 6933 24548
rect 6891 24499 6933 24508
rect 6891 23792 6933 23801
rect 6891 23752 6892 23792
rect 6932 23752 6933 23792
rect 6891 23743 6933 23752
rect 6604 22037 6644 22240
rect 6700 22828 6836 22868
rect 6603 22028 6645 22037
rect 6603 21988 6604 22028
rect 6644 21988 6645 22028
rect 6603 21979 6645 21988
rect 6507 21776 6549 21785
rect 6507 21736 6508 21776
rect 6548 21736 6549 21776
rect 6507 21727 6549 21736
rect 6452 21568 6548 21608
rect 6412 21559 6452 21568
rect 6316 21474 6356 21559
rect 6411 20936 6453 20945
rect 6411 20896 6412 20936
rect 6452 20896 6453 20936
rect 6411 20887 6453 20896
rect 6315 20768 6357 20777
rect 6315 20728 6316 20768
rect 6356 20728 6357 20768
rect 6315 20719 6357 20728
rect 6316 20634 6356 20719
rect 5932 19972 6068 20012
rect 6124 20140 6260 20180
rect 5451 18584 5493 18593
rect 5451 18544 5452 18584
rect 5492 18544 5493 18584
rect 5451 18535 5493 18544
rect 5835 18584 5877 18593
rect 5835 18544 5836 18584
rect 5876 18544 5877 18584
rect 5835 18535 5877 18544
rect 5452 18450 5492 18535
rect 5932 18341 5972 19972
rect 6027 19844 6069 19853
rect 6027 19804 6028 19844
rect 6068 19804 6069 19844
rect 6027 19795 6069 19804
rect 6028 19710 6068 19795
rect 6027 19256 6069 19265
rect 6027 19216 6028 19256
rect 6068 19216 6069 19256
rect 6027 19207 6069 19216
rect 6124 19256 6164 20140
rect 6316 20096 6356 20105
rect 6316 19517 6356 20056
rect 6412 20096 6452 20887
rect 6412 19769 6452 20056
rect 6411 19760 6453 19769
rect 6411 19720 6412 19760
rect 6452 19720 6453 19760
rect 6411 19711 6453 19720
rect 6315 19508 6357 19517
rect 6315 19468 6316 19508
rect 6356 19468 6357 19508
rect 6315 19459 6357 19468
rect 5451 18332 5493 18341
rect 5451 18292 5452 18332
rect 5492 18292 5493 18332
rect 5451 18283 5493 18292
rect 5931 18332 5973 18341
rect 5931 18292 5932 18332
rect 5972 18292 5973 18332
rect 5931 18283 5973 18292
rect 5356 17695 5396 17704
rect 5260 17536 5396 17576
rect 4587 17492 4629 17501
rect 4587 17452 4588 17492
rect 4628 17452 4629 17492
rect 4587 17443 4629 17452
rect 4588 17072 4628 17443
rect 4928 17408 5296 17417
rect 4968 17368 5010 17408
rect 5050 17368 5092 17408
rect 5132 17368 5174 17408
rect 5214 17368 5256 17408
rect 4928 17359 5296 17368
rect 4588 17023 4628 17032
rect 5068 17072 5108 17081
rect 4684 16988 4724 16999
rect 4684 16913 4724 16948
rect 4971 16988 5013 16997
rect 4971 16948 4972 16988
rect 5012 16948 5013 16988
rect 4971 16939 5013 16948
rect 4683 16904 4725 16913
rect 4683 16864 4684 16904
rect 4724 16864 4725 16904
rect 4683 16855 4725 16864
rect 4780 16316 4820 16325
rect 4972 16316 5012 16939
rect 5068 16400 5108 17032
rect 5163 17072 5205 17081
rect 5163 17032 5164 17072
rect 5204 17032 5205 17072
rect 5163 17023 5205 17032
rect 5164 16938 5204 17023
rect 5356 16904 5396 17536
rect 5452 17492 5492 18283
rect 5932 17753 5972 17838
rect 5836 17744 5876 17753
rect 5548 17660 5588 17669
rect 5836 17660 5876 17704
rect 5931 17744 5973 17753
rect 5931 17704 5932 17744
rect 5972 17704 5973 17744
rect 5931 17695 5973 17704
rect 5588 17620 5876 17660
rect 5548 17611 5588 17620
rect 6028 17576 6068 19207
rect 6124 18761 6164 19216
rect 6219 19172 6261 19181
rect 6219 19132 6220 19172
rect 6260 19132 6261 19172
rect 6219 19123 6261 19132
rect 6123 18752 6165 18761
rect 6123 18712 6124 18752
rect 6164 18712 6165 18752
rect 6123 18703 6165 18712
rect 6123 18584 6165 18593
rect 6123 18544 6124 18584
rect 6164 18544 6165 18584
rect 6123 18535 6165 18544
rect 6124 18450 6164 18535
rect 5932 17536 6068 17576
rect 5739 17492 5781 17501
rect 5452 17452 5684 17492
rect 5488 17156 5530 17165
rect 5488 17116 5489 17156
rect 5529 17116 5530 17156
rect 5488 17107 5530 17116
rect 5489 17072 5529 17107
rect 5489 17021 5529 17032
rect 5644 17072 5684 17452
rect 5739 17452 5740 17492
rect 5780 17452 5781 17492
rect 5739 17443 5781 17452
rect 5644 17023 5684 17032
rect 5740 17072 5780 17443
rect 5835 17240 5877 17249
rect 5835 17200 5836 17240
rect 5876 17200 5877 17240
rect 5835 17191 5877 17200
rect 5836 17106 5876 17191
rect 5740 17023 5780 17032
rect 5932 17072 5972 17536
rect 6220 17492 6260 19123
rect 6315 18164 6357 18173
rect 6315 18124 6316 18164
rect 6356 18124 6357 18164
rect 6315 18115 6357 18124
rect 6316 17828 6356 18115
rect 6411 17996 6453 18005
rect 6411 17956 6412 17996
rect 6452 17956 6453 17996
rect 6411 17947 6453 17956
rect 6316 17779 6356 17788
rect 6412 17828 6452 17947
rect 6412 17779 6452 17788
rect 6508 17753 6548 21568
rect 6700 20012 6740 22828
rect 6795 22700 6837 22709
rect 6795 22660 6796 22700
rect 6836 22660 6837 22700
rect 6795 22651 6837 22660
rect 6796 21776 6836 22651
rect 6892 22028 6932 23743
rect 6988 22709 7028 25759
rect 7180 24641 7220 25759
rect 7179 24632 7221 24641
rect 7179 24592 7180 24632
rect 7220 24592 7221 24632
rect 7179 24583 7221 24592
rect 6987 22700 7029 22709
rect 6987 22660 6988 22700
rect 7028 22660 7029 22700
rect 6987 22651 7029 22660
rect 6987 22532 7029 22541
rect 6987 22492 6988 22532
rect 7028 22492 7029 22532
rect 6987 22483 7029 22492
rect 6988 22364 7028 22483
rect 6988 22112 7028 22324
rect 7083 22364 7125 22373
rect 7083 22324 7084 22364
rect 7124 22324 7125 22364
rect 7083 22315 7125 22324
rect 7084 22230 7124 22315
rect 7179 22280 7221 22289
rect 7276 22280 7316 26431
rect 7371 26312 7413 26321
rect 7371 26272 7372 26312
rect 7412 26272 7413 26312
rect 7371 26263 7413 26272
rect 7372 26144 7412 26263
rect 7372 26095 7412 26104
rect 7468 26144 7508 27448
rect 7564 27404 7604 27691
rect 7564 26825 7604 27364
rect 7563 26816 7605 26825
rect 7563 26776 7564 26816
rect 7604 26776 7605 26816
rect 7563 26767 7605 26776
rect 7468 26095 7508 26104
rect 7563 25892 7605 25901
rect 7563 25852 7564 25892
rect 7604 25852 7605 25892
rect 7563 25843 7605 25852
rect 7467 25304 7509 25313
rect 7467 25264 7468 25304
rect 7508 25264 7509 25304
rect 7467 25255 7509 25264
rect 7179 22240 7180 22280
rect 7220 22240 7316 22280
rect 7179 22231 7221 22240
rect 6988 22072 7124 22112
rect 6892 21988 7028 22028
rect 6891 21776 6933 21785
rect 6796 21736 6892 21776
rect 6932 21736 6933 21776
rect 6891 21727 6933 21736
rect 6795 21608 6837 21617
rect 6795 21568 6796 21608
rect 6836 21568 6837 21608
rect 6795 21559 6837 21568
rect 6892 21608 6932 21727
rect 6892 21559 6932 21568
rect 6796 21474 6836 21559
rect 6891 21356 6933 21365
rect 6891 21316 6892 21356
rect 6932 21316 6933 21356
rect 6891 21307 6933 21316
rect 6892 21029 6932 21307
rect 6891 21020 6933 21029
rect 6891 20980 6892 21020
rect 6932 20980 6933 21020
rect 6891 20971 6933 20980
rect 6796 20012 6836 20040
rect 6700 19972 6796 20012
rect 6603 19256 6645 19265
rect 6603 19216 6604 19256
rect 6644 19216 6645 19256
rect 6603 19207 6645 19216
rect 6604 19122 6644 19207
rect 6700 18929 6740 19972
rect 6796 19963 6836 19972
rect 6892 20012 6932 20023
rect 6892 19937 6932 19972
rect 6891 19928 6933 19937
rect 6891 19888 6892 19928
rect 6932 19888 6933 19928
rect 6891 19879 6933 19888
rect 6699 18920 6741 18929
rect 6699 18880 6700 18920
rect 6740 18880 6741 18920
rect 6699 18871 6741 18880
rect 6988 18845 7028 21988
rect 7084 21617 7124 22072
rect 7083 21608 7125 21617
rect 7083 21568 7084 21608
rect 7124 21568 7125 21608
rect 7083 21559 7125 21568
rect 7083 19844 7125 19853
rect 7083 19804 7084 19844
rect 7124 19804 7125 19844
rect 7083 19795 7125 19804
rect 7084 19270 7124 19795
rect 7084 19221 7124 19230
rect 6987 18836 7029 18845
rect 6987 18796 6988 18836
rect 7028 18796 7029 18836
rect 6987 18787 7029 18796
rect 6988 18677 7028 18787
rect 6603 18668 6645 18677
rect 6603 18628 6604 18668
rect 6644 18628 6645 18668
rect 6603 18619 6645 18628
rect 6987 18668 7029 18677
rect 7180 18668 7220 22231
rect 7371 21608 7413 21617
rect 7371 21568 7372 21608
rect 7412 21568 7413 21608
rect 7371 21559 7413 21568
rect 7372 21474 7412 21559
rect 7372 20096 7412 20107
rect 7372 20021 7412 20056
rect 7371 20012 7413 20021
rect 7371 19972 7372 20012
rect 7412 19972 7413 20012
rect 7371 19963 7413 19972
rect 7468 19424 7508 25255
rect 7564 22616 7604 25843
rect 7660 25229 7700 29791
rect 7756 27656 7796 29968
rect 7852 29840 7892 30640
rect 7948 30521 7988 30640
rect 7947 30512 7989 30521
rect 7947 30472 7948 30512
rect 7988 30472 7989 30512
rect 7947 30463 7989 30472
rect 7948 30185 7988 30463
rect 7947 30176 7989 30185
rect 7947 30136 7948 30176
rect 7988 30136 7989 30176
rect 7947 30127 7989 30136
rect 8332 29849 8372 31480
rect 8428 31352 8468 31361
rect 8428 31109 8468 31312
rect 8427 31100 8469 31109
rect 8427 31060 8428 31100
rect 8468 31060 8469 31100
rect 8427 31051 8469 31060
rect 8428 30941 8468 31051
rect 8427 30932 8469 30941
rect 8427 30892 8428 30932
rect 8468 30892 8469 30932
rect 8427 30883 8469 30892
rect 8331 29840 8373 29849
rect 7852 29800 7988 29840
rect 7851 29672 7893 29681
rect 7851 29632 7852 29672
rect 7892 29632 7893 29672
rect 7851 29623 7893 29632
rect 7852 27740 7892 29623
rect 7852 27691 7892 27700
rect 7756 27607 7796 27616
rect 7948 27656 7988 29800
rect 8331 29800 8332 29840
rect 8372 29800 8373 29840
rect 8331 29791 8373 29800
rect 8523 29840 8565 29849
rect 8523 29800 8524 29840
rect 8564 29800 8565 29840
rect 8523 29791 8565 29800
rect 8427 29336 8469 29345
rect 8427 29296 8428 29336
rect 8468 29296 8469 29336
rect 8427 29287 8469 29296
rect 8236 29177 8276 29262
rect 8428 29202 8468 29287
rect 8524 29177 8564 29791
rect 8716 29681 8756 34159
rect 8812 33965 8852 34243
rect 9004 34049 9044 34336
rect 9003 34040 9045 34049
rect 9003 34000 9004 34040
rect 9044 34000 9045 34040
rect 9003 33991 9045 34000
rect 8811 33956 8853 33965
rect 8811 33916 8812 33956
rect 8852 33916 8853 33956
rect 8811 33907 8853 33916
rect 8811 33788 8853 33797
rect 8811 33748 8812 33788
rect 8852 33748 8853 33788
rect 8811 33739 8853 33748
rect 8812 32192 8852 33739
rect 9004 33293 9044 33991
rect 9003 33284 9045 33293
rect 9003 33244 9004 33284
rect 9044 33244 9045 33284
rect 9003 33235 9045 33244
rect 9003 33116 9045 33125
rect 9003 33076 9004 33116
rect 9044 33076 9045 33116
rect 9003 33067 9045 33076
rect 8812 32143 8852 32152
rect 9004 31268 9044 33067
rect 9100 31529 9140 36100
rect 9387 36056 9429 36065
rect 9387 36016 9388 36056
rect 9428 36016 9429 36056
rect 9387 36007 9429 36016
rect 9292 35972 9332 35981
rect 9196 35888 9236 35897
rect 9196 35141 9236 35848
rect 9195 35132 9237 35141
rect 9195 35092 9196 35132
rect 9236 35092 9237 35132
rect 9195 35083 9237 35092
rect 9195 34376 9237 34385
rect 9195 34336 9196 34376
rect 9236 34336 9237 34376
rect 9195 34327 9237 34336
rect 9196 34242 9236 34327
rect 9292 34049 9332 35932
rect 9388 35922 9428 36007
rect 9484 35972 9524 35981
rect 9484 35804 9524 35932
rect 9579 35888 9621 35897
rect 9579 35848 9580 35888
rect 9620 35848 9621 35888
rect 9579 35839 9621 35848
rect 9388 35764 9524 35804
rect 9388 35645 9428 35764
rect 9580 35754 9620 35839
rect 9387 35636 9429 35645
rect 9676 35636 9716 36520
rect 9387 35596 9388 35636
rect 9428 35596 9429 35636
rect 9387 35587 9429 35596
rect 9484 35596 9716 35636
rect 9387 34796 9429 34805
rect 9387 34756 9388 34796
rect 9428 34756 9429 34796
rect 9387 34747 9429 34756
rect 9291 34040 9333 34049
rect 9291 34000 9292 34040
rect 9332 34000 9333 34040
rect 9291 33991 9333 34000
rect 9388 32873 9428 34747
rect 9195 32864 9237 32873
rect 9195 32824 9196 32864
rect 9236 32824 9237 32864
rect 9195 32815 9237 32824
rect 9387 32864 9429 32873
rect 9387 32824 9388 32864
rect 9428 32824 9429 32864
rect 9387 32815 9429 32824
rect 9196 32730 9236 32815
rect 9387 32192 9429 32201
rect 9387 32152 9388 32192
rect 9428 32152 9429 32192
rect 9387 32143 9429 32152
rect 9099 31520 9141 31529
rect 9099 31480 9100 31520
rect 9140 31480 9141 31520
rect 9099 31471 9141 31480
rect 9195 31268 9237 31277
rect 9004 31228 9196 31268
rect 9236 31228 9237 31268
rect 9195 31219 9237 31228
rect 9196 30680 9236 31219
rect 9388 30848 9428 32143
rect 9388 30689 9428 30808
rect 9100 30640 9196 30680
rect 8907 30596 8949 30605
rect 8907 30556 8908 30596
rect 8948 30556 8949 30596
rect 8907 30547 8949 30556
rect 8812 29849 8852 29934
rect 8811 29840 8853 29849
rect 8811 29800 8812 29840
rect 8852 29800 8853 29840
rect 8811 29791 8853 29800
rect 8715 29672 8757 29681
rect 8908 29672 8948 30547
rect 9100 30353 9140 30640
rect 9196 30631 9236 30640
rect 9387 30680 9429 30689
rect 9387 30640 9388 30680
rect 9428 30640 9429 30680
rect 9387 30631 9429 30640
rect 9099 30344 9141 30353
rect 9099 30304 9100 30344
rect 9140 30304 9141 30344
rect 9099 30295 9141 30304
rect 9484 30185 9524 35596
rect 9772 35552 9812 36931
rect 9676 35512 9812 35552
rect 9579 35216 9621 35225
rect 9579 35176 9580 35216
rect 9620 35176 9621 35216
rect 9579 35167 9621 35176
rect 9580 35082 9620 35167
rect 9579 34628 9621 34637
rect 9579 34588 9580 34628
rect 9620 34588 9621 34628
rect 9579 34579 9621 34588
rect 9580 33713 9620 34579
rect 9579 33704 9621 33713
rect 9579 33664 9580 33704
rect 9620 33664 9621 33704
rect 9579 33655 9621 33664
rect 9676 33293 9716 35512
rect 9868 35468 9908 38191
rect 10060 38106 10100 38191
rect 9963 37988 10005 37997
rect 9963 37948 9964 37988
rect 10004 37948 10005 37988
rect 9963 37939 10005 37948
rect 9964 37854 10004 37939
rect 10059 37904 10101 37913
rect 10059 37864 10060 37904
rect 10100 37864 10101 37904
rect 10059 37855 10101 37864
rect 10060 36723 10100 37855
rect 10060 36674 10100 36683
rect 9772 35428 9908 35468
rect 9964 35888 10004 35897
rect 9772 35300 9812 35428
rect 9964 35300 10004 35848
rect 10156 35477 10196 39040
rect 10443 38996 10485 39005
rect 10443 38956 10444 38996
rect 10484 38956 10485 38996
rect 10443 38947 10485 38956
rect 10540 38996 10580 39005
rect 10580 38956 10772 38996
rect 10540 38947 10580 38956
rect 10251 38912 10293 38921
rect 10251 38872 10252 38912
rect 10292 38872 10293 38912
rect 10251 38863 10293 38872
rect 10252 38585 10292 38863
rect 10348 38744 10388 38753
rect 10444 38744 10484 38947
rect 10388 38704 10484 38744
rect 10348 38695 10388 38704
rect 10251 38576 10293 38585
rect 10251 38536 10252 38576
rect 10292 38536 10293 38576
rect 10251 38527 10293 38536
rect 10252 38240 10292 38249
rect 10252 36989 10292 38200
rect 10444 38240 10484 38249
rect 10484 38200 10580 38240
rect 10444 38191 10484 38200
rect 10444 37988 10484 37997
rect 10251 36980 10293 36989
rect 10251 36940 10252 36980
rect 10292 36940 10293 36980
rect 10251 36931 10293 36940
rect 10251 36812 10293 36821
rect 10251 36772 10252 36812
rect 10292 36772 10293 36812
rect 10251 36763 10293 36772
rect 10155 35468 10197 35477
rect 10155 35428 10156 35468
rect 10196 35428 10197 35468
rect 10155 35419 10197 35428
rect 10059 35384 10101 35393
rect 10059 35344 10060 35384
rect 10100 35344 10101 35384
rect 10059 35335 10101 35344
rect 9772 35251 9812 35260
rect 9868 35260 10004 35300
rect 9868 33797 9908 35260
rect 9964 35174 10004 35183
rect 9963 35134 9964 35141
rect 10004 35134 10005 35141
rect 9963 35132 10005 35134
rect 9963 35092 9964 35132
rect 10004 35092 10005 35132
rect 9963 35083 10005 35092
rect 9964 35039 10004 35083
rect 10060 34040 10100 35335
rect 10155 35300 10197 35309
rect 10155 35260 10156 35300
rect 10196 35260 10197 35300
rect 10155 35251 10197 35260
rect 9964 34000 10100 34040
rect 9867 33788 9909 33797
rect 9867 33748 9868 33788
rect 9908 33748 9909 33788
rect 9867 33739 9909 33748
rect 9868 33704 9908 33739
rect 9868 33545 9908 33664
rect 9867 33536 9909 33545
rect 9867 33496 9868 33536
rect 9908 33496 9909 33536
rect 9867 33487 9909 33496
rect 9675 33284 9717 33293
rect 9675 33244 9676 33284
rect 9716 33244 9717 33284
rect 9675 33235 9717 33244
rect 9580 32864 9620 32873
rect 9580 32537 9620 32824
rect 9675 32864 9717 32873
rect 9675 32824 9676 32864
rect 9716 32824 9717 32864
rect 9964 32864 10004 34000
rect 10059 33872 10101 33881
rect 10059 33832 10060 33872
rect 10100 33832 10101 33872
rect 10059 33823 10101 33832
rect 10060 33704 10100 33823
rect 10060 33655 10100 33664
rect 10059 33452 10101 33461
rect 10059 33412 10060 33452
rect 10100 33412 10101 33452
rect 10059 33403 10101 33412
rect 10060 33318 10100 33403
rect 10156 32948 10196 35251
rect 10252 33881 10292 36763
rect 10444 36737 10484 37948
rect 10540 37829 10580 38200
rect 10636 38156 10676 38165
rect 10539 37820 10581 37829
rect 10539 37780 10540 37820
rect 10580 37780 10581 37820
rect 10539 37771 10581 37780
rect 10636 36812 10676 38116
rect 10540 36772 10676 36812
rect 10443 36728 10485 36737
rect 10443 36688 10444 36728
rect 10484 36688 10485 36728
rect 10443 36679 10485 36688
rect 10347 36056 10389 36065
rect 10347 36016 10348 36056
rect 10388 36016 10389 36056
rect 10347 36007 10389 36016
rect 10251 33872 10293 33881
rect 10251 33832 10252 33872
rect 10292 33832 10293 33872
rect 10251 33823 10293 33832
rect 10252 33704 10292 33713
rect 10252 33125 10292 33664
rect 10348 33704 10388 36007
rect 10443 35132 10485 35141
rect 10443 35092 10444 35132
rect 10484 35092 10485 35132
rect 10443 35083 10485 35092
rect 10444 34376 10484 35083
rect 10444 34301 10484 34336
rect 10443 34292 10485 34301
rect 10443 34252 10444 34292
rect 10484 34252 10485 34292
rect 10443 34243 10485 34252
rect 10444 34133 10484 34243
rect 10443 34124 10485 34133
rect 10443 34084 10444 34124
rect 10484 34084 10485 34124
rect 10443 34075 10485 34084
rect 10540 33872 10580 36772
rect 10636 36644 10676 36653
rect 10636 35561 10676 36604
rect 10635 35552 10677 35561
rect 10635 35512 10636 35552
rect 10676 35512 10677 35552
rect 10635 35503 10677 35512
rect 10732 35309 10772 38956
rect 10828 38912 10868 39376
rect 10924 39257 10964 39544
rect 10923 39248 10965 39257
rect 10923 39208 10924 39248
rect 10964 39208 10965 39248
rect 10923 39199 10965 39208
rect 10923 39080 10965 39089
rect 10923 39040 10924 39080
rect 10964 39040 10965 39080
rect 10923 39031 10965 39040
rect 10828 38863 10868 38872
rect 10924 38912 10964 39031
rect 10924 38863 10964 38872
rect 11020 38744 11060 40123
rect 11212 40097 11252 42928
rect 11307 41600 11349 41609
rect 11307 41560 11308 41600
rect 11348 41560 11349 41600
rect 11307 41551 11349 41560
rect 11211 40088 11253 40097
rect 11211 40048 11212 40088
rect 11252 40048 11253 40088
rect 11211 40039 11253 40048
rect 11308 39920 11348 41551
rect 11404 39929 11444 42928
rect 11499 41012 11541 41021
rect 11499 40972 11500 41012
rect 11540 40972 11541 41012
rect 11499 40963 11541 40972
rect 11500 40438 11540 40963
rect 11500 40389 11540 40398
rect 11499 40256 11541 40265
rect 11499 40216 11500 40256
rect 11540 40216 11541 40256
rect 11499 40207 11541 40216
rect 11212 39880 11348 39920
rect 11403 39920 11445 39929
rect 11403 39880 11404 39920
rect 11444 39880 11445 39920
rect 11115 39416 11157 39425
rect 11115 39376 11116 39416
rect 11156 39376 11157 39416
rect 11115 39367 11157 39376
rect 10828 38704 11060 38744
rect 10828 38408 10868 38704
rect 11019 38576 11061 38585
rect 11019 38536 11020 38576
rect 11060 38536 11061 38576
rect 11019 38527 11061 38536
rect 10828 38359 10868 38368
rect 10923 37484 10965 37493
rect 10923 37444 10924 37484
rect 10964 37444 10965 37484
rect 10923 37435 10965 37444
rect 10827 37148 10869 37157
rect 10827 37108 10828 37148
rect 10868 37108 10869 37148
rect 10827 37099 10869 37108
rect 10828 36821 10868 37099
rect 10827 36812 10869 36821
rect 10827 36772 10828 36812
rect 10868 36772 10869 36812
rect 10827 36763 10869 36772
rect 10924 36644 10964 37435
rect 11020 37400 11060 38527
rect 11116 38240 11156 39367
rect 11212 39257 11252 39880
rect 11403 39871 11445 39880
rect 11320 39761 11360 39780
rect 11308 39752 11360 39761
rect 11403 39752 11445 39761
rect 11348 39712 11404 39752
rect 11444 39712 11445 39752
rect 11308 39703 11348 39712
rect 11403 39703 11445 39712
rect 11211 39248 11253 39257
rect 11211 39208 11212 39248
rect 11252 39208 11253 39248
rect 11211 39199 11253 39208
rect 11211 39080 11253 39089
rect 11211 39040 11212 39080
rect 11252 39040 11253 39080
rect 11211 39031 11253 39040
rect 11116 38191 11156 38200
rect 11212 38240 11252 39031
rect 11404 38996 11444 39005
rect 11500 38996 11540 40207
rect 11444 38956 11540 38996
rect 11404 38947 11444 38956
rect 11212 37913 11252 38200
rect 11308 38912 11348 38921
rect 11308 38165 11348 38872
rect 11500 38492 11540 38956
rect 11596 38669 11636 42928
rect 11691 42188 11733 42197
rect 11691 42148 11692 42188
rect 11732 42148 11733 42188
rect 11691 42139 11733 42148
rect 11692 40433 11732 42139
rect 11691 40424 11733 40433
rect 11691 40384 11692 40424
rect 11732 40384 11733 40424
rect 11788 40424 11828 42928
rect 11980 42113 12020 42928
rect 11979 42104 12021 42113
rect 11979 42064 11980 42104
rect 12020 42064 12021 42104
rect 11979 42055 12021 42064
rect 11883 41348 11925 41357
rect 11883 41308 11884 41348
rect 11924 41308 11925 41348
rect 11883 41299 11925 41308
rect 11884 41264 11924 41299
rect 11884 41213 11924 41224
rect 12172 41189 12212 42928
rect 12364 42533 12404 42928
rect 12363 42524 12405 42533
rect 12363 42484 12364 42524
rect 12404 42484 12405 42524
rect 12363 42475 12405 42484
rect 12556 41609 12596 42928
rect 12555 41600 12597 41609
rect 12555 41560 12556 41600
rect 12596 41560 12597 41600
rect 12555 41551 12597 41560
rect 12651 41432 12693 41441
rect 12651 41392 12652 41432
rect 12692 41392 12693 41432
rect 12651 41383 12693 41392
rect 12555 41348 12597 41357
rect 12555 41308 12556 41348
rect 12596 41308 12597 41348
rect 12555 41299 12597 41308
rect 12459 41264 12501 41273
rect 12459 41224 12460 41264
rect 12500 41224 12501 41264
rect 12459 41215 12501 41224
rect 12171 41180 12213 41189
rect 12171 41140 12172 41180
rect 12212 41140 12213 41180
rect 12171 41131 12213 41140
rect 12460 41130 12500 41215
rect 12076 41012 12116 41021
rect 12267 41012 12309 41021
rect 12116 40972 12212 41012
rect 12076 40963 12116 40972
rect 12076 40424 12116 40433
rect 11788 40384 11924 40424
rect 11691 40375 11733 40384
rect 11692 40256 11732 40265
rect 11732 40216 11828 40256
rect 11692 40207 11732 40216
rect 11595 38660 11637 38669
rect 11595 38620 11596 38660
rect 11636 38620 11637 38660
rect 11595 38611 11637 38620
rect 11500 38452 11732 38492
rect 11692 38240 11732 38452
rect 11307 38156 11349 38165
rect 11307 38116 11308 38156
rect 11348 38116 11349 38156
rect 11307 38107 11349 38116
rect 11595 38156 11637 38165
rect 11595 38116 11596 38156
rect 11636 38116 11637 38156
rect 11595 38107 11637 38116
rect 11596 38022 11636 38107
rect 11211 37904 11253 37913
rect 11211 37864 11212 37904
rect 11252 37864 11253 37904
rect 11211 37855 11253 37864
rect 11595 37904 11637 37913
rect 11595 37864 11596 37904
rect 11636 37864 11637 37904
rect 11595 37855 11637 37864
rect 11115 37820 11157 37829
rect 11115 37780 11116 37820
rect 11156 37780 11157 37820
rect 11115 37771 11157 37780
rect 11020 37073 11060 37360
rect 11019 37064 11061 37073
rect 11019 37024 11020 37064
rect 11060 37024 11061 37064
rect 11019 37015 11061 37024
rect 11020 36644 11060 36653
rect 10924 36604 11020 36644
rect 10827 36560 10869 36569
rect 10827 36520 10828 36560
rect 10868 36520 10869 36560
rect 10827 36511 10869 36520
rect 10828 36426 10868 36511
rect 10731 35300 10773 35309
rect 10731 35260 10732 35300
rect 10772 35260 10773 35300
rect 10731 35251 10773 35260
rect 10924 35141 10964 36604
rect 11020 36595 11060 36604
rect 11116 35561 11156 37771
rect 11596 37409 11636 37855
rect 11692 37577 11732 38200
rect 11691 37568 11733 37577
rect 11691 37528 11692 37568
rect 11732 37528 11733 37568
rect 11691 37519 11733 37528
rect 11500 37400 11540 37409
rect 11212 37360 11500 37400
rect 11212 37316 11252 37360
rect 11500 37351 11540 37360
rect 11595 37400 11637 37409
rect 11595 37360 11596 37400
rect 11636 37360 11637 37400
rect 11595 37351 11637 37360
rect 11212 37267 11252 37276
rect 11596 37266 11636 37351
rect 11211 36896 11253 36905
rect 11788 36896 11828 40216
rect 11884 39416 11924 40384
rect 11980 40384 12076 40424
rect 11980 39593 12020 40384
rect 12076 40375 12116 40384
rect 12172 40172 12212 40972
rect 12267 40972 12268 41012
rect 12308 40972 12309 41012
rect 12267 40963 12309 40972
rect 12268 40878 12308 40963
rect 12172 40132 12404 40172
rect 11979 39584 12021 39593
rect 11979 39544 11980 39584
rect 12020 39544 12021 39584
rect 11979 39535 12021 39544
rect 11884 39376 12116 39416
rect 11883 38912 11925 38921
rect 11883 38872 11884 38912
rect 11924 38872 11925 38912
rect 11883 38863 11925 38872
rect 11884 38778 11924 38863
rect 11979 38828 12021 38837
rect 11979 38788 11980 38828
rect 12020 38788 12021 38828
rect 11979 38779 12021 38788
rect 11883 38660 11925 38669
rect 11883 38620 11884 38660
rect 11924 38620 11925 38660
rect 11883 38611 11925 38620
rect 11211 36856 11212 36896
rect 11252 36856 11253 36896
rect 11211 36847 11253 36856
rect 11692 36856 11828 36896
rect 11212 36762 11252 36847
rect 11404 36644 11444 36653
rect 11211 35972 11253 35981
rect 11211 35932 11212 35972
rect 11252 35932 11253 35972
rect 11211 35923 11253 35932
rect 11212 35888 11252 35923
rect 11404 35888 11444 36604
rect 11596 36476 11636 36485
rect 11596 36065 11636 36436
rect 11595 36056 11637 36065
rect 11595 36016 11596 36056
rect 11636 36016 11637 36056
rect 11595 36007 11637 36016
rect 11212 35837 11252 35848
rect 11308 35848 11444 35888
rect 11596 35888 11636 35897
rect 11115 35552 11157 35561
rect 11115 35512 11116 35552
rect 11156 35512 11157 35552
rect 11115 35503 11157 35512
rect 11019 35384 11061 35393
rect 11019 35344 11020 35384
rect 11060 35344 11061 35384
rect 11019 35335 11061 35344
rect 10923 35132 10965 35141
rect 10923 35092 10924 35132
rect 10964 35092 10965 35132
rect 10923 35083 10965 35092
rect 10923 34544 10965 34553
rect 10923 34504 10924 34544
rect 10964 34504 10965 34544
rect 10923 34495 10965 34504
rect 10828 34376 10868 34385
rect 10828 34217 10868 34336
rect 10348 33655 10388 33664
rect 10444 33832 10580 33872
rect 10636 34208 10676 34217
rect 10251 33116 10293 33125
rect 10251 33076 10252 33116
rect 10292 33076 10293 33116
rect 10251 33067 10293 33076
rect 10347 32948 10389 32957
rect 10156 32908 10292 32948
rect 10060 32864 10100 32873
rect 9964 32824 10060 32864
rect 10252 32864 10292 32908
rect 10347 32908 10348 32948
rect 10388 32908 10389 32948
rect 10347 32899 10389 32908
rect 9675 32815 9717 32824
rect 10060 32815 10100 32824
rect 10156 32843 10196 32852
rect 9676 32730 9716 32815
rect 10252 32815 10292 32824
rect 10348 32864 10388 32899
rect 10348 32813 10388 32824
rect 9868 32696 9908 32705
rect 9772 32656 9868 32696
rect 9579 32528 9621 32537
rect 9579 32488 9580 32528
rect 9620 32488 9621 32528
rect 9579 32479 9621 32488
rect 9579 32024 9621 32033
rect 9579 31984 9580 32024
rect 9620 31984 9621 32024
rect 9579 31975 9621 31984
rect 9580 30680 9620 31975
rect 9676 31352 9716 31363
rect 9676 31277 9716 31312
rect 9675 31268 9717 31277
rect 9675 31228 9676 31268
rect 9716 31228 9717 31268
rect 9675 31219 9717 31228
rect 9580 30631 9620 30640
rect 9675 30680 9717 30689
rect 9675 30640 9676 30680
rect 9716 30640 9717 30680
rect 9772 30680 9812 32656
rect 9868 32647 9908 32656
rect 10059 32696 10101 32705
rect 10059 32656 10060 32696
rect 10100 32656 10101 32696
rect 10059 32647 10101 32656
rect 9867 32528 9909 32537
rect 9867 32488 9868 32528
rect 9908 32488 9909 32528
rect 9867 32479 9909 32488
rect 9868 31604 9908 32479
rect 10060 32192 10100 32647
rect 9868 31555 9908 31564
rect 9964 32152 10060 32192
rect 9964 31277 10004 32152
rect 10060 32143 10100 32152
rect 10059 31856 10101 31865
rect 10059 31816 10060 31856
rect 10100 31816 10101 31856
rect 10059 31807 10101 31816
rect 10060 31352 10100 31807
rect 10156 31445 10196 32803
rect 10444 32705 10484 33832
rect 10539 33704 10581 33713
rect 10539 33664 10540 33704
rect 10580 33664 10581 33704
rect 10539 33655 10581 33664
rect 10636 33704 10676 34168
rect 10827 34208 10869 34217
rect 10827 34168 10828 34208
rect 10868 34168 10869 34208
rect 10827 34159 10869 34168
rect 10636 33655 10676 33664
rect 10732 33704 10772 33713
rect 10540 32873 10580 33655
rect 10539 32864 10581 32873
rect 10636 32864 10676 32873
rect 10539 32824 10540 32864
rect 10580 32824 10636 32864
rect 10539 32815 10581 32824
rect 10636 32815 10676 32824
rect 10540 32730 10580 32815
rect 10443 32696 10485 32705
rect 10443 32656 10444 32696
rect 10484 32656 10485 32696
rect 10443 32647 10485 32656
rect 10732 32537 10772 33664
rect 10731 32528 10773 32537
rect 10731 32488 10732 32528
rect 10772 32488 10773 32528
rect 10731 32479 10773 32488
rect 10635 32360 10677 32369
rect 10635 32320 10636 32360
rect 10676 32320 10677 32360
rect 10635 32311 10677 32320
rect 10252 32276 10292 32285
rect 10292 32236 10580 32276
rect 10252 32227 10292 32236
rect 10540 32192 10580 32236
rect 10540 32143 10580 32152
rect 10636 32192 10676 32311
rect 10636 32117 10676 32152
rect 10635 32108 10677 32117
rect 10635 32068 10636 32108
rect 10676 32068 10677 32108
rect 10635 32059 10677 32068
rect 10635 31772 10677 31781
rect 10635 31732 10636 31772
rect 10676 31732 10677 31772
rect 10635 31723 10677 31732
rect 10155 31436 10197 31445
rect 10155 31396 10156 31436
rect 10196 31396 10197 31436
rect 10155 31387 10197 31396
rect 10060 31303 10100 31312
rect 9963 31268 10005 31277
rect 9963 31228 9964 31268
rect 10004 31228 10005 31268
rect 9963 31219 10005 31228
rect 10443 31268 10485 31277
rect 10443 31228 10444 31268
rect 10484 31228 10485 31268
rect 10443 31219 10485 31228
rect 9868 31184 9908 31193
rect 9868 31100 9908 31144
rect 9868 31060 10100 31100
rect 9868 30857 9908 30942
rect 9867 30848 9909 30857
rect 9867 30808 9868 30848
rect 9908 30808 9909 30848
rect 9867 30799 9909 30808
rect 10060 30689 10100 31060
rect 9868 30680 9908 30689
rect 9772 30640 9868 30680
rect 9675 30631 9717 30640
rect 9868 30631 9908 30640
rect 9964 30680 10004 30689
rect 10060 30680 10105 30689
rect 10060 30640 10065 30680
rect 9676 30546 9716 30631
rect 9483 30176 9525 30185
rect 9483 30136 9484 30176
rect 9524 30136 9525 30176
rect 9483 30127 9525 30136
rect 9964 30101 10004 30640
rect 10065 30631 10105 30640
rect 10444 30680 10484 31219
rect 10444 30521 10484 30640
rect 10443 30512 10485 30521
rect 10443 30472 10444 30512
rect 10484 30472 10485 30512
rect 10443 30463 10485 30472
rect 10155 30428 10197 30437
rect 10155 30388 10156 30428
rect 10196 30388 10197 30428
rect 10155 30379 10197 30388
rect 9099 30092 9141 30101
rect 9099 30052 9100 30092
rect 9140 30052 9141 30092
rect 9099 30043 9141 30052
rect 9963 30092 10005 30101
rect 9963 30052 9964 30092
rect 10004 30052 10005 30092
rect 9963 30043 10005 30052
rect 9004 29681 9044 29766
rect 8715 29632 8716 29672
rect 8756 29632 8757 29672
rect 8715 29623 8757 29632
rect 8812 29632 8948 29672
rect 9003 29672 9045 29681
rect 9003 29632 9004 29672
rect 9044 29632 9045 29672
rect 8715 29336 8757 29345
rect 8715 29296 8716 29336
rect 8756 29296 8757 29336
rect 8715 29287 8757 29296
rect 8812 29336 8852 29632
rect 9003 29623 9045 29632
rect 9100 29504 9140 30043
rect 9292 29968 9716 30008
rect 9195 29672 9237 29681
rect 9195 29632 9196 29672
rect 9236 29632 9237 29672
rect 9195 29623 9237 29632
rect 8812 29287 8852 29296
rect 9004 29464 9140 29504
rect 8235 29168 8277 29177
rect 8235 29128 8236 29168
rect 8276 29128 8277 29168
rect 8235 29119 8277 29128
rect 8523 29168 8565 29177
rect 8523 29128 8524 29168
rect 8564 29128 8565 29168
rect 8523 29119 8565 29128
rect 8620 29168 8660 29177
rect 8620 29000 8660 29128
rect 8236 28960 8660 29000
rect 8716 29168 8756 29287
rect 8908 29177 8948 29262
rect 8716 29000 8756 29128
rect 8907 29168 8949 29177
rect 8907 29128 8908 29168
rect 8948 29128 8949 29168
rect 8907 29119 8949 29128
rect 8716 28960 8948 29000
rect 8140 28328 8180 28337
rect 8044 28288 8140 28328
rect 8044 27833 8084 28288
rect 8140 28279 8180 28288
rect 8139 27992 8181 28001
rect 8139 27952 8140 27992
rect 8180 27952 8181 27992
rect 8139 27943 8181 27952
rect 8043 27824 8085 27833
rect 8043 27784 8044 27824
rect 8084 27784 8085 27824
rect 8043 27775 8085 27784
rect 7948 27607 7988 27616
rect 8043 27656 8085 27665
rect 8043 27616 8044 27656
rect 8084 27616 8085 27656
rect 8043 27607 8085 27616
rect 8044 27522 8084 27607
rect 7755 27488 7797 27497
rect 7755 27448 7756 27488
rect 7796 27448 7797 27488
rect 7755 27439 7797 27448
rect 7756 26144 7796 27439
rect 7852 26816 7892 26825
rect 8140 26816 8180 27943
rect 7892 26776 8180 26816
rect 8236 27656 8276 28960
rect 8811 28748 8853 28757
rect 8811 28708 8812 28748
rect 8852 28708 8853 28748
rect 8811 28699 8853 28708
rect 8715 28664 8757 28673
rect 8715 28624 8716 28664
rect 8756 28624 8757 28664
rect 8715 28615 8757 28624
rect 8427 28412 8469 28421
rect 8427 28372 8428 28412
rect 8468 28372 8469 28412
rect 8427 28363 8469 28372
rect 8332 28160 8372 28169
rect 8332 27833 8372 28120
rect 8428 28001 8468 28363
rect 8619 28328 8661 28337
rect 8619 28288 8620 28328
rect 8660 28288 8661 28328
rect 8619 28279 8661 28288
rect 8716 28328 8756 28615
rect 8716 28279 8756 28288
rect 8812 28328 8852 28699
rect 8908 28337 8948 28960
rect 8812 28279 8852 28288
rect 8907 28328 8949 28337
rect 8907 28288 8908 28328
rect 8948 28288 8949 28328
rect 8907 28279 8949 28288
rect 8523 28244 8565 28253
rect 8523 28204 8524 28244
rect 8564 28204 8565 28244
rect 8523 28195 8565 28204
rect 8524 28110 8564 28195
rect 8620 28194 8660 28279
rect 8427 27992 8469 28001
rect 8427 27952 8428 27992
rect 8468 27952 8469 27992
rect 8427 27943 8469 27952
rect 8331 27824 8373 27833
rect 8331 27784 8332 27824
rect 8372 27784 8373 27824
rect 8331 27775 8373 27784
rect 8811 27824 8853 27833
rect 8811 27784 8812 27824
rect 8852 27784 8853 27824
rect 9004 27824 9044 29464
rect 9196 29261 9236 29623
rect 9292 29336 9332 29968
rect 9388 29840 9428 29849
rect 9388 29420 9428 29800
rect 9483 29840 9525 29849
rect 9483 29800 9484 29840
rect 9524 29800 9525 29840
rect 9483 29791 9525 29800
rect 9580 29840 9620 29849
rect 9676 29840 9716 29968
rect 9868 29840 9908 29849
rect 9676 29800 9868 29840
rect 9484 29706 9524 29791
rect 9580 29420 9620 29800
rect 9868 29791 9908 29800
rect 9964 29840 10004 29849
rect 9676 29672 9716 29681
rect 9964 29672 10004 29800
rect 10156 29840 10196 30379
rect 10251 30260 10293 30269
rect 10251 30220 10252 30260
rect 10292 30220 10293 30260
rect 10251 30211 10293 30220
rect 10156 29791 10196 29800
rect 9716 29632 10004 29672
rect 10059 29672 10101 29681
rect 10059 29632 10060 29672
rect 10100 29632 10101 29672
rect 9676 29623 9716 29632
rect 10059 29623 10101 29632
rect 10060 29538 10100 29623
rect 9388 29380 9524 29420
rect 9580 29380 9716 29420
rect 9292 29287 9332 29296
rect 9195 29252 9237 29261
rect 9195 29212 9196 29252
rect 9236 29212 9237 29252
rect 9195 29203 9237 29212
rect 9100 29168 9140 29177
rect 9100 28580 9140 29128
rect 9196 29168 9236 29203
rect 9196 29118 9236 29128
rect 9388 29168 9428 29179
rect 9388 29093 9428 29128
rect 9387 29084 9429 29093
rect 9387 29044 9388 29084
rect 9428 29044 9429 29084
rect 9387 29035 9429 29044
rect 9484 28757 9524 29380
rect 9580 29093 9620 29095
rect 9579 29084 9621 29093
rect 9579 29044 9580 29084
rect 9620 29044 9621 29084
rect 9579 29035 9621 29044
rect 9580 29000 9620 29035
rect 9580 28920 9620 28960
rect 9676 28757 9716 29380
rect 9963 29252 10005 29261
rect 9963 29212 9964 29252
rect 10004 29212 10005 29252
rect 9963 29203 10005 29212
rect 9772 29168 9812 29177
rect 9772 29009 9812 29128
rect 9771 29000 9813 29009
rect 9771 28960 9772 29000
rect 9812 28960 9813 29000
rect 9771 28951 9813 28960
rect 9483 28748 9525 28757
rect 9483 28708 9484 28748
rect 9524 28708 9525 28748
rect 9483 28699 9525 28708
rect 9675 28748 9717 28757
rect 9675 28708 9676 28748
rect 9716 28708 9717 28748
rect 9675 28699 9717 28708
rect 9867 28664 9909 28673
rect 9867 28624 9868 28664
rect 9908 28624 9909 28664
rect 9867 28615 9909 28624
rect 9772 28580 9812 28589
rect 9100 28540 9772 28580
rect 9772 28531 9812 28540
rect 9387 28412 9429 28421
rect 9387 28372 9388 28412
rect 9428 28372 9429 28412
rect 9387 28363 9429 28372
rect 9099 28328 9141 28337
rect 9099 28288 9100 28328
rect 9140 28288 9141 28328
rect 9099 28279 9141 28288
rect 9388 28328 9428 28363
rect 9868 28337 9908 28615
rect 9100 28076 9140 28279
rect 9388 28277 9428 28288
rect 9483 28328 9525 28337
rect 9483 28288 9484 28328
rect 9524 28288 9525 28328
rect 9483 28279 9525 28288
rect 9867 28328 9909 28337
rect 9867 28288 9868 28328
rect 9908 28288 9909 28328
rect 9867 28279 9909 28288
rect 9964 28328 10004 29203
rect 10155 29000 10197 29009
rect 10155 28960 10156 29000
rect 10196 28960 10197 29000
rect 10155 28951 10197 28960
rect 9964 28279 10004 28288
rect 10060 28328 10100 28337
rect 9484 28194 9524 28279
rect 9100 28036 9812 28076
rect 9676 27824 9716 27833
rect 9004 27784 9140 27824
rect 8811 27775 8853 27784
rect 7852 26321 7892 26776
rect 7851 26312 7893 26321
rect 7851 26272 7852 26312
rect 7892 26272 7893 26312
rect 7851 26263 7893 26272
rect 7659 25220 7701 25229
rect 7659 25180 7660 25220
rect 7700 25180 7701 25220
rect 7659 25171 7701 25180
rect 7756 24053 7796 26104
rect 7851 26144 7893 26153
rect 7851 26104 7852 26144
rect 7892 26104 7893 26144
rect 7851 26095 7893 26104
rect 8044 26144 8084 26153
rect 7852 26010 7892 26095
rect 7852 25892 7892 25901
rect 7892 25852 7988 25892
rect 7852 25843 7892 25852
rect 7852 25304 7892 25313
rect 7755 24044 7797 24053
rect 7755 24004 7756 24044
rect 7796 24004 7797 24044
rect 7755 23995 7797 24004
rect 7852 23549 7892 25264
rect 7851 23540 7893 23549
rect 7851 23500 7852 23540
rect 7892 23500 7893 23540
rect 7851 23491 7893 23500
rect 7948 23288 7988 25852
rect 8044 25556 8084 26104
rect 8236 26060 8276 27616
rect 8332 27656 8372 27775
rect 8524 27665 8564 27750
rect 8332 26830 8372 27616
rect 8523 27656 8565 27665
rect 8523 27616 8524 27656
rect 8564 27616 8565 27656
rect 8523 27607 8565 27616
rect 8812 27656 8852 27775
rect 8907 27740 8949 27749
rect 8907 27700 8908 27740
rect 8948 27700 8949 27740
rect 8907 27691 8949 27700
rect 8812 27607 8852 27616
rect 8908 27656 8948 27691
rect 8908 27605 8948 27616
rect 9004 27656 9044 27665
rect 9004 27581 9044 27616
rect 8427 27572 8469 27581
rect 8427 27532 8428 27572
rect 8468 27532 8469 27572
rect 8427 27523 8469 27532
rect 9003 27572 9045 27581
rect 9003 27532 9004 27572
rect 9044 27532 9045 27572
rect 9003 27523 9045 27532
rect 8332 26781 8372 26790
rect 8428 26321 8468 27523
rect 8523 27488 8565 27497
rect 8523 27448 8524 27488
rect 8564 27448 8565 27488
rect 8523 27439 8565 27448
rect 8524 27354 8564 27439
rect 8619 27236 8661 27245
rect 8619 27196 8620 27236
rect 8660 27196 8661 27236
rect 8619 27187 8661 27196
rect 8524 26648 8564 26657
rect 8427 26312 8469 26321
rect 8427 26272 8428 26312
rect 8468 26272 8469 26312
rect 8427 26263 8469 26272
rect 8428 26153 8468 26263
rect 8427 26144 8469 26153
rect 8427 26104 8428 26144
rect 8468 26104 8469 26144
rect 8427 26095 8469 26104
rect 8236 26020 8372 26060
rect 8332 25976 8372 26020
rect 8332 25936 8468 25976
rect 8236 25892 8276 25903
rect 8236 25817 8276 25852
rect 8235 25808 8277 25817
rect 8235 25768 8236 25808
rect 8276 25768 8277 25808
rect 8235 25759 8277 25768
rect 8044 25507 8084 25516
rect 8332 25304 8372 25313
rect 8044 25136 8084 25145
rect 8332 25136 8372 25264
rect 8084 25096 8372 25136
rect 8044 25087 8084 25096
rect 8235 24968 8277 24977
rect 8235 24928 8236 24968
rect 8276 24928 8277 24968
rect 8235 24919 8277 24928
rect 8140 24632 8180 24641
rect 8140 24389 8180 24592
rect 8139 24380 8181 24389
rect 8139 24340 8140 24380
rect 8180 24340 8181 24380
rect 8139 24331 8181 24340
rect 8140 24221 8180 24331
rect 8139 24212 8181 24221
rect 8139 24172 8140 24212
rect 8180 24172 8181 24212
rect 8139 24163 8181 24172
rect 8140 23792 8180 23801
rect 8140 23549 8180 23752
rect 8139 23540 8181 23549
rect 8139 23500 8140 23540
rect 8180 23500 8181 23540
rect 8139 23491 8181 23500
rect 7948 23248 8084 23288
rect 8044 23129 8084 23248
rect 7948 23120 7988 23129
rect 7564 22576 7892 22616
rect 7659 22448 7701 22457
rect 7659 22408 7660 22448
rect 7700 22408 7701 22448
rect 7659 22399 7701 22408
rect 7564 22289 7604 22374
rect 7563 22280 7605 22289
rect 7563 22240 7564 22280
rect 7604 22240 7605 22280
rect 7563 22231 7605 22240
rect 7563 22112 7605 22121
rect 7563 22072 7564 22112
rect 7604 22072 7605 22112
rect 7563 22063 7605 22072
rect 7564 20768 7604 22063
rect 7564 20719 7604 20728
rect 7660 20180 7700 22399
rect 7852 22028 7892 22576
rect 7948 22205 7988 23080
rect 8043 23120 8085 23129
rect 8043 23080 8044 23120
rect 8084 23080 8085 23120
rect 8043 23071 8085 23080
rect 8140 22868 8180 22877
rect 8044 22828 8140 22868
rect 8044 22294 8084 22828
rect 8140 22819 8180 22828
rect 8236 22373 8276 24919
rect 8332 24641 8372 25096
rect 8331 24632 8373 24641
rect 8331 24592 8332 24632
rect 8372 24592 8373 24632
rect 8331 24583 8373 24592
rect 8332 23960 8372 23971
rect 8332 23885 8372 23920
rect 8331 23876 8373 23885
rect 8331 23836 8332 23876
rect 8372 23836 8373 23876
rect 8331 23827 8373 23836
rect 8332 23045 8372 23827
rect 8331 23036 8373 23045
rect 8331 22996 8332 23036
rect 8372 22996 8373 23036
rect 8331 22987 8373 22996
rect 8428 22952 8468 25936
rect 8524 24809 8564 26608
rect 8620 25472 8660 27187
rect 8811 27068 8853 27077
rect 8811 27028 8812 27068
rect 8852 27028 8853 27068
rect 8811 27019 8853 27028
rect 8812 26934 8852 27019
rect 8715 26816 8757 26825
rect 9004 26816 9044 27523
rect 9100 27077 9140 27784
rect 9387 27740 9429 27749
rect 9387 27700 9388 27740
rect 9428 27700 9429 27740
rect 9387 27691 9429 27700
rect 9388 27656 9428 27691
rect 9388 27605 9428 27616
rect 9484 27656 9524 27665
rect 9484 27497 9524 27616
rect 9483 27488 9525 27497
rect 9483 27448 9484 27488
rect 9524 27448 9525 27488
rect 9483 27439 9525 27448
rect 9196 27404 9236 27413
rect 9099 27068 9141 27077
rect 9099 27028 9100 27068
rect 9140 27028 9141 27068
rect 9099 27019 9141 27028
rect 8715 26776 8716 26816
rect 8756 26776 8757 26816
rect 8715 26767 8757 26776
rect 8908 26776 9044 26816
rect 9100 26816 9140 26825
rect 9196 26816 9236 27364
rect 9676 27320 9716 27784
rect 9772 27656 9812 28036
rect 9868 27824 9908 28279
rect 10060 28169 10100 28288
rect 10156 28328 10196 28951
rect 10156 28279 10196 28288
rect 10252 28328 10292 30211
rect 10444 29849 10484 29935
rect 10636 29849 10676 31723
rect 10828 30092 10868 30101
rect 10924 30092 10964 34495
rect 11020 34469 11060 35335
rect 11116 35048 11156 35503
rect 11212 35225 11252 35310
rect 11211 35216 11253 35225
rect 11211 35176 11212 35216
rect 11252 35176 11253 35216
rect 11211 35167 11253 35176
rect 11308 35132 11348 35848
rect 11404 35720 11444 35729
rect 11404 35216 11444 35680
rect 11596 35393 11636 35848
rect 11595 35384 11637 35393
rect 11595 35344 11596 35384
rect 11636 35344 11637 35384
rect 11595 35335 11637 35344
rect 11500 35216 11540 35225
rect 11404 35176 11500 35216
rect 11500 35167 11540 35176
rect 11595 35216 11637 35225
rect 11595 35176 11596 35216
rect 11636 35176 11637 35216
rect 11595 35167 11637 35176
rect 11308 35092 11444 35132
rect 11404 35048 11444 35092
rect 11596 35082 11636 35167
rect 11116 35008 11348 35048
rect 11404 35008 11540 35048
rect 11019 34460 11061 34469
rect 11019 34420 11020 34460
rect 11060 34420 11061 34460
rect 11019 34411 11061 34420
rect 11020 33797 11060 34411
rect 11019 33788 11061 33797
rect 11019 33748 11020 33788
rect 11060 33748 11061 33788
rect 11019 33739 11061 33748
rect 11116 33620 11156 33629
rect 11116 33461 11156 33580
rect 11211 33620 11253 33629
rect 11211 33580 11212 33620
rect 11252 33580 11253 33620
rect 11211 33571 11253 33580
rect 11212 33486 11252 33571
rect 11115 33452 11157 33461
rect 11115 33412 11116 33452
rect 11156 33412 11157 33452
rect 11115 33403 11157 33412
rect 11308 33368 11348 35008
rect 11212 33328 11348 33368
rect 11019 32780 11061 32789
rect 11019 32740 11020 32780
rect 11060 32740 11061 32780
rect 11019 32731 11061 32740
rect 11020 32192 11060 32731
rect 11020 32143 11060 32152
rect 11116 32108 11156 32117
rect 11116 31193 11156 32068
rect 11115 31184 11157 31193
rect 11115 31144 11116 31184
rect 11156 31144 11157 31184
rect 11115 31135 11157 31144
rect 11019 30176 11061 30185
rect 11019 30136 11020 30176
rect 11060 30136 11061 30176
rect 11019 30127 11061 30136
rect 10868 30052 10964 30092
rect 10828 30043 10868 30052
rect 11020 30008 11060 30127
rect 11020 29959 11060 29968
rect 10348 29840 10388 29849
rect 10348 29345 10388 29800
rect 10443 29848 10485 29849
rect 10443 29800 10444 29848
rect 10484 29800 10485 29848
rect 10443 29791 10485 29800
rect 10540 29840 10580 29849
rect 10443 29672 10485 29681
rect 10443 29632 10444 29672
rect 10484 29632 10485 29672
rect 10443 29623 10485 29632
rect 10347 29336 10389 29345
rect 10347 29296 10348 29336
rect 10388 29296 10389 29336
rect 10347 29287 10389 29296
rect 10444 29168 10484 29623
rect 10540 29261 10580 29800
rect 10635 29840 10677 29849
rect 11020 29840 11060 29849
rect 10635 29800 10636 29840
rect 10676 29800 10677 29840
rect 10635 29791 10677 29800
rect 10828 29800 11020 29840
rect 10636 29672 10676 29681
rect 10539 29252 10581 29261
rect 10539 29212 10540 29252
rect 10580 29212 10581 29252
rect 10539 29203 10581 29212
rect 10252 28279 10292 28288
rect 10348 29128 10484 29168
rect 10059 28160 10101 28169
rect 10059 28120 10060 28160
rect 10100 28120 10101 28160
rect 10059 28111 10101 28120
rect 9868 27775 9908 27784
rect 10059 27740 10101 27749
rect 10059 27700 10060 27740
rect 10100 27700 10101 27740
rect 10059 27691 10101 27700
rect 9964 27656 10004 27665
rect 9772 27616 9964 27656
rect 9964 27607 10004 27616
rect 9867 27488 9909 27497
rect 9867 27448 9868 27488
rect 9908 27448 9909 27488
rect 9867 27439 9909 27448
rect 9676 27280 9812 27320
rect 9292 26984 9332 26993
rect 9332 26944 9716 26984
rect 9292 26935 9332 26944
rect 9140 26776 9236 26816
rect 9484 26816 9524 26825
rect 8716 26682 8756 26767
rect 8811 25976 8853 25985
rect 8811 25936 8812 25976
rect 8852 25936 8853 25976
rect 8811 25927 8853 25936
rect 8812 25565 8852 25927
rect 8811 25556 8853 25565
rect 8811 25516 8812 25556
rect 8852 25516 8853 25556
rect 8811 25507 8853 25516
rect 8620 25432 8756 25472
rect 8620 25304 8660 25315
rect 8620 25229 8660 25264
rect 8716 25304 8756 25432
rect 8908 25304 8948 26776
rect 9100 26767 9140 26776
rect 9004 26648 9044 26657
rect 9004 25817 9044 26608
rect 9003 25808 9045 25817
rect 9003 25768 9004 25808
rect 9044 25768 9045 25808
rect 9003 25759 9045 25768
rect 9484 25640 9524 26776
rect 9676 26816 9716 26944
rect 9676 26767 9716 26776
rect 9772 26816 9812 27280
rect 9772 26767 9812 26776
rect 9579 26648 9621 26657
rect 9579 26608 9580 26648
rect 9620 26608 9621 26648
rect 9579 26599 9621 26608
rect 9580 26514 9620 26599
rect 9868 26573 9908 27439
rect 9963 26816 10005 26825
rect 9963 26776 9964 26816
rect 10004 26776 10005 26816
rect 9963 26767 10005 26776
rect 9964 26682 10004 26767
rect 9867 26564 9909 26573
rect 9867 26524 9868 26564
rect 9908 26524 9909 26564
rect 9867 26515 9909 26524
rect 10060 26153 10100 27691
rect 10156 27656 10196 27665
rect 10348 27656 10388 29128
rect 10540 29000 10580 29203
rect 10636 29177 10676 29632
rect 10635 29168 10677 29177
rect 10635 29128 10636 29168
rect 10676 29128 10677 29168
rect 10635 29119 10677 29128
rect 10828 29009 10868 29800
rect 11020 29791 11060 29800
rect 11019 29672 11061 29681
rect 11019 29632 11020 29672
rect 11060 29632 11061 29672
rect 11019 29623 11061 29632
rect 11020 29168 11060 29623
rect 11212 29177 11252 33328
rect 11307 32444 11349 32453
rect 11307 32404 11308 32444
rect 11348 32404 11349 32444
rect 11307 32395 11349 32404
rect 11308 32285 11348 32395
rect 11307 32276 11349 32285
rect 11307 32236 11308 32276
rect 11348 32236 11349 32276
rect 11307 32227 11349 32236
rect 11500 32201 11540 35008
rect 11595 33872 11637 33881
rect 11595 33832 11596 33872
rect 11636 33832 11637 33872
rect 11595 33823 11637 33832
rect 11596 33545 11636 33823
rect 11692 33713 11732 36856
rect 11788 36728 11828 36739
rect 11788 36653 11828 36688
rect 11787 36644 11829 36653
rect 11787 36604 11788 36644
rect 11828 36604 11829 36644
rect 11787 36595 11829 36604
rect 11884 35897 11924 38611
rect 11980 38501 12020 38779
rect 11979 38492 12021 38501
rect 11979 38452 11980 38492
rect 12020 38452 12021 38492
rect 11979 38443 12021 38452
rect 11979 38156 12021 38165
rect 11979 38116 11980 38156
rect 12020 38116 12021 38156
rect 11979 38107 12021 38116
rect 11980 37400 12020 38107
rect 12076 37745 12116 39376
rect 12364 38926 12404 40132
rect 12556 39752 12596 41299
rect 12652 40349 12692 41383
rect 12748 40424 12788 42928
rect 12940 40844 12980 42928
rect 13132 41693 13172 42928
rect 13131 41684 13173 41693
rect 13131 41644 13132 41684
rect 13172 41644 13173 41684
rect 13131 41635 13173 41644
rect 13324 41609 13364 42928
rect 13323 41600 13365 41609
rect 13323 41560 13324 41600
rect 13364 41560 13365 41600
rect 13323 41551 13365 41560
rect 13516 41525 13556 42928
rect 13708 41945 13748 42928
rect 13707 41936 13749 41945
rect 13707 41896 13708 41936
rect 13748 41896 13749 41936
rect 13707 41887 13749 41896
rect 13515 41516 13557 41525
rect 13515 41476 13516 41516
rect 13556 41476 13557 41516
rect 13515 41467 13557 41476
rect 13900 41441 13940 42928
rect 14092 41777 14132 42928
rect 14284 42365 14324 42928
rect 14379 42440 14421 42449
rect 14379 42400 14380 42440
rect 14420 42400 14421 42440
rect 14379 42391 14421 42400
rect 14283 42356 14325 42365
rect 14283 42316 14284 42356
rect 14324 42316 14325 42356
rect 14283 42307 14325 42316
rect 14091 41768 14133 41777
rect 14091 41728 14092 41768
rect 14132 41728 14133 41768
rect 14091 41719 14133 41728
rect 13899 41432 13941 41441
rect 13899 41392 13900 41432
rect 13940 41392 13941 41432
rect 13899 41383 13941 41392
rect 13707 41264 13749 41273
rect 13707 41224 13708 41264
rect 13748 41224 13749 41264
rect 13707 41215 13749 41224
rect 14092 41264 14132 41273
rect 14132 41224 14228 41264
rect 14092 41215 14132 41224
rect 13708 41130 13748 41215
rect 14188 41105 14228 41224
rect 14187 41096 14229 41105
rect 14187 41056 14188 41096
rect 14228 41056 14229 41096
rect 14187 41047 14229 41056
rect 13899 41012 13941 41021
rect 13899 40972 13900 41012
rect 13940 40972 13941 41012
rect 13899 40963 13941 40972
rect 13900 40878 13940 40963
rect 12940 40804 13172 40844
rect 13035 40676 13077 40685
rect 13035 40636 13036 40676
rect 13076 40636 13077 40676
rect 13035 40627 13077 40636
rect 12748 40384 12884 40424
rect 12651 40340 12693 40349
rect 12651 40300 12652 40340
rect 12692 40300 12693 40340
rect 12651 40291 12693 40300
rect 12556 39703 12596 39712
rect 12555 39584 12597 39593
rect 12555 39544 12556 39584
rect 12596 39544 12597 39584
rect 12555 39535 12597 39544
rect 12171 38912 12213 38921
rect 12171 38872 12172 38912
rect 12212 38872 12213 38912
rect 12556 38912 12596 39535
rect 12748 39500 12788 39509
rect 12364 38877 12404 38886
rect 12171 38863 12213 38872
rect 12460 38872 12596 38912
rect 12652 39460 12748 39500
rect 12172 38501 12212 38863
rect 12171 38492 12213 38501
rect 12171 38452 12172 38492
rect 12212 38452 12213 38492
rect 12171 38443 12213 38452
rect 12172 38240 12212 38443
rect 12172 38191 12212 38200
rect 12075 37736 12117 37745
rect 12075 37696 12076 37736
rect 12116 37696 12117 37736
rect 12075 37687 12117 37696
rect 12075 37568 12117 37577
rect 12075 37528 12076 37568
rect 12116 37528 12117 37568
rect 12075 37519 12117 37528
rect 11883 35888 11925 35897
rect 11883 35848 11884 35888
rect 11924 35848 11925 35888
rect 11883 35839 11925 35848
rect 11980 35132 12020 37360
rect 11787 34544 11829 34553
rect 11787 34504 11788 34544
rect 11828 34504 11829 34544
rect 11787 34495 11829 34504
rect 11691 33704 11733 33713
rect 11691 33664 11692 33704
rect 11732 33664 11733 33704
rect 11691 33655 11733 33664
rect 11595 33536 11637 33545
rect 11595 33496 11596 33536
rect 11636 33496 11732 33536
rect 11595 33487 11637 33496
rect 11595 33368 11637 33377
rect 11595 33328 11596 33368
rect 11636 33328 11637 33368
rect 11595 33319 11637 33328
rect 11499 32192 11541 32201
rect 11499 32152 11500 32192
rect 11540 32152 11541 32192
rect 11499 32143 11541 32152
rect 11596 32192 11636 33319
rect 11596 31781 11636 32152
rect 11595 31772 11637 31781
rect 11595 31732 11596 31772
rect 11636 31732 11637 31772
rect 11595 31723 11637 31732
rect 11692 31697 11732 33496
rect 11307 31688 11349 31697
rect 11307 31648 11308 31688
rect 11348 31648 11349 31688
rect 11307 31639 11349 31648
rect 11691 31688 11733 31697
rect 11691 31648 11692 31688
rect 11732 31648 11733 31688
rect 11691 31639 11733 31648
rect 11308 31445 11348 31639
rect 11595 31520 11637 31529
rect 11595 31480 11596 31520
rect 11636 31480 11637 31520
rect 11595 31471 11637 31480
rect 11307 31436 11349 31445
rect 11307 31396 11308 31436
rect 11348 31396 11349 31436
rect 11307 31387 11349 31396
rect 11308 31352 11348 31387
rect 11308 31301 11348 31312
rect 11500 31184 11540 31193
rect 11403 30512 11445 30521
rect 11403 30472 11404 30512
rect 11444 30472 11445 30512
rect 11403 30463 11445 30472
rect 11307 30344 11349 30353
rect 11307 30304 11308 30344
rect 11348 30304 11349 30344
rect 11307 30295 11349 30304
rect 11308 29261 11348 30295
rect 11404 29756 11444 30463
rect 11500 29840 11540 31144
rect 11596 30680 11636 31471
rect 11691 31352 11733 31361
rect 11691 31312 11692 31352
rect 11732 31312 11733 31352
rect 11691 31303 11733 31312
rect 11692 31109 11732 31303
rect 11691 31100 11733 31109
rect 11691 31060 11692 31100
rect 11732 31060 11733 31100
rect 11691 31051 11733 31060
rect 11692 30680 11732 30689
rect 11596 30640 11692 30680
rect 11596 30521 11636 30640
rect 11692 30631 11732 30640
rect 11595 30512 11637 30521
rect 11595 30472 11596 30512
rect 11636 30472 11637 30512
rect 11595 30463 11637 30472
rect 11691 30008 11733 30017
rect 11691 29968 11692 30008
rect 11732 29968 11733 30008
rect 11691 29959 11733 29968
rect 11596 29840 11636 29849
rect 11500 29800 11596 29840
rect 11596 29791 11636 29800
rect 11692 29840 11732 29959
rect 11404 29716 11540 29756
rect 11307 29252 11349 29261
rect 11307 29212 11308 29252
rect 11348 29212 11349 29252
rect 11307 29203 11349 29212
rect 11020 29119 11060 29128
rect 11211 29168 11253 29177
rect 11211 29128 11212 29168
rect 11252 29128 11253 29168
rect 11211 29119 11253 29128
rect 11212 29034 11252 29119
rect 10827 29000 10869 29009
rect 10540 28960 10676 29000
rect 10539 28580 10581 28589
rect 10539 28540 10540 28580
rect 10580 28540 10581 28580
rect 10539 28531 10581 28540
rect 10443 28328 10485 28337
rect 10443 28288 10444 28328
rect 10484 28288 10485 28328
rect 10443 28279 10485 28288
rect 10540 28328 10580 28531
rect 10636 28328 10676 28960
rect 10827 28960 10828 29000
rect 10868 28960 10869 29000
rect 10827 28951 10869 28960
rect 10827 28832 10869 28841
rect 10827 28792 10828 28832
rect 10868 28792 10869 28832
rect 10827 28783 10869 28792
rect 10731 28748 10773 28757
rect 10731 28708 10732 28748
rect 10772 28708 10773 28748
rect 10731 28699 10773 28708
rect 10732 28580 10772 28699
rect 10732 28531 10772 28540
rect 10732 28328 10772 28337
rect 10636 28288 10732 28328
rect 10540 28279 10580 28288
rect 10732 28279 10772 28288
rect 10444 28194 10484 28279
rect 10828 28160 10868 28783
rect 10923 28496 10965 28505
rect 10923 28456 10924 28496
rect 10964 28456 10965 28496
rect 10923 28447 10965 28456
rect 10924 28341 10964 28447
rect 10924 28292 10964 28301
rect 11116 28328 11156 28337
rect 10196 27616 10388 27656
rect 10732 28120 10868 28160
rect 11020 28160 11060 28169
rect 9676 26144 9716 26153
rect 9676 25985 9716 26104
rect 9867 26144 9909 26153
rect 9867 26104 9868 26144
rect 9908 26104 9909 26144
rect 9867 26095 9909 26104
rect 10059 26144 10101 26153
rect 10059 26104 10060 26144
rect 10100 26104 10101 26144
rect 10059 26095 10101 26104
rect 9868 25985 9908 26095
rect 9675 25976 9717 25985
rect 9675 25936 9676 25976
rect 9716 25936 9717 25976
rect 9675 25927 9717 25936
rect 9867 25976 9909 25985
rect 9867 25936 9868 25976
rect 9908 25936 9909 25976
rect 9867 25927 9909 25936
rect 9484 25600 9812 25640
rect 9004 25472 9044 25481
rect 9388 25472 9428 25481
rect 9044 25432 9332 25472
rect 9004 25423 9044 25432
rect 9292 25388 9332 25432
rect 9292 25339 9332 25348
rect 9196 25304 9236 25313
rect 8908 25264 9140 25304
rect 8619 25220 8661 25229
rect 8619 25180 8620 25220
rect 8660 25180 8661 25220
rect 8619 25171 8661 25180
rect 8619 24968 8661 24977
rect 8619 24928 8620 24968
rect 8660 24928 8661 24968
rect 8619 24919 8661 24928
rect 8523 24800 8565 24809
rect 8523 24760 8524 24800
rect 8564 24760 8565 24800
rect 8523 24751 8565 24760
rect 8523 24632 8565 24641
rect 8523 24592 8524 24632
rect 8564 24592 8565 24632
rect 8523 24583 8565 24592
rect 8524 23792 8564 24583
rect 8524 23743 8564 23752
rect 8524 23129 8564 23214
rect 8523 23120 8565 23129
rect 8523 23080 8524 23120
rect 8564 23080 8565 23120
rect 8523 23071 8565 23080
rect 8620 23036 8660 24919
rect 8716 24809 8756 25264
rect 8715 24800 8757 24809
rect 8715 24760 8716 24800
rect 8756 24760 8757 24800
rect 8715 24751 8757 24760
rect 8812 24632 8852 24641
rect 8716 24592 8812 24632
rect 8716 24221 8756 24592
rect 8812 24583 8852 24592
rect 8908 24632 8948 24641
rect 8908 24305 8948 24592
rect 9003 24632 9045 24641
rect 9003 24592 9004 24632
rect 9044 24592 9045 24632
rect 9003 24583 9045 24592
rect 8907 24296 8949 24305
rect 8907 24256 8908 24296
rect 8948 24256 8949 24296
rect 8907 24247 8949 24256
rect 8715 24212 8757 24221
rect 8715 24172 8716 24212
rect 8756 24172 8757 24212
rect 8715 24163 8757 24172
rect 9004 24128 9044 24583
rect 8812 24088 9044 24128
rect 8716 23969 8756 24054
rect 8715 23960 8757 23969
rect 8715 23920 8716 23960
rect 8756 23920 8757 23960
rect 8715 23911 8757 23920
rect 8715 23792 8757 23801
rect 8715 23752 8716 23792
rect 8756 23752 8757 23792
rect 8715 23743 8757 23752
rect 8716 23633 8756 23743
rect 8812 23708 8852 24088
rect 8908 23960 8948 23969
rect 8948 23920 9044 23960
rect 8908 23911 8948 23920
rect 8812 23668 8948 23708
rect 8715 23624 8757 23633
rect 8715 23584 8716 23624
rect 8756 23584 8757 23624
rect 8715 23575 8757 23584
rect 8812 23045 8852 23130
rect 8908 23120 8948 23668
rect 8908 23071 8948 23080
rect 8620 22987 8660 22996
rect 8811 23036 8853 23045
rect 8811 22996 8812 23036
rect 8852 22996 8853 23036
rect 8811 22987 8853 22996
rect 8715 22952 8757 22961
rect 8428 22912 8564 22952
rect 8331 22868 8373 22877
rect 8331 22828 8332 22868
rect 8372 22828 8373 22868
rect 8331 22819 8373 22828
rect 8235 22364 8277 22373
rect 8235 22324 8236 22364
rect 8276 22324 8277 22364
rect 8235 22315 8277 22324
rect 8044 22245 8084 22254
rect 7947 22196 7989 22205
rect 7947 22156 7948 22196
rect 7988 22156 7989 22196
rect 7947 22147 7989 22156
rect 8235 22112 8277 22121
rect 8235 22072 8236 22112
rect 8276 22072 8277 22112
rect 8235 22063 8277 22072
rect 7852 21988 8180 22028
rect 8044 21692 8084 21701
rect 7852 21594 7892 21603
rect 7756 21020 7796 21029
rect 7852 21020 7892 21554
rect 8044 21533 8084 21652
rect 8043 21524 8085 21533
rect 8043 21484 8044 21524
rect 8084 21484 8085 21524
rect 8043 21475 8085 21484
rect 7796 20980 7892 21020
rect 7756 20971 7796 20980
rect 8044 20180 8084 20220
rect 7660 20140 7796 20180
rect 7659 19760 7701 19769
rect 7659 19720 7660 19760
rect 7700 19720 7701 19760
rect 7659 19711 7701 19720
rect 7372 19384 7508 19424
rect 7660 19424 7700 19711
rect 7275 19088 7317 19097
rect 7275 19048 7276 19088
rect 7316 19048 7317 19088
rect 7275 19039 7317 19048
rect 7276 18954 7316 19039
rect 7372 18761 7412 19384
rect 7660 19375 7700 19384
rect 7564 19340 7604 19349
rect 7468 19256 7508 19265
rect 7371 18752 7413 18761
rect 7371 18712 7372 18752
rect 7412 18712 7413 18752
rect 7371 18703 7413 18712
rect 6987 18628 6988 18668
rect 7028 18628 7029 18668
rect 6987 18619 7029 18628
rect 7084 18628 7220 18668
rect 6507 17744 6549 17753
rect 6507 17704 6508 17744
rect 6548 17704 6549 17744
rect 6507 17695 6549 17704
rect 6315 17660 6357 17669
rect 6315 17620 6316 17660
rect 6356 17620 6357 17660
rect 6315 17611 6357 17620
rect 5932 17023 5972 17032
rect 6028 17452 6260 17492
rect 6028 17072 6068 17452
rect 6220 17072 6260 17081
rect 6028 17023 6068 17032
rect 6124 17032 6220 17072
rect 5356 16864 5492 16904
rect 5068 16360 5396 16400
rect 4972 16276 5108 16316
rect 4588 16064 4628 16073
rect 4588 15149 4628 16024
rect 4683 16064 4725 16073
rect 4683 16024 4684 16064
rect 4724 16024 4725 16064
rect 4683 16015 4725 16024
rect 4587 15140 4629 15149
rect 4587 15100 4588 15140
rect 4628 15100 4629 15140
rect 4587 15091 4629 15100
rect 4107 14636 4149 14645
rect 4107 14596 4108 14636
rect 4148 14596 4149 14636
rect 4107 14587 4149 14596
rect 4107 14300 4149 14309
rect 4107 14260 4108 14300
rect 4148 14260 4149 14300
rect 4107 14251 4149 14260
rect 3819 14048 3861 14057
rect 3819 14008 3820 14048
rect 3860 14008 3861 14048
rect 3819 13999 3861 14008
rect 3724 13964 3764 13973
rect 3532 13924 3724 13964
rect 3532 13637 3572 13924
rect 3724 13915 3764 13924
rect 3820 13914 3860 13999
rect 3531 13628 3573 13637
rect 3531 13588 3532 13628
rect 3572 13588 3573 13628
rect 3531 13579 3573 13588
rect 3688 13628 4056 13637
rect 3728 13588 3770 13628
rect 3810 13588 3852 13628
rect 3892 13588 3934 13628
rect 3974 13588 4016 13628
rect 3688 13579 4056 13588
rect 3627 13376 3669 13385
rect 3532 13336 3628 13376
rect 3668 13336 3669 13376
rect 3532 13303 3572 13336
rect 3627 13327 3669 13336
rect 3532 13254 3572 13263
rect 3916 13292 3956 13301
rect 3724 13040 3764 13049
rect 3724 12797 3764 13000
rect 3723 12788 3765 12797
rect 3723 12748 3724 12788
rect 3764 12748 3765 12788
rect 3723 12739 3765 12748
rect 3532 12545 3572 12630
rect 3531 12536 3573 12545
rect 3531 12496 3532 12536
rect 3572 12496 3573 12536
rect 3531 12487 3573 12496
rect 3916 12293 3956 13252
rect 4011 12620 4053 12629
rect 4011 12580 4012 12620
rect 4052 12580 4053 12620
rect 4011 12571 4053 12580
rect 4012 12536 4052 12571
rect 4012 12485 4052 12496
rect 4108 12536 4148 14251
rect 4203 14048 4245 14057
rect 4203 14008 4204 14048
rect 4244 14008 4245 14048
rect 4203 13999 4245 14008
rect 4300 14048 4340 14057
rect 4204 13914 4244 13999
rect 4300 13889 4340 14008
rect 4299 13880 4341 13889
rect 4299 13840 4300 13880
rect 4340 13840 4341 13880
rect 4299 13831 4341 13840
rect 4299 13628 4341 13637
rect 4299 13588 4300 13628
rect 4340 13588 4341 13628
rect 4299 13579 4341 13588
rect 4300 13208 4340 13579
rect 4300 13159 4340 13168
rect 4492 13040 4532 14680
rect 4684 14048 4724 16015
rect 4780 15737 4820 16276
rect 5068 16232 5108 16276
rect 4972 16073 5012 16158
rect 4971 16064 5013 16073
rect 4971 16024 4972 16064
rect 5012 16024 5013 16064
rect 5068 16064 5108 16192
rect 5260 16232 5300 16243
rect 5260 16157 5300 16192
rect 5259 16148 5301 16157
rect 5259 16108 5260 16148
rect 5300 16108 5301 16148
rect 5259 16099 5301 16108
rect 5163 16064 5205 16073
rect 5068 16024 5164 16064
rect 5204 16024 5205 16064
rect 4971 16015 5013 16024
rect 5163 16015 5205 16024
rect 4928 15896 5296 15905
rect 4968 15856 5010 15896
rect 5050 15856 5092 15896
rect 5132 15856 5174 15896
rect 5214 15856 5256 15896
rect 4928 15847 5296 15856
rect 4779 15728 4821 15737
rect 4779 15688 4780 15728
rect 4820 15688 4821 15728
rect 4779 15679 4821 15688
rect 5163 15728 5205 15737
rect 5163 15688 5164 15728
rect 5204 15688 5205 15728
rect 5163 15679 5205 15688
rect 4972 14725 5012 14734
rect 4972 14561 5012 14685
rect 5164 14636 5204 15679
rect 5164 14587 5204 14596
rect 4971 14552 5013 14561
rect 4971 14512 4972 14552
rect 5012 14512 5013 14552
rect 4971 14503 5013 14512
rect 4779 14468 4821 14477
rect 4779 14428 4780 14468
rect 4820 14428 4821 14468
rect 4779 14419 4821 14428
rect 4587 13460 4629 13469
rect 4587 13420 4588 13460
rect 4628 13420 4629 13460
rect 4587 13411 4629 13420
rect 4588 13217 4628 13411
rect 4587 13208 4629 13217
rect 4587 13168 4588 13208
rect 4628 13168 4629 13208
rect 4587 13159 4629 13168
rect 3915 12284 3957 12293
rect 3915 12244 3916 12284
rect 3956 12244 3957 12284
rect 3915 12235 3957 12244
rect 3688 12116 4056 12125
rect 3728 12076 3770 12116
rect 3810 12076 3852 12116
rect 3892 12076 3934 12116
rect 3974 12076 4016 12116
rect 3688 12067 4056 12076
rect 3435 11444 3477 11453
rect 3435 11404 3436 11444
rect 3476 11404 3477 11444
rect 3435 11395 3477 11404
rect 3435 11108 3477 11117
rect 3435 11068 3436 11108
rect 3476 11068 3477 11108
rect 3435 11059 3477 11068
rect 3436 11024 3476 11059
rect 3436 10973 3476 10984
rect 3819 11024 3861 11033
rect 3819 10984 3820 11024
rect 3860 10984 3861 11024
rect 3819 10975 3861 10984
rect 3820 10890 3860 10975
rect 3628 10772 3668 10781
rect 3436 10732 3628 10772
rect 2955 9596 2997 9605
rect 2955 9556 2956 9596
rect 2996 9556 2997 9596
rect 2955 9547 2997 9556
rect 3244 9596 3284 9605
rect 2860 9442 2900 9451
rect 2859 9344 2901 9353
rect 2859 9304 2860 9344
rect 2900 9304 2901 9344
rect 2859 9295 2901 9304
rect 2860 8345 2900 9295
rect 2956 8756 2996 9547
rect 3244 8933 3284 9556
rect 3339 9596 3381 9605
rect 3339 9556 3340 9596
rect 3380 9556 3381 9596
rect 3339 9547 3381 9556
rect 3436 9507 3476 10732
rect 3628 10723 3668 10732
rect 3688 10604 4056 10613
rect 3728 10564 3770 10604
rect 3810 10564 3852 10604
rect 3892 10564 3934 10604
rect 3974 10564 4016 10604
rect 3688 10555 4056 10564
rect 3531 10352 3573 10361
rect 3531 10312 3532 10352
rect 3572 10312 3573 10352
rect 3531 10303 3573 10312
rect 3436 9458 3476 9467
rect 3435 9260 3477 9269
rect 3435 9220 3436 9260
rect 3476 9220 3477 9260
rect 3435 9211 3477 9220
rect 3339 9008 3381 9017
rect 3339 8968 3340 9008
rect 3380 8968 3381 9008
rect 3339 8959 3381 8968
rect 3243 8924 3285 8933
rect 3243 8884 3244 8924
rect 3284 8884 3285 8924
rect 3243 8875 3285 8884
rect 2956 8513 2996 8716
rect 3052 8672 3092 8681
rect 2955 8504 2997 8513
rect 2955 8464 2956 8504
rect 2996 8464 2997 8504
rect 2955 8455 2997 8464
rect 3052 8345 3092 8632
rect 3147 8672 3189 8681
rect 3147 8632 3148 8672
rect 3188 8632 3189 8672
rect 3147 8623 3189 8632
rect 2859 8336 2901 8345
rect 2859 8296 2860 8336
rect 2900 8296 2901 8336
rect 2859 8287 2901 8296
rect 3051 8336 3093 8345
rect 3051 8296 3052 8336
rect 3092 8296 3093 8336
rect 3051 8287 3093 8296
rect 2763 8168 2805 8177
rect 2763 8128 2764 8168
rect 2804 8128 2805 8168
rect 2763 8119 2805 8128
rect 3051 8168 3093 8177
rect 3051 8128 3052 8168
rect 3092 8128 3093 8168
rect 3051 8119 3093 8128
rect 3052 8034 3092 8119
rect 2955 8000 2997 8009
rect 2860 7979 2956 8000
rect 2900 7960 2956 7979
rect 2996 7960 2997 8000
rect 2955 7951 2997 7960
rect 2860 7930 2900 7939
rect 2763 7916 2805 7925
rect 2763 7876 2764 7916
rect 2804 7876 2805 7916
rect 2763 7867 2805 7876
rect 2764 7412 2804 7867
rect 2764 7363 2804 7372
rect 3052 7160 3092 7169
rect 2956 7120 3052 7160
rect 2859 6992 2901 7001
rect 2859 6952 2860 6992
rect 2900 6952 2901 6992
rect 2859 6943 2901 6952
rect 2763 6656 2805 6665
rect 2763 6616 2764 6656
rect 2804 6616 2805 6656
rect 2763 6607 2805 6616
rect 2764 6488 2804 6607
rect 2860 6497 2900 6943
rect 2764 6439 2804 6448
rect 2859 6488 2901 6497
rect 2859 6448 2860 6488
rect 2900 6448 2901 6488
rect 2859 6439 2901 6448
rect 2668 6280 2804 6320
rect 2571 6271 2613 6280
rect 2668 5816 2708 5825
rect 2476 5776 2668 5816
rect 2668 5767 2708 5776
rect 2475 5648 2517 5657
rect 2475 5608 2476 5648
rect 2516 5608 2517 5648
rect 2475 5599 2517 5608
rect 2284 4852 2420 4892
rect 2091 4843 2133 4852
rect 2092 4758 2132 4843
rect 2283 4724 2325 4733
rect 2283 4684 2284 4724
rect 2324 4684 2325 4724
rect 2283 4675 2325 4684
rect 2284 4590 2324 4675
rect 2380 4649 2420 4852
rect 2476 4724 2516 5599
rect 2667 5564 2709 5573
rect 2667 5524 2668 5564
rect 2708 5524 2709 5564
rect 2667 5515 2709 5524
rect 2571 5060 2613 5069
rect 2571 5020 2572 5060
rect 2612 5020 2613 5060
rect 2571 5011 2613 5020
rect 2572 4976 2612 5011
rect 2572 4925 2612 4936
rect 2668 4976 2708 5515
rect 2476 4684 2612 4724
rect 2379 4640 2421 4649
rect 2379 4600 2380 4640
rect 2420 4600 2421 4640
rect 2379 4591 2421 4600
rect 2283 4388 2325 4397
rect 2283 4348 2284 4388
rect 2324 4348 2325 4388
rect 2283 4339 2325 4348
rect 1996 3760 2132 3800
rect 1995 3632 2037 3641
rect 1995 3592 1996 3632
rect 2036 3592 2037 3632
rect 1995 3583 2037 3592
rect 1996 3498 2036 3583
rect 1804 3296 1844 3305
rect 1804 2885 1844 3256
rect 1803 2876 1845 2885
rect 1803 2836 1804 2876
rect 1844 2836 1845 2876
rect 1803 2827 1845 2836
rect 2092 2717 2132 3760
rect 2188 3473 2228 3554
rect 2187 3464 2229 3473
rect 2187 3419 2188 3464
rect 2228 3419 2229 3464
rect 2187 3415 2229 3419
rect 2188 3410 2228 3415
rect 2091 2708 2133 2717
rect 2091 2668 2092 2708
rect 2132 2668 2133 2708
rect 2091 2659 2133 2668
rect 1899 2204 1941 2213
rect 1899 2164 1900 2204
rect 1940 2164 1941 2204
rect 1899 2155 1941 2164
rect 1612 1457 1652 1828
rect 1804 1700 1844 1709
rect 1611 1448 1653 1457
rect 1611 1408 1612 1448
rect 1652 1408 1653 1448
rect 1611 1399 1653 1408
rect 1804 1373 1844 1660
rect 1803 1364 1845 1373
rect 1803 1324 1804 1364
rect 1844 1324 1845 1364
rect 1803 1315 1845 1324
rect 1900 1112 1940 2155
rect 1995 1868 2037 1877
rect 1995 1828 1996 1868
rect 2036 1828 2037 1868
rect 1995 1819 2037 1828
rect 1996 1734 2036 1819
rect 2187 1700 2229 1709
rect 2187 1660 2188 1700
rect 2228 1660 2229 1700
rect 2187 1651 2229 1660
rect 2188 1566 2228 1651
rect 2284 1448 2324 4339
rect 2572 4136 2612 4684
rect 2572 3296 2612 4096
rect 2668 3977 2708 4936
rect 2764 4388 2804 6280
rect 2860 5825 2900 6439
rect 2859 5816 2901 5825
rect 2859 5776 2860 5816
rect 2900 5776 2901 5816
rect 2859 5767 2901 5776
rect 2860 5648 2900 5657
rect 2860 5237 2900 5608
rect 2859 5228 2901 5237
rect 2859 5188 2860 5228
rect 2900 5188 2901 5228
rect 2859 5179 2901 5188
rect 2956 4808 2996 7120
rect 3052 7111 3092 7120
rect 3148 7160 3188 8623
rect 3243 8588 3285 8597
rect 3243 8548 3244 8588
rect 3284 8548 3285 8588
rect 3243 8539 3285 8548
rect 3148 7111 3188 7120
rect 3244 6992 3284 8539
rect 3052 6952 3284 6992
rect 3052 5657 3092 6952
rect 3147 5900 3189 5909
rect 3147 5860 3148 5900
rect 3188 5860 3189 5900
rect 3147 5851 3189 5860
rect 3148 5766 3188 5851
rect 3340 5657 3380 8959
rect 3436 8000 3476 9211
rect 3532 8924 3572 10303
rect 4108 9596 4148 12496
rect 4300 13000 4532 13040
rect 4203 12284 4245 12293
rect 4203 12244 4204 12284
rect 4244 12244 4245 12284
rect 4203 12235 4245 12244
rect 4012 9556 4148 9596
rect 3916 9512 3956 9521
rect 3916 9269 3956 9472
rect 4012 9437 4052 9556
rect 4011 9428 4053 9437
rect 4011 9388 4012 9428
rect 4052 9388 4053 9428
rect 4011 9379 4053 9388
rect 4107 9344 4149 9353
rect 4107 9304 4108 9344
rect 4148 9304 4149 9344
rect 4107 9295 4149 9304
rect 3915 9260 3957 9269
rect 3915 9220 3916 9260
rect 3956 9220 3957 9260
rect 3915 9211 3957 9220
rect 3688 9092 4056 9101
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 3688 9043 4056 9052
rect 3532 8884 3668 8924
rect 3532 8672 3572 8681
rect 3532 8429 3572 8632
rect 3531 8420 3573 8429
rect 3531 8380 3532 8420
rect 3572 8380 3573 8420
rect 3531 8371 3573 8380
rect 3436 7951 3476 7960
rect 3628 8000 3668 8884
rect 4108 8840 4148 9295
rect 3916 8800 4148 8840
rect 3819 8756 3861 8765
rect 3819 8716 3820 8756
rect 3860 8716 3861 8756
rect 3819 8707 3861 8716
rect 3628 7951 3668 7960
rect 3820 8000 3860 8707
rect 3916 8177 3956 8800
rect 4204 8743 4244 12235
rect 4300 10781 4340 13000
rect 4395 12872 4437 12881
rect 4395 12832 4396 12872
rect 4436 12832 4437 12872
rect 4395 12823 4437 12832
rect 4396 12531 4436 12823
rect 4492 12536 4532 12545
rect 4491 12531 4492 12536
rect 4396 12496 4492 12531
rect 4396 12491 4532 12496
rect 4492 12487 4532 12491
rect 4587 12536 4629 12545
rect 4587 12496 4588 12536
rect 4628 12496 4629 12536
rect 4587 12487 4629 12496
rect 4588 12402 4628 12487
rect 4684 12125 4724 14008
rect 4780 14048 4820 14419
rect 4928 14384 5296 14393
rect 4968 14344 5010 14384
rect 5050 14344 5092 14384
rect 5132 14344 5174 14384
rect 5214 14344 5256 14384
rect 4928 14335 5296 14344
rect 5356 14309 5396 16360
rect 5452 15149 5492 16864
rect 5739 16652 5781 16661
rect 5739 16612 5740 16652
rect 5780 16612 5781 16652
rect 5739 16603 5781 16612
rect 5643 16400 5685 16409
rect 5643 16360 5644 16400
rect 5684 16360 5685 16400
rect 5643 16351 5685 16360
rect 5644 15560 5684 16351
rect 5644 15511 5684 15520
rect 5451 15140 5493 15149
rect 5451 15100 5452 15140
rect 5492 15100 5493 15140
rect 5451 15091 5493 15100
rect 5740 14972 5780 16603
rect 5931 16316 5973 16325
rect 5931 16276 5932 16316
rect 5972 16276 5973 16316
rect 5931 16267 5973 16276
rect 5835 15728 5877 15737
rect 5835 15688 5836 15728
rect 5876 15688 5877 15728
rect 5835 15679 5877 15688
rect 5836 15594 5876 15679
rect 5932 15653 5972 16267
rect 6027 15812 6069 15821
rect 6027 15772 6028 15812
rect 6068 15772 6069 15812
rect 6027 15763 6069 15772
rect 5931 15644 5973 15653
rect 5931 15604 5932 15644
rect 5972 15604 5973 15644
rect 5931 15595 5973 15604
rect 5835 15392 5877 15401
rect 5835 15352 5836 15392
rect 5876 15352 5877 15392
rect 5835 15343 5877 15352
rect 5644 14932 5780 14972
rect 5644 14813 5684 14932
rect 5643 14804 5685 14813
rect 5643 14764 5644 14804
rect 5684 14764 5685 14804
rect 5643 14755 5685 14764
rect 5548 14720 5588 14729
rect 5452 14552 5492 14561
rect 5355 14300 5397 14309
rect 5355 14260 5356 14300
rect 5396 14260 5397 14300
rect 5355 14251 5397 14260
rect 5452 14225 5492 14512
rect 4971 14216 5013 14225
rect 4971 14176 4972 14216
rect 5012 14176 5013 14216
rect 4971 14167 5013 14176
rect 5451 14216 5493 14225
rect 5451 14176 5452 14216
rect 5492 14176 5493 14216
rect 5451 14167 5493 14176
rect 4780 13999 4820 14008
rect 4972 14048 5012 14167
rect 4972 13999 5012 14008
rect 5164 14048 5204 14057
rect 4972 13796 5012 13805
rect 4780 13756 4972 13796
rect 4780 12536 4820 13756
rect 4972 13747 5012 13756
rect 5164 13040 5204 14008
rect 5260 14048 5300 14057
rect 5260 13217 5300 14008
rect 5356 14048 5396 14057
rect 5259 13208 5301 13217
rect 5259 13168 5260 13208
rect 5300 13168 5301 13208
rect 5259 13159 5301 13168
rect 5356 13124 5396 14008
rect 5452 14048 5492 14057
rect 5548 14048 5588 14680
rect 5644 14720 5684 14755
rect 5644 14669 5684 14680
rect 5740 14720 5780 14729
rect 5740 14477 5780 14680
rect 5739 14468 5781 14477
rect 5739 14428 5740 14468
rect 5780 14428 5781 14468
rect 5739 14419 5781 14428
rect 5740 14225 5780 14419
rect 5739 14216 5781 14225
rect 5739 14176 5740 14216
rect 5780 14176 5781 14216
rect 5739 14167 5781 14176
rect 5740 14048 5780 14057
rect 5492 14008 5740 14048
rect 5452 13999 5492 14008
rect 5643 13460 5685 13469
rect 5643 13420 5644 13460
rect 5684 13420 5685 13460
rect 5643 13411 5685 13420
rect 5740 13460 5780 14008
rect 5836 14048 5876 15343
rect 5932 14729 5972 15595
rect 6028 15560 6068 15763
rect 6028 15511 6068 15520
rect 6027 14972 6069 14981
rect 6027 14932 6028 14972
rect 6068 14932 6069 14972
rect 6027 14923 6069 14932
rect 6028 14838 6068 14923
rect 5931 14720 5973 14729
rect 5931 14680 5932 14720
rect 5972 14680 5973 14720
rect 5931 14671 5973 14680
rect 5932 14586 5972 14671
rect 6027 14132 6069 14141
rect 6027 14092 6028 14132
rect 6068 14092 6069 14132
rect 6027 14083 6069 14092
rect 5836 13999 5876 14008
rect 6028 13973 6068 14083
rect 6027 13964 6069 13973
rect 6027 13924 6028 13964
rect 6068 13924 6069 13964
rect 6027 13915 6069 13924
rect 5740 13411 5780 13420
rect 5547 13208 5589 13217
rect 5547 13168 5548 13208
rect 5588 13168 5589 13208
rect 5547 13159 5589 13168
rect 5356 13084 5492 13124
rect 5164 13000 5396 13040
rect 4928 12872 5296 12881
rect 4968 12832 5010 12872
rect 5050 12832 5092 12872
rect 5132 12832 5174 12872
rect 5214 12832 5256 12872
rect 4928 12823 5296 12832
rect 5356 12704 5396 13000
rect 5068 12664 5396 12704
rect 5068 12547 5108 12664
rect 5452 12620 5492 13084
rect 5548 13074 5588 13159
rect 5452 12571 5492 12580
rect 4876 12536 4916 12545
rect 4780 12496 4876 12536
rect 4876 12487 4916 12496
rect 4971 12536 5013 12545
rect 4971 12496 4972 12536
rect 5012 12496 5013 12536
rect 5068 12498 5108 12507
rect 5163 12536 5205 12545
rect 5260 12536 5300 12545
rect 4971 12487 5013 12496
rect 5163 12496 5164 12536
rect 5204 12496 5260 12536
rect 5163 12487 5205 12496
rect 5260 12487 5300 12496
rect 5356 12536 5396 12545
rect 4779 12368 4821 12377
rect 4779 12328 4780 12368
rect 4820 12328 4821 12368
rect 4779 12319 4821 12328
rect 4683 12116 4725 12125
rect 4683 12076 4684 12116
rect 4724 12076 4725 12116
rect 4683 12067 4725 12076
rect 4588 11864 4628 11873
rect 4683 11864 4725 11873
rect 4628 11824 4684 11864
rect 4724 11824 4725 11864
rect 4588 11815 4628 11824
rect 4683 11815 4725 11824
rect 4396 11701 4436 11705
rect 4396 11696 4532 11701
rect 4436 11661 4532 11696
rect 4396 11647 4436 11656
rect 4492 11537 4532 11661
rect 4780 11696 4820 12319
rect 4780 11647 4820 11656
rect 4972 11696 5012 12487
rect 5356 12293 5396 12496
rect 5548 12536 5588 12545
rect 5644 12536 5684 13411
rect 5932 13208 5972 13217
rect 5932 12797 5972 13168
rect 6027 13208 6069 13217
rect 6027 13168 6028 13208
rect 6068 13168 6069 13208
rect 6027 13159 6069 13168
rect 5931 12788 5973 12797
rect 5931 12748 5932 12788
rect 5972 12748 5973 12788
rect 5931 12739 5973 12748
rect 5588 12496 5684 12536
rect 5548 12487 5588 12496
rect 5932 12461 5972 12546
rect 5931 12452 5973 12461
rect 5931 12412 5932 12452
rect 5972 12412 5973 12452
rect 5931 12403 5973 12412
rect 5068 12284 5108 12293
rect 5355 12284 5397 12293
rect 5108 12244 5204 12284
rect 5068 12235 5108 12244
rect 5067 12116 5109 12125
rect 5067 12076 5068 12116
rect 5108 12076 5109 12116
rect 5067 12067 5109 12076
rect 4972 11621 5012 11656
rect 5068 11696 5108 12067
rect 5164 11957 5204 12244
rect 5355 12244 5356 12284
rect 5396 12244 5397 12284
rect 5355 12235 5397 12244
rect 5643 12284 5685 12293
rect 5643 12244 5644 12284
rect 5684 12244 5685 12284
rect 5643 12235 5685 12244
rect 5740 12284 5780 12293
rect 5163 11948 5205 11957
rect 5163 11908 5164 11948
rect 5204 11908 5205 11948
rect 5163 11899 5205 11908
rect 5068 11647 5108 11656
rect 5356 11696 5396 11705
rect 4971 11612 5013 11621
rect 4971 11572 4972 11612
rect 5012 11572 5013 11612
rect 4971 11563 5013 11572
rect 4491 11528 4533 11537
rect 4876 11528 4916 11537
rect 4491 11488 4492 11528
rect 4532 11488 4533 11528
rect 4491 11479 4533 11488
rect 4780 11488 4876 11528
rect 4395 11276 4437 11285
rect 4395 11236 4396 11276
rect 4436 11236 4437 11276
rect 4395 11227 4437 11236
rect 4299 10772 4341 10781
rect 4299 10732 4300 10772
rect 4340 10732 4341 10772
rect 4299 10723 4341 10732
rect 4299 10520 4341 10529
rect 4299 10480 4300 10520
rect 4340 10480 4341 10520
rect 4299 10471 4341 10480
rect 4300 8840 4340 10471
rect 4396 9932 4436 11227
rect 4492 10865 4532 11479
rect 4491 10856 4533 10865
rect 4491 10816 4492 10856
rect 4532 10816 4533 10856
rect 4491 10807 4533 10816
rect 4587 10772 4629 10781
rect 4587 10732 4588 10772
rect 4628 10732 4629 10772
rect 4587 10723 4629 10732
rect 4492 10184 4532 10195
rect 4492 10109 4532 10144
rect 4491 10100 4533 10109
rect 4491 10060 4492 10100
rect 4532 10060 4533 10100
rect 4491 10051 4533 10060
rect 4396 9892 4532 9932
rect 4492 9512 4532 9892
rect 4395 9428 4437 9437
rect 4395 9388 4396 9428
rect 4436 9388 4437 9428
rect 4395 9379 4437 9388
rect 4396 9294 4436 9379
rect 4492 9101 4532 9472
rect 4491 9092 4533 9101
rect 4491 9052 4492 9092
rect 4532 9052 4533 9092
rect 4491 9043 4533 9052
rect 4588 8924 4628 10723
rect 4684 10361 4724 10446
rect 4683 10352 4725 10361
rect 4683 10312 4684 10352
rect 4724 10312 4725 10352
rect 4683 10303 4725 10312
rect 4683 10184 4725 10193
rect 4683 10144 4684 10184
rect 4724 10144 4725 10184
rect 4780 10184 4820 11488
rect 4876 11479 4916 11488
rect 4928 11360 5296 11369
rect 4968 11320 5010 11360
rect 5050 11320 5092 11360
rect 5132 11320 5174 11360
rect 5214 11320 5256 11360
rect 4928 11311 5296 11320
rect 5260 11192 5300 11201
rect 5356 11192 5396 11656
rect 5452 11696 5492 11705
rect 5452 11285 5492 11656
rect 5547 11360 5589 11369
rect 5547 11320 5548 11360
rect 5588 11320 5589 11360
rect 5547 11311 5589 11320
rect 5451 11276 5493 11285
rect 5451 11236 5452 11276
rect 5492 11236 5493 11276
rect 5451 11227 5493 11236
rect 5300 11152 5396 11192
rect 5260 11143 5300 11152
rect 5067 11108 5109 11117
rect 5067 11068 5068 11108
rect 5108 11068 5109 11108
rect 5067 11059 5109 11068
rect 5068 11024 5108 11059
rect 5068 10973 5108 10984
rect 5548 11024 5588 11311
rect 5644 11192 5684 12235
rect 5740 11360 5780 12244
rect 5835 12032 5877 12041
rect 5835 11992 5836 12032
rect 5876 11992 5877 12032
rect 5835 11983 5877 11992
rect 5836 11780 5876 11983
rect 5836 11705 5876 11740
rect 5931 11780 5973 11789
rect 5931 11740 5932 11780
rect 5972 11740 5973 11780
rect 5931 11731 5973 11740
rect 5835 11696 5877 11705
rect 5835 11656 5836 11696
rect 5876 11656 5877 11696
rect 5835 11647 5877 11656
rect 5836 11616 5876 11647
rect 5932 11646 5972 11731
rect 5931 11528 5973 11537
rect 5931 11488 5932 11528
rect 5972 11488 5973 11528
rect 5931 11479 5973 11488
rect 5932 11360 5972 11479
rect 6028 11360 6068 13159
rect 6124 11957 6164 17032
rect 6220 17023 6260 17032
rect 6316 16904 6356 17611
rect 6412 17072 6452 17081
rect 6604 17072 6644 18619
rect 6891 18332 6933 18341
rect 6891 18292 6892 18332
rect 6932 18292 6933 18332
rect 6891 18283 6933 18292
rect 6892 17744 6932 18283
rect 6892 17669 6932 17704
rect 6891 17660 6933 17669
rect 6891 17620 6892 17660
rect 6932 17620 6933 17660
rect 6891 17611 6933 17620
rect 6452 17032 6548 17072
rect 6412 17023 6452 17032
rect 6220 16864 6356 16904
rect 6220 16325 6260 16864
rect 6412 16820 6452 16829
rect 6219 16316 6261 16325
rect 6219 16276 6220 16316
rect 6260 16276 6261 16316
rect 6219 16267 6261 16276
rect 6315 16232 6357 16241
rect 6315 16192 6316 16232
rect 6356 16192 6357 16232
rect 6315 16183 6357 16192
rect 6219 14720 6261 14729
rect 6219 14680 6220 14720
rect 6260 14680 6261 14720
rect 6219 14671 6261 14680
rect 6220 14586 6260 14671
rect 6316 13973 6356 16183
rect 6220 13964 6260 13973
rect 6220 12788 6260 13924
rect 6315 13964 6357 13973
rect 6315 13924 6316 13964
rect 6356 13924 6357 13964
rect 6315 13915 6357 13924
rect 6316 13830 6356 13915
rect 6220 12748 6356 12788
rect 6220 12545 6260 12630
rect 6219 12536 6261 12545
rect 6219 12496 6220 12536
rect 6260 12496 6261 12536
rect 6219 12487 6261 12496
rect 6316 12377 6356 12748
rect 6412 12461 6452 16780
rect 6508 16400 6548 17032
rect 6604 17023 6644 17032
rect 7084 16661 7124 18628
rect 7372 18584 7412 18593
rect 7180 18544 7372 18584
rect 7180 17081 7220 18544
rect 7372 18535 7412 18544
rect 7468 18080 7508 19216
rect 7564 19181 7604 19300
rect 7756 19340 7796 20140
rect 8044 20105 8084 20140
rect 8043 20096 8085 20105
rect 7900 20054 7940 20063
rect 8043 20056 8044 20096
rect 8084 20056 8085 20096
rect 8043 20047 8085 20056
rect 8044 20045 8084 20047
rect 7900 20012 7940 20014
rect 7900 19972 7988 20012
rect 7851 19424 7893 19433
rect 7851 19384 7852 19424
rect 7892 19384 7893 19424
rect 7851 19375 7893 19384
rect 7756 19291 7796 19300
rect 7852 19256 7892 19375
rect 7852 19207 7892 19216
rect 7563 19172 7605 19181
rect 7563 19132 7564 19172
rect 7604 19132 7605 19172
rect 7563 19123 7605 19132
rect 7564 18752 7604 18761
rect 7948 18752 7988 19972
rect 7604 18712 7988 18752
rect 7564 18703 7604 18712
rect 8140 18668 8180 21988
rect 8236 21978 8276 22063
rect 7852 18628 8180 18668
rect 8236 21608 8276 21617
rect 8332 21608 8372 22819
rect 8427 22112 8469 22121
rect 8427 22072 8428 22112
rect 8468 22072 8469 22112
rect 8427 22063 8469 22072
rect 8428 21978 8468 22063
rect 8276 21568 8372 21608
rect 7755 18584 7797 18593
rect 7755 18544 7756 18584
rect 7796 18544 7797 18584
rect 7755 18535 7797 18544
rect 7756 18450 7796 18535
rect 7276 18040 7508 18080
rect 7276 17249 7316 18040
rect 7755 17912 7797 17921
rect 7755 17872 7756 17912
rect 7796 17872 7797 17912
rect 7755 17863 7797 17872
rect 7756 17778 7796 17863
rect 7372 17749 7412 17758
rect 7275 17240 7317 17249
rect 7275 17200 7276 17240
rect 7316 17200 7317 17240
rect 7275 17191 7317 17200
rect 7179 17072 7221 17081
rect 7179 17032 7180 17072
rect 7220 17032 7221 17072
rect 7179 17023 7221 17032
rect 7083 16652 7125 16661
rect 7083 16612 7084 16652
rect 7124 16612 7125 16652
rect 7083 16603 7125 16612
rect 7180 16409 7220 17023
rect 7179 16400 7221 16409
rect 6508 16360 6644 16400
rect 6507 16232 6549 16241
rect 6507 16192 6508 16232
rect 6548 16192 6549 16232
rect 6507 16183 6549 16192
rect 6508 16098 6548 16183
rect 6507 14552 6549 14561
rect 6507 14512 6508 14552
rect 6548 14512 6549 14552
rect 6507 14503 6549 14512
rect 6411 12452 6453 12461
rect 6411 12412 6412 12452
rect 6452 12412 6453 12452
rect 6411 12403 6453 12412
rect 6315 12368 6357 12377
rect 6315 12328 6316 12368
rect 6356 12328 6357 12368
rect 6315 12319 6357 12328
rect 6123 11948 6165 11957
rect 6123 11908 6124 11948
rect 6164 11908 6165 11948
rect 6123 11899 6165 11908
rect 6316 11789 6356 12319
rect 6508 11948 6548 14503
rect 6604 12032 6644 16360
rect 7179 16360 7180 16400
rect 7220 16360 7221 16400
rect 7179 16351 7221 16360
rect 7084 16241 7124 16246
rect 6891 16232 6933 16241
rect 6796 16192 6892 16232
rect 6932 16192 6933 16232
rect 6700 16148 6740 16157
rect 6796 16148 6836 16192
rect 6891 16183 6933 16192
rect 7083 16237 7125 16241
rect 7083 16192 7084 16237
rect 7124 16192 7125 16237
rect 7083 16183 7125 16192
rect 6740 16108 6836 16148
rect 6700 16099 6740 16108
rect 7084 16102 7124 16183
rect 6891 16064 6933 16073
rect 6891 16024 6892 16064
rect 6932 16024 6933 16064
rect 6891 16015 6933 16024
rect 6892 15930 6932 16015
rect 7180 14729 7220 16351
rect 7275 15896 7317 15905
rect 7275 15856 7276 15896
rect 7316 15856 7317 15896
rect 7275 15847 7317 15856
rect 7276 15560 7316 15847
rect 7276 15511 7316 15520
rect 7179 14720 7221 14729
rect 7179 14680 7180 14720
rect 7220 14680 7221 14720
rect 7179 14671 7221 14680
rect 6795 14048 6837 14057
rect 6795 14008 6796 14048
rect 6836 14008 6837 14048
rect 6795 13999 6837 14008
rect 6987 14048 7029 14057
rect 6987 14008 6988 14048
rect 7028 14008 7029 14048
rect 6987 13999 7029 14008
rect 6699 13964 6741 13973
rect 6699 13924 6700 13964
rect 6740 13924 6741 13964
rect 6699 13915 6741 13924
rect 6700 12629 6740 13915
rect 6796 13914 6836 13999
rect 6795 13544 6837 13553
rect 6795 13504 6796 13544
rect 6836 13504 6837 13544
rect 6795 13495 6837 13504
rect 6699 12620 6741 12629
rect 6699 12580 6700 12620
rect 6740 12580 6741 12620
rect 6699 12571 6741 12580
rect 6700 12209 6740 12571
rect 6796 12545 6836 13495
rect 6795 12536 6837 12545
rect 6795 12496 6796 12536
rect 6836 12496 6837 12536
rect 6795 12487 6837 12496
rect 6699 12200 6741 12209
rect 6699 12160 6700 12200
rect 6740 12160 6741 12200
rect 6699 12151 6741 12160
rect 6891 12032 6933 12041
rect 6604 11992 6892 12032
rect 6932 11992 6933 12032
rect 6891 11983 6933 11992
rect 6508 11908 6644 11948
rect 6315 11780 6357 11789
rect 6315 11740 6316 11780
rect 6356 11740 6357 11780
rect 6315 11731 6357 11740
rect 6507 11780 6549 11789
rect 6507 11740 6508 11780
rect 6548 11740 6549 11780
rect 6507 11731 6549 11740
rect 6412 11696 6452 11705
rect 6412 11612 6452 11656
rect 5740 11320 5876 11360
rect 5740 11192 5780 11201
rect 5644 11152 5740 11192
rect 5740 11143 5780 11152
rect 5548 10975 5588 10984
rect 5451 10856 5493 10865
rect 5451 10816 5452 10856
rect 5492 10816 5493 10856
rect 5451 10807 5493 10816
rect 5452 10722 5492 10807
rect 5836 10613 5876 11320
rect 5932 11320 6068 11360
rect 6316 11572 6452 11612
rect 5932 11024 5972 11320
rect 6219 11276 6261 11285
rect 6219 11236 6220 11276
rect 6260 11236 6261 11276
rect 6219 11227 6261 11236
rect 6027 11192 6069 11201
rect 6027 11152 6028 11192
rect 6068 11152 6069 11192
rect 6027 11143 6069 11152
rect 5835 10604 5877 10613
rect 5835 10564 5836 10604
rect 5876 10564 5877 10604
rect 5835 10555 5877 10564
rect 5068 10436 5108 10445
rect 5108 10396 5780 10436
rect 5068 10387 5108 10396
rect 5259 10268 5301 10277
rect 5259 10228 5260 10268
rect 5300 10228 5301 10268
rect 5259 10219 5301 10228
rect 4876 10184 4916 10193
rect 4780 10144 4876 10184
rect 4683 10135 4725 10144
rect 4876 10135 4916 10144
rect 4684 10050 4724 10135
rect 5260 10134 5300 10219
rect 5451 10184 5493 10193
rect 5451 10144 5452 10184
rect 5492 10144 5493 10184
rect 5451 10135 5493 10144
rect 5452 10050 5492 10135
rect 5643 10016 5685 10025
rect 5643 9976 5644 10016
rect 5684 9976 5685 10016
rect 5643 9967 5685 9976
rect 4928 9848 5296 9857
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 4928 9799 5296 9808
rect 4779 9596 4821 9605
rect 4779 9556 4780 9596
rect 4820 9556 4821 9596
rect 4779 9547 4821 9556
rect 4588 8884 4724 8924
rect 4396 8840 4436 8849
rect 4300 8800 4396 8840
rect 4396 8791 4436 8800
rect 4108 8703 4244 8743
rect 4577 8767 4617 8776
rect 4684 8743 4724 8884
rect 4780 8849 4820 9547
rect 4876 9512 4916 9521
rect 4779 8840 4821 8849
rect 4779 8800 4780 8840
rect 4820 8800 4821 8840
rect 4876 8840 4916 9472
rect 4971 9512 5013 9521
rect 4971 9472 4972 9512
rect 5012 9472 5013 9512
rect 4971 9463 5013 9472
rect 5356 9512 5396 9521
rect 5547 9512 5589 9521
rect 5396 9472 5492 9512
rect 5356 9463 5396 9472
rect 4972 9378 5012 9463
rect 5356 9260 5396 9269
rect 5164 9220 5356 9260
rect 4876 8800 5108 8840
rect 4779 8791 4821 8800
rect 4012 8677 4052 8686
rect 3915 8168 3957 8177
rect 3915 8128 3916 8168
rect 3956 8128 3957 8168
rect 3915 8119 3957 8128
rect 3820 7951 3860 7960
rect 4012 7925 4052 8637
rect 3532 7916 3572 7925
rect 3532 7673 3572 7876
rect 4011 7916 4053 7925
rect 4011 7876 4012 7916
rect 4052 7876 4053 7916
rect 4011 7867 4053 7876
rect 3531 7664 3573 7673
rect 3531 7624 3532 7664
rect 3572 7624 3573 7664
rect 3531 7615 3573 7624
rect 3688 7580 4056 7589
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 3688 7531 4056 7540
rect 4108 7421 4148 8703
rect 4577 8677 4617 8727
rect 4492 8637 4617 8677
rect 4666 8703 4724 8743
rect 4204 8588 4244 8597
rect 4492 8588 4532 8637
rect 4666 8588 4706 8703
rect 5068 8681 5108 8800
rect 4972 8672 5012 8681
rect 4244 8548 4532 8588
rect 4588 8548 4706 8588
rect 4780 8632 4972 8672
rect 4204 8539 4244 8548
rect 4299 8336 4341 8345
rect 4299 8296 4300 8336
rect 4340 8296 4341 8336
rect 4299 8287 4341 8296
rect 4203 8168 4245 8177
rect 4203 8128 4204 8168
rect 4244 8128 4245 8168
rect 4203 8119 4245 8128
rect 4107 7412 4149 7421
rect 4107 7372 4108 7412
rect 4148 7372 4149 7412
rect 4107 7363 4149 7372
rect 3531 7244 3573 7253
rect 3531 7204 3532 7244
rect 3572 7204 3573 7244
rect 3531 7195 3573 7204
rect 3532 7110 3572 7195
rect 3628 7160 3668 7169
rect 3435 6320 3477 6329
rect 3435 6280 3436 6320
rect 3476 6280 3477 6320
rect 3435 6271 3477 6280
rect 3051 5648 3093 5657
rect 3051 5608 3052 5648
rect 3092 5608 3093 5648
rect 3051 5599 3093 5608
rect 3148 5648 3188 5657
rect 3148 5321 3188 5608
rect 3339 5648 3381 5657
rect 3339 5608 3340 5648
rect 3380 5608 3381 5648
rect 3339 5599 3381 5608
rect 3436 5648 3476 6271
rect 3628 6236 3668 7120
rect 4108 7160 4148 7169
rect 4204 7160 4244 8119
rect 4148 7120 4244 7160
rect 4108 7111 4148 7120
rect 4204 6665 4244 6750
rect 4203 6656 4245 6665
rect 4203 6616 4204 6656
rect 4244 6616 4245 6656
rect 4203 6607 4245 6616
rect 4300 6497 4340 8287
rect 4588 7328 4628 8548
rect 4492 7288 4628 7328
rect 4395 6572 4437 6581
rect 4395 6532 4396 6572
rect 4436 6532 4437 6572
rect 4395 6523 4437 6532
rect 4011 6488 4053 6497
rect 4011 6448 4012 6488
rect 4052 6448 4053 6488
rect 4011 6439 4053 6448
rect 4299 6488 4341 6497
rect 4299 6448 4300 6488
rect 4340 6448 4341 6488
rect 4299 6439 4341 6448
rect 4012 6354 4052 6439
rect 4396 6438 4436 6523
rect 3532 6196 3668 6236
rect 3532 5900 3572 6196
rect 4203 6152 4245 6161
rect 4203 6112 4204 6152
rect 4244 6112 4245 6152
rect 4203 6103 4245 6112
rect 3688 6068 4056 6077
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 3688 6019 4056 6028
rect 3532 5860 3668 5900
rect 3628 5816 3668 5860
rect 3819 5816 3861 5825
rect 3628 5776 3764 5816
rect 3532 5657 3572 5742
rect 3340 5480 3380 5489
rect 3147 5312 3189 5321
rect 3147 5272 3148 5312
rect 3188 5272 3189 5312
rect 3147 5263 3189 5272
rect 2764 4339 2804 4348
rect 2860 4768 2996 4808
rect 3052 4892 3092 4901
rect 2667 3968 2709 3977
rect 2667 3928 2668 3968
rect 2708 3928 2709 3968
rect 2667 3919 2709 3928
rect 2667 3548 2709 3557
rect 2667 3508 2668 3548
rect 2708 3508 2709 3548
rect 2667 3499 2709 3508
rect 2668 3464 2708 3499
rect 2668 3413 2708 3424
rect 2667 3296 2709 3305
rect 2572 3256 2668 3296
rect 2708 3256 2709 3296
rect 2667 3247 2709 3256
rect 2668 2624 2708 3247
rect 2763 3212 2805 3221
rect 2763 3172 2764 3212
rect 2804 3172 2805 3212
rect 2763 3163 2805 3172
rect 2668 2575 2708 2584
rect 2379 2372 2421 2381
rect 2379 2332 2380 2372
rect 2420 2332 2421 2372
rect 2379 2323 2421 2332
rect 2380 1952 2420 2323
rect 2380 1903 2420 1912
rect 2667 1952 2709 1961
rect 2667 1912 2668 1952
rect 2708 1912 2709 1952
rect 2667 1903 2709 1912
rect 1460 1072 1556 1112
rect 1804 1072 1940 1112
rect 2188 1408 2324 1448
rect 1420 1063 1460 1072
rect 1035 356 1077 365
rect 1035 316 1036 356
rect 1076 316 1077 356
rect 1035 307 1077 316
rect 1804 80 1844 1072
rect 1995 1028 2037 1037
rect 1995 988 1996 1028
rect 2036 988 2037 1028
rect 1995 979 2037 988
rect 1996 80 2036 979
rect 2188 80 2228 1408
rect 2571 1280 2613 1289
rect 2571 1240 2572 1280
rect 2612 1240 2613 1280
rect 2571 1231 2613 1240
rect 2379 440 2421 449
rect 2379 400 2380 440
rect 2420 400 2421 440
rect 2379 391 2421 400
rect 2380 80 2420 391
rect 2572 80 2612 1231
rect 2668 1112 2708 1903
rect 2668 1063 2708 1072
rect 2764 80 2804 3163
rect 2860 2876 2900 4768
rect 3052 4229 3092 4852
rect 3148 4892 3188 4901
rect 3148 4649 3188 4852
rect 3147 4640 3189 4649
rect 3147 4600 3148 4640
rect 3188 4600 3189 4640
rect 3147 4591 3189 4600
rect 3340 4388 3380 5440
rect 3436 5153 3476 5608
rect 3531 5648 3573 5657
rect 3531 5608 3532 5648
rect 3572 5608 3573 5648
rect 3531 5599 3573 5608
rect 3628 5648 3668 5657
rect 3531 5480 3573 5489
rect 3531 5440 3532 5480
rect 3572 5440 3573 5480
rect 3531 5431 3573 5440
rect 3435 5144 3477 5153
rect 3435 5104 3436 5144
rect 3476 5104 3477 5144
rect 3435 5095 3477 5104
rect 3148 4348 3380 4388
rect 3051 4220 3093 4229
rect 3051 4180 3052 4220
rect 3092 4180 3093 4220
rect 3051 4171 3093 4180
rect 2956 4136 2996 4145
rect 2956 3809 2996 4096
rect 3148 4052 3188 4348
rect 3339 4220 3381 4229
rect 3339 4180 3340 4220
rect 3380 4180 3381 4220
rect 3339 4171 3381 4180
rect 3052 4012 3188 4052
rect 2955 3800 2997 3809
rect 2955 3760 2956 3800
rect 2996 3760 2997 3800
rect 2955 3751 2997 3760
rect 2955 3632 2997 3641
rect 2955 3592 2956 3632
rect 2996 3592 2997 3632
rect 2955 3583 2997 3592
rect 2860 2827 2900 2836
rect 2859 2624 2901 2633
rect 2859 2584 2860 2624
rect 2900 2584 2901 2624
rect 2859 2575 2901 2584
rect 2860 1280 2900 2575
rect 2860 1231 2900 1240
rect 2956 80 2996 3583
rect 3052 2624 3092 4012
rect 3243 3884 3285 3893
rect 3243 3844 3244 3884
rect 3284 3844 3285 3884
rect 3243 3835 3285 3844
rect 3244 3464 3284 3835
rect 3244 3415 3284 3424
rect 3148 3380 3188 3389
rect 3148 3221 3188 3340
rect 3147 3212 3189 3221
rect 3147 3172 3148 3212
rect 3188 3172 3189 3212
rect 3147 3163 3189 3172
rect 3340 3137 3380 4171
rect 3435 3800 3477 3809
rect 3435 3760 3436 3800
rect 3476 3760 3477 3800
rect 3435 3751 3477 3760
rect 3339 3128 3381 3137
rect 3339 3088 3340 3128
rect 3380 3088 3381 3128
rect 3339 3079 3381 3088
rect 3243 2792 3285 2801
rect 3243 2752 3244 2792
rect 3284 2752 3285 2792
rect 3243 2743 3285 2752
rect 3147 2708 3189 2717
rect 3147 2668 3148 2708
rect 3188 2668 3189 2708
rect 3147 2659 3189 2668
rect 3052 2575 3092 2584
rect 3148 2574 3188 2659
rect 3244 2624 3284 2743
rect 3244 2575 3284 2584
rect 3436 2540 3476 3751
rect 3532 2801 3572 5431
rect 3628 5405 3668 5608
rect 3627 5396 3669 5405
rect 3627 5356 3628 5396
rect 3668 5356 3669 5396
rect 3627 5347 3669 5356
rect 3724 5237 3764 5776
rect 3819 5776 3820 5816
rect 3860 5776 3861 5816
rect 3819 5767 3861 5776
rect 3820 5648 3860 5767
rect 3820 5599 3860 5608
rect 3915 5648 3957 5657
rect 3915 5608 3916 5648
rect 3956 5608 3957 5648
rect 3915 5599 3957 5608
rect 3723 5228 3765 5237
rect 3723 5188 3724 5228
rect 3764 5188 3765 5228
rect 3723 5179 3765 5188
rect 3627 4976 3669 4985
rect 3916 4976 3956 5599
rect 3627 4936 3628 4976
rect 3668 4936 3956 4976
rect 4108 4962 4148 4971
rect 3627 4927 3669 4936
rect 3628 4842 3668 4927
rect 3688 4556 4056 4565
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 3688 4507 4056 4516
rect 4108 3893 4148 4922
rect 4204 4808 4244 6103
rect 4492 5993 4532 7288
rect 4588 7165 4628 7174
rect 4780 7160 4820 8632
rect 4972 8623 5012 8632
rect 5067 8672 5109 8681
rect 5067 8632 5068 8672
rect 5108 8632 5109 8672
rect 5067 8623 5109 8632
rect 5164 8672 5204 9220
rect 5356 9211 5396 9220
rect 5356 8681 5396 8766
rect 5164 8623 5204 8632
rect 5355 8672 5397 8681
rect 5355 8632 5356 8672
rect 5396 8632 5397 8672
rect 5355 8623 5397 8632
rect 5068 8504 5108 8513
rect 5108 8464 5396 8504
rect 5068 8455 5108 8464
rect 4928 8336 5296 8345
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 4928 8287 5296 8296
rect 5259 8168 5301 8177
rect 5259 8128 5260 8168
rect 5300 8128 5301 8168
rect 5259 8119 5301 8128
rect 5260 8034 5300 8119
rect 5067 8000 5109 8009
rect 5067 7960 5068 8000
rect 5108 7960 5109 8000
rect 5067 7951 5109 7960
rect 5068 7866 5108 7951
rect 5164 7421 5204 7506
rect 5163 7412 5205 7421
rect 5163 7372 5164 7412
rect 5204 7372 5205 7412
rect 5163 7363 5205 7372
rect 5163 7244 5205 7253
rect 5163 7204 5164 7244
rect 5204 7204 5205 7244
rect 5163 7195 5205 7204
rect 4588 6665 4628 7125
rect 4684 7120 4820 7160
rect 4971 7160 5013 7169
rect 4971 7120 4972 7160
rect 5012 7120 5013 7160
rect 4587 6656 4629 6665
rect 4587 6616 4588 6656
rect 4628 6616 4629 6656
rect 4587 6607 4629 6616
rect 4684 6581 4724 7120
rect 4971 7111 5013 7120
rect 5164 7160 5204 7195
rect 5356 7169 5396 8464
rect 5452 8261 5492 9472
rect 5547 9472 5548 9512
rect 5588 9472 5589 9512
rect 5547 9463 5589 9472
rect 5644 9510 5684 9967
rect 5451 8252 5493 8261
rect 5451 8212 5452 8252
rect 5492 8212 5493 8252
rect 5451 8203 5493 8212
rect 5548 8177 5588 9463
rect 5644 9461 5684 9470
rect 5740 8504 5780 10396
rect 5932 9680 5972 10984
rect 6028 10865 6068 11143
rect 6027 10856 6069 10865
rect 6027 10816 6028 10856
rect 6068 10816 6069 10856
rect 6027 10807 6069 10816
rect 6027 10436 6069 10445
rect 6027 10396 6028 10436
rect 6068 10396 6069 10436
rect 6027 10387 6069 10396
rect 5644 8464 5780 8504
rect 5836 9640 5972 9680
rect 5547 8168 5589 8177
rect 5547 8128 5548 8168
rect 5588 8128 5589 8168
rect 5547 8119 5589 8128
rect 5451 8000 5493 8009
rect 5451 7960 5452 8000
rect 5492 7960 5493 8000
rect 5451 7951 5493 7960
rect 5452 7866 5492 7951
rect 4972 7026 5012 7111
rect 5164 7109 5204 7120
rect 5355 7160 5397 7169
rect 5355 7120 5356 7160
rect 5396 7120 5397 7160
rect 5355 7111 5397 7120
rect 5452 7160 5492 7169
rect 5452 7001 5492 7120
rect 5548 7160 5588 7169
rect 4780 6992 4820 7001
rect 4780 6833 4820 6952
rect 5451 6992 5493 7001
rect 5451 6952 5452 6992
rect 5492 6952 5493 6992
rect 5451 6943 5493 6952
rect 5548 6833 5588 7120
rect 5644 7085 5684 8464
rect 5739 8252 5781 8261
rect 5739 8212 5740 8252
rect 5780 8212 5781 8252
rect 5739 8203 5781 8212
rect 5643 7076 5685 7085
rect 5643 7036 5644 7076
rect 5684 7036 5685 7076
rect 5643 7027 5685 7036
rect 4779 6824 4821 6833
rect 4779 6784 4780 6824
rect 4820 6784 4821 6824
rect 4779 6775 4821 6784
rect 4928 6824 5296 6833
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 4928 6775 5296 6784
rect 5547 6824 5589 6833
rect 5547 6784 5548 6824
rect 5588 6784 5589 6824
rect 5547 6775 5589 6784
rect 5643 6740 5685 6749
rect 5643 6700 5644 6740
rect 5684 6700 5685 6740
rect 5643 6691 5685 6700
rect 5067 6656 5109 6665
rect 5067 6616 5068 6656
rect 5108 6616 5109 6656
rect 5067 6607 5109 6616
rect 4683 6572 4725 6581
rect 4683 6532 4684 6572
rect 4724 6532 4725 6572
rect 4683 6523 4725 6532
rect 5068 6488 5108 6607
rect 4588 6474 4628 6483
rect 5068 6439 5108 6448
rect 5547 6488 5589 6497
rect 5547 6448 5548 6488
rect 5588 6448 5589 6488
rect 5547 6439 5589 6448
rect 5644 6488 5684 6691
rect 5644 6439 5684 6448
rect 4491 5984 4533 5993
rect 4491 5944 4492 5984
rect 4532 5944 4533 5984
rect 4491 5935 4533 5944
rect 4395 5900 4437 5909
rect 4395 5860 4396 5900
rect 4436 5860 4437 5900
rect 4395 5851 4437 5860
rect 4300 5060 4340 5071
rect 4300 4985 4340 5020
rect 4299 4976 4341 4985
rect 4299 4936 4300 4976
rect 4340 4936 4341 4976
rect 4299 4927 4341 4936
rect 4204 4768 4340 4808
rect 4203 4220 4245 4229
rect 4203 4180 4204 4220
rect 4244 4180 4245 4220
rect 4203 4171 4245 4180
rect 4204 4136 4244 4171
rect 4204 4085 4244 4096
rect 4300 3968 4340 4768
rect 4396 4640 4436 5851
rect 4492 5657 4532 5935
rect 4491 5648 4533 5657
rect 4491 5608 4492 5648
rect 4532 5608 4533 5648
rect 4491 5599 4533 5608
rect 4588 5405 4628 6434
rect 5548 6354 5588 6439
rect 5740 6329 5780 8203
rect 5836 7925 5876 9640
rect 5931 9512 5973 9521
rect 5931 9472 5932 9512
rect 5972 9472 5973 9512
rect 5931 9463 5973 9472
rect 6028 9512 6068 10387
rect 6220 10361 6260 11227
rect 6219 10352 6261 10361
rect 6219 10312 6220 10352
rect 6260 10312 6261 10352
rect 6219 10303 6261 10312
rect 6219 10100 6261 10109
rect 6219 10060 6220 10100
rect 6260 10060 6261 10100
rect 6219 10051 6261 10060
rect 6028 9463 6068 9472
rect 5932 9378 5972 9463
rect 6123 8672 6165 8681
rect 6123 8632 6124 8672
rect 6164 8632 6165 8672
rect 6123 8623 6165 8632
rect 5835 7916 5877 7925
rect 5835 7876 5836 7916
rect 5876 7876 5877 7916
rect 5835 7867 5877 7876
rect 6124 7757 6164 8623
rect 6123 7748 6165 7757
rect 6123 7708 6124 7748
rect 6164 7708 6165 7748
rect 6123 7699 6165 7708
rect 5835 7580 5877 7589
rect 5835 7540 5836 7580
rect 5876 7540 5877 7580
rect 5835 7531 5877 7540
rect 5836 6665 5876 7531
rect 5931 7160 5973 7169
rect 5931 7120 5932 7160
rect 5972 7120 5973 7160
rect 5931 7111 5973 7120
rect 6028 7160 6068 7171
rect 5932 7026 5972 7111
rect 6028 7085 6068 7120
rect 6027 7076 6069 7085
rect 6027 7036 6028 7076
rect 6068 7036 6069 7076
rect 6027 7027 6069 7036
rect 5835 6656 5877 6665
rect 5835 6616 5836 6656
rect 5876 6616 5877 6656
rect 5835 6607 5877 6616
rect 6027 6488 6069 6497
rect 6027 6448 6028 6488
rect 6068 6448 6069 6488
rect 6027 6439 6069 6448
rect 6124 6488 6164 6497
rect 5835 6404 5877 6413
rect 5835 6364 5836 6404
rect 5876 6364 5877 6404
rect 5835 6355 5877 6364
rect 5739 6320 5781 6329
rect 5739 6280 5740 6320
rect 5780 6280 5781 6320
rect 5739 6271 5781 6280
rect 5643 6236 5685 6245
rect 5643 6196 5644 6236
rect 5684 6196 5685 6236
rect 5643 6187 5685 6196
rect 5259 6152 5301 6161
rect 5259 6112 5260 6152
rect 5300 6112 5301 6152
rect 5259 6103 5301 6112
rect 5260 5900 5300 6103
rect 5260 5851 5300 5860
rect 4683 5648 4725 5657
rect 4683 5608 4684 5648
rect 4724 5608 4725 5648
rect 4683 5599 4725 5608
rect 5067 5648 5109 5657
rect 5067 5608 5068 5648
rect 5108 5608 5109 5648
rect 5067 5599 5109 5608
rect 5452 5648 5492 5657
rect 4587 5396 4629 5405
rect 4587 5356 4588 5396
rect 4628 5356 4629 5396
rect 4587 5347 4629 5356
rect 4491 5144 4533 5153
rect 4491 5104 4492 5144
rect 4532 5104 4533 5144
rect 4491 5095 4533 5104
rect 4492 5010 4532 5095
rect 4684 4976 4724 5599
rect 5068 5514 5108 5599
rect 4928 5312 5296 5321
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 4928 5263 5296 5272
rect 4396 4600 4532 4640
rect 4395 4472 4437 4481
rect 4395 4432 4396 4472
rect 4436 4432 4437 4472
rect 4395 4423 4437 4432
rect 4396 4388 4436 4423
rect 4396 4337 4436 4348
rect 4395 4052 4437 4061
rect 4395 4012 4396 4052
rect 4436 4012 4437 4052
rect 4395 4003 4437 4012
rect 4204 3928 4340 3968
rect 4107 3884 4149 3893
rect 4107 3844 4108 3884
rect 4148 3844 4149 3884
rect 4107 3835 4149 3844
rect 3915 3800 3957 3809
rect 3915 3760 3916 3800
rect 3956 3760 3957 3800
rect 3915 3751 3957 3760
rect 3723 3548 3765 3557
rect 3723 3508 3724 3548
rect 3764 3508 3765 3548
rect 3916 3548 3956 3751
rect 4012 3548 4052 3557
rect 3916 3508 4012 3548
rect 3723 3499 3765 3508
rect 4012 3499 4052 3508
rect 3628 3464 3668 3475
rect 3628 3389 3668 3424
rect 3724 3464 3764 3499
rect 3724 3413 3764 3424
rect 3627 3380 3669 3389
rect 3627 3340 3628 3380
rect 3668 3340 3669 3380
rect 3627 3331 3669 3340
rect 3688 3044 4056 3053
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 3688 2995 4056 3004
rect 4204 2876 4244 3928
rect 4396 3884 4436 4003
rect 4300 3844 4436 3884
rect 4300 3632 4340 3844
rect 4395 3716 4437 3725
rect 4395 3676 4396 3716
rect 4436 3676 4437 3716
rect 4395 3667 4437 3676
rect 4300 3583 4340 3592
rect 4396 3464 4436 3667
rect 4396 3415 4436 3424
rect 4299 3044 4341 3053
rect 4299 3004 4300 3044
rect 4340 3004 4341 3044
rect 4299 2995 4341 3004
rect 4204 2836 4254 2876
rect 3531 2792 3573 2801
rect 3531 2752 3532 2792
rect 3572 2752 3573 2792
rect 3531 2743 3573 2752
rect 3819 2792 3861 2801
rect 3819 2752 3820 2792
rect 3860 2752 3861 2792
rect 3819 2743 3861 2752
rect 3627 2708 3669 2717
rect 3627 2668 3628 2708
rect 3668 2668 3669 2708
rect 3627 2659 3669 2668
rect 3628 2574 3668 2659
rect 3820 2658 3860 2743
rect 4214 2717 4254 2836
rect 4204 2708 4254 2717
rect 4244 2668 4254 2708
rect 4204 2659 4244 2668
rect 3340 2500 3476 2540
rect 3147 1280 3189 1289
rect 3147 1240 3148 1280
rect 3188 1240 3189 1280
rect 3147 1231 3189 1240
rect 3052 1112 3092 1121
rect 3052 197 3092 1072
rect 3051 188 3093 197
rect 3051 148 3052 188
rect 3092 148 3093 188
rect 3051 139 3093 148
rect 3148 80 3188 1231
rect 3340 80 3380 2500
rect 4011 2456 4053 2465
rect 4011 2416 4012 2456
rect 4052 2416 4053 2456
rect 4011 2407 4053 2416
rect 4012 2322 4052 2407
rect 4107 2288 4149 2297
rect 4107 2248 4108 2288
rect 4148 2248 4149 2288
rect 4107 2239 4149 2248
rect 3820 2036 3860 2045
rect 3860 1996 3956 2036
rect 3820 1987 3860 1996
rect 3627 1952 3669 1961
rect 3627 1912 3628 1952
rect 3668 1912 3669 1952
rect 3916 1952 3956 1996
rect 4011 1952 4053 1961
rect 3916 1912 4012 1952
rect 4052 1912 4053 1952
rect 3627 1903 3669 1912
rect 4011 1903 4053 1912
rect 4108 1952 4148 2239
rect 4300 2120 4340 2995
rect 4395 2960 4437 2969
rect 4395 2920 4396 2960
rect 4436 2920 4437 2960
rect 4395 2911 4437 2920
rect 4396 2792 4436 2911
rect 4396 2743 4436 2752
rect 4395 2204 4437 2213
rect 4395 2164 4396 2204
rect 4436 2164 4437 2204
rect 4395 2155 4437 2164
rect 4300 2071 4340 2080
rect 3628 1818 3668 1903
rect 4012 1818 4052 1903
rect 3688 1532 4056 1541
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 3688 1483 4056 1492
rect 4108 1289 4148 1912
rect 4396 1709 4436 2155
rect 4395 1700 4437 1709
rect 4395 1660 4396 1700
rect 4436 1660 4437 1700
rect 4395 1651 4437 1660
rect 3723 1280 3765 1289
rect 3723 1240 3724 1280
rect 3764 1240 3765 1280
rect 3723 1231 3765 1240
rect 4107 1280 4149 1289
rect 4107 1240 4108 1280
rect 4148 1240 4149 1280
rect 4107 1231 4149 1240
rect 4492 1280 4532 4600
rect 4684 4229 4724 4936
rect 4683 4220 4725 4229
rect 4683 4180 4684 4220
rect 4724 4180 4725 4220
rect 4683 4171 4725 4180
rect 4587 4136 4629 4145
rect 4587 4096 4588 4136
rect 4628 4096 4629 4136
rect 4587 4087 4629 4096
rect 4588 4002 4628 4087
rect 5355 4052 5397 4061
rect 5355 4012 5356 4052
rect 5396 4012 5397 4052
rect 5355 4003 5397 4012
rect 4928 3800 5296 3809
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 4928 3751 5296 3760
rect 4587 3548 4629 3557
rect 4587 3508 4588 3548
rect 4628 3508 4629 3548
rect 4587 3499 4629 3508
rect 4588 3414 4628 3499
rect 4780 3464 4820 3473
rect 4780 3305 4820 3424
rect 5356 3389 5396 4003
rect 5355 3380 5397 3389
rect 5355 3340 5356 3380
rect 5396 3340 5397 3380
rect 5355 3331 5397 3340
rect 4779 3296 4821 3305
rect 4779 3256 4780 3296
rect 4820 3256 4821 3296
rect 4779 3247 4821 3256
rect 4683 2876 4725 2885
rect 4683 2836 4684 2876
rect 4724 2836 4725 2876
rect 4683 2827 4725 2836
rect 4684 2624 4724 2827
rect 4684 2213 4724 2584
rect 5068 2624 5108 2633
rect 5068 2456 5108 2584
rect 5164 2624 5204 2633
rect 5356 2624 5396 3331
rect 5204 2584 5396 2624
rect 5164 2575 5204 2584
rect 5068 2416 5396 2456
rect 4928 2288 5296 2297
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 4928 2239 5296 2248
rect 4683 2204 4725 2213
rect 4683 2164 4684 2204
rect 4724 2164 4725 2204
rect 4683 2155 4725 2164
rect 4684 1868 4724 2155
rect 4684 1819 4724 1828
rect 5067 1868 5109 1877
rect 5067 1828 5068 1868
rect 5108 1828 5109 1868
rect 5067 1819 5109 1828
rect 4875 1784 4917 1793
rect 4875 1744 4876 1784
rect 4916 1744 4917 1784
rect 4875 1735 4917 1744
rect 4876 1650 4916 1735
rect 5068 1734 5108 1819
rect 5260 1700 5300 1709
rect 4492 1231 4532 1240
rect 3531 1196 3573 1205
rect 3531 1156 3532 1196
rect 3572 1156 3573 1196
rect 3531 1147 3573 1156
rect 3532 80 3572 1147
rect 3724 80 3764 1231
rect 5068 1196 5108 1205
rect 4107 1112 4149 1121
rect 4107 1072 4108 1112
rect 4148 1072 4149 1112
rect 4107 1063 4149 1072
rect 4300 1112 4340 1121
rect 4340 1072 4436 1112
rect 4300 1063 4340 1072
rect 3915 608 3957 617
rect 3915 568 3916 608
rect 3956 568 3957 608
rect 3915 559 3957 568
rect 3916 80 3956 559
rect 4108 80 4148 1063
rect 4299 944 4341 953
rect 4299 904 4300 944
rect 4340 904 4341 944
rect 4299 895 4341 904
rect 4300 80 4340 895
rect 4396 701 4436 1072
rect 4876 1037 4916 1122
rect 5068 1037 5108 1156
rect 5260 1121 5300 1660
rect 5259 1112 5301 1121
rect 5259 1072 5260 1112
rect 5300 1072 5301 1112
rect 5356 1112 5396 2416
rect 5452 2120 5492 5608
rect 5644 5648 5684 6187
rect 5836 6152 5876 6355
rect 6028 6354 6068 6439
rect 6124 6245 6164 6448
rect 6123 6236 6165 6245
rect 6123 6196 6124 6236
rect 6164 6196 6165 6236
rect 6123 6187 6165 6196
rect 5547 5480 5589 5489
rect 5547 5440 5548 5480
rect 5588 5440 5589 5480
rect 5547 5431 5589 5440
rect 5548 5346 5588 5431
rect 5644 4481 5684 5608
rect 5740 6112 5876 6152
rect 5740 5648 5780 6112
rect 6220 6068 6260 10051
rect 6316 9353 6356 11572
rect 6412 9437 6452 9522
rect 6411 9428 6453 9437
rect 6411 9388 6412 9428
rect 6452 9388 6453 9428
rect 6411 9379 6453 9388
rect 6508 9428 6548 11731
rect 6604 10109 6644 11908
rect 6795 11780 6837 11789
rect 6795 11740 6796 11780
rect 6836 11740 6837 11780
rect 6795 11731 6837 11740
rect 6796 11621 6836 11731
rect 6892 11701 6932 11710
rect 6795 11612 6837 11621
rect 6795 11572 6796 11612
rect 6836 11572 6837 11612
rect 6795 11563 6837 11572
rect 6699 11108 6741 11117
rect 6699 11068 6700 11108
rect 6740 11068 6741 11108
rect 6699 11059 6741 11068
rect 6700 10184 6740 11059
rect 6700 10135 6740 10144
rect 6603 10100 6645 10109
rect 6603 10060 6604 10100
rect 6644 10060 6645 10100
rect 6603 10051 6645 10060
rect 6315 9344 6357 9353
rect 6315 9304 6316 9344
rect 6356 9304 6357 9344
rect 6315 9295 6357 9304
rect 6411 9260 6453 9269
rect 6411 9220 6412 9260
rect 6452 9220 6453 9260
rect 6411 9211 6453 9220
rect 6315 9092 6357 9101
rect 6315 9052 6316 9092
rect 6356 9052 6357 9092
rect 6315 9043 6357 9052
rect 6316 7085 6356 9043
rect 6412 7160 6452 9211
rect 6508 9017 6548 9388
rect 6603 9428 6645 9437
rect 6603 9388 6604 9428
rect 6644 9388 6645 9428
rect 6603 9379 6645 9388
rect 6604 9101 6644 9379
rect 6796 9176 6836 11563
rect 6892 10436 6932 11661
rect 6988 11117 7028 13999
rect 7180 13208 7220 14671
rect 7275 14216 7317 14225
rect 7275 14176 7276 14216
rect 7316 14176 7317 14216
rect 7275 14167 7317 14176
rect 7276 14043 7316 14167
rect 7276 13994 7316 14003
rect 7372 13460 7412 17709
rect 7467 17744 7509 17753
rect 7467 17704 7468 17744
rect 7508 17704 7509 17744
rect 7467 17695 7509 17704
rect 7468 15728 7508 17695
rect 7563 17660 7605 17669
rect 7563 17620 7564 17660
rect 7604 17620 7605 17660
rect 7563 17611 7605 17620
rect 7564 17526 7604 17611
rect 7852 17249 7892 18628
rect 8139 18500 8181 18509
rect 8139 18460 8140 18500
rect 8180 18460 8181 18500
rect 8139 18451 8181 18460
rect 8043 17912 8085 17921
rect 8043 17872 8044 17912
rect 8084 17872 8085 17912
rect 8043 17863 8085 17872
rect 7948 17828 7988 17837
rect 7851 17240 7893 17249
rect 7756 17200 7852 17240
rect 7892 17200 7893 17240
rect 7564 16325 7604 16356
rect 7563 16316 7605 16325
rect 7563 16276 7564 16316
rect 7604 16276 7605 16316
rect 7563 16267 7605 16276
rect 7564 16232 7604 16267
rect 7564 16157 7604 16192
rect 7563 16148 7605 16157
rect 7563 16108 7564 16148
rect 7604 16108 7605 16148
rect 7563 16099 7605 16108
rect 7468 15679 7508 15688
rect 7564 15653 7604 16099
rect 7756 16073 7796 17200
rect 7851 17191 7893 17200
rect 7852 17072 7892 17081
rect 7755 16064 7797 16073
rect 7755 16024 7756 16064
rect 7796 16024 7797 16064
rect 7755 16015 7797 16024
rect 7852 15905 7892 17032
rect 7948 16409 7988 17788
rect 8044 17240 8084 17863
rect 8044 17191 8084 17200
rect 8140 17072 8180 18451
rect 8236 17492 8276 21568
rect 8331 19256 8373 19265
rect 8331 19216 8332 19256
rect 8372 19216 8373 19256
rect 8331 19207 8373 19216
rect 8332 17921 8372 19207
rect 8427 19172 8469 19181
rect 8427 19132 8428 19172
rect 8468 19132 8469 19172
rect 8427 19123 8469 19132
rect 8331 17912 8373 17921
rect 8331 17872 8332 17912
rect 8372 17872 8373 17912
rect 8331 17863 8373 17872
rect 8331 17744 8373 17753
rect 8331 17704 8332 17744
rect 8372 17704 8373 17744
rect 8331 17695 8373 17704
rect 8428 17744 8468 19123
rect 8332 17610 8372 17695
rect 8236 17452 8372 17492
rect 8235 17240 8277 17249
rect 8235 17200 8236 17240
rect 8276 17200 8277 17240
rect 8235 17191 8277 17200
rect 8044 17032 8180 17072
rect 8236 17072 8276 17191
rect 7947 16400 7989 16409
rect 7947 16360 7948 16400
rect 7988 16360 7989 16400
rect 7947 16351 7989 16360
rect 8044 16316 8084 17032
rect 8236 17023 8276 17032
rect 8235 16652 8277 16661
rect 8235 16612 8236 16652
rect 8276 16612 8277 16652
rect 8235 16603 8277 16612
rect 8044 16267 8084 16276
rect 8140 16232 8180 16241
rect 8140 16148 8180 16192
rect 8044 16108 8180 16148
rect 7851 15896 7893 15905
rect 7851 15856 7852 15896
rect 7892 15856 7893 15896
rect 7851 15847 7893 15856
rect 7563 15644 7605 15653
rect 7563 15604 7564 15644
rect 7604 15604 7605 15644
rect 7563 15595 7605 15604
rect 7660 15560 7700 15569
rect 7948 15560 7988 15569
rect 7700 15520 7796 15560
rect 7660 15511 7700 15520
rect 7660 15308 7700 15317
rect 7564 15268 7660 15308
rect 7467 14720 7509 14729
rect 7467 14680 7468 14720
rect 7508 14680 7509 14720
rect 7467 14671 7509 14680
rect 7468 14586 7508 14671
rect 7372 13411 7412 13420
rect 7468 14132 7508 14141
rect 7180 13159 7220 13168
rect 7468 12704 7508 14092
rect 7564 13469 7604 15268
rect 7660 15259 7700 15268
rect 7659 15140 7701 15149
rect 7659 15100 7660 15140
rect 7700 15100 7701 15140
rect 7659 15091 7701 15100
rect 7660 14972 7700 15091
rect 7660 14923 7700 14932
rect 7659 14468 7701 14477
rect 7659 14428 7660 14468
rect 7700 14428 7701 14468
rect 7659 14419 7701 14428
rect 7660 14048 7700 14419
rect 7756 14225 7796 15520
rect 7852 15520 7948 15560
rect 7755 14216 7797 14225
rect 7755 14176 7756 14216
rect 7796 14176 7797 14216
rect 7755 14167 7797 14176
rect 7756 14048 7796 14057
rect 7660 14008 7756 14048
rect 7756 13637 7796 14008
rect 7755 13628 7797 13637
rect 7755 13588 7756 13628
rect 7796 13588 7797 13628
rect 7755 13579 7797 13588
rect 7563 13460 7605 13469
rect 7563 13420 7564 13460
rect 7604 13420 7605 13460
rect 7563 13411 7605 13420
rect 7852 13385 7892 15520
rect 7948 15511 7988 15520
rect 8044 15401 8084 16108
rect 8236 15728 8276 16603
rect 8140 15688 8276 15728
rect 8043 15392 8085 15401
rect 8043 15352 8044 15392
rect 8084 15352 8085 15392
rect 8043 15343 8085 15352
rect 8140 14981 8180 15688
rect 8235 15560 8277 15569
rect 8332 15560 8372 17452
rect 8235 15520 8236 15560
rect 8276 15520 8372 15560
rect 8235 15511 8277 15520
rect 8236 15426 8276 15511
rect 8428 15392 8468 17704
rect 8524 16661 8564 22912
rect 8715 22912 8716 22952
rect 8756 22912 8757 22952
rect 8715 22903 8757 22912
rect 8619 22868 8661 22877
rect 8619 22828 8620 22868
rect 8660 22828 8661 22868
rect 8619 22819 8661 22828
rect 8620 19013 8660 22819
rect 8716 22818 8756 22903
rect 9004 22868 9044 23920
rect 9100 23624 9140 25264
rect 9196 25061 9236 25264
rect 9195 25052 9237 25061
rect 9195 25012 9196 25052
rect 9236 25012 9237 25052
rect 9195 25003 9237 25012
rect 9388 24977 9428 25432
rect 9484 25388 9524 25397
rect 9387 24968 9429 24977
rect 9387 24928 9388 24968
rect 9428 24928 9429 24968
rect 9484 24968 9524 25348
rect 9580 25304 9620 25313
rect 9620 25264 9716 25304
rect 9580 25255 9620 25264
rect 9484 24928 9620 24968
rect 9387 24919 9429 24928
rect 9484 24800 9524 24809
rect 9292 24760 9484 24800
rect 9292 24641 9332 24760
rect 9484 24751 9524 24760
rect 9291 24632 9333 24641
rect 9291 24592 9292 24632
rect 9332 24592 9333 24632
rect 9580 24632 9620 24928
rect 9291 24583 9333 24592
rect 9422 24617 9462 24626
rect 9196 24464 9236 24473
rect 9422 24464 9462 24577
rect 9236 24424 9462 24464
rect 9196 24415 9236 24424
rect 9580 24380 9620 24592
rect 9484 24340 9620 24380
rect 9676 24632 9716 25264
rect 9195 24296 9237 24305
rect 9195 24256 9196 24296
rect 9236 24256 9237 24296
rect 9195 24247 9237 24256
rect 9196 23792 9236 24247
rect 9291 24212 9333 24221
rect 9291 24172 9292 24212
rect 9332 24172 9333 24212
rect 9291 24163 9333 24172
rect 9196 23743 9236 23752
rect 9292 23792 9332 24163
rect 9387 24044 9429 24053
rect 9387 24004 9388 24044
rect 9428 24004 9429 24044
rect 9387 23995 9429 24004
rect 9100 23584 9236 23624
rect 9099 23120 9141 23129
rect 9099 23080 9100 23120
rect 9140 23080 9141 23120
rect 9099 23071 9141 23080
rect 9100 22986 9140 23071
rect 8812 22828 9044 22868
rect 8715 22700 8757 22709
rect 8715 22660 8716 22700
rect 8756 22660 8757 22700
rect 8715 22651 8757 22660
rect 8716 22280 8756 22651
rect 8812 22364 8852 22828
rect 9003 22700 9045 22709
rect 9003 22660 9004 22700
rect 9044 22660 9045 22700
rect 9003 22651 9045 22660
rect 8812 22315 8852 22324
rect 8908 22448 8948 22457
rect 8716 22231 8756 22240
rect 8715 22112 8757 22121
rect 8715 22072 8716 22112
rect 8756 22072 8757 22112
rect 8715 22063 8757 22072
rect 8619 19004 8661 19013
rect 8619 18964 8620 19004
rect 8660 18964 8661 19004
rect 8619 18955 8661 18964
rect 8523 16652 8565 16661
rect 8523 16612 8524 16652
rect 8564 16612 8565 16652
rect 8523 16603 8565 16612
rect 8620 16484 8660 18955
rect 8524 16444 8660 16484
rect 8524 16232 8564 16444
rect 8524 15989 8564 16192
rect 8620 16232 8660 16241
rect 8523 15980 8565 15989
rect 8523 15940 8524 15980
rect 8564 15940 8565 15980
rect 8523 15931 8565 15940
rect 8620 15737 8660 16192
rect 8619 15728 8661 15737
rect 8619 15688 8620 15728
rect 8660 15688 8661 15728
rect 8619 15679 8661 15688
rect 8619 15560 8661 15569
rect 8619 15520 8620 15560
rect 8660 15520 8661 15560
rect 8619 15511 8661 15520
rect 8332 15352 8468 15392
rect 8139 14972 8181 14981
rect 8139 14932 8140 14972
rect 8180 14932 8181 14972
rect 8139 14923 8181 14932
rect 7948 14720 7988 14729
rect 7851 13376 7893 13385
rect 7851 13336 7852 13376
rect 7892 13336 7893 13376
rect 7851 13327 7893 13336
rect 7372 12664 7508 12704
rect 7564 13208 7604 13217
rect 7275 11864 7317 11873
rect 7275 11824 7276 11864
rect 7316 11824 7317 11864
rect 7275 11815 7317 11824
rect 7276 11696 7316 11815
rect 7372 11696 7412 12664
rect 7468 12536 7508 12547
rect 7468 12461 7508 12496
rect 7467 12452 7509 12461
rect 7467 12412 7468 12452
rect 7508 12412 7509 12452
rect 7467 12403 7509 12412
rect 7564 12452 7604 13168
rect 7756 13208 7796 13217
rect 7659 13040 7701 13049
rect 7659 13000 7660 13040
rect 7700 13000 7701 13040
rect 7659 12991 7701 13000
rect 7660 12906 7700 12991
rect 7756 12629 7796 13168
rect 7852 13208 7892 13217
rect 7755 12620 7797 12629
rect 7755 12580 7756 12620
rect 7796 12580 7797 12620
rect 7755 12571 7797 12580
rect 7852 12545 7892 13168
rect 7851 12536 7893 12545
rect 7851 12496 7852 12536
rect 7892 12496 7893 12536
rect 7851 12487 7893 12496
rect 7564 12412 7796 12452
rect 7467 12032 7509 12041
rect 7467 11992 7468 12032
rect 7508 11992 7509 12032
rect 7467 11983 7509 11992
rect 7468 11948 7508 11983
rect 7468 11897 7508 11908
rect 7468 11696 7508 11705
rect 7372 11656 7468 11696
rect 7276 11647 7316 11656
rect 7468 11647 7508 11656
rect 7084 11528 7124 11537
rect 6987 11108 7029 11117
rect 6987 11068 6988 11108
rect 7028 11068 7029 11108
rect 6987 11059 7029 11068
rect 6892 10387 6932 10396
rect 6891 10268 6933 10277
rect 6891 10228 6892 10268
rect 6932 10228 6933 10268
rect 6891 10219 6933 10228
rect 6700 9136 6836 9176
rect 6603 9092 6645 9101
rect 6603 9052 6604 9092
rect 6644 9052 6645 9092
rect 6603 9043 6645 9052
rect 6507 9008 6549 9017
rect 6507 8968 6508 9008
rect 6548 8968 6549 9008
rect 6507 8959 6549 8968
rect 6700 8840 6740 9136
rect 6795 9008 6837 9017
rect 6795 8968 6796 9008
rect 6836 8968 6837 9008
rect 6795 8959 6837 8968
rect 6796 8924 6836 8959
rect 6796 8873 6836 8884
rect 6508 8800 6740 8840
rect 6508 7337 6548 8800
rect 6604 8672 6644 8681
rect 6699 8672 6741 8681
rect 6644 8632 6700 8672
rect 6740 8632 6741 8672
rect 6604 8623 6644 8632
rect 6699 8623 6741 8632
rect 6603 8168 6645 8177
rect 6603 8128 6604 8168
rect 6644 8128 6645 8168
rect 6603 8119 6645 8128
rect 6507 7328 6549 7337
rect 6507 7288 6508 7328
rect 6548 7288 6549 7328
rect 6507 7279 6549 7288
rect 6508 7160 6548 7169
rect 6412 7120 6508 7160
rect 6315 7076 6357 7085
rect 6315 7036 6316 7076
rect 6356 7036 6357 7076
rect 6315 7027 6357 7036
rect 6316 6749 6356 7027
rect 6315 6740 6357 6749
rect 6315 6700 6316 6740
rect 6356 6700 6357 6740
rect 6315 6691 6357 6700
rect 6412 6665 6452 7120
rect 6508 7111 6548 7120
rect 6507 6824 6549 6833
rect 6507 6784 6508 6824
rect 6548 6784 6549 6824
rect 6507 6775 6549 6784
rect 6411 6656 6453 6665
rect 6411 6616 6412 6656
rect 6452 6616 6453 6656
rect 6411 6607 6453 6616
rect 6508 6656 6548 6775
rect 6508 6607 6548 6616
rect 6412 6488 6452 6497
rect 6604 6488 6644 8119
rect 6700 8000 6740 8623
rect 6700 7925 6740 7960
rect 6796 8504 6836 8513
rect 6699 7916 6741 7925
rect 6699 7876 6700 7916
rect 6740 7876 6741 7916
rect 6699 7867 6741 7876
rect 6796 7505 6836 8464
rect 6892 7925 6932 10219
rect 6988 9512 7028 11059
rect 7084 10529 7124 11488
rect 7564 11453 7604 12412
rect 7756 12368 7796 12412
rect 7852 12368 7892 12377
rect 7756 12328 7852 12368
rect 7852 12319 7892 12328
rect 7660 12284 7700 12293
rect 7660 12116 7700 12244
rect 7948 12116 7988 14680
rect 8044 14720 8084 14729
rect 8332 14720 8372 15352
rect 8084 14680 8372 14720
rect 8044 14671 8084 14680
rect 8139 13796 8181 13805
rect 8139 13756 8140 13796
rect 8180 13756 8181 13796
rect 8139 13747 8181 13756
rect 8140 13208 8180 13747
rect 8140 13133 8180 13168
rect 8139 13124 8181 13133
rect 8139 13084 8140 13124
rect 8180 13084 8181 13124
rect 8139 13075 8181 13084
rect 8140 13044 8180 13075
rect 8235 12620 8277 12629
rect 8235 12580 8236 12620
rect 8276 12580 8277 12620
rect 8235 12571 8277 12580
rect 8044 12536 8084 12545
rect 8084 12496 8180 12536
rect 8044 12487 8084 12496
rect 7660 12076 7988 12116
rect 7659 11948 7701 11957
rect 7659 11908 7660 11948
rect 7700 11908 7701 11948
rect 7659 11899 7701 11908
rect 7660 11814 7700 11899
rect 7852 11696 7892 11705
rect 7660 11528 7700 11537
rect 7563 11444 7605 11453
rect 7563 11404 7564 11444
rect 7604 11404 7605 11444
rect 7563 11395 7605 11404
rect 7179 11360 7221 11369
rect 7179 11320 7180 11360
rect 7220 11320 7221 11360
rect 7179 11311 7221 11320
rect 7180 11024 7220 11311
rect 7180 10975 7220 10984
rect 7371 11024 7413 11033
rect 7371 10984 7372 11024
rect 7412 10984 7413 11024
rect 7371 10975 7413 10984
rect 7372 10890 7412 10975
rect 7083 10520 7125 10529
rect 7083 10480 7084 10520
rect 7124 10480 7125 10520
rect 7083 10471 7125 10480
rect 7179 10352 7221 10361
rect 7179 10312 7180 10352
rect 7220 10312 7221 10352
rect 7179 10303 7221 10312
rect 7180 10184 7220 10303
rect 7467 10268 7509 10277
rect 7467 10228 7468 10268
rect 7508 10228 7509 10268
rect 7467 10219 7509 10228
rect 7180 10135 7220 10144
rect 7276 10184 7316 10193
rect 7276 10109 7316 10144
rect 7372 10184 7412 10193
rect 7275 10100 7317 10109
rect 7275 10060 7276 10100
rect 7316 10060 7317 10100
rect 7275 10051 7317 10060
rect 6988 9269 7028 9472
rect 7083 9512 7125 9521
rect 7083 9472 7084 9512
rect 7124 9472 7125 9512
rect 7083 9463 7125 9472
rect 6987 9260 7029 9269
rect 6987 9220 6988 9260
rect 7028 9220 7029 9260
rect 6987 9211 7029 9220
rect 6988 8924 7028 8933
rect 7084 8924 7124 9463
rect 7028 8884 7124 8924
rect 6988 8875 7028 8884
rect 7276 8840 7316 10051
rect 7084 8800 7316 8840
rect 6988 8504 7028 8513
rect 6891 7916 6933 7925
rect 6891 7876 6892 7916
rect 6932 7876 6933 7916
rect 6891 7867 6933 7876
rect 6988 7832 7028 8464
rect 7084 8000 7124 8800
rect 7179 8672 7221 8681
rect 7179 8632 7180 8672
rect 7220 8632 7221 8672
rect 7179 8623 7221 8632
rect 7180 8538 7220 8623
rect 7276 8168 7316 8177
rect 7372 8168 7412 10144
rect 7468 10184 7508 10219
rect 7660 10184 7700 11488
rect 7852 11285 7892 11656
rect 7947 11444 7989 11453
rect 7947 11404 7948 11444
rect 7988 11404 7989 11444
rect 7947 11395 7989 11404
rect 7851 11276 7893 11285
rect 7851 11236 7852 11276
rect 7892 11236 7893 11276
rect 7851 11227 7893 11236
rect 7852 10613 7892 11227
rect 7851 10604 7893 10613
rect 7851 10564 7852 10604
rect 7892 10564 7893 10604
rect 7851 10555 7893 10564
rect 7948 10352 7988 11395
rect 8140 11285 8180 12496
rect 8236 12041 8276 12571
rect 8235 12032 8277 12041
rect 8235 11992 8236 12032
rect 8276 11992 8277 12032
rect 8235 11983 8277 11992
rect 8139 11276 8181 11285
rect 8139 11236 8140 11276
rect 8180 11236 8181 11276
rect 8139 11227 8181 11236
rect 8139 10772 8181 10781
rect 8139 10732 8140 10772
rect 8180 10732 8181 10772
rect 8139 10723 8181 10732
rect 8140 10529 8180 10723
rect 8139 10520 8181 10529
rect 8139 10480 8140 10520
rect 8180 10480 8181 10520
rect 8139 10471 8181 10480
rect 7948 10312 8084 10352
rect 7468 10133 7508 10144
rect 7564 10144 7660 10184
rect 7468 9498 7508 9507
rect 7468 9017 7508 9458
rect 7467 9008 7509 9017
rect 7467 8968 7468 9008
rect 7508 8968 7509 9008
rect 7467 8959 7509 8968
rect 7564 8840 7604 10144
rect 7660 10135 7700 10144
rect 7756 10184 7796 10193
rect 7756 9764 7796 10144
rect 7947 10184 7989 10193
rect 7947 10144 7948 10184
rect 7988 10144 7989 10184
rect 7947 10135 7989 10144
rect 7948 10016 7988 10135
rect 7948 9967 7988 9976
rect 8044 9773 8084 10312
rect 8140 10184 8180 10471
rect 8332 10361 8372 14680
rect 8428 14720 8468 14729
rect 8428 14561 8468 14680
rect 8524 14720 8564 14731
rect 8524 14645 8564 14680
rect 8523 14636 8565 14645
rect 8523 14596 8524 14636
rect 8564 14596 8565 14636
rect 8523 14587 8565 14596
rect 8427 14552 8469 14561
rect 8427 14512 8428 14552
rect 8468 14512 8469 14552
rect 8427 14503 8469 14512
rect 8428 14057 8468 14503
rect 8523 14384 8565 14393
rect 8523 14344 8524 14384
rect 8564 14344 8565 14384
rect 8523 14335 8565 14344
rect 8427 14048 8469 14057
rect 8427 14008 8428 14048
rect 8468 14008 8469 14048
rect 8427 13999 8469 14008
rect 8427 13124 8469 13133
rect 8427 13084 8428 13124
rect 8468 13084 8469 13124
rect 8427 13075 8469 13084
rect 8331 10352 8373 10361
rect 8331 10312 8332 10352
rect 8372 10312 8373 10352
rect 8331 10303 8373 10312
rect 8140 10135 8180 10144
rect 8331 9932 8373 9941
rect 8331 9892 8332 9932
rect 8372 9892 8373 9932
rect 8331 9883 8373 9892
rect 8043 9764 8085 9773
rect 7756 9724 7988 9764
rect 7660 9596 7700 9605
rect 7700 9556 7892 9596
rect 7660 9547 7700 9556
rect 7852 9512 7892 9556
rect 7852 9463 7892 9472
rect 7659 9428 7701 9437
rect 7659 9388 7660 9428
rect 7700 9388 7701 9428
rect 7659 9379 7701 9388
rect 7316 8128 7412 8168
rect 7468 8800 7604 8840
rect 7276 8119 7316 8128
rect 7180 8009 7220 8094
rect 7084 7951 7124 7960
rect 7179 8000 7221 8009
rect 7179 7960 7180 8000
rect 7220 7960 7221 8000
rect 7179 7951 7221 7960
rect 7372 8000 7412 8009
rect 7468 8000 7508 8800
rect 7660 8756 7700 9379
rect 7948 9344 7988 9724
rect 8043 9724 8044 9764
rect 8084 9724 8085 9764
rect 8043 9715 8085 9724
rect 8044 9521 8084 9606
rect 8043 9512 8085 9521
rect 8043 9472 8044 9512
rect 8084 9472 8085 9512
rect 8043 9463 8085 9472
rect 8236 9344 8276 9353
rect 7948 9304 8236 9344
rect 8236 9295 8276 9304
rect 7412 7960 7508 8000
rect 7564 8716 7700 8756
rect 7852 9260 7892 9269
rect 7564 8000 7604 8716
rect 7372 7951 7412 7960
rect 7564 7951 7604 7960
rect 7179 7832 7221 7841
rect 6988 7792 7124 7832
rect 6892 7748 6932 7757
rect 6932 7708 7028 7748
rect 6892 7699 6932 7708
rect 6795 7496 6837 7505
rect 6795 7456 6796 7496
rect 6836 7456 6837 7496
rect 6795 7447 6837 7456
rect 6699 7328 6741 7337
rect 6699 7288 6700 7328
rect 6740 7288 6741 7328
rect 6699 7279 6741 7288
rect 6700 7169 6740 7279
rect 6988 7174 7028 7708
rect 6699 7160 6741 7169
rect 6699 7120 6700 7160
rect 6740 7120 6741 7160
rect 6988 7125 7028 7134
rect 6699 7111 6741 7120
rect 6028 6028 6260 6068
rect 6316 6448 6412 6488
rect 5835 5732 5877 5741
rect 5835 5692 5836 5732
rect 5876 5692 5877 5732
rect 5835 5683 5877 5692
rect 5740 5599 5780 5608
rect 5739 5396 5781 5405
rect 5739 5356 5740 5396
rect 5780 5356 5781 5396
rect 5739 5347 5781 5356
rect 5643 4472 5685 4481
rect 5643 4432 5644 4472
rect 5684 4432 5685 4472
rect 5643 4423 5685 4432
rect 5644 3389 5684 4423
rect 5740 3968 5780 5347
rect 5836 4976 5876 5683
rect 5932 5648 5972 5657
rect 5932 5489 5972 5608
rect 5931 5480 5973 5489
rect 5931 5440 5932 5480
rect 5972 5440 5973 5480
rect 5931 5431 5973 5440
rect 5932 4976 5972 4985
rect 5836 4936 5932 4976
rect 5932 4927 5972 4936
rect 5835 4388 5877 4397
rect 5835 4348 5836 4388
rect 5876 4348 5877 4388
rect 5835 4339 5877 4348
rect 5836 4229 5876 4339
rect 5835 4220 5877 4229
rect 5835 4180 5836 4220
rect 5876 4180 5877 4220
rect 5835 4171 5877 4180
rect 5836 4136 5876 4171
rect 6028 4136 6068 6028
rect 6220 5900 6260 5909
rect 6316 5900 6356 6448
rect 6412 6439 6452 6448
rect 6508 6448 6604 6488
rect 6508 6320 6548 6448
rect 6604 6439 6644 6448
rect 6700 6488 6740 7111
rect 7084 7076 7124 7792
rect 7179 7792 7180 7832
rect 7220 7792 7221 7832
rect 7179 7783 7221 7792
rect 6988 7036 7124 7076
rect 7180 7076 7220 7783
rect 7275 7496 7317 7505
rect 7275 7456 7276 7496
rect 7316 7456 7317 7496
rect 7275 7447 7317 7456
rect 6891 6572 6933 6581
rect 6891 6532 6892 6572
rect 6932 6532 6933 6572
rect 6891 6523 6933 6532
rect 6700 6439 6740 6448
rect 6892 6438 6932 6523
rect 6988 6488 7028 7036
rect 7180 7027 7220 7036
rect 7276 6908 7316 7447
rect 7852 7253 7892 9220
rect 8332 9008 8372 9883
rect 8044 8968 8372 9008
rect 7851 7244 7893 7253
rect 7851 7204 7852 7244
rect 7892 7204 7893 7244
rect 7851 7195 7893 7204
rect 7467 7160 7509 7169
rect 7467 7120 7468 7160
rect 7508 7120 7509 7160
rect 7372 7085 7412 7116
rect 7467 7111 7509 7120
rect 7564 7160 7604 7169
rect 7371 7076 7413 7085
rect 7371 7036 7372 7076
rect 7412 7036 7413 7076
rect 7371 7027 7413 7036
rect 7180 6868 7316 6908
rect 7372 6992 7412 7027
rect 7083 6824 7125 6833
rect 7083 6784 7084 6824
rect 7124 6784 7125 6824
rect 7083 6775 7125 6784
rect 6988 6439 7028 6448
rect 7084 6488 7124 6775
rect 7084 6439 7124 6448
rect 7180 6488 7220 6868
rect 7372 6749 7412 6952
rect 7468 6833 7508 7111
rect 7467 6824 7509 6833
rect 7467 6784 7468 6824
rect 7508 6784 7509 6824
rect 7467 6775 7509 6784
rect 7564 6749 7604 7120
rect 7659 7160 7701 7169
rect 7659 7120 7660 7160
rect 7700 7120 7701 7160
rect 7659 7111 7701 7120
rect 7371 6740 7413 6749
rect 7371 6700 7372 6740
rect 7412 6700 7413 6740
rect 7371 6691 7413 6700
rect 7563 6740 7605 6749
rect 7563 6700 7564 6740
rect 7604 6700 7605 6740
rect 7563 6691 7605 6700
rect 7275 6656 7317 6665
rect 7275 6616 7276 6656
rect 7316 6616 7317 6656
rect 7275 6607 7317 6616
rect 7180 6320 7220 6448
rect 6260 5860 6356 5900
rect 6412 6280 6548 6320
rect 6604 6280 7220 6320
rect 6220 5851 6260 5860
rect 6220 5648 6260 5657
rect 6412 5648 6452 6280
rect 6507 5984 6549 5993
rect 6507 5944 6508 5984
rect 6548 5944 6549 5984
rect 6507 5935 6549 5944
rect 6260 5608 6412 5648
rect 6220 5599 6260 5608
rect 6412 5599 6452 5608
rect 6508 5648 6548 5935
rect 6508 5599 6548 5608
rect 6604 5648 6644 6280
rect 6699 6152 6741 6161
rect 6699 6112 6700 6152
rect 6740 6112 6741 6152
rect 6699 6103 6741 6112
rect 6891 6152 6933 6161
rect 7276 6152 7316 6607
rect 7467 6572 7509 6581
rect 7372 6532 7468 6572
rect 7508 6532 7509 6572
rect 7372 6488 7412 6532
rect 7467 6523 7509 6532
rect 7372 6439 7412 6448
rect 7467 6404 7509 6413
rect 7467 6364 7468 6404
rect 7508 6364 7509 6404
rect 7467 6355 7509 6364
rect 7660 6404 7700 7111
rect 7947 6572 7989 6581
rect 7947 6532 7948 6572
rect 7988 6532 7989 6572
rect 7947 6523 7989 6532
rect 7756 6488 7796 6497
rect 7796 6448 7892 6488
rect 7756 6439 7796 6448
rect 7660 6355 7700 6364
rect 7371 6320 7413 6329
rect 7371 6280 7372 6320
rect 7412 6280 7413 6320
rect 7371 6271 7413 6280
rect 6891 6112 6892 6152
rect 6932 6112 6933 6152
rect 6891 6103 6933 6112
rect 6988 6112 7316 6152
rect 6604 5599 6644 5608
rect 6700 5648 6740 6103
rect 6795 6068 6837 6077
rect 6795 6028 6796 6068
rect 6836 6028 6837 6068
rect 6795 6019 6837 6028
rect 6700 5599 6740 5608
rect 6411 5480 6453 5489
rect 6411 5440 6412 5480
rect 6452 5440 6453 5480
rect 6411 5431 6453 5440
rect 6699 5480 6741 5489
rect 6699 5440 6700 5480
rect 6740 5440 6741 5480
rect 6699 5431 6741 5440
rect 6123 5060 6165 5069
rect 6123 5020 6124 5060
rect 6164 5020 6165 5060
rect 6123 5011 6165 5020
rect 6124 4926 6164 5011
rect 6316 4976 6356 4985
rect 6316 4817 6356 4936
rect 6315 4808 6357 4817
rect 6315 4768 6316 4808
rect 6356 4768 6357 4808
rect 6315 4759 6357 4768
rect 6220 4145 6260 4230
rect 6315 4220 6357 4229
rect 6315 4180 6316 4220
rect 6356 4180 6357 4220
rect 6315 4171 6357 4180
rect 6219 4136 6261 4145
rect 6028 4096 6164 4136
rect 5836 4086 5876 4096
rect 6028 3968 6068 3977
rect 5740 3928 6028 3968
rect 6124 3968 6164 4096
rect 6219 4096 6220 4136
rect 6260 4096 6261 4136
rect 6219 4087 6261 4096
rect 6316 4136 6356 4171
rect 6316 4085 6356 4096
rect 6412 4136 6452 5431
rect 6603 5228 6645 5237
rect 6603 5188 6604 5228
rect 6644 5188 6645 5228
rect 6603 5179 6645 5188
rect 6507 4388 6549 4397
rect 6507 4348 6508 4388
rect 6548 4348 6549 4388
rect 6507 4339 6549 4348
rect 6412 4087 6452 4096
rect 6508 4136 6548 4339
rect 6508 4087 6548 4096
rect 6604 3968 6644 5179
rect 6124 3928 6260 3968
rect 5739 3800 5781 3809
rect 5739 3760 5740 3800
rect 5780 3760 5781 3800
rect 5739 3751 5781 3760
rect 5643 3380 5685 3389
rect 5643 3340 5644 3380
rect 5684 3340 5685 3380
rect 5643 3331 5685 3340
rect 5548 2633 5588 2718
rect 5644 2708 5684 2717
rect 5740 2708 5780 3751
rect 5684 2668 5780 2708
rect 5644 2659 5684 2668
rect 5547 2624 5589 2633
rect 5547 2584 5548 2624
rect 5588 2584 5589 2624
rect 5547 2575 5589 2584
rect 5836 2540 5876 3928
rect 6028 3919 6068 3928
rect 6027 3800 6069 3809
rect 6027 3760 6028 3800
rect 6068 3760 6069 3800
rect 6027 3751 6069 3760
rect 6028 3464 6068 3751
rect 5931 3380 5973 3389
rect 5931 3340 5932 3380
rect 5972 3340 5973 3380
rect 5931 3331 5973 3340
rect 5644 2500 5876 2540
rect 5644 2456 5684 2500
rect 5932 2456 5972 3331
rect 5452 2071 5492 2080
rect 5548 2416 5684 2456
rect 5740 2416 5972 2456
rect 5548 1952 5588 2416
rect 5643 2288 5685 2297
rect 5643 2248 5644 2288
rect 5684 2248 5685 2288
rect 5643 2239 5685 2248
rect 5548 1903 5588 1912
rect 5644 1952 5684 2239
rect 5644 1903 5684 1912
rect 5740 1952 5780 2416
rect 6028 2381 6068 3424
rect 6124 2633 6164 2718
rect 6123 2624 6165 2633
rect 6123 2584 6124 2624
rect 6164 2584 6165 2624
rect 6123 2575 6165 2584
rect 6027 2372 6069 2381
rect 6027 2332 6028 2372
rect 6068 2332 6069 2372
rect 6027 2323 6069 2332
rect 5740 1903 5780 1912
rect 5931 1952 5973 1961
rect 5931 1912 5932 1952
rect 5972 1912 5973 1952
rect 5931 1903 5973 1912
rect 5932 1818 5972 1903
rect 5739 1532 5781 1541
rect 5739 1492 5740 1532
rect 5780 1492 5781 1532
rect 5739 1483 5781 1492
rect 5643 1196 5685 1205
rect 5643 1156 5644 1196
rect 5684 1156 5685 1196
rect 5643 1147 5685 1156
rect 5356 1072 5588 1112
rect 5259 1063 5301 1072
rect 4875 1028 4917 1037
rect 4875 988 4876 1028
rect 4916 988 4917 1028
rect 4875 979 4917 988
rect 5067 1028 5109 1037
rect 5067 988 5068 1028
rect 5108 988 5109 1028
rect 5067 979 5109 988
rect 5260 944 5300 953
rect 5451 944 5493 953
rect 5300 904 5396 944
rect 5260 895 5300 904
rect 5356 785 5396 904
rect 5451 904 5452 944
rect 5492 904 5493 944
rect 5451 895 5493 904
rect 5452 810 5492 895
rect 4683 776 4725 785
rect 4683 736 4684 776
rect 4724 736 4725 776
rect 4683 727 4725 736
rect 4928 776 5296 785
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 4928 727 5296 736
rect 5355 776 5397 785
rect 5355 736 5356 776
rect 5396 736 5397 776
rect 5355 727 5397 736
rect 4395 692 4437 701
rect 4395 652 4396 692
rect 4436 652 4437 692
rect 4395 643 4437 652
rect 4491 272 4533 281
rect 4491 232 4492 272
rect 4532 232 4533 272
rect 4491 223 4533 232
rect 4492 80 4532 223
rect 4684 80 4724 727
rect 5067 608 5109 617
rect 5067 568 5068 608
rect 5108 568 5109 608
rect 5067 559 5109 568
rect 4875 356 4917 365
rect 4875 316 4876 356
rect 4916 316 4917 356
rect 4875 307 4917 316
rect 4876 80 4916 307
rect 5068 80 5108 559
rect 5548 533 5588 1072
rect 5644 1062 5684 1147
rect 5740 944 5780 1483
rect 5835 1280 5877 1289
rect 5835 1240 5836 1280
rect 5876 1240 5877 1280
rect 5835 1231 5877 1240
rect 5836 1146 5876 1231
rect 6123 1196 6165 1205
rect 6123 1156 6124 1196
rect 6164 1156 6165 1196
rect 6123 1147 6165 1156
rect 6124 1112 6164 1147
rect 6124 1061 6164 1072
rect 5644 904 5780 944
rect 5547 524 5589 533
rect 5547 484 5548 524
rect 5588 484 5589 524
rect 5547 475 5589 484
rect 5451 272 5493 281
rect 5451 232 5452 272
rect 5492 232 5493 272
rect 5451 223 5493 232
rect 5259 188 5301 197
rect 5259 148 5260 188
rect 5300 148 5301 188
rect 5259 139 5301 148
rect 5260 80 5300 139
rect 5452 80 5492 223
rect 5644 80 5684 904
rect 5835 860 5877 869
rect 5835 820 5836 860
rect 5876 820 5877 860
rect 5835 811 5877 820
rect 5836 80 5876 811
rect 6027 104 6069 113
rect 6027 80 6028 104
rect 1784 0 1864 80
rect 1976 0 2056 80
rect 2168 0 2248 80
rect 2360 0 2440 80
rect 2552 0 2632 80
rect 2744 0 2824 80
rect 2936 0 3016 80
rect 3128 0 3208 80
rect 3320 0 3400 80
rect 3512 0 3592 80
rect 3704 0 3784 80
rect 3896 0 3976 80
rect 4088 0 4168 80
rect 4280 0 4360 80
rect 4472 0 4552 80
rect 4664 0 4744 80
rect 4856 0 4936 80
rect 5048 0 5128 80
rect 5240 0 5320 80
rect 5432 0 5512 80
rect 5624 0 5704 80
rect 5816 0 5896 80
rect 6008 64 6028 80
rect 6068 80 6069 104
rect 6220 80 6260 3928
rect 6316 3928 6644 3968
rect 6316 3464 6356 3928
rect 6412 3632 6452 3641
rect 6700 3632 6740 5431
rect 6796 5237 6836 6019
rect 6892 5648 6932 6103
rect 6892 5599 6932 5608
rect 6795 5228 6837 5237
rect 6795 5188 6796 5228
rect 6836 5188 6837 5228
rect 6795 5179 6837 5188
rect 6988 5060 7028 6112
rect 7275 5984 7317 5993
rect 7275 5944 7276 5984
rect 7316 5944 7317 5984
rect 7275 5935 7317 5944
rect 7179 5564 7221 5573
rect 7179 5524 7180 5564
rect 7220 5524 7221 5564
rect 7179 5515 7221 5524
rect 6796 5020 7028 5060
rect 6796 4397 6836 5020
rect 6891 4892 6933 4901
rect 6891 4852 6892 4892
rect 6932 4852 6933 4892
rect 6891 4843 6933 4852
rect 6795 4388 6837 4397
rect 6795 4348 6796 4388
rect 6836 4348 6837 4388
rect 6795 4339 6837 4348
rect 6452 3592 6740 3632
rect 6796 4136 6836 4145
rect 6412 3583 6452 3592
rect 6316 3415 6356 3424
rect 6508 3464 6548 3475
rect 6508 3389 6548 3424
rect 6604 3464 6644 3473
rect 6796 3464 6836 4096
rect 6892 4136 6932 4843
rect 7083 4808 7125 4817
rect 7083 4768 7084 4808
rect 7124 4768 7125 4808
rect 7083 4759 7125 4768
rect 6987 4640 7029 4649
rect 6987 4600 6988 4640
rect 7028 4600 7029 4640
rect 6987 4591 7029 4600
rect 6892 4087 6932 4096
rect 6892 3464 6932 3473
rect 6796 3424 6892 3464
rect 6507 3380 6549 3389
rect 6507 3340 6508 3380
rect 6548 3340 6549 3380
rect 6507 3331 6549 3340
rect 6604 3380 6644 3424
rect 6699 3380 6741 3389
rect 6604 3340 6700 3380
rect 6740 3340 6741 3380
rect 6604 3137 6644 3340
rect 6699 3331 6741 3340
rect 6603 3128 6645 3137
rect 6603 3088 6604 3128
rect 6644 3088 6645 3128
rect 6603 3079 6645 3088
rect 6604 2633 6644 2719
rect 6603 2629 6645 2633
rect 6603 2584 6604 2629
rect 6644 2584 6645 2629
rect 6603 2575 6645 2584
rect 6795 2540 6837 2549
rect 6795 2500 6796 2540
rect 6836 2500 6837 2540
rect 6795 2491 6837 2500
rect 6796 2406 6836 2491
rect 6892 1938 6932 3424
rect 6988 3464 7028 4591
rect 6988 3415 7028 3424
rect 7084 3305 7124 4759
rect 7083 3296 7125 3305
rect 7083 3256 7084 3296
rect 7124 3256 7125 3296
rect 7083 3247 7125 3256
rect 7180 3128 7220 5515
rect 7084 3088 7220 3128
rect 7276 4220 7316 5935
rect 6987 2708 7029 2717
rect 6987 2668 6988 2708
rect 7028 2668 7029 2708
rect 6987 2659 7029 2668
rect 6988 2574 7028 2659
rect 7084 2204 7124 3088
rect 7179 2456 7221 2465
rect 7179 2416 7180 2456
rect 7220 2416 7221 2456
rect 7179 2407 7221 2416
rect 7180 2322 7220 2407
rect 7276 2297 7316 4180
rect 7372 4220 7412 6271
rect 7468 6270 7508 6355
rect 7852 6329 7892 6448
rect 7947 6474 7987 6523
rect 7947 6434 7988 6474
rect 7563 6320 7605 6329
rect 7563 6280 7564 6320
rect 7604 6280 7605 6320
rect 7563 6271 7605 6280
rect 7851 6320 7893 6329
rect 7851 6280 7852 6320
rect 7892 6280 7893 6320
rect 7851 6271 7893 6280
rect 7948 6320 7988 6434
rect 7948 6271 7988 6280
rect 7564 6186 7604 6271
rect 7659 6152 7701 6161
rect 7659 6112 7660 6152
rect 7700 6112 7701 6152
rect 7659 6103 7701 6112
rect 7467 5984 7509 5993
rect 7467 5944 7468 5984
rect 7508 5944 7509 5984
rect 7467 5935 7509 5944
rect 7372 4171 7412 4180
rect 7371 3968 7413 3977
rect 7371 3928 7372 3968
rect 7412 3928 7413 3968
rect 7371 3919 7413 3928
rect 7372 3380 7412 3919
rect 7372 3137 7412 3340
rect 7468 3464 7508 5935
rect 7660 5405 7700 6103
rect 8044 5648 8084 8968
rect 8428 8840 8468 13075
rect 8524 11705 8564 14335
rect 8523 11696 8565 11705
rect 8523 11656 8524 11696
rect 8564 11656 8565 11696
rect 8523 11647 8565 11656
rect 8524 10436 8564 11647
rect 8620 11360 8660 15511
rect 8716 12629 8756 22063
rect 8811 21608 8853 21617
rect 8811 21568 8812 21608
rect 8852 21568 8853 21608
rect 8811 21559 8853 21568
rect 8812 17921 8852 21559
rect 8908 21533 8948 22408
rect 9004 22364 9044 22651
rect 9099 22616 9141 22625
rect 9099 22576 9100 22616
rect 9140 22576 9141 22616
rect 9099 22567 9141 22576
rect 9004 22315 9044 22324
rect 9100 22280 9140 22567
rect 9100 22231 9140 22240
rect 9196 21953 9236 23584
rect 9292 23381 9332 23752
rect 9291 23372 9333 23381
rect 9291 23332 9292 23372
rect 9332 23332 9333 23372
rect 9291 23323 9333 23332
rect 9291 22448 9333 22457
rect 9291 22408 9292 22448
rect 9332 22408 9333 22448
rect 9291 22399 9333 22408
rect 9292 22280 9332 22399
rect 9195 21944 9237 21953
rect 9195 21904 9196 21944
rect 9236 21904 9237 21944
rect 9195 21895 9237 21904
rect 8907 21524 8949 21533
rect 8907 21484 8908 21524
rect 8948 21484 8949 21524
rect 8907 21475 8949 21484
rect 9099 20936 9141 20945
rect 9292 20936 9332 22240
rect 9388 21440 9428 23995
rect 9484 23633 9524 24340
rect 9676 23969 9716 24592
rect 9772 24473 9812 25600
rect 9868 25304 9908 25313
rect 9868 24893 9908 25264
rect 10059 25052 10101 25061
rect 10059 25012 10060 25052
rect 10100 25012 10101 25052
rect 10059 25003 10101 25012
rect 9867 24884 9909 24893
rect 9867 24844 9868 24884
rect 9908 24844 9909 24884
rect 9867 24835 9909 24844
rect 9867 24632 9909 24641
rect 9867 24592 9868 24632
rect 9908 24592 9909 24632
rect 9867 24583 9909 24592
rect 9964 24632 10004 24641
rect 9771 24464 9813 24473
rect 9771 24424 9772 24464
rect 9812 24424 9813 24464
rect 9771 24415 9813 24424
rect 9868 24137 9908 24583
rect 9867 24128 9909 24137
rect 9867 24088 9868 24128
rect 9908 24088 9909 24128
rect 9867 24079 9909 24088
rect 9964 23969 10004 24592
rect 9675 23960 9717 23969
rect 9675 23920 9676 23960
rect 9716 23920 9717 23960
rect 9675 23911 9717 23920
rect 9840 23960 9882 23969
rect 9963 23960 10005 23969
rect 9840 23920 9841 23960
rect 9881 23920 9908 23960
rect 9840 23911 9908 23920
rect 9963 23920 9964 23960
rect 10004 23920 10005 23960
rect 9963 23911 10005 23920
rect 9580 23792 9620 23801
rect 9483 23624 9525 23633
rect 9483 23584 9484 23624
rect 9524 23584 9525 23624
rect 9483 23575 9525 23584
rect 9580 22280 9620 23752
rect 9771 23792 9813 23801
rect 9771 23752 9772 23792
rect 9812 23752 9813 23792
rect 9771 23743 9813 23752
rect 9868 23792 9908 23911
rect 10060 23885 10100 25003
rect 10156 24380 10196 27616
rect 10539 26228 10581 26237
rect 10539 26188 10540 26228
rect 10580 26188 10581 26228
rect 10539 26179 10581 26188
rect 10348 24632 10388 24643
rect 10348 24557 10388 24592
rect 10443 24632 10485 24641
rect 10443 24592 10444 24632
rect 10484 24592 10485 24632
rect 10443 24583 10485 24592
rect 10347 24548 10389 24557
rect 10347 24508 10348 24548
rect 10388 24508 10389 24548
rect 10347 24499 10389 24508
rect 10444 24498 10484 24583
rect 10156 24340 10388 24380
rect 10059 23876 10101 23885
rect 10059 23836 10060 23876
rect 10100 23836 10101 23876
rect 10059 23827 10101 23836
rect 9868 23743 9908 23752
rect 9964 23792 10004 23801
rect 9675 22280 9717 22289
rect 9580 22240 9676 22280
rect 9716 22240 9717 22280
rect 9675 22231 9717 22240
rect 9579 21944 9621 21953
rect 9579 21904 9580 21944
rect 9620 21904 9621 21944
rect 9579 21895 9621 21904
rect 9484 21617 9524 21702
rect 9483 21608 9525 21617
rect 9483 21568 9484 21608
rect 9524 21568 9525 21608
rect 9580 21608 9620 21895
rect 9676 21776 9716 22231
rect 9772 22037 9812 23743
rect 9867 23624 9909 23633
rect 9867 23584 9868 23624
rect 9908 23584 9909 23624
rect 9867 23575 9909 23584
rect 9771 22028 9813 22037
rect 9771 21988 9772 22028
rect 9812 21988 9813 22028
rect 9771 21979 9813 21988
rect 9676 21727 9716 21736
rect 9580 21568 9812 21608
rect 9483 21559 9525 21568
rect 9388 21400 9524 21440
rect 9099 20896 9100 20936
rect 9140 20896 9332 20936
rect 9099 20887 9141 20896
rect 9387 20852 9429 20861
rect 9387 20812 9388 20852
rect 9428 20812 9429 20852
rect 9387 20803 9429 20812
rect 9003 20768 9045 20777
rect 9003 20728 9004 20768
rect 9044 20728 9045 20768
rect 9003 20719 9045 20728
rect 9388 20768 9428 20803
rect 9004 18584 9044 20719
rect 9388 20693 9428 20728
rect 9387 20684 9429 20693
rect 9387 20644 9388 20684
rect 9428 20644 9429 20684
rect 9387 20635 9429 20644
rect 9388 20604 9428 20635
rect 9292 20096 9332 20105
rect 9099 19256 9141 19265
rect 9099 19216 9100 19256
rect 9140 19216 9141 19256
rect 9099 19207 9141 19216
rect 9196 19256 9236 19267
rect 9100 19122 9140 19207
rect 9196 19181 9236 19216
rect 9195 19172 9237 19181
rect 9195 19132 9196 19172
rect 9236 19132 9237 19172
rect 9195 19123 9237 19132
rect 9099 19004 9141 19013
rect 9099 18964 9100 19004
rect 9140 18964 9141 19004
rect 9099 18955 9141 18964
rect 9100 18584 9140 18955
rect 9196 18752 9236 18761
rect 9292 18752 9332 20056
rect 9388 20096 9428 20105
rect 9388 19181 9428 20056
rect 9387 19172 9429 19181
rect 9387 19132 9388 19172
rect 9428 19132 9429 19172
rect 9387 19123 9429 19132
rect 9236 18712 9332 18752
rect 9387 18752 9429 18761
rect 9387 18712 9388 18752
rect 9428 18712 9429 18752
rect 9196 18703 9236 18712
rect 9387 18703 9429 18712
rect 9388 18584 9428 18703
rect 9100 18544 9236 18584
rect 8811 17912 8853 17921
rect 8811 17872 8812 17912
rect 8852 17872 8853 17912
rect 8811 17863 8853 17872
rect 8812 17744 8852 17753
rect 8812 17585 8852 17704
rect 8908 17744 8948 17755
rect 8908 17669 8948 17704
rect 8907 17660 8949 17669
rect 8907 17620 8908 17660
rect 8948 17620 8949 17660
rect 8907 17611 8949 17620
rect 8811 17576 8853 17585
rect 8811 17536 8812 17576
rect 8852 17536 8853 17576
rect 8811 17527 8853 17536
rect 8812 14561 8852 17527
rect 8907 16064 8949 16073
rect 8907 16024 8908 16064
rect 8948 16024 8949 16064
rect 8907 16015 8949 16024
rect 8908 15930 8948 16015
rect 9004 14888 9044 18544
rect 8908 14848 9044 14888
rect 9100 16316 9140 16325
rect 8811 14552 8853 14561
rect 8811 14512 8812 14552
rect 8852 14512 8853 14552
rect 8811 14503 8853 14512
rect 8715 12620 8757 12629
rect 8715 12580 8716 12620
rect 8756 12580 8757 12620
rect 8715 12571 8757 12580
rect 8620 11320 8756 11360
rect 8620 11024 8660 11033
rect 8620 10613 8660 10984
rect 8619 10604 8661 10613
rect 8619 10564 8620 10604
rect 8660 10564 8661 10604
rect 8619 10555 8661 10564
rect 8716 10445 8756 11320
rect 8812 10772 8852 10781
rect 8715 10436 8757 10445
rect 8524 10396 8660 10436
rect 8524 9512 8564 9521
rect 8524 9353 8564 9472
rect 8620 9512 8660 10396
rect 8715 10396 8716 10436
rect 8756 10396 8757 10436
rect 8715 10387 8757 10396
rect 8620 9463 8660 9472
rect 8523 9344 8565 9353
rect 8523 9304 8524 9344
rect 8564 9304 8565 9344
rect 8523 9295 8565 9304
rect 8716 9017 8756 10387
rect 8812 10109 8852 10732
rect 8811 10100 8853 10109
rect 8811 10060 8812 10100
rect 8852 10060 8853 10100
rect 8811 10051 8853 10060
rect 8908 9773 8948 14848
rect 9003 14720 9045 14729
rect 9003 14680 9004 14720
rect 9044 14680 9045 14720
rect 9003 14671 9045 14680
rect 9004 14586 9044 14671
rect 9004 14048 9044 14057
rect 9004 13973 9044 14008
rect 9003 13964 9045 13973
rect 9003 13924 9004 13964
rect 9044 13924 9045 13964
rect 9003 13915 9045 13924
rect 9004 12293 9044 13915
rect 9100 12788 9140 16276
rect 9196 15728 9236 18544
rect 9388 18425 9428 18544
rect 9387 18416 9429 18425
rect 9387 18376 9388 18416
rect 9428 18376 9429 18416
rect 9387 18367 9429 18376
rect 9291 17912 9333 17921
rect 9291 17872 9292 17912
rect 9332 17872 9333 17912
rect 9291 17863 9333 17872
rect 9292 16232 9332 17863
rect 9387 17744 9429 17753
rect 9387 17704 9388 17744
rect 9428 17704 9429 17744
rect 9387 17695 9429 17704
rect 9388 17610 9428 17695
rect 9484 17240 9524 21400
rect 9772 20180 9812 21568
rect 9868 21449 9908 23575
rect 9964 23381 10004 23752
rect 10156 23792 10196 23801
rect 10196 23752 10292 23792
rect 10156 23743 10196 23752
rect 10156 23624 10196 23633
rect 10060 23584 10156 23624
rect 9963 23372 10005 23381
rect 9963 23332 9964 23372
rect 10004 23332 10005 23372
rect 9963 23323 10005 23332
rect 10060 21692 10100 23584
rect 10156 23575 10196 23584
rect 10155 23456 10197 23465
rect 10155 23416 10156 23456
rect 10196 23416 10197 23456
rect 10155 23407 10197 23416
rect 10156 22877 10196 23407
rect 10155 22868 10197 22877
rect 10155 22828 10156 22868
rect 10196 22828 10197 22868
rect 10155 22819 10197 22828
rect 10155 22364 10197 22373
rect 10155 22324 10156 22364
rect 10196 22324 10197 22364
rect 10155 22315 10197 22324
rect 10156 22205 10196 22315
rect 10252 22289 10292 23752
rect 10348 23624 10388 24340
rect 10443 24128 10485 24137
rect 10443 24088 10444 24128
rect 10484 24088 10485 24128
rect 10443 24079 10485 24088
rect 10444 23792 10484 24079
rect 10540 23969 10580 26179
rect 10732 24305 10772 28120
rect 11020 27665 11060 28120
rect 11116 27833 11156 28288
rect 11115 27824 11157 27833
rect 11115 27784 11116 27824
rect 11156 27784 11157 27824
rect 11115 27775 11157 27784
rect 11019 27656 11061 27665
rect 11019 27616 11020 27656
rect 11060 27616 11061 27656
rect 11019 27607 11061 27616
rect 11019 26816 11061 26825
rect 11019 26776 11020 26816
rect 11060 26776 11061 26816
rect 11019 26767 11061 26776
rect 11211 26816 11253 26825
rect 11308 26816 11348 29203
rect 11403 29000 11445 29009
rect 11403 28960 11404 29000
rect 11444 28960 11445 29000
rect 11403 28951 11445 28960
rect 11404 28328 11444 28951
rect 11404 28253 11444 28288
rect 11403 28244 11445 28253
rect 11403 28204 11404 28244
rect 11444 28204 11445 28244
rect 11403 28195 11445 28204
rect 11403 27740 11445 27749
rect 11403 27700 11404 27740
rect 11444 27700 11445 27740
rect 11403 27691 11445 27700
rect 11404 27656 11444 27691
rect 11404 27605 11444 27616
rect 11403 26984 11445 26993
rect 11403 26944 11404 26984
rect 11444 26944 11445 26984
rect 11403 26935 11445 26944
rect 11404 26850 11444 26935
rect 11211 26776 11212 26816
rect 11252 26776 11348 26816
rect 11211 26767 11253 26776
rect 10923 24632 10965 24641
rect 10923 24592 10924 24632
rect 10964 24592 10965 24632
rect 10923 24583 10965 24592
rect 10828 24548 10868 24557
rect 10731 24296 10773 24305
rect 10731 24256 10732 24296
rect 10772 24256 10773 24296
rect 10731 24247 10773 24256
rect 10828 24044 10868 24508
rect 10924 24498 10964 24583
rect 11020 24221 11060 26767
rect 11212 26682 11252 26767
rect 11500 26564 11540 29716
rect 11596 27404 11636 27413
rect 11596 26900 11636 27364
rect 11692 26984 11732 29800
rect 11788 27068 11828 34495
rect 11884 32873 11924 32958
rect 11883 32864 11925 32873
rect 11883 32824 11884 32864
rect 11924 32824 11925 32864
rect 11883 32815 11925 32824
rect 11883 32696 11925 32705
rect 11883 32656 11884 32696
rect 11924 32656 11925 32696
rect 11883 32647 11925 32656
rect 11884 31100 11924 32647
rect 11980 31184 12020 35092
rect 12076 37400 12116 37519
rect 12076 35132 12116 37360
rect 12460 37325 12500 38872
rect 12556 38744 12596 38755
rect 12556 38669 12596 38704
rect 12555 38660 12597 38669
rect 12555 38620 12556 38660
rect 12596 38620 12597 38660
rect 12555 38611 12597 38620
rect 12555 38492 12597 38501
rect 12555 38452 12556 38492
rect 12596 38452 12597 38492
rect 12555 38443 12597 38452
rect 12556 37400 12596 38443
rect 12652 38235 12692 39460
rect 12748 39451 12788 39460
rect 12844 39257 12884 40384
rect 12939 39752 12981 39761
rect 12939 39712 12940 39752
rect 12980 39712 12981 39752
rect 12939 39703 12981 39712
rect 12940 39618 12980 39703
rect 12939 39500 12981 39509
rect 12939 39460 12940 39500
rect 12980 39460 12981 39500
rect 12939 39451 12981 39460
rect 12843 39248 12885 39257
rect 12843 39208 12844 39248
rect 12884 39208 12885 39248
rect 12843 39199 12885 39208
rect 12940 38912 12980 39451
rect 13036 39341 13076 40627
rect 13035 39332 13077 39341
rect 13035 39292 13036 39332
rect 13076 39292 13077 39332
rect 13035 39283 13077 39292
rect 13035 38996 13077 39005
rect 13035 38956 13036 38996
rect 13076 38956 13077 38996
rect 13035 38947 13077 38956
rect 12940 38837 12980 38872
rect 12939 38828 12981 38837
rect 12939 38788 12940 38828
rect 12980 38788 12981 38828
rect 12939 38779 12981 38788
rect 12747 38744 12789 38753
rect 12747 38704 12748 38744
rect 12788 38704 12789 38744
rect 12747 38695 12789 38704
rect 12748 38610 12788 38695
rect 12844 38324 12884 38333
rect 12652 38186 12692 38195
rect 12748 38284 12844 38324
rect 12748 37577 12788 38284
rect 12844 38275 12884 38284
rect 12940 38156 12980 38779
rect 13036 38744 13076 38947
rect 13132 38921 13172 40804
rect 14283 40676 14325 40685
rect 14283 40636 14284 40676
rect 14324 40636 14325 40676
rect 14283 40627 14325 40636
rect 14284 40542 14324 40627
rect 13324 40445 13364 40454
rect 13324 39836 13364 40405
rect 13611 40424 13653 40433
rect 13742 40431 13782 40440
rect 13611 40384 13612 40424
rect 13652 40384 13653 40424
rect 13611 40375 13653 40384
rect 13708 40391 13742 40424
rect 13708 40382 13782 40391
rect 13899 40424 13941 40433
rect 13899 40384 13900 40424
rect 13940 40384 13941 40424
rect 13515 40340 13557 40349
rect 13515 40300 13516 40340
rect 13556 40300 13557 40340
rect 13515 40291 13557 40300
rect 13516 40206 13556 40291
rect 13324 39796 13460 39836
rect 13323 39668 13365 39677
rect 13323 39628 13324 39668
rect 13364 39628 13365 39668
rect 13323 39619 13365 39628
rect 13131 38912 13173 38921
rect 13131 38872 13132 38912
rect 13172 38872 13173 38912
rect 13131 38863 13173 38872
rect 13036 38704 13172 38744
rect 12844 38116 12980 38156
rect 13036 38145 13076 38154
rect 12747 37568 12789 37577
rect 12747 37528 12748 37568
rect 12788 37528 12789 37568
rect 12747 37519 12789 37528
rect 12459 37316 12501 37325
rect 12459 37276 12460 37316
rect 12500 37276 12501 37316
rect 12459 37267 12501 37276
rect 12171 36308 12213 36317
rect 12171 36268 12172 36308
rect 12212 36268 12213 36308
rect 12171 36259 12213 36268
rect 12076 34553 12116 35092
rect 12075 34544 12117 34553
rect 12075 34504 12076 34544
rect 12116 34504 12117 34544
rect 12075 34495 12117 34504
rect 12076 34376 12116 34385
rect 12076 34301 12116 34336
rect 12075 34292 12117 34301
rect 12075 34252 12076 34292
rect 12116 34252 12117 34292
rect 12075 34243 12117 34252
rect 12076 34133 12116 34243
rect 12075 34124 12117 34133
rect 12075 34084 12076 34124
rect 12116 34084 12117 34124
rect 12075 34075 12117 34084
rect 12172 33788 12212 36259
rect 12363 35300 12405 35309
rect 12363 35260 12364 35300
rect 12404 35260 12405 35300
rect 12363 35251 12405 35260
rect 12076 33748 12212 33788
rect 12268 34208 12308 34217
rect 12076 33536 12116 33748
rect 12268 33704 12308 34168
rect 12364 33872 12404 35251
rect 12556 35216 12596 37360
rect 12651 37400 12693 37409
rect 12651 37360 12652 37400
rect 12692 37360 12693 37400
rect 12651 37351 12693 37360
rect 12460 34460 12500 34471
rect 12460 34385 12500 34420
rect 12459 34376 12501 34385
rect 12459 34336 12460 34376
rect 12500 34336 12501 34376
rect 12459 34327 12501 34336
rect 12364 33823 12404 33832
rect 12556 33788 12596 35176
rect 12652 34376 12692 37351
rect 12747 37316 12789 37325
rect 12747 37276 12748 37316
rect 12788 37276 12789 37316
rect 12747 37267 12789 37276
rect 12748 34460 12788 37267
rect 12844 35981 12884 38116
rect 12939 37904 12981 37913
rect 12939 37864 12940 37904
rect 12980 37864 12981 37904
rect 12939 37855 12981 37864
rect 12843 35972 12885 35981
rect 12843 35932 12844 35972
rect 12884 35932 12885 35972
rect 12843 35923 12885 35932
rect 12844 35888 12884 35923
rect 12844 35838 12884 35848
rect 12844 34460 12884 34469
rect 12748 34420 12844 34460
rect 12652 34336 12788 34376
rect 12652 34208 12692 34219
rect 12652 34133 12692 34168
rect 12651 34124 12693 34133
rect 12651 34084 12652 34124
rect 12692 34084 12693 34124
rect 12651 34075 12693 34084
rect 12556 33748 12692 33788
rect 12220 33694 12308 33704
rect 12260 33664 12308 33694
rect 12220 33645 12260 33654
rect 12556 33662 12596 33671
rect 12556 33620 12596 33622
rect 12364 33580 12596 33620
rect 12364 33536 12404 33580
rect 12076 33496 12404 33536
rect 12076 32696 12116 32705
rect 12076 32187 12116 32656
rect 12076 32138 12116 32147
rect 12172 31361 12212 33496
rect 12652 33368 12692 33748
rect 12556 33328 12692 33368
rect 12459 32780 12501 32789
rect 12459 32740 12460 32780
rect 12500 32740 12501 32780
rect 12459 32731 12501 32740
rect 12460 32646 12500 32731
rect 12459 32360 12501 32369
rect 12459 32320 12460 32360
rect 12500 32320 12501 32360
rect 12459 32311 12501 32320
rect 12267 32276 12309 32285
rect 12267 32236 12268 32276
rect 12308 32236 12309 32276
rect 12267 32227 12309 32236
rect 12268 32142 12308 32227
rect 12460 32226 12500 32311
rect 12363 32192 12405 32201
rect 12363 32152 12364 32192
rect 12404 32152 12405 32192
rect 12363 32143 12405 32152
rect 12364 31613 12404 32143
rect 12459 31688 12501 31697
rect 12459 31648 12460 31688
rect 12500 31648 12501 31688
rect 12459 31639 12501 31648
rect 12363 31604 12405 31613
rect 12363 31564 12364 31604
rect 12404 31564 12405 31604
rect 12363 31555 12405 31564
rect 12171 31352 12213 31361
rect 12171 31312 12172 31352
rect 12212 31312 12213 31352
rect 12171 31303 12213 31312
rect 12363 31184 12405 31193
rect 11980 31144 12308 31184
rect 11884 31060 12020 31100
rect 11980 30857 12020 31060
rect 11979 30848 12021 30857
rect 11979 30808 11980 30848
rect 12020 30808 12021 30848
rect 11979 30799 12021 30808
rect 11883 30764 11925 30773
rect 11883 30724 11884 30764
rect 11924 30724 11925 30764
rect 11883 30715 11925 30724
rect 11884 30630 11924 30715
rect 11883 27656 11925 27665
rect 11883 27616 11884 27656
rect 11924 27616 11925 27656
rect 11883 27607 11925 27616
rect 11884 27522 11924 27607
rect 11788 27028 11924 27068
rect 11692 26944 11828 26984
rect 11596 26860 11732 26900
rect 11692 26835 11732 26860
rect 11692 26786 11732 26795
rect 11788 26796 11828 26944
rect 11691 26732 11733 26741
rect 11788 26732 11828 26756
rect 11691 26692 11692 26732
rect 11732 26692 11828 26732
rect 11691 26683 11733 26692
rect 11884 26648 11924 27028
rect 11788 26608 11924 26648
rect 11500 26524 11732 26564
rect 11115 26312 11157 26321
rect 11115 26272 11116 26312
rect 11156 26272 11157 26312
rect 11115 26263 11157 26272
rect 11499 26312 11541 26321
rect 11499 26272 11500 26312
rect 11540 26272 11541 26312
rect 11499 26263 11541 26272
rect 11116 26144 11156 26263
rect 11500 26178 11540 26263
rect 11116 25304 11156 26104
rect 11308 25892 11348 25901
rect 11019 24212 11061 24221
rect 11019 24172 11020 24212
rect 11060 24172 11061 24212
rect 11019 24163 11061 24172
rect 10732 24004 10868 24044
rect 10539 23960 10581 23969
rect 10539 23920 10540 23960
rect 10580 23920 10581 23960
rect 10539 23911 10581 23920
rect 10444 23743 10484 23752
rect 10540 23792 10580 23803
rect 10540 23717 10580 23752
rect 10539 23708 10581 23717
rect 10539 23668 10540 23708
rect 10580 23668 10581 23708
rect 10539 23659 10581 23668
rect 10348 23584 10484 23624
rect 10348 23213 10388 23244
rect 10347 23204 10389 23213
rect 10347 23164 10348 23204
rect 10388 23164 10389 23204
rect 10347 23155 10389 23164
rect 10348 23120 10388 23155
rect 10348 22373 10388 23080
rect 10347 22364 10389 22373
rect 10347 22324 10348 22364
rect 10388 22324 10389 22364
rect 10347 22315 10389 22324
rect 10251 22280 10293 22289
rect 10251 22240 10252 22280
rect 10292 22240 10293 22280
rect 10251 22231 10293 22240
rect 10155 22196 10197 22205
rect 10155 22156 10156 22196
rect 10196 22156 10197 22196
rect 10155 22147 10197 22156
rect 10251 22028 10293 22037
rect 10251 21988 10252 22028
rect 10292 21988 10293 22028
rect 10444 22028 10484 23584
rect 10732 23465 10772 24004
rect 10923 23960 10965 23969
rect 10923 23920 10924 23960
rect 10964 23920 10965 23960
rect 10923 23911 10965 23920
rect 10924 23876 10964 23911
rect 10924 23825 10964 23836
rect 11020 23801 11060 23886
rect 11116 23885 11156 25264
rect 11212 25852 11308 25892
rect 11212 24137 11252 25852
rect 11308 25843 11348 25852
rect 11596 25397 11636 25482
rect 11595 25388 11637 25397
rect 11595 25348 11596 25388
rect 11636 25348 11637 25388
rect 11595 25339 11637 25348
rect 11308 25136 11348 25145
rect 11308 24557 11348 25096
rect 11404 24632 11444 24641
rect 11307 24548 11349 24557
rect 11307 24508 11308 24548
rect 11348 24508 11349 24548
rect 11307 24499 11349 24508
rect 11211 24128 11253 24137
rect 11211 24088 11212 24128
rect 11252 24088 11253 24128
rect 11211 24079 11253 24088
rect 11404 24053 11444 24592
rect 11403 24044 11445 24053
rect 11403 24004 11404 24044
rect 11444 24004 11445 24044
rect 11403 23995 11445 24004
rect 11115 23876 11157 23885
rect 11115 23836 11116 23876
rect 11156 23836 11157 23876
rect 11115 23827 11157 23836
rect 11019 23792 11061 23801
rect 11500 23792 11540 23801
rect 11019 23752 11020 23792
rect 11060 23752 11061 23792
rect 11019 23743 11061 23752
rect 11404 23752 11500 23792
rect 10731 23456 10773 23465
rect 10731 23416 10732 23456
rect 10772 23416 10773 23456
rect 10731 23407 10773 23416
rect 10539 23372 10581 23381
rect 10539 23332 10540 23372
rect 10580 23332 10581 23372
rect 10539 23323 10581 23332
rect 10828 23332 10964 23372
rect 10540 23288 10580 23323
rect 10828 23288 10868 23332
rect 10540 23237 10580 23248
rect 10636 23248 10868 23288
rect 10924 23288 10964 23332
rect 10539 22364 10581 22373
rect 10539 22324 10540 22364
rect 10580 22324 10581 22364
rect 10539 22315 10581 22324
rect 10540 22280 10580 22315
rect 10540 22229 10580 22240
rect 10444 21988 10580 22028
rect 10251 21979 10293 21988
rect 9964 21652 10100 21692
rect 9964 21608 10004 21652
rect 9964 21559 10004 21568
rect 10059 21524 10101 21533
rect 10059 21484 10060 21524
rect 10100 21484 10101 21524
rect 10059 21475 10101 21484
rect 10252 21524 10292 21979
rect 10347 21944 10389 21953
rect 10347 21904 10348 21944
rect 10388 21904 10389 21944
rect 10347 21895 10389 21904
rect 10348 21608 10388 21895
rect 10540 21617 10580 21988
rect 10636 21953 10676 23248
rect 10924 23239 10964 23248
rect 11116 23213 11156 23244
rect 11115 23204 11157 23213
rect 11115 23164 11116 23204
rect 11156 23164 11157 23204
rect 11115 23155 11157 23164
rect 10732 23120 10772 23129
rect 11020 23120 11060 23129
rect 10876 23110 10916 23119
rect 10732 22532 10772 23080
rect 10855 23070 10876 23110
rect 10855 23061 10916 23070
rect 10855 23045 10895 23061
rect 10827 23036 10895 23045
rect 10827 22996 10828 23036
rect 10868 22996 10895 23036
rect 10827 22987 10869 22996
rect 11020 22625 11060 23080
rect 11116 23120 11156 23155
rect 11116 22709 11156 23080
rect 11273 23105 11313 23114
rect 11273 23045 11313 23065
rect 11273 23036 11349 23045
rect 11273 22996 11308 23036
rect 11348 22996 11349 23036
rect 11307 22987 11349 22996
rect 11307 22868 11349 22877
rect 11307 22828 11308 22868
rect 11348 22828 11349 22868
rect 11307 22819 11349 22828
rect 11115 22700 11157 22709
rect 11115 22660 11116 22700
rect 11156 22660 11157 22700
rect 11115 22651 11157 22660
rect 11019 22616 11061 22625
rect 11019 22576 11020 22616
rect 11060 22576 11061 22616
rect 11019 22567 11061 22576
rect 10732 22483 10772 22492
rect 11019 22280 11061 22289
rect 11019 22240 11020 22280
rect 11060 22240 11061 22280
rect 11019 22231 11061 22240
rect 11308 22280 11348 22819
rect 11404 22364 11444 23752
rect 11500 23743 11540 23752
rect 11499 23372 11541 23381
rect 11499 23332 11500 23372
rect 11540 23332 11541 23372
rect 11499 23323 11541 23332
rect 11500 23120 11540 23323
rect 11692 23297 11732 26524
rect 11788 26144 11828 26608
rect 11883 26312 11925 26321
rect 11883 26272 11884 26312
rect 11924 26272 11925 26312
rect 11883 26263 11925 26272
rect 11884 26178 11924 26263
rect 11788 24893 11828 26104
rect 11787 24884 11829 24893
rect 11787 24844 11788 24884
rect 11828 24844 11829 24884
rect 11787 24835 11829 24844
rect 11980 24716 12020 30799
rect 12171 30764 12213 30773
rect 12171 30724 12172 30764
rect 12212 30724 12213 30764
rect 12171 30715 12213 30724
rect 12172 30680 12212 30715
rect 12172 30629 12212 30640
rect 12268 30680 12308 31144
rect 12363 31144 12364 31184
rect 12404 31144 12405 31184
rect 12363 31135 12405 31144
rect 12268 30605 12308 30640
rect 12267 30596 12309 30605
rect 12267 30556 12268 30596
rect 12308 30556 12309 30596
rect 12267 30547 12309 30556
rect 12075 30092 12117 30101
rect 12075 30052 12076 30092
rect 12116 30052 12117 30092
rect 12075 30043 12117 30052
rect 12076 29840 12116 30043
rect 12171 29924 12213 29933
rect 12171 29884 12172 29924
rect 12212 29884 12213 29924
rect 12171 29875 12213 29884
rect 12076 29681 12116 29800
rect 12172 29790 12212 29875
rect 12075 29672 12117 29681
rect 12364 29672 12404 31135
rect 12460 30092 12500 31639
rect 12556 30691 12596 33328
rect 12651 33200 12693 33209
rect 12651 33160 12652 33200
rect 12692 33160 12693 33200
rect 12651 33151 12693 33160
rect 12652 33116 12692 33151
rect 12652 33065 12692 33076
rect 12748 32696 12788 34336
rect 12844 33965 12884 34420
rect 12843 33956 12885 33965
rect 12843 33916 12844 33956
rect 12884 33916 12885 33956
rect 12843 33907 12885 33916
rect 12844 33797 12884 33907
rect 12843 33788 12885 33797
rect 12843 33748 12844 33788
rect 12884 33748 12885 33788
rect 12843 33739 12885 33748
rect 12843 33452 12885 33461
rect 12843 33412 12844 33452
rect 12884 33412 12885 33452
rect 12843 33403 12885 33412
rect 12844 32864 12884 33403
rect 12844 32815 12884 32824
rect 12748 32656 12884 32696
rect 12747 32444 12789 32453
rect 12747 32404 12748 32444
rect 12788 32404 12789 32444
rect 12747 32395 12789 32404
rect 12748 32192 12788 32395
rect 12748 30941 12788 32152
rect 12747 30932 12789 30941
rect 12747 30892 12748 30932
rect 12788 30892 12789 30932
rect 12747 30883 12789 30892
rect 12556 30680 12692 30691
rect 12556 30651 12652 30680
rect 12652 30631 12692 30640
rect 12747 30596 12789 30605
rect 12747 30556 12748 30596
rect 12788 30556 12789 30596
rect 12747 30547 12789 30556
rect 12748 30462 12788 30547
rect 12460 30052 12596 30092
rect 12459 29924 12501 29933
rect 12459 29884 12460 29924
rect 12500 29884 12501 29924
rect 12459 29875 12501 29884
rect 12075 29632 12076 29672
rect 12116 29632 12117 29672
rect 12075 29623 12117 29632
rect 12172 29632 12404 29672
rect 12172 27917 12212 29632
rect 12460 29588 12500 29875
rect 12268 29548 12500 29588
rect 12171 27908 12213 27917
rect 12171 27868 12172 27908
rect 12212 27868 12213 27908
rect 12171 27859 12213 27868
rect 12075 26984 12117 26993
rect 12075 26944 12076 26984
rect 12116 26944 12117 26984
rect 12075 26935 12117 26944
rect 12076 26396 12116 26935
rect 12172 26900 12212 27859
rect 12172 26851 12212 26860
rect 12268 26816 12308 29548
rect 12556 29504 12596 30052
rect 12076 26356 12212 26396
rect 12075 26228 12117 26237
rect 12075 26188 12076 26228
rect 12116 26188 12117 26228
rect 12075 26179 12117 26188
rect 12076 26094 12116 26179
rect 12172 25304 12212 26356
rect 12268 25649 12308 26776
rect 12364 29464 12596 29504
rect 12652 29840 12692 29849
rect 12364 26312 12404 29464
rect 12459 29252 12501 29261
rect 12459 29212 12460 29252
rect 12500 29212 12501 29252
rect 12459 29203 12501 29212
rect 12460 29168 12500 29203
rect 12460 28328 12500 29128
rect 12652 29084 12692 29800
rect 12844 29513 12884 32656
rect 12940 31697 12980 37855
rect 13036 37829 13076 38105
rect 13035 37820 13077 37829
rect 13035 37780 13036 37820
rect 13076 37780 13077 37820
rect 13035 37771 13077 37780
rect 13132 37568 13172 38704
rect 13227 38492 13269 38501
rect 13227 38452 13228 38492
rect 13268 38452 13269 38492
rect 13227 38443 13269 38452
rect 13228 38408 13268 38443
rect 13228 38357 13268 38368
rect 13324 37820 13364 39619
rect 13420 39593 13460 39796
rect 13419 39584 13461 39593
rect 13419 39544 13420 39584
rect 13460 39544 13461 39584
rect 13419 39535 13461 39544
rect 13612 39080 13652 40375
rect 13708 39761 13748 40382
rect 13899 40375 13941 40384
rect 13996 40424 14036 40433
rect 14188 40431 14228 40433
rect 13900 40290 13940 40375
rect 13803 40256 13845 40265
rect 13803 40216 13804 40256
rect 13844 40216 13845 40256
rect 13803 40207 13845 40216
rect 13707 39752 13749 39761
rect 13707 39712 13708 39752
rect 13748 39712 13749 39752
rect 13707 39703 13749 39712
rect 13516 39040 13652 39080
rect 13419 38156 13461 38165
rect 13419 38116 13420 38156
rect 13460 38116 13461 38156
rect 13419 38107 13461 38116
rect 13420 38022 13460 38107
rect 13324 37780 13460 37820
rect 13132 37528 13364 37568
rect 13084 37409 13124 37418
rect 13124 37369 13172 37400
rect 13084 37360 13172 37369
rect 13035 37064 13077 37073
rect 13035 37024 13036 37064
rect 13076 37024 13077 37064
rect 13035 37015 13077 37024
rect 13036 36728 13076 37015
rect 13132 36896 13172 37360
rect 13227 37316 13269 37325
rect 13227 37276 13228 37316
rect 13268 37276 13269 37316
rect 13227 37267 13269 37276
rect 13228 37182 13268 37267
rect 13324 37064 13364 37528
rect 13420 37409 13460 37780
rect 13419 37400 13461 37409
rect 13419 37360 13420 37400
rect 13460 37360 13461 37400
rect 13419 37351 13461 37360
rect 13420 37266 13460 37351
rect 13419 37064 13461 37073
rect 13324 37024 13420 37064
rect 13460 37024 13461 37064
rect 13419 37015 13461 37024
rect 13228 36896 13268 36905
rect 13132 36856 13228 36896
rect 13228 36847 13268 36856
rect 13323 36812 13365 36821
rect 13323 36772 13324 36812
rect 13364 36772 13365 36812
rect 13323 36763 13365 36772
rect 13036 36679 13076 36688
rect 13324 36056 13364 36763
rect 13420 36728 13460 37015
rect 13420 36679 13460 36688
rect 13516 36569 13556 39040
rect 13611 38744 13653 38753
rect 13611 38704 13612 38744
rect 13652 38704 13653 38744
rect 13611 38695 13653 38704
rect 13612 38408 13652 38695
rect 13707 38660 13749 38669
rect 13707 38620 13708 38660
rect 13748 38620 13749 38660
rect 13707 38611 13749 38620
rect 13612 38359 13652 38368
rect 13708 38165 13748 38611
rect 13804 38240 13844 40207
rect 13996 39929 14036 40384
rect 14092 40424 14228 40431
rect 14092 40391 14188 40424
rect 14092 40349 14132 40391
rect 14188 40375 14228 40384
rect 14284 40424 14324 40433
rect 14091 40340 14133 40349
rect 14091 40300 14092 40340
rect 14132 40300 14133 40340
rect 14091 40291 14133 40300
rect 14284 40265 14324 40384
rect 14283 40256 14325 40265
rect 14283 40216 14284 40256
rect 14324 40216 14325 40256
rect 14283 40207 14325 40216
rect 14380 40088 14420 42391
rect 14476 41693 14516 42928
rect 14571 42608 14613 42617
rect 14571 42568 14572 42608
rect 14612 42568 14613 42608
rect 14571 42559 14613 42568
rect 14475 41684 14517 41693
rect 14475 41644 14476 41684
rect 14516 41644 14517 41684
rect 14475 41635 14517 41644
rect 14572 40769 14612 42559
rect 14668 42029 14708 42928
rect 14667 42020 14709 42029
rect 14667 41980 14668 42020
rect 14708 41980 14709 42020
rect 14667 41971 14709 41980
rect 14763 41852 14805 41861
rect 14763 41812 14764 41852
rect 14804 41812 14805 41852
rect 14763 41803 14805 41812
rect 14571 40760 14613 40769
rect 14571 40720 14572 40760
rect 14612 40720 14613 40760
rect 14571 40711 14613 40720
rect 14571 40592 14613 40601
rect 14571 40552 14572 40592
rect 14612 40552 14613 40592
rect 14571 40543 14613 40552
rect 14572 40458 14612 40543
rect 14284 40048 14420 40088
rect 14476 40424 14516 40433
rect 13995 39920 14037 39929
rect 13995 39880 13996 39920
rect 14036 39880 14037 39920
rect 13995 39871 14037 39880
rect 14188 39752 14228 39761
rect 14188 39593 14228 39712
rect 14187 39584 14229 39593
rect 14187 39544 14188 39584
rect 14228 39544 14229 39584
rect 14187 39535 14229 39544
rect 14091 39500 14133 39509
rect 14091 39460 14092 39500
rect 14132 39460 14133 39500
rect 14091 39451 14133 39460
rect 13707 38156 13749 38165
rect 13707 38116 13708 38156
rect 13748 38116 13749 38156
rect 13707 38107 13749 38116
rect 13708 37820 13748 38107
rect 13612 37780 13748 37820
rect 13515 36560 13557 36569
rect 13515 36520 13516 36560
rect 13556 36520 13557 36560
rect 13515 36511 13557 36520
rect 13132 36016 13364 36056
rect 13036 35720 13076 35729
rect 13036 35211 13076 35680
rect 13036 35162 13076 35171
rect 13036 34628 13076 34637
rect 13132 34628 13172 36016
rect 13323 35888 13365 35897
rect 13323 35848 13324 35888
rect 13364 35848 13365 35888
rect 13323 35839 13365 35848
rect 13227 35804 13269 35813
rect 13227 35764 13228 35804
rect 13268 35764 13269 35804
rect 13227 35755 13269 35764
rect 13228 35426 13268 35755
rect 13324 35754 13364 35839
rect 13323 35636 13365 35645
rect 13323 35596 13324 35636
rect 13364 35596 13365 35636
rect 13323 35587 13365 35596
rect 13228 35377 13268 35386
rect 13324 35300 13364 35587
rect 13076 34588 13172 34628
rect 13228 35260 13364 35300
rect 13036 34579 13076 34588
rect 13131 34376 13173 34385
rect 13131 34336 13132 34376
rect 13172 34336 13173 34376
rect 13131 34327 13173 34336
rect 12939 31688 12981 31697
rect 12939 31648 12940 31688
rect 12980 31648 12981 31688
rect 12939 31639 12981 31648
rect 13132 31520 13172 34327
rect 13132 31480 13179 31520
rect 12940 31361 12980 31446
rect 13139 31361 13179 31480
rect 12939 31352 12981 31361
rect 12939 31312 12940 31352
rect 12980 31312 12981 31352
rect 12939 31303 12981 31312
rect 13131 31352 13179 31361
rect 13131 31312 13132 31352
rect 13172 31312 13179 31352
rect 13131 31303 13173 31312
rect 12939 31184 12981 31193
rect 12939 31144 12940 31184
rect 12980 31144 12981 31184
rect 12939 31135 12981 31144
rect 13132 31184 13172 31193
rect 12843 29504 12885 29513
rect 12843 29464 12844 29504
rect 12884 29464 12885 29504
rect 12843 29455 12885 29464
rect 12843 29168 12885 29177
rect 12843 29128 12844 29168
rect 12884 29128 12885 29168
rect 12843 29119 12885 29128
rect 12556 29044 12692 29084
rect 12556 28664 12596 29044
rect 12844 29034 12884 29119
rect 12651 28916 12693 28925
rect 12651 28876 12652 28916
rect 12692 28876 12693 28916
rect 12651 28867 12693 28876
rect 12652 28782 12692 28867
rect 12556 28624 12692 28664
rect 12652 28505 12692 28624
rect 12843 28580 12885 28589
rect 12843 28540 12844 28580
rect 12884 28540 12885 28580
rect 12843 28531 12885 28540
rect 12651 28496 12693 28505
rect 12651 28456 12652 28496
rect 12692 28456 12693 28496
rect 12651 28447 12693 28456
rect 12844 28446 12884 28531
rect 12652 28328 12692 28337
rect 12460 28288 12652 28328
rect 12652 27833 12692 28288
rect 12843 28328 12885 28337
rect 12843 28288 12844 28328
rect 12884 28288 12885 28328
rect 12843 28279 12885 28288
rect 12651 27824 12693 27833
rect 12651 27784 12652 27824
rect 12692 27784 12693 27824
rect 12651 27775 12693 27784
rect 12844 27413 12884 28279
rect 12843 27404 12885 27413
rect 12843 27364 12844 27404
rect 12884 27364 12885 27404
rect 12843 27355 12885 27364
rect 12843 27236 12885 27245
rect 12843 27196 12844 27236
rect 12884 27196 12885 27236
rect 12843 27187 12885 27196
rect 12747 26816 12789 26825
rect 12747 26776 12748 26816
rect 12788 26776 12789 26816
rect 12747 26767 12789 26776
rect 12748 26682 12788 26767
rect 12364 26272 12596 26312
rect 12364 26144 12404 26153
rect 12364 25817 12404 26104
rect 12363 25808 12405 25817
rect 12363 25768 12364 25808
rect 12404 25768 12405 25808
rect 12363 25759 12405 25768
rect 12267 25640 12309 25649
rect 12267 25600 12268 25640
rect 12308 25600 12309 25640
rect 12267 25591 12309 25600
rect 12364 25397 12404 25759
rect 12363 25388 12405 25397
rect 12363 25348 12364 25388
rect 12404 25348 12405 25388
rect 12363 25339 12405 25348
rect 12172 25255 12212 25264
rect 12267 25304 12309 25313
rect 12267 25264 12268 25304
rect 12308 25264 12309 25304
rect 12267 25255 12309 25264
rect 12268 25170 12308 25255
rect 11788 24676 12020 24716
rect 12076 24716 12116 24725
rect 12116 24676 12500 24716
rect 11691 23288 11733 23297
rect 11691 23248 11692 23288
rect 11732 23248 11733 23288
rect 11691 23239 11733 23248
rect 11595 23204 11637 23213
rect 11595 23164 11596 23204
rect 11636 23164 11637 23204
rect 11595 23155 11637 23164
rect 11500 23071 11540 23080
rect 11596 23070 11636 23155
rect 11691 23036 11733 23045
rect 11691 22996 11692 23036
rect 11732 22996 11733 23036
rect 11691 22987 11733 22996
rect 11692 22532 11732 22987
rect 11692 22483 11732 22492
rect 11788 22364 11828 24676
rect 12076 24667 12116 24676
rect 11884 24618 11924 24627
rect 11884 24137 11924 24578
rect 11979 24548 12021 24557
rect 11979 24508 11980 24548
rect 12020 24508 12021 24548
rect 11979 24499 12021 24508
rect 11883 24128 11925 24137
rect 11883 24088 11884 24128
rect 11924 24088 11925 24128
rect 11883 24079 11925 24088
rect 11980 23806 12020 24499
rect 12364 23960 12404 23969
rect 11980 23757 12020 23766
rect 12076 23920 12364 23960
rect 11980 23120 12020 23129
rect 12076 23120 12116 23920
rect 12364 23911 12404 23920
rect 12460 23792 12500 24676
rect 12556 23960 12596 26272
rect 12747 25388 12789 25397
rect 12747 25348 12748 25388
rect 12788 25348 12789 25388
rect 12747 25339 12789 25348
rect 12652 25304 12692 25313
rect 12652 24389 12692 25264
rect 12651 24380 12693 24389
rect 12651 24340 12652 24380
rect 12692 24340 12693 24380
rect 12651 24331 12693 24340
rect 12556 23920 12692 23960
rect 12268 23752 12500 23792
rect 12555 23792 12597 23801
rect 12555 23752 12556 23792
rect 12596 23752 12597 23792
rect 12020 23080 12116 23120
rect 12172 23624 12212 23633
rect 12172 23120 12212 23584
rect 12268 23288 12308 23752
rect 12555 23743 12597 23752
rect 12556 23658 12596 23743
rect 12652 23540 12692 23920
rect 12748 23801 12788 25339
rect 12844 24221 12884 27187
rect 12940 24464 12980 31135
rect 13035 31016 13077 31025
rect 13035 30976 13036 31016
rect 13076 30976 13077 31016
rect 13035 30967 13077 30976
rect 13036 29420 13076 30967
rect 13132 29854 13172 31144
rect 13228 31025 13268 35260
rect 13419 35216 13461 35225
rect 13419 35176 13420 35216
rect 13460 35176 13461 35216
rect 13419 35167 13461 35176
rect 13420 35145 13460 35167
rect 13323 35132 13365 35141
rect 13323 35092 13324 35132
rect 13364 35092 13365 35132
rect 13323 35083 13365 35092
rect 13612 35132 13652 37780
rect 13707 35468 13749 35477
rect 13707 35428 13708 35468
rect 13748 35428 13749 35468
rect 13707 35419 13749 35428
rect 13324 34460 13364 35083
rect 13420 35081 13460 35105
rect 13516 35092 13652 35132
rect 13420 34460 13460 34469
rect 13324 34420 13420 34460
rect 13227 31016 13269 31025
rect 13227 30976 13228 31016
rect 13268 30976 13269 31016
rect 13227 30967 13269 30976
rect 13227 30764 13269 30773
rect 13227 30724 13228 30764
rect 13268 30724 13269 30764
rect 13227 30715 13269 30724
rect 13228 30680 13268 30715
rect 13228 29933 13268 30640
rect 13324 30101 13364 34420
rect 13420 34411 13460 34420
rect 13516 34040 13556 35092
rect 13612 34964 13652 34973
rect 13708 34964 13748 35419
rect 13804 35309 13844 38200
rect 13995 37736 14037 37745
rect 13995 37696 13996 37736
rect 14036 37696 14037 37736
rect 13995 37687 14037 37696
rect 13899 35888 13941 35897
rect 13899 35848 13900 35888
rect 13940 35848 13941 35888
rect 13899 35839 13941 35848
rect 13900 35561 13940 35839
rect 13899 35552 13941 35561
rect 13899 35512 13900 35552
rect 13940 35512 13941 35552
rect 13899 35503 13941 35512
rect 13803 35300 13845 35309
rect 13803 35260 13804 35300
rect 13844 35260 13845 35300
rect 13803 35251 13845 35260
rect 13652 34924 13748 34964
rect 13804 35132 13844 35141
rect 13612 34915 13652 34924
rect 13707 34544 13749 34553
rect 13707 34504 13708 34544
rect 13748 34504 13749 34544
rect 13707 34495 13749 34504
rect 13804 34544 13844 35092
rect 13804 34495 13844 34504
rect 13611 34208 13653 34217
rect 13611 34168 13612 34208
rect 13652 34168 13653 34208
rect 13611 34159 13653 34168
rect 13612 34074 13652 34159
rect 13708 34133 13748 34495
rect 13900 34376 13940 35503
rect 13996 35225 14036 37687
rect 13995 35216 14037 35225
rect 13995 35176 13996 35216
rect 14036 35176 14037 35216
rect 13995 35167 14037 35176
rect 13996 35048 14036 35057
rect 14092 35048 14132 39451
rect 14188 38912 14228 38921
rect 14188 37829 14228 38872
rect 14187 37820 14229 37829
rect 14187 37780 14188 37820
rect 14228 37780 14229 37820
rect 14284 37820 14324 40048
rect 14380 39836 14420 39847
rect 14380 39761 14420 39796
rect 14379 39752 14421 39761
rect 14379 39712 14380 39752
rect 14420 39712 14421 39752
rect 14379 39703 14421 39712
rect 14379 39332 14421 39341
rect 14379 39292 14380 39332
rect 14420 39292 14421 39332
rect 14379 39283 14421 39292
rect 14380 38912 14420 39283
rect 14380 38863 14420 38872
rect 14476 38417 14516 40384
rect 14764 40424 14804 41803
rect 14860 41189 14900 42928
rect 14955 42860 14997 42869
rect 14955 42820 14956 42860
rect 14996 42820 14997 42860
rect 14955 42811 14997 42820
rect 14859 41180 14901 41189
rect 14859 41140 14860 41180
rect 14900 41140 14901 41180
rect 14859 41131 14901 41140
rect 14956 41105 14996 42811
rect 15052 42113 15092 42928
rect 15244 42533 15284 42928
rect 15243 42524 15285 42533
rect 15243 42484 15244 42524
rect 15284 42484 15285 42524
rect 15243 42475 15285 42484
rect 15051 42104 15093 42113
rect 15051 42064 15052 42104
rect 15092 42064 15093 42104
rect 15051 42055 15093 42064
rect 15436 41432 15476 42928
rect 15244 41392 15476 41432
rect 14955 41096 14997 41105
rect 14955 41056 14956 41096
rect 14996 41056 14997 41096
rect 14955 41047 14997 41056
rect 14764 40375 14804 40384
rect 14955 40424 14997 40433
rect 14955 40384 14956 40424
rect 14996 40384 14997 40424
rect 14955 40375 14997 40384
rect 14571 40256 14613 40265
rect 14571 40216 14572 40256
rect 14612 40216 14613 40256
rect 14571 40207 14613 40216
rect 14763 40256 14805 40265
rect 14763 40216 14764 40256
rect 14804 40216 14805 40256
rect 14763 40207 14805 40216
rect 14572 39920 14612 40207
rect 14668 39920 14708 39929
rect 14572 39880 14668 39920
rect 14668 39871 14708 39880
rect 14572 39752 14612 39761
rect 14572 39089 14612 39712
rect 14764 39752 14804 40207
rect 14764 39703 14804 39712
rect 14859 39752 14901 39761
rect 14859 39712 14860 39752
rect 14900 39712 14901 39752
rect 14859 39703 14901 39712
rect 14860 39618 14900 39703
rect 14763 39500 14805 39509
rect 14763 39460 14764 39500
rect 14804 39460 14805 39500
rect 14763 39451 14805 39460
rect 14571 39080 14613 39089
rect 14571 39040 14572 39080
rect 14612 39040 14613 39080
rect 14571 39031 14613 39040
rect 14475 38408 14517 38417
rect 14475 38368 14476 38408
rect 14516 38368 14517 38408
rect 14475 38359 14517 38368
rect 14667 38240 14709 38249
rect 14667 38200 14668 38240
rect 14708 38200 14709 38240
rect 14667 38191 14709 38200
rect 14284 37780 14420 37820
rect 14187 37771 14229 37780
rect 14283 35636 14325 35645
rect 14283 35596 14284 35636
rect 14324 35596 14325 35636
rect 14283 35587 14325 35596
rect 14036 35008 14132 35048
rect 14188 35132 14228 35141
rect 13996 34999 14036 35008
rect 13900 34336 14036 34376
rect 13900 34208 13940 34217
rect 13707 34124 13749 34133
rect 13707 34084 13708 34124
rect 13748 34084 13749 34124
rect 13707 34075 13749 34084
rect 13900 34049 13940 34168
rect 13420 34000 13556 34040
rect 13899 34040 13941 34049
rect 13899 34000 13900 34040
rect 13940 34000 13941 34040
rect 13420 31361 13460 34000
rect 13899 33991 13941 34000
rect 13803 33956 13845 33965
rect 13803 33916 13804 33956
rect 13844 33916 13845 33956
rect 13803 33907 13845 33916
rect 13804 33704 13844 33907
rect 13804 33461 13844 33664
rect 13996 33620 14036 34336
rect 14188 34208 14228 35092
rect 14188 34133 14228 34168
rect 14187 34124 14229 34133
rect 14187 34084 14188 34124
rect 14228 34084 14229 34124
rect 14187 34075 14229 34084
rect 14284 33956 14324 35587
rect 14380 35048 14420 37780
rect 14668 37493 14708 38191
rect 14667 37484 14709 37493
rect 14667 37444 14668 37484
rect 14708 37444 14709 37484
rect 14667 37435 14709 37444
rect 14668 37400 14708 37435
rect 14668 37349 14708 37360
rect 14668 36728 14708 36737
rect 14572 36688 14668 36728
rect 14572 35981 14612 36688
rect 14668 36679 14708 36688
rect 14764 36560 14804 39451
rect 14859 38072 14901 38081
rect 14859 38032 14860 38072
rect 14900 38032 14901 38072
rect 14859 38023 14901 38032
rect 14860 37652 14900 38023
rect 14860 37409 14900 37612
rect 14859 37400 14901 37409
rect 14859 37360 14860 37400
rect 14900 37360 14901 37400
rect 14859 37351 14901 37360
rect 14859 36980 14901 36989
rect 14859 36940 14860 36980
rect 14900 36940 14901 36980
rect 14859 36931 14901 36940
rect 14860 36896 14900 36931
rect 14860 36569 14900 36856
rect 14668 36520 14804 36560
rect 14859 36560 14901 36569
rect 14859 36520 14860 36560
rect 14900 36520 14901 36560
rect 14571 35972 14613 35981
rect 14571 35932 14572 35972
rect 14612 35932 14613 35972
rect 14571 35923 14613 35932
rect 14572 35888 14612 35923
rect 14572 35837 14612 35848
rect 14668 35309 14708 36520
rect 14859 36511 14901 36520
rect 14763 36392 14805 36401
rect 14763 36352 14764 36392
rect 14804 36352 14805 36392
rect 14763 36343 14805 36352
rect 14764 36140 14804 36343
rect 14764 36091 14804 36100
rect 14956 36056 14996 40375
rect 15244 40265 15284 41392
rect 15339 41264 15381 41273
rect 15339 41224 15340 41264
rect 15380 41224 15381 41264
rect 15339 41215 15381 41224
rect 15340 41130 15380 41215
rect 15532 41012 15572 41021
rect 15436 40972 15532 41012
rect 15243 40256 15285 40265
rect 15243 40216 15244 40256
rect 15284 40216 15285 40256
rect 15243 40207 15285 40216
rect 15147 40088 15189 40097
rect 15147 40048 15148 40088
rect 15188 40048 15189 40088
rect 15147 40039 15189 40048
rect 15051 39752 15093 39761
rect 15051 39712 15052 39752
rect 15092 39712 15093 39752
rect 15051 39703 15093 39712
rect 15148 39752 15188 40039
rect 15339 39920 15381 39929
rect 15339 39880 15340 39920
rect 15380 39880 15381 39920
rect 15339 39871 15381 39880
rect 15340 39786 15380 39871
rect 15148 39703 15188 39712
rect 15052 39618 15092 39703
rect 15051 38912 15093 38921
rect 15051 38872 15052 38912
rect 15092 38872 15093 38912
rect 15051 38863 15093 38872
rect 15052 38249 15092 38863
rect 15051 38240 15093 38249
rect 15051 38200 15052 38240
rect 15092 38200 15093 38240
rect 15051 38191 15093 38200
rect 15052 38106 15092 38191
rect 15244 37988 15284 37997
rect 15244 37829 15284 37948
rect 15243 37820 15285 37829
rect 15243 37780 15244 37820
rect 15284 37780 15285 37820
rect 15243 37771 15285 37780
rect 15436 37661 15476 40972
rect 15532 40963 15572 40972
rect 15628 40433 15668 42928
rect 15724 41264 15764 41273
rect 15627 40424 15669 40433
rect 15627 40384 15628 40424
rect 15668 40384 15669 40424
rect 15627 40375 15669 40384
rect 15724 39836 15764 41224
rect 15820 40685 15860 42928
rect 16012 42197 16052 42928
rect 16011 42188 16053 42197
rect 16011 42148 16012 42188
rect 16052 42148 16053 42188
rect 16011 42139 16053 42148
rect 15819 40676 15861 40685
rect 15819 40636 15820 40676
rect 15860 40636 15861 40676
rect 15819 40627 15861 40636
rect 15628 39796 15764 39836
rect 16012 40424 16052 40433
rect 16204 40424 16244 42928
rect 16396 41180 16436 42928
rect 16588 41768 16628 42928
rect 16588 41728 16724 41768
rect 16587 41600 16629 41609
rect 16587 41560 16588 41600
rect 16628 41560 16629 41600
rect 16587 41551 16629 41560
rect 16300 41140 16436 41180
rect 16300 40928 16340 41140
rect 16300 40888 16532 40928
rect 16204 40384 16340 40424
rect 15531 39500 15573 39509
rect 15531 39460 15532 39500
rect 15572 39460 15573 39500
rect 15531 39451 15573 39460
rect 15532 39366 15572 39451
rect 15628 38921 15668 39796
rect 15723 39668 15765 39677
rect 15723 39628 15724 39668
rect 15764 39628 15765 39668
rect 15723 39619 15765 39628
rect 15724 39534 15764 39619
rect 16012 39089 16052 40384
rect 16204 40256 16244 40265
rect 16108 40216 16204 40256
rect 16108 39752 16148 40216
rect 16204 40207 16244 40216
rect 16300 40013 16340 40384
rect 16396 40256 16436 40265
rect 16396 40097 16436 40216
rect 16395 40088 16437 40097
rect 16395 40048 16396 40088
rect 16436 40048 16437 40088
rect 16395 40039 16437 40048
rect 16299 40004 16341 40013
rect 16299 39964 16300 40004
rect 16340 39964 16341 40004
rect 16299 39955 16341 39964
rect 16108 39703 16148 39712
rect 16203 39752 16245 39761
rect 16203 39712 16204 39752
rect 16244 39712 16245 39752
rect 16203 39703 16245 39712
rect 16204 39618 16244 39703
rect 16299 39332 16341 39341
rect 16299 39292 16300 39332
rect 16340 39292 16341 39332
rect 16299 39283 16341 39292
rect 16011 39080 16053 39089
rect 16011 39040 16012 39080
rect 16052 39040 16053 39080
rect 16011 39031 16053 39040
rect 15627 38912 15669 38921
rect 15627 38872 15628 38912
rect 15668 38872 15669 38912
rect 15627 38863 15669 38872
rect 16300 38912 16340 39283
rect 15628 38778 15668 38863
rect 16300 38837 16340 38872
rect 16299 38828 16341 38837
rect 16299 38788 16300 38828
rect 16340 38788 16341 38828
rect 16299 38779 16341 38788
rect 15820 38744 15860 38753
rect 15532 38240 15572 38249
rect 15820 38240 15860 38704
rect 16012 38744 16052 38753
rect 16012 38417 16052 38704
rect 16011 38408 16053 38417
rect 16011 38368 16012 38408
rect 16052 38368 16053 38408
rect 16011 38359 16053 38368
rect 15915 38240 15957 38249
rect 15572 38200 15668 38240
rect 15820 38200 15916 38240
rect 15956 38200 15957 38240
rect 15532 38191 15572 38200
rect 15531 38072 15573 38081
rect 15531 38032 15532 38072
rect 15572 38032 15573 38072
rect 15531 38023 15573 38032
rect 15532 37938 15572 38023
rect 15628 37913 15668 38200
rect 15915 38191 15957 38200
rect 16012 38240 16052 38249
rect 15916 38106 15956 38191
rect 15724 37988 15764 37997
rect 15627 37904 15669 37913
rect 15627 37864 15628 37904
rect 15668 37864 15669 37904
rect 15627 37855 15669 37864
rect 15051 37652 15093 37661
rect 15051 37612 15052 37652
rect 15092 37612 15093 37652
rect 15051 37603 15093 37612
rect 15435 37652 15477 37661
rect 15435 37612 15436 37652
rect 15476 37612 15477 37652
rect 15435 37603 15477 37612
rect 15052 37148 15092 37603
rect 15531 37568 15573 37577
rect 15531 37528 15532 37568
rect 15572 37528 15573 37568
rect 15531 37519 15573 37528
rect 15147 37400 15189 37409
rect 15147 37360 15148 37400
rect 15188 37360 15189 37400
rect 15147 37351 15189 37360
rect 15435 37400 15477 37409
rect 15435 37360 15436 37400
rect 15476 37360 15477 37400
rect 15435 37351 15477 37360
rect 15532 37400 15572 37519
rect 15148 37266 15188 37351
rect 15436 37266 15476 37351
rect 15532 37241 15572 37360
rect 15531 37232 15573 37241
rect 15531 37192 15532 37232
rect 15572 37192 15573 37232
rect 15531 37183 15573 37192
rect 15052 37108 15188 37148
rect 15148 36844 15188 37108
rect 15052 36737 15092 36822
rect 15148 36737 15196 36844
rect 15051 36728 15093 36737
rect 15051 36688 15052 36728
rect 15092 36688 15093 36728
rect 15051 36679 15093 36688
rect 15148 36728 15197 36737
rect 15148 36688 15156 36728
rect 15196 36688 15197 36728
rect 15148 36686 15197 36688
rect 15188 36679 15197 36686
rect 15436 36728 15476 36737
rect 15532 36728 15572 37183
rect 15627 37148 15669 37157
rect 15627 37108 15628 37148
rect 15668 37108 15669 37148
rect 15627 37099 15669 37108
rect 15476 36688 15572 36728
rect 15436 36679 15476 36688
rect 15148 36637 15188 36646
rect 15340 36644 15380 36653
rect 15051 36560 15093 36569
rect 15051 36520 15052 36560
rect 15092 36520 15093 36560
rect 15051 36511 15093 36520
rect 15244 36560 15284 36569
rect 14860 36016 14996 36056
rect 14764 35720 14804 35731
rect 14764 35645 14804 35680
rect 14763 35636 14805 35645
rect 14763 35596 14764 35636
rect 14804 35596 14805 35636
rect 14763 35587 14805 35596
rect 14667 35300 14709 35309
rect 14667 35260 14668 35300
rect 14708 35260 14709 35300
rect 14667 35251 14709 35260
rect 14475 35216 14517 35225
rect 14475 35176 14476 35216
rect 14516 35176 14517 35216
rect 14475 35167 14517 35176
rect 14380 34999 14420 35008
rect 14476 34385 14516 35167
rect 14571 35132 14613 35141
rect 14571 35092 14572 35132
rect 14612 35092 14613 35132
rect 14571 35083 14613 35092
rect 14572 34998 14612 35083
rect 14668 34805 14708 35251
rect 14860 35048 14900 36016
rect 14956 35888 14996 35897
rect 14956 35309 14996 35848
rect 14955 35300 14997 35309
rect 14955 35260 14956 35300
rect 14996 35260 14997 35300
rect 14955 35251 14997 35260
rect 15052 35216 15092 36511
rect 15052 35132 15092 35176
rect 15244 35141 15284 36520
rect 15340 36485 15380 36604
rect 15435 36560 15477 36569
rect 15435 36520 15436 36560
rect 15476 36520 15477 36560
rect 15628 36560 15668 37099
rect 15724 36737 15764 37948
rect 15915 37988 15957 37997
rect 15915 37948 15916 37988
rect 15956 37948 15957 37988
rect 15915 37939 15957 37948
rect 15820 37568 15860 37577
rect 15820 36905 15860 37528
rect 15916 37409 15956 37939
rect 15915 37400 15957 37409
rect 15915 37360 15916 37400
rect 15956 37360 15957 37400
rect 15915 37351 15957 37360
rect 16012 37232 16052 38200
rect 16108 38240 16148 38249
rect 16108 37829 16148 38200
rect 16204 38240 16244 38249
rect 16396 38240 16436 38249
rect 16244 38200 16396 38240
rect 16204 38191 16244 38200
rect 16396 38191 16436 38200
rect 16395 38072 16437 38081
rect 16395 38032 16396 38072
rect 16436 38032 16437 38072
rect 16395 38023 16437 38032
rect 16396 37938 16436 38023
rect 16492 37829 16532 40888
rect 16588 40508 16628 41551
rect 16684 40769 16724 41728
rect 16780 41609 16820 42928
rect 16875 41684 16917 41693
rect 16875 41644 16876 41684
rect 16916 41644 16917 41684
rect 16875 41635 16917 41644
rect 16779 41600 16821 41609
rect 16779 41560 16780 41600
rect 16820 41560 16821 41600
rect 16779 41551 16821 41560
rect 16779 41348 16821 41357
rect 16779 41308 16780 41348
rect 16820 41308 16821 41348
rect 16779 41299 16821 41308
rect 16683 40760 16725 40769
rect 16683 40720 16684 40760
rect 16724 40720 16725 40760
rect 16683 40711 16725 40720
rect 16780 40592 16820 41299
rect 16876 40676 16916 41635
rect 16972 41609 17012 42928
rect 16971 41600 17013 41609
rect 16971 41560 16972 41600
rect 17012 41560 17013 41600
rect 16971 41551 17013 41560
rect 17164 41357 17204 42928
rect 17356 41861 17396 42928
rect 17548 42281 17588 42928
rect 17740 42281 17780 42928
rect 17835 42356 17877 42365
rect 17835 42316 17836 42356
rect 17876 42316 17877 42356
rect 17835 42307 17877 42316
rect 17547 42272 17589 42281
rect 17547 42232 17548 42272
rect 17588 42232 17589 42272
rect 17547 42223 17589 42232
rect 17739 42272 17781 42281
rect 17739 42232 17740 42272
rect 17780 42232 17781 42272
rect 17739 42223 17781 42232
rect 17739 41936 17781 41945
rect 17739 41896 17740 41936
rect 17780 41896 17781 41936
rect 17739 41887 17781 41896
rect 17355 41852 17397 41861
rect 17355 41812 17356 41852
rect 17396 41812 17397 41852
rect 17355 41803 17397 41812
rect 17259 41768 17301 41777
rect 17259 41728 17260 41768
rect 17300 41728 17301 41768
rect 17259 41719 17301 41728
rect 17163 41348 17205 41357
rect 17163 41308 17164 41348
rect 17204 41308 17205 41348
rect 17163 41299 17205 41308
rect 16972 41264 17012 41273
rect 16972 40853 17012 41224
rect 17163 41012 17205 41021
rect 17163 40972 17164 41012
rect 17204 40972 17205 41012
rect 17163 40963 17205 40972
rect 17164 40878 17204 40963
rect 16971 40844 17013 40853
rect 16971 40804 16972 40844
rect 17012 40804 17013 40844
rect 16971 40795 17013 40804
rect 16876 40636 17012 40676
rect 16588 40459 16628 40468
rect 16684 40552 16820 40592
rect 16684 40349 16724 40552
rect 16972 40508 17012 40636
rect 17163 40592 17205 40601
rect 17163 40552 17164 40592
rect 17204 40552 17205 40592
rect 17163 40543 17205 40552
rect 16972 40459 17012 40468
rect 17164 40458 17204 40543
rect 17260 40508 17300 41719
rect 17355 41516 17397 41525
rect 17355 41476 17356 41516
rect 17396 41476 17397 41516
rect 17355 41467 17397 41476
rect 17356 41180 17396 41467
rect 17643 41348 17685 41357
rect 17643 41308 17644 41348
rect 17684 41308 17685 41348
rect 17643 41299 17685 41308
rect 17356 41131 17396 41140
rect 17547 41012 17589 41021
rect 17547 40972 17548 41012
rect 17588 40972 17589 41012
rect 17547 40963 17589 40972
rect 17548 40878 17588 40963
rect 17547 40592 17589 40601
rect 17547 40552 17548 40592
rect 17588 40552 17589 40592
rect 17547 40543 17589 40552
rect 17356 40508 17396 40517
rect 17260 40468 17356 40508
rect 17356 40459 17396 40468
rect 17548 40458 17588 40543
rect 17644 40508 17684 41299
rect 17740 41180 17780 41887
rect 17836 41180 17876 42307
rect 17932 41525 17972 42928
rect 18124 41609 18164 42928
rect 18316 41777 18356 42928
rect 18411 42272 18453 42281
rect 18411 42232 18412 42272
rect 18452 42232 18453 42272
rect 18411 42223 18453 42232
rect 18315 41768 18357 41777
rect 18315 41728 18316 41768
rect 18356 41728 18357 41768
rect 18315 41719 18357 41728
rect 18123 41600 18165 41609
rect 18123 41560 18124 41600
rect 18164 41560 18165 41600
rect 18123 41551 18165 41560
rect 17931 41516 17973 41525
rect 17931 41476 17932 41516
rect 17972 41476 17973 41516
rect 17931 41467 17973 41476
rect 18219 41516 18261 41525
rect 18219 41476 18220 41516
rect 18260 41476 18261 41516
rect 18219 41467 18261 41476
rect 18124 41180 18164 41189
rect 17836 41140 18124 41180
rect 17740 41131 17780 41140
rect 18124 41131 18164 41140
rect 17931 41012 17973 41021
rect 17931 40972 17932 41012
rect 17972 40972 17973 41012
rect 17931 40963 17973 40972
rect 17932 40878 17972 40963
rect 18123 40928 18165 40937
rect 18123 40888 18124 40928
rect 18164 40888 18165 40928
rect 18123 40879 18165 40888
rect 17931 40592 17973 40601
rect 17931 40552 17932 40592
rect 17972 40552 17973 40592
rect 17931 40543 17973 40552
rect 17740 40508 17780 40517
rect 17644 40468 17740 40508
rect 17740 40459 17780 40468
rect 17932 40458 17972 40543
rect 18124 40508 18164 40879
rect 18220 40760 18260 41467
rect 18315 41012 18357 41021
rect 18315 40972 18316 41012
rect 18356 40972 18357 41012
rect 18315 40963 18357 40972
rect 18316 40878 18356 40963
rect 18220 40720 18356 40760
rect 18124 40459 18164 40468
rect 16683 40340 16725 40349
rect 16683 40300 16684 40340
rect 16724 40300 16725 40340
rect 16683 40291 16725 40300
rect 17163 40340 17205 40349
rect 17163 40300 17164 40340
rect 17204 40300 17205 40340
rect 17163 40291 17205 40300
rect 16780 40256 16820 40265
rect 16780 39929 16820 40216
rect 16779 39920 16821 39929
rect 17164 39920 17204 40291
rect 17259 40172 17301 40181
rect 17259 40132 17260 40172
rect 17300 40132 17301 40172
rect 17259 40123 17301 40132
rect 16779 39880 16780 39920
rect 16820 39880 16821 39920
rect 16779 39871 16821 39880
rect 16972 39880 17204 39920
rect 16587 39668 16629 39677
rect 16587 39628 16588 39668
rect 16628 39628 16629 39668
rect 16587 39619 16629 39628
rect 16684 39668 16724 39677
rect 16588 39534 16628 39619
rect 16684 38501 16724 39628
rect 16683 38492 16725 38501
rect 16683 38452 16684 38492
rect 16724 38452 16725 38492
rect 16683 38443 16725 38452
rect 16587 38408 16629 38417
rect 16587 38368 16588 38408
rect 16628 38368 16629 38408
rect 16587 38359 16629 38368
rect 16588 38226 16628 38359
rect 16684 38240 16724 38249
rect 16875 38240 16917 38249
rect 16724 38200 16820 38235
rect 16684 38195 16820 38200
rect 16684 38191 16724 38195
rect 16588 38177 16628 38186
rect 16107 37820 16149 37829
rect 16107 37780 16108 37820
rect 16148 37780 16149 37820
rect 16107 37771 16149 37780
rect 16491 37820 16533 37829
rect 16491 37780 16492 37820
rect 16532 37780 16533 37820
rect 16491 37771 16533 37780
rect 16108 37652 16148 37771
rect 16683 37736 16725 37745
rect 16683 37696 16684 37736
rect 16724 37696 16725 37736
rect 16683 37687 16725 37696
rect 16587 37652 16629 37661
rect 16108 37612 16244 37652
rect 16108 37409 16148 37494
rect 16204 37493 16244 37612
rect 16587 37612 16588 37652
rect 16628 37612 16629 37652
rect 16587 37603 16629 37612
rect 16203 37484 16245 37493
rect 16203 37444 16204 37484
rect 16244 37444 16245 37484
rect 16203 37435 16245 37444
rect 16107 37400 16149 37409
rect 16107 37360 16108 37400
rect 16148 37360 16149 37400
rect 16107 37351 16149 37360
rect 16396 37400 16436 37409
rect 16012 37192 16340 37232
rect 16107 36980 16149 36989
rect 16107 36940 16108 36980
rect 16148 36940 16149 36980
rect 16107 36931 16149 36940
rect 15819 36896 15861 36905
rect 15819 36856 15820 36896
rect 15860 36856 15861 36896
rect 15819 36847 15861 36856
rect 15723 36728 15765 36737
rect 15723 36688 15724 36728
rect 15764 36688 15765 36728
rect 15723 36679 15765 36688
rect 15820 36728 15860 36737
rect 15820 36569 15860 36688
rect 15916 36728 15956 36737
rect 15819 36560 15861 36569
rect 15628 36520 15820 36560
rect 15860 36520 15861 36560
rect 15435 36511 15477 36520
rect 15819 36511 15861 36520
rect 15339 36476 15381 36485
rect 15339 36436 15340 36476
rect 15380 36436 15381 36476
rect 15339 36427 15381 36436
rect 15339 35636 15381 35645
rect 15339 35596 15340 35636
rect 15380 35596 15381 35636
rect 15339 35587 15381 35596
rect 15340 35216 15380 35587
rect 15243 35132 15285 35141
rect 15052 35092 15188 35132
rect 14860 35008 15092 35048
rect 14763 34964 14805 34973
rect 14763 34924 14764 34964
rect 14804 34924 14805 34964
rect 14763 34915 14805 34924
rect 14764 34830 14804 34915
rect 14667 34796 14709 34805
rect 14667 34756 14668 34796
rect 14708 34756 14709 34796
rect 14667 34747 14709 34756
rect 14571 34712 14613 34721
rect 14571 34672 14572 34712
rect 14612 34672 14613 34712
rect 14571 34663 14613 34672
rect 14475 34376 14517 34385
rect 14475 34336 14476 34376
rect 14516 34336 14517 34376
rect 14475 34327 14517 34336
rect 14476 34208 14516 34217
rect 13900 33580 14036 33620
rect 14092 33916 14324 33956
rect 14380 34168 14476 34208
rect 13803 33452 13845 33461
rect 13803 33412 13804 33452
rect 13844 33412 13845 33452
rect 13803 33403 13845 33412
rect 13803 32948 13845 32957
rect 13803 32908 13804 32948
rect 13844 32908 13845 32948
rect 13803 32899 13845 32908
rect 13804 32285 13844 32899
rect 13900 32696 13940 33580
rect 13996 33452 14036 33461
rect 14092 33452 14132 33916
rect 14188 33704 14228 33715
rect 14188 33629 14228 33664
rect 14283 33704 14325 33713
rect 14283 33664 14284 33704
rect 14324 33664 14325 33704
rect 14283 33655 14325 33664
rect 14187 33620 14229 33629
rect 14187 33580 14188 33620
rect 14228 33580 14229 33620
rect 14187 33571 14229 33580
rect 14284 33570 14324 33655
rect 14380 33629 14420 34168
rect 14476 34159 14516 34168
rect 14476 33704 14516 33713
rect 14379 33620 14421 33629
rect 14379 33580 14380 33620
rect 14420 33580 14421 33620
rect 14379 33571 14421 33580
rect 14379 33452 14421 33461
rect 14092 33412 14324 33452
rect 13996 32873 14036 33412
rect 14187 33284 14229 33293
rect 14187 33244 14188 33284
rect 14228 33244 14229 33284
rect 14187 33235 14229 33244
rect 13995 32864 14037 32873
rect 13995 32824 13996 32864
rect 14036 32824 14037 32864
rect 13995 32815 14037 32824
rect 14092 32864 14132 32873
rect 14092 32696 14132 32824
rect 13900 32656 14132 32696
rect 13803 32276 13845 32285
rect 13803 32236 13804 32276
rect 13844 32236 13845 32276
rect 13803 32227 13845 32236
rect 13996 32192 14036 32201
rect 14188 32192 14228 33235
rect 13900 32152 13996 32192
rect 14036 32152 14228 32192
rect 13900 31688 13940 32152
rect 13996 32143 14036 32152
rect 13612 31648 13940 31688
rect 14188 31940 14228 31949
rect 13612 31529 13652 31648
rect 14188 31529 14228 31900
rect 14284 31856 14324 33412
rect 14379 33412 14380 33452
rect 14420 33412 14421 33452
rect 14379 33403 14421 33412
rect 14380 32948 14420 33403
rect 14476 33125 14516 33664
rect 14572 33704 14612 34663
rect 14668 34376 14708 34385
rect 14668 34049 14708 34336
rect 14955 34124 14997 34133
rect 14955 34084 14956 34124
rect 14996 34084 14997 34124
rect 14955 34075 14997 34084
rect 14667 34040 14709 34049
rect 14667 34000 14668 34040
rect 14708 34000 14709 34040
rect 14667 33991 14709 34000
rect 14668 33872 14708 33881
rect 14859 33872 14901 33881
rect 14708 33832 14804 33872
rect 14668 33823 14708 33832
rect 14572 33545 14612 33664
rect 14673 33704 14713 33713
rect 14571 33536 14613 33545
rect 14571 33496 14572 33536
rect 14612 33496 14613 33536
rect 14571 33487 14613 33496
rect 14673 33368 14713 33664
rect 14572 33328 14713 33368
rect 14475 33116 14517 33125
rect 14475 33076 14476 33116
rect 14516 33076 14517 33116
rect 14475 33067 14517 33076
rect 14476 32948 14516 32957
rect 14380 32908 14476 32948
rect 14476 32201 14516 32908
rect 14475 32192 14517 32201
rect 14475 32152 14476 32192
rect 14516 32152 14517 32192
rect 14475 32143 14517 32152
rect 14380 32024 14420 32033
rect 14572 32024 14612 33328
rect 14667 33032 14709 33041
rect 14667 32992 14668 33032
rect 14708 32992 14709 33032
rect 14667 32983 14709 32992
rect 14668 32898 14708 32983
rect 14667 32696 14709 32705
rect 14667 32656 14668 32696
rect 14708 32656 14709 32696
rect 14667 32647 14709 32656
rect 14420 31984 14612 32024
rect 14668 32192 14708 32647
rect 14764 32369 14804 33832
rect 14859 33832 14860 33872
rect 14900 33832 14901 33872
rect 14859 33823 14901 33832
rect 14860 32948 14900 33823
rect 14860 32899 14900 32908
rect 14956 33536 14996 34075
rect 14763 32360 14805 32369
rect 14956 32360 14996 33496
rect 15052 33116 15092 35008
rect 15148 34889 15188 35092
rect 15243 35092 15244 35132
rect 15284 35092 15285 35132
rect 15243 35083 15285 35092
rect 15147 34880 15189 34889
rect 15147 34840 15148 34880
rect 15188 34840 15189 34880
rect 15147 34831 15189 34840
rect 15340 34133 15380 35176
rect 15436 35216 15476 36511
rect 15531 36476 15573 36485
rect 15531 36436 15532 36476
rect 15572 36436 15764 36476
rect 15531 36427 15573 36436
rect 15531 36224 15573 36233
rect 15531 36184 15532 36224
rect 15572 36184 15573 36224
rect 15531 36175 15573 36184
rect 15339 34124 15381 34133
rect 15339 34084 15340 34124
rect 15380 34084 15381 34124
rect 15339 34075 15381 34084
rect 15436 34049 15476 35176
rect 15532 35057 15572 36175
rect 15627 35300 15669 35309
rect 15627 35260 15628 35300
rect 15668 35260 15669 35300
rect 15627 35251 15669 35260
rect 15531 35048 15573 35057
rect 15531 35008 15532 35048
rect 15572 35008 15573 35048
rect 15531 34999 15573 35008
rect 15435 34040 15477 34049
rect 15435 34000 15436 34040
rect 15476 34000 15477 34040
rect 15435 33991 15477 34000
rect 15531 33704 15573 33713
rect 15531 33664 15532 33704
rect 15572 33664 15573 33704
rect 15531 33655 15573 33664
rect 15628 33704 15668 35251
rect 15724 35216 15764 36436
rect 15820 36426 15860 36511
rect 15916 36485 15956 36688
rect 16108 36728 16148 36931
rect 16300 36896 16340 37192
rect 16396 36989 16436 37360
rect 16491 37316 16533 37325
rect 16491 37276 16492 37316
rect 16532 37276 16533 37316
rect 16491 37267 16533 37276
rect 16492 37182 16532 37267
rect 16395 36980 16437 36989
rect 16588 36980 16628 37603
rect 16395 36940 16396 36980
rect 16436 36940 16437 36980
rect 16395 36931 16437 36940
rect 16492 36940 16628 36980
rect 16300 36847 16340 36856
rect 16396 36749 16436 36758
rect 16108 36679 16148 36688
rect 16299 36728 16341 36737
rect 16299 36688 16300 36728
rect 16340 36709 16396 36728
rect 16340 36688 16436 36709
rect 16492 36728 16532 36940
rect 16299 36679 16341 36688
rect 16492 36644 16532 36688
rect 16396 36604 16532 36644
rect 16588 36728 16628 36737
rect 15915 36476 15957 36485
rect 15915 36436 15916 36476
rect 15956 36436 15957 36476
rect 15915 36427 15957 36436
rect 16108 36476 16148 36485
rect 16011 36392 16053 36401
rect 16011 36352 16012 36392
rect 16052 36352 16053 36392
rect 16011 36343 16053 36352
rect 15724 35176 15956 35216
rect 15723 35048 15765 35057
rect 15723 35008 15724 35048
rect 15764 35008 15765 35048
rect 15723 34999 15765 35008
rect 15916 35048 15956 35176
rect 15916 34999 15956 35008
rect 15724 34914 15764 34999
rect 15723 34712 15765 34721
rect 15723 34672 15724 34712
rect 15764 34672 15765 34712
rect 15723 34663 15765 34672
rect 15628 33655 15668 33664
rect 15147 33620 15189 33629
rect 15147 33580 15148 33620
rect 15188 33580 15189 33620
rect 15147 33571 15189 33580
rect 15052 33067 15092 33076
rect 15051 32864 15093 32873
rect 15051 32824 15052 32864
rect 15092 32824 15093 32864
rect 15051 32815 15093 32824
rect 14763 32320 14764 32360
rect 14804 32320 14805 32360
rect 14763 32311 14805 32320
rect 14860 32320 14996 32360
rect 14860 32276 14900 32320
rect 14857 32236 14900 32276
rect 14380 31975 14420 31984
rect 14284 31816 14516 31856
rect 14283 31688 14325 31697
rect 14283 31648 14284 31688
rect 14324 31648 14325 31688
rect 14283 31639 14325 31648
rect 13611 31520 13653 31529
rect 13516 31445 13556 31487
rect 13611 31480 13612 31520
rect 13652 31480 13653 31520
rect 13611 31471 13653 31480
rect 13803 31520 13845 31529
rect 13803 31480 13804 31520
rect 13844 31480 13845 31520
rect 13803 31471 13845 31480
rect 14187 31520 14229 31529
rect 14187 31480 14188 31520
rect 14228 31480 14229 31520
rect 14187 31471 14229 31480
rect 13515 31436 13557 31445
rect 13515 31396 13516 31436
rect 13556 31396 13557 31436
rect 13515 31392 13557 31396
rect 13515 31387 13516 31392
rect 13419 31352 13461 31361
rect 13419 31312 13420 31352
rect 13460 31312 13461 31352
rect 13556 31387 13557 31392
rect 13516 31343 13556 31352
rect 13612 31352 13652 31361
rect 13419 31303 13461 31312
rect 13420 31184 13460 31193
rect 13323 30092 13365 30101
rect 13323 30052 13324 30092
rect 13364 30052 13365 30092
rect 13323 30043 13365 30052
rect 13227 29924 13269 29933
rect 13227 29884 13228 29924
rect 13268 29884 13269 29924
rect 13227 29875 13269 29884
rect 13420 29849 13460 31144
rect 13612 30773 13652 31312
rect 13708 31352 13748 31361
rect 13708 31109 13748 31312
rect 13707 31100 13749 31109
rect 13707 31060 13708 31100
rect 13748 31060 13749 31100
rect 13707 31051 13749 31060
rect 13611 30764 13653 30773
rect 13611 30724 13612 30764
rect 13652 30724 13653 30764
rect 13611 30715 13653 30724
rect 13804 30680 13844 31471
rect 13995 31436 14037 31445
rect 13995 31396 13996 31436
rect 14036 31396 14037 31436
rect 13995 31387 14037 31396
rect 13900 31352 13940 31361
rect 13900 30932 13940 31312
rect 13996 31268 14036 31387
rect 13996 31219 14036 31228
rect 14092 31352 14132 31361
rect 14092 31193 14132 31312
rect 14187 31352 14229 31361
rect 14187 31312 14188 31352
rect 14228 31312 14229 31352
rect 14187 31303 14229 31312
rect 14188 31218 14228 31303
rect 14091 31184 14133 31193
rect 14091 31144 14092 31184
rect 14132 31144 14133 31184
rect 14091 31135 14133 31144
rect 13900 30892 14036 30932
rect 13899 30764 13941 30773
rect 13899 30724 13900 30764
rect 13940 30724 13941 30764
rect 13899 30715 13941 30724
rect 13756 30670 13844 30680
rect 13796 30640 13844 30670
rect 13900 30630 13940 30715
rect 13756 30621 13796 30630
rect 13996 30521 14036 30892
rect 14092 30596 14132 31135
rect 14187 31016 14229 31025
rect 14187 30976 14188 31016
rect 14228 30976 14229 31016
rect 14187 30967 14229 30976
rect 14188 30691 14228 30967
rect 14188 30642 14228 30651
rect 14092 30556 14228 30596
rect 13707 30512 13749 30521
rect 13707 30472 13708 30512
rect 13748 30472 13749 30512
rect 13707 30463 13749 30472
rect 13995 30512 14037 30521
rect 13995 30472 13996 30512
rect 14036 30472 14037 30512
rect 13995 30463 14037 30472
rect 13611 30092 13653 30101
rect 13611 30052 13612 30092
rect 13652 30052 13653 30092
rect 13611 30043 13653 30052
rect 13612 29933 13652 30043
rect 13611 29924 13653 29933
rect 13611 29884 13612 29924
rect 13652 29884 13653 29924
rect 13611 29875 13653 29884
rect 13132 29805 13172 29814
rect 13419 29840 13461 29849
rect 13419 29800 13420 29840
rect 13460 29800 13461 29840
rect 13419 29791 13461 29800
rect 13708 29840 13748 30463
rect 14092 30428 14132 30437
rect 13995 30344 14037 30353
rect 14092 30344 14132 30388
rect 13995 30304 13996 30344
rect 14036 30304 14132 30344
rect 13995 30295 14037 30304
rect 14188 30260 14228 30556
rect 14092 30220 14228 30260
rect 14092 29924 14132 30220
rect 13996 29884 14132 29924
rect 14187 29924 14229 29933
rect 14187 29884 14188 29924
rect 14228 29884 14229 29924
rect 13708 29791 13748 29800
rect 13804 29840 13844 29851
rect 13804 29765 13844 29800
rect 13899 29840 13941 29849
rect 13899 29800 13900 29840
rect 13940 29800 13941 29840
rect 13899 29791 13941 29800
rect 13996 29840 14036 29884
rect 14187 29875 14229 29884
rect 13996 29791 14036 29800
rect 14188 29840 14228 29875
rect 13323 29756 13365 29765
rect 13323 29716 13324 29756
rect 13364 29716 13365 29756
rect 13323 29707 13365 29716
rect 13803 29756 13845 29765
rect 13803 29716 13804 29756
rect 13844 29716 13845 29756
rect 13803 29707 13845 29716
rect 13324 29622 13364 29707
rect 13900 29706 13940 29791
rect 13611 29504 13653 29513
rect 13611 29464 13612 29504
rect 13652 29464 13653 29504
rect 13611 29455 13653 29464
rect 13323 29420 13365 29429
rect 13036 29380 13324 29420
rect 13364 29380 13365 29420
rect 13323 29371 13365 29380
rect 13036 29296 13268 29336
rect 13036 29168 13076 29296
rect 13036 29119 13076 29128
rect 13132 29168 13172 29177
rect 13036 29000 13076 29009
rect 13036 28328 13076 28960
rect 13132 28589 13172 29128
rect 13228 28925 13268 29296
rect 13323 29168 13365 29177
rect 13323 29128 13324 29168
rect 13364 29128 13365 29168
rect 13323 29119 13365 29128
rect 13612 29168 13652 29455
rect 13803 29420 13845 29429
rect 13803 29380 13804 29420
rect 13844 29380 13845 29420
rect 13803 29371 13845 29380
rect 13612 29119 13652 29128
rect 13324 29034 13364 29119
rect 13804 29000 13844 29371
rect 13995 29168 14037 29177
rect 13995 29128 13996 29168
rect 14036 29128 14037 29168
rect 13995 29119 14037 29128
rect 13612 28960 13844 29000
rect 13227 28916 13269 28925
rect 13227 28876 13228 28916
rect 13268 28876 13269 28916
rect 13227 28867 13269 28876
rect 13420 28916 13460 28925
rect 13131 28580 13173 28589
rect 13131 28540 13132 28580
rect 13172 28540 13173 28580
rect 13131 28531 13173 28540
rect 13036 28279 13076 28288
rect 13132 28328 13172 28337
rect 13228 28328 13268 28867
rect 13172 28288 13268 28328
rect 13323 28328 13365 28337
rect 13323 28288 13324 28328
rect 13364 28288 13365 28328
rect 13132 28279 13172 28288
rect 13323 28279 13365 28288
rect 13420 28328 13460 28876
rect 13520 28580 13562 28589
rect 13520 28540 13521 28580
rect 13561 28540 13562 28580
rect 13520 28531 13562 28540
rect 13420 28279 13460 28288
rect 13521 28328 13561 28531
rect 13324 28194 13364 28279
rect 13035 28160 13077 28169
rect 13035 28120 13036 28160
rect 13076 28120 13077 28160
rect 13035 28111 13077 28120
rect 13420 28160 13460 28169
rect 13036 24884 13076 28111
rect 13131 27656 13173 27665
rect 13131 27616 13132 27656
rect 13172 27616 13173 27656
rect 13131 27607 13173 27616
rect 13132 27522 13172 27607
rect 13420 27413 13460 28120
rect 13521 28076 13561 28288
rect 13612 28169 13652 28960
rect 13707 28328 13749 28337
rect 13707 28288 13708 28328
rect 13748 28288 13749 28328
rect 13707 28279 13749 28288
rect 13996 28328 14036 29119
rect 14188 29093 14228 29800
rect 14284 29597 14324 31639
rect 14379 31520 14421 31529
rect 14379 31480 14380 31520
rect 14420 31480 14421 31520
rect 14379 31471 14421 31480
rect 14380 31184 14420 31471
rect 14380 30941 14420 31144
rect 14379 30932 14421 30941
rect 14379 30892 14380 30932
rect 14420 30892 14421 30932
rect 14379 30883 14421 30892
rect 14380 30848 14420 30883
rect 14380 30768 14420 30808
rect 14379 29840 14421 29849
rect 14379 29800 14380 29840
rect 14420 29800 14421 29840
rect 14379 29791 14421 29800
rect 14283 29588 14325 29597
rect 14283 29548 14284 29588
rect 14324 29548 14325 29588
rect 14283 29539 14325 29548
rect 14283 29252 14325 29261
rect 14283 29212 14284 29252
rect 14324 29212 14325 29252
rect 14283 29203 14325 29212
rect 14187 29084 14229 29093
rect 14187 29044 14188 29084
rect 14228 29044 14229 29084
rect 14187 29035 14229 29044
rect 13611 28160 13653 28169
rect 13611 28120 13612 28160
rect 13652 28120 13653 28160
rect 13611 28111 13653 28120
rect 13516 28036 13561 28076
rect 13516 27656 13556 28036
rect 13708 27992 13748 28279
rect 13804 28169 13844 28254
rect 13803 28160 13845 28169
rect 13803 28120 13804 28160
rect 13844 28120 13940 28160
rect 13803 28111 13845 28120
rect 13708 27952 13844 27992
rect 13707 27824 13749 27833
rect 13707 27784 13708 27824
rect 13748 27784 13749 27824
rect 13707 27775 13749 27784
rect 13804 27824 13844 27952
rect 13804 27775 13844 27784
rect 13611 27740 13653 27749
rect 13611 27700 13612 27740
rect 13652 27700 13653 27740
rect 13611 27691 13653 27700
rect 13516 27607 13556 27616
rect 13612 27656 13652 27691
rect 13612 27605 13652 27616
rect 13515 27488 13557 27497
rect 13708 27488 13748 27775
rect 13803 27572 13845 27581
rect 13803 27532 13804 27572
rect 13844 27532 13845 27572
rect 13803 27523 13845 27532
rect 13515 27448 13516 27488
rect 13556 27448 13557 27488
rect 13515 27439 13557 27448
rect 13612 27448 13748 27488
rect 13324 27404 13364 27413
rect 13324 26835 13364 27364
rect 13419 27404 13461 27413
rect 13419 27364 13420 27404
rect 13460 27364 13461 27404
rect 13419 27355 13461 27364
rect 13298 26834 13364 26835
rect 13276 26825 13364 26834
rect 13420 26825 13460 27355
rect 13316 26795 13364 26825
rect 13419 26816 13461 26825
rect 13316 26785 13338 26795
rect 13276 26776 13316 26785
rect 13419 26776 13420 26816
rect 13460 26776 13461 26816
rect 13419 26767 13461 26776
rect 13227 26648 13269 26657
rect 13227 26608 13228 26648
rect 13268 26608 13269 26648
rect 13227 26599 13269 26608
rect 13419 26648 13461 26657
rect 13419 26608 13420 26648
rect 13460 26608 13461 26648
rect 13419 26599 13461 26608
rect 13228 25304 13268 26599
rect 13420 26514 13460 26599
rect 13036 24844 13172 24884
rect 13036 24641 13076 24726
rect 13035 24632 13077 24641
rect 13035 24592 13036 24632
rect 13076 24592 13077 24632
rect 13035 24583 13077 24592
rect 12940 24424 13076 24464
rect 12843 24212 12885 24221
rect 12843 24172 12844 24212
rect 12884 24172 12885 24212
rect 12843 24163 12885 24172
rect 12843 24044 12885 24053
rect 12843 24004 12844 24044
rect 12884 24004 12885 24044
rect 12843 23995 12885 24004
rect 12747 23792 12789 23801
rect 12747 23752 12748 23792
rect 12788 23752 12789 23792
rect 12747 23743 12789 23752
rect 12556 23500 12692 23540
rect 12459 23288 12501 23297
rect 12268 23248 12404 23288
rect 12364 23204 12404 23248
rect 12459 23248 12460 23288
rect 12500 23248 12501 23288
rect 12459 23239 12501 23248
rect 12364 23155 12404 23164
rect 12268 23120 12308 23129
rect 12172 23080 12268 23120
rect 11980 23071 12020 23080
rect 12268 23071 12308 23080
rect 11883 22700 11925 22709
rect 11883 22660 11884 22700
rect 11924 22660 11925 22700
rect 11883 22651 11925 22660
rect 11404 22324 11540 22364
rect 11308 22231 11348 22240
rect 11020 22146 11060 22231
rect 11403 22196 11445 22205
rect 11403 22156 11404 22196
rect 11444 22156 11445 22196
rect 11403 22147 11445 22156
rect 10732 22112 10772 22123
rect 10732 22037 10772 22072
rect 11404 22062 11444 22147
rect 10731 22028 10773 22037
rect 10731 21988 10732 22028
rect 10772 21988 10773 22028
rect 10731 21979 10773 21988
rect 11500 21953 11540 22324
rect 11596 22324 11828 22364
rect 10635 21944 10677 21953
rect 10635 21904 10636 21944
rect 10676 21904 10677 21944
rect 10635 21895 10677 21904
rect 11499 21944 11541 21953
rect 11499 21904 11500 21944
rect 11540 21904 11541 21944
rect 11499 21895 11541 21904
rect 11019 21860 11061 21869
rect 11019 21820 11020 21860
rect 11060 21820 11061 21860
rect 11019 21811 11061 21820
rect 10348 21559 10388 21568
rect 10539 21608 10581 21617
rect 10539 21568 10540 21608
rect 10580 21568 10581 21608
rect 10539 21559 10581 21568
rect 10252 21475 10292 21484
rect 9867 21440 9909 21449
rect 9867 21400 9868 21440
rect 9908 21400 9909 21440
rect 9867 21391 9909 21400
rect 10060 21390 10100 21475
rect 10156 21440 10196 21449
rect 10156 20945 10196 21400
rect 10443 21272 10485 21281
rect 10443 21232 10444 21272
rect 10484 21232 10485 21272
rect 10443 21223 10485 21232
rect 10251 21188 10293 21197
rect 10251 21148 10252 21188
rect 10292 21148 10293 21188
rect 10251 21139 10293 21148
rect 10155 20936 10197 20945
rect 10155 20896 10156 20936
rect 10196 20896 10197 20936
rect 10155 20887 10197 20896
rect 9772 20140 10100 20180
rect 9772 20012 9812 20021
rect 9772 19424 9812 19972
rect 9867 20012 9909 20021
rect 9867 19972 9868 20012
rect 9908 19972 9909 20012
rect 9867 19963 9909 19972
rect 9868 19878 9908 19963
rect 9580 19384 9812 19424
rect 9580 19256 9620 19384
rect 9580 17585 9620 19216
rect 9675 19256 9717 19265
rect 9675 19216 9676 19256
rect 9716 19216 9717 19256
rect 9675 19207 9717 19216
rect 9676 17669 9716 19207
rect 9771 18500 9813 18509
rect 9771 18460 9772 18500
rect 9812 18460 9813 18500
rect 9771 18451 9813 18460
rect 9675 17660 9717 17669
rect 9675 17620 9676 17660
rect 9716 17620 9717 17660
rect 9675 17611 9717 17620
rect 9579 17576 9621 17585
rect 9579 17536 9580 17576
rect 9620 17536 9621 17576
rect 9579 17527 9621 17536
rect 9772 17417 9812 18451
rect 9868 17749 9908 17758
rect 9771 17408 9813 17417
rect 9771 17368 9772 17408
rect 9812 17368 9813 17408
rect 9771 17359 9813 17368
rect 9388 17200 9524 17240
rect 9675 17240 9717 17249
rect 9675 17200 9676 17240
rect 9716 17200 9717 17240
rect 9388 16409 9428 17200
rect 9675 17191 9717 17200
rect 9676 17106 9716 17191
rect 9483 17072 9525 17081
rect 9868 17072 9908 17709
rect 10060 17660 10100 20140
rect 10155 20096 10197 20105
rect 10155 20056 10156 20096
rect 10196 20056 10197 20096
rect 10155 20047 10197 20056
rect 10156 19256 10196 20047
rect 10156 17753 10196 19216
rect 10155 17744 10197 17753
rect 10155 17704 10156 17744
rect 10196 17704 10197 17744
rect 10155 17695 10197 17704
rect 9963 17324 10005 17333
rect 9963 17284 9964 17324
rect 10004 17284 10005 17324
rect 9963 17275 10005 17284
rect 9964 17240 10004 17275
rect 9964 17189 10004 17200
rect 9483 17032 9484 17072
rect 9524 17032 9525 17072
rect 9483 17023 9525 17032
rect 9772 17032 9908 17072
rect 9484 16938 9524 17023
rect 9387 16400 9429 16409
rect 9387 16360 9388 16400
rect 9428 16360 9429 16400
rect 9387 16351 9429 16360
rect 9484 16316 9524 16325
rect 9524 16276 9620 16316
rect 9484 16267 9524 16276
rect 9292 16192 9428 16232
rect 9291 16064 9333 16073
rect 9291 16024 9292 16064
rect 9332 16024 9333 16064
rect 9291 16015 9333 16024
rect 9292 15930 9332 16015
rect 9196 15688 9332 15728
rect 9195 14216 9237 14225
rect 9195 14176 9196 14216
rect 9236 14176 9237 14216
rect 9195 14167 9237 14176
rect 9196 14082 9236 14167
rect 9100 12748 9236 12788
rect 9099 12620 9141 12629
rect 9099 12580 9100 12620
rect 9140 12580 9141 12620
rect 9099 12571 9141 12580
rect 9003 12284 9045 12293
rect 9003 12244 9004 12284
rect 9044 12244 9045 12284
rect 9003 12235 9045 12244
rect 9100 11948 9140 12571
rect 9004 11908 9140 11948
rect 9004 11360 9044 11908
rect 9099 11696 9141 11705
rect 9099 11656 9100 11696
rect 9140 11656 9141 11696
rect 9099 11647 9141 11656
rect 9100 11562 9140 11647
rect 9004 11320 9140 11360
rect 9100 11024 9140 11320
rect 9003 10100 9045 10109
rect 9100 10100 9140 10984
rect 9003 10060 9004 10100
rect 9044 10060 9140 10100
rect 9003 10051 9045 10060
rect 8907 9764 8949 9773
rect 8907 9724 8908 9764
rect 8948 9724 8949 9764
rect 8907 9715 8949 9724
rect 9004 9596 9044 10051
rect 9196 10016 9236 12748
rect 9292 12704 9332 15688
rect 9388 13376 9428 16192
rect 9483 15560 9525 15569
rect 9483 15520 9484 15560
rect 9524 15520 9525 15560
rect 9483 15511 9525 15520
rect 9484 15426 9524 15511
rect 9484 14725 9524 14734
rect 9484 14309 9524 14685
rect 9483 14300 9525 14309
rect 9483 14260 9484 14300
rect 9524 14260 9525 14300
rect 9483 14251 9525 14260
rect 9580 14225 9620 16276
rect 9676 15728 9716 15737
rect 9772 15728 9812 17032
rect 10060 16913 10100 17620
rect 9868 16904 9908 16913
rect 9868 16241 9908 16864
rect 10059 16904 10101 16913
rect 10059 16864 10060 16904
rect 10100 16864 10101 16904
rect 10059 16855 10101 16864
rect 10059 16400 10101 16409
rect 10059 16360 10060 16400
rect 10100 16360 10101 16400
rect 10059 16351 10101 16360
rect 9867 16232 9909 16241
rect 9867 16192 9868 16232
rect 9908 16192 9909 16232
rect 9867 16183 9909 16192
rect 9964 16232 10004 16241
rect 9716 15688 9812 15728
rect 9868 15728 9908 16183
rect 9676 15679 9716 15688
rect 9868 14888 9908 15688
rect 9964 15149 10004 16192
rect 10060 16232 10100 16351
rect 10060 16183 10100 16192
rect 9963 15140 10005 15149
rect 9963 15100 9964 15140
rect 10004 15100 10005 15140
rect 9963 15091 10005 15100
rect 9868 14839 9908 14848
rect 10156 14729 10196 17695
rect 10252 16325 10292 21139
rect 10347 20684 10389 20693
rect 10347 20644 10348 20684
rect 10388 20644 10389 20684
rect 10347 20635 10389 20644
rect 10348 20273 10388 20635
rect 10347 20264 10389 20273
rect 10347 20224 10348 20264
rect 10388 20224 10389 20264
rect 10347 20215 10389 20224
rect 10347 20096 10389 20105
rect 10347 20056 10348 20096
rect 10388 20056 10389 20096
rect 10347 20047 10389 20056
rect 10348 19962 10388 20047
rect 10444 16400 10484 21223
rect 11020 20936 11060 21811
rect 11115 21776 11157 21785
rect 11115 21736 11116 21776
rect 11156 21736 11157 21776
rect 11115 21727 11157 21736
rect 10732 20896 11060 20936
rect 10635 20768 10677 20777
rect 10635 20728 10636 20768
rect 10676 20728 10677 20768
rect 10635 20719 10677 20728
rect 10636 20634 10676 20719
rect 10732 20180 10772 20896
rect 11020 20768 11060 20779
rect 11020 20693 11060 20728
rect 11019 20684 11061 20693
rect 11019 20644 11020 20684
rect 11060 20644 11061 20684
rect 11019 20635 11061 20644
rect 10540 20140 10772 20180
rect 10828 20600 10868 20609
rect 10540 16484 10580 20140
rect 10828 20091 10868 20560
rect 11020 20180 11060 20189
rect 11116 20180 11156 21727
rect 11307 21608 11349 21617
rect 11307 21568 11308 21608
rect 11348 21568 11349 21608
rect 11307 21559 11349 21568
rect 11060 20140 11156 20180
rect 11020 20131 11060 20140
rect 10828 20042 10868 20051
rect 10827 19340 10869 19349
rect 10827 19300 10828 19340
rect 10868 19300 10869 19340
rect 10827 19291 10869 19300
rect 10684 19265 10724 19274
rect 10724 19225 10772 19256
rect 10684 19216 10772 19225
rect 10635 18752 10677 18761
rect 10635 18712 10636 18752
rect 10676 18712 10677 18752
rect 10732 18752 10772 19216
rect 10828 19172 10868 19291
rect 10828 19123 10868 19132
rect 10828 18752 10868 18761
rect 10732 18712 10828 18752
rect 10635 18703 10677 18712
rect 10828 18703 10868 18712
rect 10636 18584 10676 18703
rect 10636 18509 10676 18544
rect 11020 18584 11060 18593
rect 10635 18500 10677 18509
rect 11020 18500 11060 18544
rect 10635 18460 10636 18500
rect 10676 18460 10677 18500
rect 10635 18451 10677 18460
rect 10924 18460 11060 18500
rect 10924 18416 10964 18460
rect 10855 18376 10964 18416
rect 10855 18332 10895 18376
rect 10732 18292 10895 18332
rect 11019 18332 11061 18341
rect 11019 18292 11020 18332
rect 11060 18292 11061 18332
rect 10540 16444 10676 16484
rect 10348 16360 10484 16400
rect 10251 16316 10293 16325
rect 10251 16276 10252 16316
rect 10292 16276 10293 16316
rect 10251 16267 10293 16276
rect 10252 15569 10292 15654
rect 10251 15560 10293 15569
rect 10251 15520 10252 15560
rect 10292 15520 10293 15560
rect 10251 15511 10293 15520
rect 10348 15392 10388 16360
rect 10539 16316 10581 16325
rect 10539 16276 10540 16316
rect 10580 16276 10581 16316
rect 10539 16267 10581 16276
rect 10443 16232 10485 16241
rect 10443 16192 10444 16232
rect 10484 16192 10485 16232
rect 10443 16183 10485 16192
rect 10444 16098 10484 16183
rect 10540 15989 10580 16267
rect 10539 15980 10581 15989
rect 10539 15940 10540 15980
rect 10580 15940 10581 15980
rect 10539 15931 10581 15940
rect 10443 15896 10485 15905
rect 10443 15856 10444 15896
rect 10484 15856 10485 15896
rect 10443 15847 10485 15856
rect 10444 15569 10484 15847
rect 10443 15560 10485 15569
rect 10443 15520 10444 15560
rect 10484 15520 10485 15560
rect 10443 15511 10485 15520
rect 10252 15352 10388 15392
rect 9963 14720 10005 14729
rect 9963 14680 9964 14720
rect 10004 14680 10005 14720
rect 9963 14671 10005 14680
rect 10155 14720 10197 14729
rect 10155 14680 10156 14720
rect 10196 14680 10197 14720
rect 10155 14671 10197 14680
rect 9676 14552 9716 14561
rect 9676 14393 9716 14512
rect 9675 14384 9717 14393
rect 9675 14344 9676 14384
rect 9716 14344 9717 14384
rect 9675 14335 9717 14344
rect 9579 14216 9621 14225
rect 9579 14176 9580 14216
rect 9620 14176 9621 14216
rect 9579 14167 9621 14176
rect 9867 14216 9909 14225
rect 9867 14176 9868 14216
rect 9908 14176 9909 14216
rect 9867 14167 9909 14176
rect 9484 14048 9524 14057
rect 9484 13460 9524 14008
rect 9579 14048 9621 14057
rect 9579 14008 9580 14048
rect 9620 14008 9621 14048
rect 9579 13999 9621 14008
rect 9580 13914 9620 13999
rect 9868 13796 9908 14167
rect 9964 14048 10004 14671
rect 9964 13999 10004 14008
rect 10059 14048 10101 14057
rect 10059 14008 10060 14048
rect 10100 14008 10196 14048
rect 10059 13999 10101 14008
rect 10060 13914 10100 13999
rect 9868 13756 10004 13796
rect 9580 13460 9620 13469
rect 9484 13420 9580 13460
rect 9580 13411 9620 13420
rect 9771 13376 9813 13385
rect 9388 13336 9524 13376
rect 9388 13208 9428 13219
rect 9388 13133 9428 13168
rect 9387 13124 9429 13133
rect 9387 13084 9388 13124
rect 9428 13084 9429 13124
rect 9387 13075 9429 13084
rect 9388 12881 9428 13075
rect 9387 12872 9429 12881
rect 9387 12832 9388 12872
rect 9428 12832 9429 12872
rect 9387 12823 9429 12832
rect 9484 12704 9524 13336
rect 9771 13336 9772 13376
rect 9812 13336 9813 13376
rect 9771 13327 9813 13336
rect 9772 12881 9812 13327
rect 9867 13208 9909 13217
rect 9867 13168 9868 13208
rect 9908 13168 9909 13208
rect 9867 13159 9909 13168
rect 9868 13074 9908 13159
rect 9771 12872 9813 12881
rect 9771 12832 9772 12872
rect 9812 12832 9813 12872
rect 9771 12823 9813 12832
rect 9292 12664 9428 12704
rect 9484 12664 9716 12704
rect 9292 12536 9332 12547
rect 9292 12461 9332 12496
rect 9291 12452 9333 12461
rect 9291 12412 9292 12452
rect 9332 12412 9333 12452
rect 9291 12403 9333 12412
rect 9388 12377 9428 12664
rect 9483 12536 9525 12545
rect 9483 12496 9484 12536
rect 9524 12496 9525 12536
rect 9483 12487 9525 12496
rect 9387 12368 9429 12377
rect 9387 12328 9388 12368
rect 9428 12328 9429 12368
rect 9387 12319 9429 12328
rect 9484 12368 9524 12487
rect 9484 12319 9524 12328
rect 9291 12284 9333 12293
rect 9291 12244 9292 12284
rect 9332 12244 9333 12284
rect 9291 12235 9333 12244
rect 9292 10436 9332 12235
rect 9388 11705 9428 12319
rect 9387 11696 9429 11705
rect 9387 11656 9388 11696
rect 9428 11656 9429 11696
rect 9387 11647 9429 11656
rect 9579 11696 9621 11705
rect 9579 11656 9580 11696
rect 9620 11656 9621 11696
rect 9579 11647 9621 11656
rect 9580 11562 9620 11647
rect 9676 11537 9716 12664
rect 9772 12620 9812 12823
rect 9772 12571 9812 12580
rect 9868 12536 9908 12545
rect 9868 12209 9908 12496
rect 9867 12200 9909 12209
rect 9867 12160 9868 12200
rect 9908 12160 9909 12200
rect 9867 12151 9909 12160
rect 9771 11948 9813 11957
rect 9771 11908 9772 11948
rect 9812 11908 9813 11948
rect 9771 11899 9813 11908
rect 9675 11528 9717 11537
rect 9675 11488 9676 11528
rect 9716 11488 9717 11528
rect 9675 11479 9717 11488
rect 9387 11276 9429 11285
rect 9387 11236 9388 11276
rect 9428 11236 9429 11276
rect 9387 11227 9429 11236
rect 9388 11024 9428 11227
rect 9484 11108 9524 11117
rect 9676 11108 9716 11479
rect 9524 11068 9716 11108
rect 9484 11059 9524 11068
rect 9388 10604 9428 10984
rect 9772 10856 9812 11899
rect 9868 11873 9908 12151
rect 9867 11864 9909 11873
rect 9867 11824 9868 11864
rect 9908 11824 9909 11864
rect 9867 11815 9909 11824
rect 9964 11780 10004 13756
rect 10156 12788 10196 14008
rect 10252 13133 10292 15352
rect 10347 14720 10389 14729
rect 10347 14680 10348 14720
rect 10388 14680 10389 14720
rect 10347 14671 10389 14680
rect 10348 14586 10388 14671
rect 10444 14468 10484 15511
rect 10348 14428 10484 14468
rect 10251 13124 10293 13133
rect 10251 13084 10252 13124
rect 10292 13084 10293 13124
rect 10251 13075 10293 13084
rect 10156 12748 10292 12788
rect 10059 12536 10101 12545
rect 10059 12496 10060 12536
rect 10100 12527 10196 12536
rect 10100 12496 10156 12527
rect 10059 12487 10101 12496
rect 10156 12478 10196 12487
rect 10252 12368 10292 12748
rect 10348 12545 10388 14428
rect 10540 14048 10580 14059
rect 10636 14057 10676 16444
rect 10732 14645 10772 18292
rect 11019 18283 11061 18292
rect 10923 18248 10965 18257
rect 10923 18208 10924 18248
rect 10964 18208 10965 18248
rect 10923 18199 10965 18208
rect 10828 17744 10868 17753
rect 10828 17249 10868 17704
rect 10924 17744 10964 18199
rect 10924 17695 10964 17704
rect 10827 17240 10869 17249
rect 10827 17200 10828 17240
rect 10868 17200 10869 17240
rect 10827 17191 10869 17200
rect 11020 16400 11060 18283
rect 11116 16661 11156 20140
rect 11211 20180 11253 20189
rect 11211 20140 11212 20180
rect 11252 20140 11253 20180
rect 11211 20131 11253 20140
rect 11115 16652 11157 16661
rect 11115 16612 11116 16652
rect 11156 16612 11157 16652
rect 11115 16603 11157 16612
rect 10828 16360 11060 16400
rect 10828 14897 10868 16360
rect 11115 16316 11157 16325
rect 11115 16276 11116 16316
rect 11156 16276 11157 16316
rect 11115 16267 11157 16276
rect 11019 16232 11061 16241
rect 11019 16192 11020 16232
rect 11060 16192 11061 16232
rect 11019 16183 11061 16192
rect 11020 16098 11060 16183
rect 11116 15905 11156 16267
rect 11115 15896 11157 15905
rect 11115 15856 11116 15896
rect 11156 15856 11157 15896
rect 11115 15847 11157 15856
rect 11212 15653 11252 20131
rect 11308 18341 11348 21559
rect 11403 20516 11445 20525
rect 11403 20476 11404 20516
rect 11444 20476 11445 20516
rect 11403 20467 11445 20476
rect 11404 18929 11444 20467
rect 11596 19433 11636 22324
rect 11884 22280 11924 22651
rect 11979 22616 12021 22625
rect 11979 22576 11980 22616
rect 12020 22576 12021 22616
rect 11979 22567 12021 22576
rect 11980 22364 12020 22567
rect 11980 22315 12020 22324
rect 11884 22231 11924 22240
rect 12075 22280 12117 22289
rect 12075 22240 12076 22280
rect 12116 22240 12117 22280
rect 12075 22231 12117 22240
rect 12268 22280 12308 22289
rect 12460 22280 12500 23239
rect 12308 22240 12500 22280
rect 12268 22231 12308 22240
rect 11691 22196 11733 22205
rect 11691 22156 11692 22196
rect 11732 22156 11733 22196
rect 11691 22147 11733 22156
rect 11595 19424 11637 19433
rect 11595 19384 11596 19424
rect 11636 19384 11637 19424
rect 11595 19375 11637 19384
rect 11596 19256 11636 19265
rect 11403 18920 11445 18929
rect 11403 18880 11404 18920
rect 11444 18880 11445 18920
rect 11403 18871 11445 18880
rect 11307 18332 11349 18341
rect 11307 18292 11308 18332
rect 11348 18292 11349 18332
rect 11307 18283 11349 18292
rect 11307 18080 11349 18089
rect 11307 18040 11308 18080
rect 11348 18040 11349 18080
rect 11307 18031 11349 18040
rect 11308 17828 11348 18031
rect 11308 17779 11348 17788
rect 11404 17828 11444 18871
rect 11596 18845 11636 19216
rect 11595 18836 11637 18845
rect 11595 18796 11596 18836
rect 11636 18796 11637 18836
rect 11595 18787 11637 18796
rect 11404 17779 11444 17788
rect 11596 17669 11636 18787
rect 11595 17660 11637 17669
rect 11595 17620 11596 17660
rect 11636 17620 11637 17660
rect 11595 17611 11637 17620
rect 11692 17240 11732 22147
rect 12076 22146 12116 22231
rect 11787 22028 11829 22037
rect 11787 21988 11788 22028
rect 11828 21988 11829 22028
rect 11787 21979 11829 21988
rect 11788 21608 11828 21979
rect 11980 21692 12020 21701
rect 12020 21652 12308 21692
rect 11980 21643 12020 21652
rect 11788 21559 11828 21568
rect 12268 21608 12308 21652
rect 12268 21559 12308 21568
rect 12364 21608 12404 21619
rect 12364 21533 12404 21568
rect 12075 21524 12117 21533
rect 12075 21484 12076 21524
rect 12116 21484 12117 21524
rect 12075 21475 12117 21484
rect 12363 21524 12405 21533
rect 12363 21484 12364 21524
rect 12404 21484 12405 21524
rect 12363 21475 12405 21484
rect 11787 21440 11829 21449
rect 11787 21400 11788 21440
rect 11828 21400 11829 21440
rect 11787 21391 11829 21400
rect 11596 17200 11732 17240
rect 11403 16568 11445 16577
rect 11403 16528 11404 16568
rect 11444 16528 11445 16568
rect 11403 16519 11445 16528
rect 11404 16157 11444 16519
rect 11596 16400 11636 17200
rect 11692 17072 11732 17081
rect 11692 16661 11732 17032
rect 11691 16652 11733 16661
rect 11691 16612 11692 16652
rect 11732 16612 11733 16652
rect 11691 16603 11733 16612
rect 11788 16577 11828 21391
rect 11979 21272 12021 21281
rect 11979 21232 11980 21272
rect 12020 21232 12021 21272
rect 11979 21223 12021 21232
rect 11883 19424 11925 19433
rect 11883 19384 11884 19424
rect 11924 19384 11925 19424
rect 11883 19375 11925 19384
rect 11884 17744 11924 19375
rect 11787 16568 11829 16577
rect 11787 16528 11788 16568
rect 11828 16528 11829 16568
rect 11787 16519 11829 16528
rect 11596 16360 11828 16400
rect 11548 16274 11625 16316
rect 11588 16234 11625 16274
rect 11548 16232 11625 16234
rect 11548 16225 11636 16232
rect 11585 16192 11636 16225
rect 11403 16148 11445 16157
rect 11403 16108 11404 16148
rect 11444 16108 11445 16148
rect 11403 16099 11445 16108
rect 11596 15728 11636 16192
rect 11691 16064 11733 16073
rect 11691 16024 11692 16064
rect 11732 16024 11733 16064
rect 11691 16015 11733 16024
rect 11692 15930 11732 16015
rect 11692 15728 11732 15737
rect 11596 15688 11692 15728
rect 11692 15679 11732 15688
rect 10923 15644 10965 15653
rect 10923 15604 10924 15644
rect 10964 15604 10965 15644
rect 10923 15595 10965 15604
rect 11211 15644 11253 15653
rect 11211 15604 11212 15644
rect 11252 15604 11253 15644
rect 11211 15595 11253 15604
rect 10827 14888 10869 14897
rect 10827 14848 10828 14888
rect 10868 14848 10869 14888
rect 10827 14839 10869 14848
rect 10731 14636 10773 14645
rect 10731 14596 10732 14636
rect 10772 14596 10773 14636
rect 10731 14587 10773 14596
rect 10540 13973 10580 14008
rect 10635 14048 10677 14057
rect 10635 14008 10636 14048
rect 10676 14008 10677 14048
rect 10635 13999 10677 14008
rect 10539 13964 10581 13973
rect 10539 13924 10540 13964
rect 10580 13924 10581 13964
rect 10539 13915 10581 13924
rect 10827 13040 10869 13049
rect 10827 13000 10828 13040
rect 10868 13000 10869 13040
rect 10827 12991 10869 13000
rect 10347 12536 10389 12545
rect 10347 12496 10348 12536
rect 10388 12496 10389 12536
rect 10347 12487 10389 12496
rect 10444 12536 10484 12545
rect 10636 12536 10676 12545
rect 10484 12496 10580 12536
rect 10444 12487 10484 12496
rect 10252 12328 10388 12368
rect 10155 12284 10197 12293
rect 10155 12244 10156 12284
rect 10196 12244 10197 12284
rect 10155 12235 10197 12244
rect 9964 11740 10100 11780
rect 9868 11696 9908 11705
rect 9868 11612 9908 11656
rect 9964 11612 10004 11623
rect 9868 11572 9909 11612
rect 9869 11528 9909 11572
rect 9964 11537 10004 11572
rect 9868 11488 9909 11528
rect 9963 11528 10005 11537
rect 9963 11488 9964 11528
rect 10004 11488 10005 11528
rect 9868 11369 9908 11488
rect 9963 11479 10005 11488
rect 9867 11360 9909 11369
rect 10060 11360 10100 11740
rect 9867 11320 9868 11360
rect 9908 11320 9909 11360
rect 9867 11311 9909 11320
rect 9964 11320 10100 11360
rect 9772 10807 9812 10816
rect 9675 10688 9717 10697
rect 9675 10648 9676 10688
rect 9716 10648 9717 10688
rect 9675 10639 9717 10648
rect 9388 10564 9524 10604
rect 9292 10396 9428 10436
rect 8908 9556 9044 9596
rect 9100 9976 9236 10016
rect 9388 10184 9428 10396
rect 8908 9512 8948 9556
rect 8908 9463 8948 9472
rect 9003 9428 9045 9437
rect 9003 9388 9004 9428
rect 9044 9388 9045 9428
rect 9003 9379 9045 9388
rect 8907 9092 8949 9101
rect 8812 9052 8908 9092
rect 8948 9052 8949 9092
rect 8715 9008 8757 9017
rect 8715 8968 8716 9008
rect 8756 8968 8757 9008
rect 8715 8959 8757 8968
rect 8428 8800 8564 8840
rect 8428 8672 8468 8681
rect 8428 8177 8468 8632
rect 8427 8168 8469 8177
rect 8427 8128 8428 8168
rect 8468 8128 8469 8168
rect 8427 8119 8469 8128
rect 8139 7412 8181 7421
rect 8139 7372 8140 7412
rect 8180 7372 8181 7412
rect 8139 7363 8181 7372
rect 8140 6749 8180 7363
rect 8427 6992 8469 7001
rect 8427 6952 8428 6992
rect 8468 6952 8469 6992
rect 8427 6943 8469 6952
rect 8139 6740 8181 6749
rect 8139 6700 8140 6740
rect 8180 6700 8181 6740
rect 8139 6691 8181 6700
rect 8331 6740 8373 6749
rect 8331 6700 8332 6740
rect 8372 6700 8373 6740
rect 8331 6691 8373 6700
rect 8428 6714 8468 6943
rect 8041 5608 8084 5648
rect 8140 5648 8180 6691
rect 8235 6656 8277 6665
rect 8235 6616 8236 6656
rect 8276 6616 8277 6656
rect 8235 6607 8277 6616
rect 8236 6488 8276 6607
rect 8332 6497 8372 6691
rect 8428 6665 8468 6674
rect 8236 6439 8276 6448
rect 8331 6488 8373 6497
rect 8331 6448 8332 6488
rect 8372 6448 8373 6488
rect 8331 6439 8373 6448
rect 8524 6320 8564 8800
rect 8812 8756 8852 9052
rect 8907 9043 8949 9052
rect 9004 9008 9044 9379
rect 9004 8968 9055 9008
rect 8812 8716 8940 8756
rect 8900 8686 8940 8716
rect 9015 8686 9055 8968
rect 8716 8672 8756 8681
rect 8900 8672 8948 8686
rect 8716 8597 8756 8632
rect 8811 8657 8853 8666
rect 8811 8611 8812 8657
rect 8852 8611 8853 8657
rect 8900 8646 8908 8672
rect 8908 8623 8948 8632
rect 9004 8672 9055 8686
rect 9044 8646 9055 8672
rect 9100 8686 9140 9976
rect 9388 9521 9428 10144
rect 9195 9512 9237 9521
rect 9195 9472 9196 9512
rect 9236 9472 9237 9512
rect 9195 9463 9237 9472
rect 9387 9512 9429 9521
rect 9387 9472 9388 9512
rect 9428 9472 9429 9512
rect 9387 9463 9429 9472
rect 9196 9378 9236 9463
rect 9291 9008 9333 9017
rect 9291 8968 9292 9008
rect 9332 8968 9333 9008
rect 9291 8959 9333 8968
rect 9100 8646 9236 8686
rect 9004 8623 9044 8632
rect 8811 8608 8853 8611
rect 8715 8588 8757 8597
rect 8715 8548 8716 8588
rect 8756 8548 8757 8588
rect 8715 8539 8757 8548
rect 8716 8084 8756 8539
rect 8812 8522 8852 8608
rect 9196 8504 9236 8646
rect 9292 8672 9332 8959
rect 9484 8840 9524 10564
rect 9580 10016 9620 10025
rect 9580 9017 9620 9976
rect 9676 9353 9716 10639
rect 9964 10352 10004 11320
rect 10059 10772 10101 10781
rect 10059 10732 10060 10772
rect 10100 10732 10101 10772
rect 10059 10723 10101 10732
rect 10060 10638 10100 10723
rect 9964 10303 10004 10312
rect 9867 10268 9909 10277
rect 9867 10228 9868 10268
rect 9908 10228 9909 10268
rect 9867 10219 9909 10228
rect 10059 10268 10101 10277
rect 10059 10228 10060 10268
rect 10100 10228 10101 10268
rect 10059 10219 10101 10228
rect 9771 10184 9813 10193
rect 9771 10144 9772 10184
rect 9812 10144 9813 10184
rect 9771 10135 9813 10144
rect 9772 10050 9812 10135
rect 9868 10134 9908 10219
rect 9963 10184 10005 10193
rect 9963 10144 9964 10184
rect 10004 10144 10005 10184
rect 9963 10135 10005 10144
rect 9675 9344 9717 9353
rect 9675 9304 9676 9344
rect 9716 9304 9717 9344
rect 9675 9295 9717 9304
rect 9579 9008 9621 9017
rect 9579 8968 9580 9008
rect 9620 8968 9621 9008
rect 9579 8959 9621 8968
rect 9484 8800 9716 8840
rect 9292 8623 9332 8632
rect 9388 8672 9428 8681
rect 9388 8588 9428 8632
rect 9388 8548 9620 8588
rect 9196 8464 9524 8504
rect 8041 5564 8081 5608
rect 8140 5573 8180 5608
rect 8236 6280 8564 6320
rect 8620 8044 8756 8084
rect 8139 5564 8181 5573
rect 8041 5524 8084 5564
rect 7659 5396 7701 5405
rect 7659 5356 7660 5396
rect 7700 5356 7701 5396
rect 7659 5347 7701 5356
rect 7564 4976 7604 4987
rect 7564 4901 7604 4936
rect 7948 4976 7988 4985
rect 7563 4892 7605 4901
rect 7563 4852 7564 4892
rect 7604 4852 7605 4892
rect 7563 4843 7605 4852
rect 7948 4733 7988 4936
rect 7756 4724 7796 4733
rect 7659 3968 7701 3977
rect 7659 3928 7660 3968
rect 7700 3928 7701 3968
rect 7659 3919 7701 3928
rect 7660 3725 7700 3919
rect 7659 3716 7701 3725
rect 7659 3676 7660 3716
rect 7700 3676 7701 3716
rect 7659 3667 7701 3676
rect 7756 3473 7796 4684
rect 7947 4724 7989 4733
rect 7947 4684 7948 4724
rect 7988 4684 7989 4724
rect 7947 4675 7989 4684
rect 7851 4220 7893 4229
rect 7851 4180 7852 4220
rect 7892 4180 7893 4220
rect 7851 4171 7893 4180
rect 7852 4136 7892 4171
rect 7852 4085 7892 4096
rect 7947 3632 7989 3641
rect 7947 3592 7948 3632
rect 7988 3592 7989 3632
rect 7947 3583 7989 3592
rect 7468 3221 7508 3424
rect 7755 3464 7797 3473
rect 7755 3424 7756 3464
rect 7796 3424 7797 3464
rect 7755 3415 7797 3424
rect 7948 3464 7988 3583
rect 7948 3415 7988 3424
rect 7467 3212 7509 3221
rect 7467 3172 7468 3212
rect 7508 3172 7509 3212
rect 7467 3163 7509 3172
rect 7371 3128 7413 3137
rect 7371 3088 7372 3128
rect 7412 3088 7413 3128
rect 7371 3079 7413 3088
rect 7371 2960 7413 2969
rect 7371 2920 7372 2960
rect 7412 2920 7413 2960
rect 7371 2911 7413 2920
rect 7372 2708 7412 2911
rect 7372 2659 7412 2668
rect 7755 2708 7797 2717
rect 7755 2668 7756 2708
rect 7796 2668 7797 2708
rect 7755 2659 7797 2668
rect 7756 2624 7796 2659
rect 7756 2573 7796 2584
rect 8044 2549 8084 5524
rect 8139 5524 8140 5564
rect 8180 5524 8181 5564
rect 8139 5515 8181 5524
rect 8139 5228 8181 5237
rect 8139 5188 8140 5228
rect 8180 5188 8181 5228
rect 8139 5179 8181 5188
rect 8140 3977 8180 5179
rect 8139 3968 8181 3977
rect 8139 3928 8140 3968
rect 8180 3928 8181 3968
rect 8139 3919 8181 3928
rect 8043 2540 8085 2549
rect 8043 2500 8044 2540
rect 8084 2500 8085 2540
rect 8043 2491 8085 2500
rect 7467 2456 7509 2465
rect 7467 2416 7468 2456
rect 7508 2416 7509 2456
rect 7467 2407 7509 2416
rect 7564 2456 7604 2465
rect 7275 2288 7317 2297
rect 7275 2248 7276 2288
rect 7316 2248 7317 2288
rect 7275 2239 7317 2248
rect 7084 2164 7220 2204
rect 7180 1952 7220 2164
rect 6892 1898 7124 1938
rect 7180 1903 7220 1912
rect 7084 1784 7124 1898
rect 7372 1784 7412 1793
rect 7084 1744 7372 1784
rect 7372 1735 7412 1744
rect 6411 1280 6453 1289
rect 6411 1240 6412 1280
rect 6452 1240 6453 1280
rect 6411 1231 6453 1240
rect 6795 1280 6837 1289
rect 6795 1240 6796 1280
rect 6836 1240 6837 1280
rect 6795 1231 6837 1240
rect 6987 1280 7029 1289
rect 6987 1240 6988 1280
rect 7028 1240 7029 1280
rect 6987 1231 7029 1240
rect 7179 1280 7221 1289
rect 7179 1240 7180 1280
rect 7220 1240 7221 1280
rect 7179 1231 7221 1240
rect 6412 80 6452 1231
rect 6603 356 6645 365
rect 6603 316 6604 356
rect 6644 316 6645 356
rect 6603 307 6645 316
rect 6604 80 6644 307
rect 6796 80 6836 1231
rect 6988 80 7028 1231
rect 7180 80 7220 1231
rect 7372 1112 7412 1121
rect 7276 1072 7372 1112
rect 7276 701 7316 1072
rect 7372 1063 7412 1072
rect 7371 944 7413 953
rect 7371 904 7372 944
rect 7412 904 7413 944
rect 7371 895 7413 904
rect 7275 692 7317 701
rect 7275 652 7276 692
rect 7316 652 7317 692
rect 7275 643 7317 652
rect 7276 281 7316 643
rect 7275 272 7317 281
rect 7275 232 7276 272
rect 7316 232 7317 272
rect 7275 223 7317 232
rect 7372 80 7412 895
rect 7468 869 7508 2407
rect 7564 2288 7604 2416
rect 7564 2248 7892 2288
rect 7563 2120 7605 2129
rect 7563 2080 7564 2120
rect 7604 2080 7605 2120
rect 7563 2071 7605 2080
rect 7564 1952 7604 2071
rect 7564 1903 7604 1912
rect 7659 1952 7701 1961
rect 7659 1912 7660 1952
rect 7700 1912 7701 1952
rect 7659 1903 7701 1912
rect 7660 1784 7700 1903
rect 7564 1744 7700 1784
rect 7564 1280 7604 1744
rect 7852 1532 7892 2248
rect 7564 1231 7604 1240
rect 7660 1492 7892 1532
rect 7563 1112 7605 1121
rect 7563 1072 7564 1112
rect 7604 1072 7605 1112
rect 7563 1063 7605 1072
rect 7467 860 7509 869
rect 7467 820 7468 860
rect 7508 820 7509 860
rect 7467 811 7509 820
rect 7564 80 7604 1063
rect 7660 617 7700 1492
rect 7755 1280 7797 1289
rect 7755 1240 7756 1280
rect 7796 1240 7797 1280
rect 7755 1231 7797 1240
rect 8139 1280 8181 1289
rect 8139 1240 8140 1280
rect 8180 1240 8181 1280
rect 8139 1231 8181 1240
rect 7756 1112 7796 1231
rect 7796 1072 7892 1112
rect 7756 1063 7796 1072
rect 7755 944 7797 953
rect 7755 904 7756 944
rect 7796 904 7797 944
rect 7852 944 7892 1072
rect 8043 944 8085 953
rect 7852 904 8044 944
rect 8084 904 8085 944
rect 7755 895 7797 904
rect 8043 895 8085 904
rect 7659 608 7701 617
rect 7659 568 7660 608
rect 7700 568 7701 608
rect 7659 559 7701 568
rect 7756 80 7796 895
rect 7947 692 7989 701
rect 7947 652 7948 692
rect 7988 652 7989 692
rect 7947 643 7989 652
rect 7948 80 7988 643
rect 8140 80 8180 1231
rect 8236 953 8276 6280
rect 8620 6236 8660 8044
rect 8812 8000 8852 8009
rect 8716 7960 8812 8000
rect 8716 7421 8756 7960
rect 8812 7589 8852 7960
rect 9099 8000 9141 8009
rect 9099 7960 9100 8000
rect 9140 7960 9141 8000
rect 9099 7951 9141 7960
rect 9196 8000 9236 8011
rect 9003 7748 9045 7757
rect 9003 7708 9004 7748
rect 9044 7708 9045 7748
rect 9003 7699 9045 7708
rect 9004 7614 9044 7699
rect 8811 7580 8853 7589
rect 8811 7540 8812 7580
rect 8852 7540 8853 7580
rect 8811 7531 8853 7540
rect 8715 7412 8757 7421
rect 8715 7372 8716 7412
rect 8756 7372 8757 7412
rect 8715 7363 8757 7372
rect 8715 7160 8757 7169
rect 8812 7160 8852 7169
rect 8715 7120 8716 7160
rect 8756 7120 8812 7160
rect 8715 7111 8757 7120
rect 8812 7111 8852 7120
rect 9004 7160 9044 7169
rect 9004 7001 9044 7120
rect 9100 7160 9140 7951
rect 9196 7925 9236 7960
rect 9484 7925 9524 8464
rect 9195 7916 9237 7925
rect 9195 7876 9196 7916
rect 9236 7876 9237 7916
rect 9195 7867 9237 7876
rect 9483 7916 9525 7925
rect 9483 7876 9484 7916
rect 9524 7876 9525 7916
rect 9483 7867 9525 7876
rect 9580 7328 9620 8548
rect 9676 8261 9716 8800
rect 9772 8672 9812 8681
rect 9675 8252 9717 8261
rect 9675 8212 9676 8252
rect 9716 8212 9717 8252
rect 9675 8203 9717 8212
rect 9772 8000 9812 8632
rect 9867 8672 9909 8681
rect 9867 8632 9868 8672
rect 9908 8632 9909 8672
rect 9867 8623 9909 8632
rect 9868 8538 9908 8623
rect 9964 8177 10004 10135
rect 10060 10134 10100 10219
rect 10156 10184 10196 12235
rect 10252 11864 10292 11873
rect 10252 11192 10292 11824
rect 10348 11369 10388 12328
rect 10443 12284 10485 12293
rect 10443 12244 10444 12284
rect 10484 12244 10485 12284
rect 10443 12235 10485 12244
rect 10444 12150 10484 12235
rect 10443 11864 10485 11873
rect 10443 11824 10444 11864
rect 10484 11824 10485 11864
rect 10443 11815 10485 11824
rect 10444 11696 10484 11815
rect 10444 11647 10484 11656
rect 10347 11360 10389 11369
rect 10347 11320 10348 11360
rect 10388 11320 10389 11360
rect 10347 11311 10389 11320
rect 10540 11201 10580 12496
rect 10636 12041 10676 12496
rect 10732 12536 10772 12545
rect 10635 12032 10677 12041
rect 10635 11992 10636 12032
rect 10676 11992 10677 12032
rect 10635 11983 10677 11992
rect 10732 11957 10772 12496
rect 10731 11948 10773 11957
rect 10731 11908 10732 11948
rect 10772 11908 10773 11948
rect 10731 11899 10773 11908
rect 10731 11780 10773 11789
rect 10731 11740 10732 11780
rect 10772 11740 10773 11780
rect 10731 11731 10773 11740
rect 10539 11192 10581 11201
rect 10252 11152 10388 11192
rect 10252 11024 10292 11033
rect 10252 10613 10292 10984
rect 10251 10604 10293 10613
rect 10251 10564 10252 10604
rect 10292 10564 10293 10604
rect 10348 10604 10388 11152
rect 10539 11152 10540 11192
rect 10580 11152 10581 11192
rect 10539 11143 10581 11152
rect 10348 10564 10580 10604
rect 10251 10555 10293 10564
rect 10252 10361 10292 10555
rect 10347 10436 10389 10445
rect 10347 10396 10348 10436
rect 10388 10396 10389 10436
rect 10347 10387 10389 10396
rect 10251 10352 10293 10361
rect 10251 10312 10252 10352
rect 10292 10312 10293 10352
rect 10251 10303 10293 10312
rect 10156 10135 10196 10144
rect 10251 10184 10293 10193
rect 10251 10144 10252 10184
rect 10292 10144 10293 10184
rect 10251 10135 10293 10144
rect 10348 10184 10388 10387
rect 10252 8513 10292 10135
rect 10348 9941 10388 10144
rect 10347 9932 10389 9941
rect 10347 9892 10348 9932
rect 10388 9892 10389 9932
rect 10347 9883 10389 9892
rect 10443 9512 10485 9521
rect 10443 9472 10444 9512
rect 10484 9472 10485 9512
rect 10443 9463 10485 9472
rect 10347 8840 10389 8849
rect 10347 8800 10348 8840
rect 10388 8800 10389 8840
rect 10347 8791 10389 8800
rect 10348 8672 10388 8791
rect 10251 8504 10293 8513
rect 10251 8464 10252 8504
rect 10292 8464 10293 8504
rect 10251 8455 10293 8464
rect 9963 8168 10005 8177
rect 9963 8128 9964 8168
rect 10004 8128 10005 8168
rect 9963 8119 10005 8128
rect 9772 7960 10100 8000
rect 9771 7748 9813 7757
rect 9771 7708 9772 7748
rect 9812 7708 9813 7748
rect 9771 7699 9813 7708
rect 9388 7288 9620 7328
rect 8715 6992 8757 7001
rect 8715 6952 8716 6992
rect 8756 6952 8757 6992
rect 8715 6943 8757 6952
rect 9003 6992 9045 7001
rect 9003 6952 9004 6992
rect 9044 6952 9045 6992
rect 9003 6943 9045 6952
rect 8716 6497 8756 6943
rect 9100 6917 9140 7120
rect 9292 7160 9332 7171
rect 9292 7085 9332 7120
rect 9291 7076 9333 7085
rect 9291 7036 9292 7076
rect 9332 7036 9333 7076
rect 9291 7027 9333 7036
rect 9388 7001 9428 7288
rect 9675 7244 9717 7253
rect 9675 7204 9676 7244
rect 9716 7204 9717 7244
rect 9675 7195 9717 7204
rect 9484 7160 9524 7169
rect 9196 6992 9236 7001
rect 9099 6908 9141 6917
rect 9099 6868 9100 6908
rect 9140 6868 9141 6908
rect 9099 6859 9141 6868
rect 9003 6824 9045 6833
rect 9003 6784 9004 6824
rect 9044 6784 9045 6824
rect 9003 6775 9045 6784
rect 8811 6572 8853 6581
rect 8811 6532 8812 6572
rect 8852 6532 8853 6572
rect 8811 6523 8853 6532
rect 8715 6488 8757 6497
rect 8715 6448 8716 6488
rect 8756 6448 8757 6488
rect 8715 6439 8757 6448
rect 8716 6354 8756 6439
rect 8428 6196 8660 6236
rect 8331 6152 8373 6161
rect 8331 6112 8332 6152
rect 8372 6112 8373 6152
rect 8331 6103 8373 6112
rect 8332 5993 8372 6103
rect 8331 5984 8373 5993
rect 8331 5944 8332 5984
rect 8372 5944 8373 5984
rect 8331 5935 8373 5944
rect 8332 5480 8372 5489
rect 8332 5237 8372 5440
rect 8331 5228 8373 5237
rect 8331 5188 8332 5228
rect 8372 5188 8373 5228
rect 8331 5179 8373 5188
rect 8428 4649 8468 6196
rect 8715 6152 8757 6161
rect 8812 6152 8852 6523
rect 9004 6488 9044 6775
rect 9099 6572 9141 6581
rect 9099 6532 9100 6572
rect 9140 6532 9141 6572
rect 9099 6523 9141 6532
rect 9004 6439 9044 6448
rect 9100 6438 9140 6523
rect 8715 6112 8716 6152
rect 8756 6112 8852 6152
rect 8715 6103 8757 6112
rect 8800 6028 8852 6112
rect 8619 5900 8661 5909
rect 8619 5860 8620 5900
rect 8660 5860 8661 5900
rect 8619 5851 8661 5860
rect 8811 5900 8853 5909
rect 8811 5860 8812 5900
rect 8852 5860 8853 5900
rect 8811 5851 8853 5860
rect 8620 5648 8660 5851
rect 8620 5599 8660 5608
rect 8523 5564 8565 5573
rect 8523 5524 8524 5564
rect 8564 5524 8565 5564
rect 8523 5515 8565 5524
rect 8427 4640 8469 4649
rect 8427 4600 8428 4640
rect 8468 4600 8469 4640
rect 8427 4591 8469 4600
rect 8380 4145 8420 4154
rect 8420 4105 8468 4136
rect 8380 4096 8468 4105
rect 8428 3450 8468 4096
rect 8524 4052 8564 5515
rect 8812 4985 8852 5851
rect 8908 5648 8948 5657
rect 8811 4976 8853 4985
rect 8811 4936 8812 4976
rect 8852 4936 8853 4976
rect 8811 4927 8853 4936
rect 8811 4808 8853 4817
rect 8811 4768 8812 4808
rect 8852 4768 8853 4808
rect 8811 4759 8853 4768
rect 8715 4388 8757 4397
rect 8715 4348 8716 4388
rect 8756 4348 8757 4388
rect 8715 4339 8757 4348
rect 8716 4229 8756 4339
rect 8715 4220 8757 4229
rect 8715 4180 8716 4220
rect 8756 4180 8757 4220
rect 8715 4171 8757 4180
rect 8812 4136 8852 4759
rect 8812 4087 8852 4096
rect 8524 4003 8564 4012
rect 8908 3968 8948 5608
rect 9003 5564 9045 5573
rect 9003 5524 9004 5564
rect 9044 5524 9045 5564
rect 9003 5515 9045 5524
rect 9004 5430 9044 5515
rect 9196 5228 9236 6952
rect 9387 6992 9429 7001
rect 9387 6952 9388 6992
rect 9428 6952 9429 6992
rect 9387 6943 9429 6952
rect 9484 6824 9524 7120
rect 9580 7160 9620 7171
rect 9580 7085 9620 7120
rect 9579 7076 9621 7085
rect 9579 7036 9580 7076
rect 9620 7036 9621 7076
rect 9579 7027 9621 7036
rect 9676 7076 9716 7195
rect 9772 7160 9812 7699
rect 9812 7120 9908 7160
rect 9772 7111 9812 7120
rect 9676 7027 9716 7036
rect 9388 6784 9524 6824
rect 9388 6698 9428 6784
rect 9291 6656 9333 6665
rect 9291 6616 9292 6656
rect 9332 6616 9333 6656
rect 9388 6649 9428 6658
rect 9580 6656 9620 7027
rect 9291 6607 9333 6616
rect 9484 6616 9620 6656
rect 9292 5900 9332 6607
rect 9484 6320 9524 6616
rect 9580 6488 9620 6497
rect 9868 6488 9908 7120
rect 10060 6740 10100 7960
rect 10155 7748 10197 7757
rect 10155 7708 10156 7748
rect 10196 7708 10197 7748
rect 10155 7699 10197 7708
rect 10156 7160 10196 7699
rect 10348 7253 10388 8632
rect 10444 8168 10484 9463
rect 10540 8597 10580 10564
rect 10636 9260 10676 9269
rect 10636 8765 10676 9220
rect 10635 8756 10677 8765
rect 10635 8716 10636 8756
rect 10676 8716 10677 8756
rect 10635 8707 10677 8716
rect 10539 8588 10581 8597
rect 10539 8548 10540 8588
rect 10580 8548 10581 8588
rect 10539 8539 10581 8548
rect 10444 8128 10580 8168
rect 10443 8000 10485 8009
rect 10443 7960 10444 8000
rect 10484 7960 10485 8000
rect 10443 7951 10485 7960
rect 10444 7866 10484 7951
rect 10347 7244 10389 7253
rect 10347 7204 10348 7244
rect 10388 7204 10389 7244
rect 10347 7195 10389 7204
rect 10156 7111 10196 7120
rect 10252 7160 10292 7169
rect 10252 6740 10292 7120
rect 10060 6700 10292 6740
rect 10347 6740 10389 6749
rect 10347 6700 10348 6740
rect 10388 6700 10389 6740
rect 9620 6448 9716 6488
rect 9580 6439 9620 6448
rect 9292 5851 9332 5860
rect 9388 6280 9524 6320
rect 9579 6320 9621 6329
rect 9579 6280 9580 6320
rect 9620 6280 9621 6320
rect 9388 5648 9428 6280
rect 9579 6271 9621 6280
rect 9580 6186 9620 6271
rect 9676 5816 9716 6448
rect 9868 6439 9908 6448
rect 10060 6488 10100 6499
rect 10060 6413 10100 6448
rect 10059 6404 10101 6413
rect 10059 6364 10060 6404
rect 10100 6364 10101 6404
rect 10059 6355 10101 6364
rect 10060 6236 10100 6245
rect 9676 5767 9716 5776
rect 9772 6196 10060 6236
rect 9484 5648 9524 5657
rect 9388 5608 9484 5648
rect 9484 5599 9524 5608
rect 9675 5648 9717 5657
rect 9675 5608 9676 5648
rect 9716 5608 9717 5648
rect 9675 5599 9717 5608
rect 9772 5648 9812 6196
rect 10060 6187 10100 6196
rect 10156 6068 10196 6700
rect 10347 6691 10389 6700
rect 10348 6572 10388 6691
rect 10252 6532 10388 6572
rect 10252 6487 10292 6532
rect 10444 6488 10484 6497
rect 10252 6438 10292 6447
rect 10348 6448 10444 6488
rect 10251 6320 10293 6329
rect 10251 6280 10252 6320
rect 10292 6280 10293 6320
rect 10251 6271 10293 6280
rect 9772 5599 9812 5608
rect 10060 6028 10196 6068
rect 9676 5514 9716 5599
rect 9100 5188 9236 5228
rect 9003 4724 9045 4733
rect 9003 4684 9004 4724
rect 9044 4684 9045 4724
rect 9003 4675 9045 4684
rect 8812 3928 8948 3968
rect 8812 3800 8852 3928
rect 8620 3760 8852 3800
rect 8907 3800 8949 3809
rect 8907 3760 8908 3800
rect 8948 3760 8949 3800
rect 8620 3632 8660 3760
rect 8907 3751 8949 3760
rect 8620 3583 8660 3592
rect 8812 3632 8852 3641
rect 8908 3632 8948 3751
rect 8852 3592 8948 3632
rect 8812 3583 8852 3592
rect 8428 1961 8468 3410
rect 9004 3464 9044 4675
rect 9100 4145 9140 5188
rect 9196 5069 9236 5100
rect 9195 5060 9237 5069
rect 9195 5020 9196 5060
rect 9236 5020 9237 5060
rect 9195 5011 9237 5020
rect 9196 4976 9236 5011
rect 9580 4976 9620 4985
rect 9099 4136 9141 4145
rect 9099 4096 9100 4136
rect 9140 4096 9141 4136
rect 9099 4087 9141 4096
rect 9004 3389 9044 3424
rect 9003 3380 9045 3389
rect 9003 3340 9004 3380
rect 9044 3340 9045 3380
rect 9003 3331 9045 3340
rect 9196 3212 9236 4936
rect 8908 3172 9236 3212
rect 9292 4936 9580 4976
rect 8715 2792 8757 2801
rect 8715 2752 8716 2792
rect 8756 2752 8757 2792
rect 8715 2743 8757 2752
rect 8427 1952 8469 1961
rect 8427 1912 8428 1952
rect 8468 1912 8469 1952
rect 8427 1903 8469 1912
rect 8331 1280 8373 1289
rect 8331 1240 8332 1280
rect 8372 1240 8373 1280
rect 8331 1231 8373 1240
rect 8523 1280 8565 1289
rect 8523 1240 8524 1280
rect 8564 1240 8565 1280
rect 8523 1231 8565 1240
rect 8235 944 8277 953
rect 8235 904 8236 944
rect 8276 904 8277 944
rect 8235 895 8277 904
rect 8332 80 8372 1231
rect 8524 80 8564 1231
rect 8716 80 8756 2743
rect 8811 2456 8853 2465
rect 8811 2416 8812 2456
rect 8852 2416 8853 2456
rect 8811 2407 8853 2416
rect 8812 1952 8852 2407
rect 8908 2129 8948 3172
rect 9196 2876 9236 2885
rect 9292 2876 9332 4936
rect 9580 4927 9620 4936
rect 9675 4976 9717 4985
rect 9675 4936 9676 4976
rect 9716 4936 9717 4976
rect 9675 4927 9717 4936
rect 9676 4842 9716 4927
rect 10060 4892 10100 6028
rect 10156 5648 10196 5657
rect 10252 5648 10292 6271
rect 10348 6077 10388 6448
rect 10444 6439 10484 6448
rect 10443 6320 10485 6329
rect 10443 6280 10444 6320
rect 10484 6280 10485 6320
rect 10443 6271 10485 6280
rect 10347 6068 10389 6077
rect 10347 6028 10348 6068
rect 10388 6028 10389 6068
rect 10347 6019 10389 6028
rect 10348 5825 10388 6019
rect 10347 5816 10389 5825
rect 10347 5776 10348 5816
rect 10388 5776 10389 5816
rect 10347 5767 10389 5776
rect 10196 5608 10292 5648
rect 10156 5599 10196 5608
rect 10155 4976 10197 4985
rect 10155 4936 10156 4976
rect 10196 4936 10197 4976
rect 10155 4927 10197 4936
rect 10060 4724 10100 4852
rect 10156 4842 10196 4927
rect 10251 4892 10293 4901
rect 10251 4852 10252 4892
rect 10292 4852 10293 4892
rect 10251 4843 10293 4852
rect 10060 4684 10196 4724
rect 10059 4220 10101 4229
rect 10059 4180 10060 4220
rect 10100 4180 10101 4220
rect 10059 4171 10101 4180
rect 10060 4136 10100 4171
rect 10060 4085 10100 4096
rect 10156 3968 10196 4684
rect 10252 4388 10292 4843
rect 10252 4339 10292 4348
rect 10347 4220 10389 4229
rect 10347 4180 10348 4220
rect 10388 4180 10389 4220
rect 10347 4171 10389 4180
rect 10060 3928 10196 3968
rect 9675 3464 9717 3473
rect 9675 3424 9676 3464
rect 9716 3424 9717 3464
rect 9675 3415 9717 3424
rect 9483 3212 9525 3221
rect 9483 3172 9484 3212
rect 9524 3172 9525 3212
rect 9483 3163 9525 3172
rect 9236 2836 9332 2876
rect 9196 2827 9236 2836
rect 9387 2708 9429 2717
rect 9387 2668 9388 2708
rect 9428 2668 9429 2708
rect 9387 2659 9429 2668
rect 9004 2624 9044 2633
rect 9004 2465 9044 2584
rect 9388 2624 9428 2659
rect 9099 2540 9141 2549
rect 9099 2500 9100 2540
rect 9140 2500 9141 2540
rect 9099 2491 9141 2500
rect 9003 2456 9045 2465
rect 9003 2416 9004 2456
rect 9044 2416 9045 2456
rect 9003 2407 9045 2416
rect 9003 2204 9045 2213
rect 9003 2164 9004 2204
rect 9044 2164 9045 2204
rect 9003 2155 9045 2164
rect 8907 2120 8949 2129
rect 8907 2080 8908 2120
rect 8948 2080 8949 2120
rect 8907 2071 8949 2080
rect 9004 2120 9044 2155
rect 9004 2069 9044 2080
rect 8812 1903 8852 1912
rect 9003 1952 9045 1961
rect 9003 1912 9004 1952
rect 9044 1912 9045 1952
rect 9003 1903 9045 1912
rect 9004 1112 9044 1903
rect 9100 1280 9140 2491
rect 9291 2120 9333 2129
rect 9291 2080 9292 2120
rect 9332 2080 9333 2120
rect 9291 2071 9333 2080
rect 9292 1986 9332 2071
rect 9388 1961 9428 2584
rect 9484 2604 9524 3163
rect 9676 2792 9716 3415
rect 9964 2885 10004 2970
rect 9963 2876 10005 2885
rect 9963 2836 9964 2876
rect 10004 2836 10005 2876
rect 9963 2827 10005 2836
rect 9676 2743 9716 2752
rect 9771 2708 9813 2717
rect 9771 2668 9772 2708
rect 9812 2668 9813 2708
rect 9771 2659 9813 2668
rect 9580 2624 9620 2633
rect 9484 2584 9580 2604
rect 9484 2564 9620 2584
rect 9676 2624 9716 2633
rect 9484 2381 9524 2564
rect 9483 2372 9525 2381
rect 9483 2332 9484 2372
rect 9524 2332 9525 2372
rect 9483 2323 9525 2332
rect 9676 2297 9716 2584
rect 9675 2288 9717 2297
rect 9675 2248 9676 2288
rect 9716 2248 9717 2288
rect 9675 2239 9717 2248
rect 9483 2120 9525 2129
rect 9483 2080 9484 2120
rect 9524 2080 9525 2120
rect 9483 2071 9525 2080
rect 9387 1952 9429 1961
rect 9387 1912 9388 1952
rect 9428 1912 9429 1952
rect 9387 1903 9429 1912
rect 9388 1709 9428 1903
rect 9484 1868 9524 2071
rect 9676 1877 9716 2239
rect 9484 1819 9524 1828
rect 9675 1868 9717 1877
rect 9675 1828 9676 1868
rect 9716 1828 9717 1868
rect 9675 1819 9717 1828
rect 9387 1700 9429 1709
rect 9387 1660 9388 1700
rect 9428 1660 9429 1700
rect 9387 1651 9429 1660
rect 9675 1700 9717 1709
rect 9675 1660 9676 1700
rect 9716 1660 9717 1700
rect 9675 1651 9717 1660
rect 9676 1566 9716 1651
rect 9387 1364 9429 1373
rect 9387 1324 9388 1364
rect 9428 1324 9429 1364
rect 9387 1315 9429 1324
rect 9100 1240 9332 1280
rect 8907 692 8949 701
rect 8907 652 8908 692
rect 8948 652 8949 692
rect 8907 643 8949 652
rect 8908 80 8948 643
rect 9004 365 9044 1072
rect 9099 1112 9141 1121
rect 9099 1072 9100 1112
rect 9140 1072 9141 1112
rect 9099 1063 9141 1072
rect 9003 356 9045 365
rect 9003 316 9004 356
rect 9044 316 9045 356
rect 9003 307 9045 316
rect 9100 80 9140 1063
rect 9195 1028 9237 1037
rect 9195 988 9196 1028
rect 9236 988 9237 1028
rect 9195 979 9237 988
rect 9196 894 9236 979
rect 9292 80 9332 1240
rect 9388 1121 9428 1315
rect 9772 1280 9812 2659
rect 10060 2549 10100 3928
rect 10155 3800 10197 3809
rect 10155 3760 10156 3800
rect 10196 3760 10197 3800
rect 10155 3751 10197 3760
rect 10156 2708 10196 3751
rect 10251 3548 10293 3557
rect 10251 3508 10252 3548
rect 10292 3508 10293 3548
rect 10251 3499 10293 3508
rect 10252 3464 10292 3499
rect 10252 3413 10292 3424
rect 10348 3296 10388 4171
rect 10444 4136 10484 6271
rect 10540 4313 10580 8128
rect 10636 7757 10676 7842
rect 10635 7748 10677 7757
rect 10635 7708 10636 7748
rect 10676 7708 10677 7748
rect 10635 7699 10677 7708
rect 10635 7244 10677 7253
rect 10635 7204 10636 7244
rect 10676 7204 10677 7244
rect 10635 7195 10677 7204
rect 10732 7244 10772 11731
rect 10828 10277 10868 12991
rect 10924 11612 10964 15595
rect 11499 15560 11541 15569
rect 11499 15520 11500 15560
rect 11540 15520 11541 15560
rect 11499 15511 11541 15520
rect 11500 15426 11540 15511
rect 11596 14720 11636 14729
rect 11788 14720 11828 16360
rect 11884 16073 11924 17704
rect 11980 16997 12020 21223
rect 12076 20684 12116 21475
rect 12267 21440 12309 21449
rect 12267 21400 12268 21440
rect 12308 21400 12309 21440
rect 12267 21391 12309 21400
rect 12268 20768 12308 21391
rect 12460 21281 12500 22240
rect 12556 22205 12596 23500
rect 12844 23120 12884 23995
rect 12844 23071 12884 23080
rect 12651 22868 12693 22877
rect 12651 22828 12652 22868
rect 12692 22828 12693 22868
rect 12651 22819 12693 22828
rect 12652 22734 12692 22819
rect 12747 22616 12789 22625
rect 12747 22576 12748 22616
rect 12788 22576 12789 22616
rect 12747 22567 12789 22576
rect 12555 22196 12597 22205
rect 12555 22156 12556 22196
rect 12596 22156 12597 22196
rect 12555 22147 12597 22156
rect 12748 21608 12788 22567
rect 12748 21559 12788 21568
rect 12843 21608 12885 21617
rect 12843 21568 12844 21608
rect 12884 21568 12980 21608
rect 12843 21559 12885 21568
rect 12844 21474 12884 21559
rect 12459 21272 12501 21281
rect 12459 21232 12460 21272
rect 12500 21232 12501 21272
rect 12459 21223 12501 21232
rect 12651 21188 12693 21197
rect 12651 21148 12652 21188
rect 12692 21148 12693 21188
rect 12651 21139 12693 21148
rect 12652 21029 12692 21139
rect 12651 21020 12693 21029
rect 12651 20980 12652 21020
rect 12692 20980 12693 21020
rect 12651 20971 12693 20980
rect 12308 20728 12596 20768
rect 12268 20719 12308 20728
rect 12076 20644 12212 20684
rect 12075 19676 12117 19685
rect 12075 19636 12076 19676
rect 12116 19636 12117 19676
rect 12075 19627 12117 19636
rect 11979 16988 12021 16997
rect 11979 16948 11980 16988
rect 12020 16948 12021 16988
rect 11979 16939 12021 16948
rect 11883 16064 11925 16073
rect 11883 16024 11884 16064
rect 11924 16024 11925 16064
rect 11883 16015 11925 16024
rect 11883 15896 11925 15905
rect 11883 15856 11884 15896
rect 11924 15856 11925 15896
rect 11883 15847 11925 15856
rect 11500 14680 11596 14720
rect 11211 14384 11253 14393
rect 11211 14344 11212 14384
rect 11252 14344 11253 14384
rect 11211 14335 11253 14344
rect 11212 14216 11252 14335
rect 11308 14225 11348 14244
rect 11212 14167 11252 14176
rect 11307 14216 11349 14225
rect 11404 14216 11444 14225
rect 11307 14176 11308 14216
rect 11348 14176 11404 14216
rect 11307 14167 11349 14176
rect 11404 14167 11444 14176
rect 11068 14038 11108 14047
rect 11108 13998 11348 14034
rect 11068 13994 11348 13998
rect 11068 13989 11108 13994
rect 11308 13460 11348 13994
rect 11500 13469 11540 14680
rect 11596 14671 11636 14680
rect 11692 14680 11828 14720
rect 11692 14393 11732 14680
rect 11787 14552 11829 14561
rect 11787 14512 11788 14552
rect 11828 14512 11829 14552
rect 11787 14503 11829 14512
rect 11788 14418 11828 14503
rect 11691 14384 11733 14393
rect 11691 14344 11692 14384
rect 11732 14344 11733 14384
rect 11691 14335 11733 14344
rect 11595 14216 11637 14225
rect 11884 14216 11924 15847
rect 11980 15560 12020 16939
rect 12076 15905 12116 19627
rect 12075 15896 12117 15905
rect 12075 15856 12076 15896
rect 12116 15856 12117 15896
rect 12075 15847 12117 15856
rect 11980 15511 12020 15520
rect 12172 15056 12212 20644
rect 12460 20600 12500 20609
rect 12268 20096 12308 20105
rect 12268 19844 12308 20056
rect 12363 20096 12405 20105
rect 12363 20056 12364 20096
rect 12404 20056 12405 20096
rect 12363 20047 12405 20056
rect 12364 19962 12404 20047
rect 12460 19844 12500 20560
rect 12268 19804 12500 19844
rect 12556 18593 12596 20728
rect 12652 20105 12692 20971
rect 12651 20096 12693 20105
rect 12651 20056 12652 20096
rect 12692 20056 12693 20096
rect 12651 20047 12693 20056
rect 12747 20012 12789 20021
rect 12747 19972 12748 20012
rect 12788 19972 12789 20012
rect 12747 19963 12789 19972
rect 12844 20012 12884 20023
rect 12748 19878 12788 19963
rect 12844 19937 12884 19972
rect 12843 19928 12885 19937
rect 12843 19888 12844 19928
rect 12884 19888 12885 19928
rect 12843 19879 12885 19888
rect 12843 19592 12885 19601
rect 12843 19552 12844 19592
rect 12884 19552 12885 19592
rect 12843 19543 12885 19552
rect 12844 19256 12884 19543
rect 12844 19207 12884 19216
rect 12267 18584 12309 18593
rect 12267 18544 12268 18584
rect 12308 18544 12309 18584
rect 12267 18535 12309 18544
rect 12555 18584 12597 18593
rect 12555 18544 12556 18584
rect 12596 18544 12597 18584
rect 12555 18535 12597 18544
rect 12652 18584 12692 18593
rect 12268 17081 12308 18535
rect 12652 18509 12692 18544
rect 12651 18500 12693 18509
rect 12651 18460 12652 18500
rect 12692 18460 12693 18500
rect 12651 18451 12693 18460
rect 12460 18332 12500 18341
rect 12460 17828 12500 18292
rect 12412 17788 12500 17828
rect 12412 17786 12452 17788
rect 12652 17753 12692 18451
rect 12412 17737 12452 17746
rect 12651 17744 12693 17753
rect 12651 17704 12652 17744
rect 12692 17704 12693 17744
rect 12651 17695 12693 17704
rect 12363 17576 12405 17585
rect 12363 17536 12364 17576
rect 12404 17536 12405 17576
rect 12363 17527 12405 17536
rect 12556 17576 12596 17585
rect 12651 17576 12693 17585
rect 12596 17536 12652 17576
rect 12692 17536 12693 17576
rect 12556 17527 12596 17536
rect 12651 17527 12693 17536
rect 12267 17072 12309 17081
rect 12267 17032 12268 17072
rect 12308 17032 12309 17072
rect 12267 17023 12309 17032
rect 12268 15569 12308 17023
rect 12364 15821 12404 17527
rect 12940 17408 12980 21568
rect 13036 19340 13076 24424
rect 13132 21617 13172 24844
rect 13228 22625 13268 25264
rect 13419 24296 13461 24305
rect 13419 24256 13420 24296
rect 13460 24256 13461 24296
rect 13419 24247 13461 24256
rect 13323 24212 13365 24221
rect 13323 24172 13324 24212
rect 13364 24172 13365 24212
rect 13323 24163 13365 24172
rect 13227 22616 13269 22625
rect 13227 22576 13228 22616
rect 13268 22576 13269 22616
rect 13227 22567 13269 22576
rect 13131 21608 13173 21617
rect 13324 21608 13364 24163
rect 13131 21568 13132 21608
rect 13172 21568 13173 21608
rect 13131 21559 13173 21568
rect 13228 21568 13324 21608
rect 13228 19517 13268 21568
rect 13324 21559 13364 21568
rect 13420 21440 13460 24247
rect 13516 22541 13556 27439
rect 13612 26144 13652 27448
rect 13708 27068 13748 27077
rect 13804 27068 13844 27523
rect 13748 27028 13844 27068
rect 13708 27019 13748 27028
rect 13900 26825 13940 28120
rect 13996 27572 14036 28288
rect 14188 27572 14228 27581
rect 14284 27572 14324 29203
rect 13996 27532 14132 27572
rect 14092 27488 14132 27532
rect 14228 27532 14324 27572
rect 14188 27523 14228 27532
rect 14092 27448 14137 27488
rect 13996 27404 14036 27413
rect 14097 27404 14137 27448
rect 14097 27364 14228 27404
rect 13996 27236 14036 27364
rect 13996 27196 14132 27236
rect 13996 26993 14036 27078
rect 14092 27077 14132 27196
rect 14091 27068 14133 27077
rect 14091 27028 14092 27068
rect 14132 27028 14133 27068
rect 14091 27019 14133 27028
rect 13995 26984 14037 26993
rect 13995 26944 13996 26984
rect 14036 26944 14037 26984
rect 13995 26935 14037 26944
rect 13803 26816 13845 26825
rect 13803 26776 13804 26816
rect 13844 26776 13845 26816
rect 13900 26816 14132 26825
rect 13900 26785 14092 26816
rect 13803 26767 13845 26776
rect 14092 26767 14132 26776
rect 13804 26682 13844 26767
rect 13612 26095 13652 26104
rect 13995 26144 14037 26153
rect 13995 26104 13996 26144
rect 14036 26104 14037 26144
rect 13995 26095 14037 26104
rect 13996 26010 14036 26095
rect 13804 25892 13844 25901
rect 13708 25852 13804 25892
rect 13708 25318 13748 25852
rect 13804 25843 13844 25852
rect 13899 25640 13941 25649
rect 13899 25600 13900 25640
rect 13940 25600 13941 25640
rect 13899 25591 13941 25600
rect 13708 25269 13748 25278
rect 13900 25220 13940 25591
rect 13995 25556 14037 25565
rect 13995 25516 13996 25556
rect 14036 25516 14037 25556
rect 13995 25507 14037 25516
rect 13900 25171 13940 25180
rect 13996 25145 14036 25507
rect 14092 25304 14132 25315
rect 14092 25229 14132 25264
rect 14091 25220 14133 25229
rect 14091 25180 14092 25220
rect 14132 25180 14133 25220
rect 14091 25171 14133 25180
rect 13995 25136 14037 25145
rect 13995 25096 13996 25136
rect 14036 25096 14037 25136
rect 13995 25087 14037 25096
rect 14188 24968 14228 27364
rect 14380 27161 14420 29791
rect 14379 27152 14421 27161
rect 14379 27112 14380 27152
rect 14420 27112 14421 27152
rect 14379 27103 14421 27112
rect 14379 26984 14421 26993
rect 14379 26944 14380 26984
rect 14420 26944 14421 26984
rect 14379 26935 14421 26944
rect 14283 26900 14325 26909
rect 14283 26860 14284 26900
rect 14324 26860 14325 26900
rect 14283 26851 14325 26860
rect 14284 26766 14324 26851
rect 14380 26816 14420 26935
rect 14476 26825 14516 31816
rect 14571 31688 14613 31697
rect 14668 31688 14708 32152
rect 14571 31648 14572 31688
rect 14612 31648 14708 31688
rect 14764 32192 14804 32201
rect 14857 32192 14897 32236
rect 14804 32152 14897 32192
rect 15052 32192 15092 32815
rect 15148 32696 15188 33571
rect 15532 33570 15572 33655
rect 15244 33452 15284 33461
rect 15284 33412 15572 33452
rect 15244 33403 15284 33412
rect 15339 33284 15381 33293
rect 15339 33244 15340 33284
rect 15380 33244 15381 33284
rect 15339 33235 15381 33244
rect 15244 32873 15284 32958
rect 15243 32864 15285 32873
rect 15243 32824 15244 32864
rect 15284 32824 15285 32864
rect 15340 32864 15380 33235
rect 15435 33116 15477 33125
rect 15435 33076 15436 33116
rect 15476 33076 15477 33116
rect 15435 33067 15477 33076
rect 15436 32982 15476 33067
rect 15436 32864 15476 32873
rect 15340 32824 15436 32864
rect 15243 32815 15285 32824
rect 15340 32696 15380 32705
rect 15148 32656 15284 32696
rect 14571 31639 14613 31648
rect 14764 31604 14804 32152
rect 15052 32143 15092 32152
rect 14955 32024 14997 32033
rect 15147 32024 15189 32033
rect 14955 31984 14956 32024
rect 14996 31984 15092 32024
rect 14955 31975 14997 31984
rect 14676 31564 14804 31604
rect 14676 31529 14716 31564
rect 14667 31520 14716 31529
rect 14859 31520 14901 31529
rect 14667 31480 14668 31520
rect 14708 31480 14716 31520
rect 14764 31480 14860 31520
rect 14900 31480 14901 31520
rect 14667 31471 14709 31480
rect 14764 31436 14804 31480
rect 14859 31471 14901 31480
rect 14764 31387 14804 31396
rect 14668 31352 14708 31361
rect 14668 30857 14708 31312
rect 14955 31184 14997 31193
rect 14955 31144 14956 31184
rect 14996 31144 14997 31184
rect 14955 31135 14997 31144
rect 14956 31050 14996 31135
rect 14667 30848 14709 30857
rect 14667 30808 14668 30848
rect 14708 30808 14709 30848
rect 14667 30799 14709 30808
rect 14668 30680 14708 30689
rect 14572 30640 14668 30680
rect 14572 30269 14612 30640
rect 14668 30631 14708 30640
rect 14859 30680 14901 30689
rect 14859 30640 14860 30680
rect 14900 30640 14901 30680
rect 14859 30631 14901 30640
rect 15052 30680 15092 31984
rect 15147 31984 15148 32024
rect 15188 31984 15189 32024
rect 15147 31975 15189 31984
rect 15148 31697 15188 31975
rect 15147 31688 15189 31697
rect 15147 31648 15148 31688
rect 15188 31648 15189 31688
rect 15147 31639 15189 31648
rect 15148 31352 15188 31639
rect 15148 31303 15188 31312
rect 15244 31184 15284 32656
rect 15340 32192 15380 32656
rect 15340 32143 15380 32152
rect 15436 32108 15476 32824
rect 15532 32528 15572 33412
rect 15628 32705 15668 32790
rect 15627 32696 15669 32705
rect 15627 32656 15628 32696
rect 15668 32656 15669 32696
rect 15627 32647 15669 32656
rect 15532 32488 15668 32528
rect 15436 32059 15476 32068
rect 15628 32108 15668 32488
rect 15724 32369 15764 34663
rect 15915 34376 15957 34385
rect 16012 34376 16052 36343
rect 16108 35309 16148 36436
rect 16396 36233 16436 36604
rect 16588 36569 16628 36688
rect 16587 36560 16629 36569
rect 16587 36520 16588 36560
rect 16628 36520 16629 36560
rect 16587 36511 16629 36520
rect 16491 36476 16533 36485
rect 16491 36436 16492 36476
rect 16532 36436 16533 36476
rect 16491 36427 16533 36436
rect 16395 36224 16437 36233
rect 16395 36184 16396 36224
rect 16436 36184 16437 36224
rect 16395 36175 16437 36184
rect 16204 35981 16244 36012
rect 16203 35972 16245 35981
rect 16203 35932 16204 35972
rect 16244 35932 16245 35972
rect 16203 35923 16245 35932
rect 16204 35888 16244 35923
rect 16204 35645 16244 35848
rect 16396 35720 16436 35729
rect 16203 35636 16245 35645
rect 16203 35596 16204 35636
rect 16244 35596 16245 35636
rect 16203 35587 16245 35596
rect 16299 35384 16341 35393
rect 16299 35344 16300 35384
rect 16340 35344 16341 35384
rect 16299 35335 16341 35344
rect 16107 35300 16149 35309
rect 16107 35260 16108 35300
rect 16148 35260 16149 35300
rect 16107 35251 16149 35260
rect 16204 35216 16244 35225
rect 16204 35048 16244 35176
rect 16300 35216 16340 35335
rect 16396 35225 16436 35680
rect 16300 35167 16340 35176
rect 16395 35216 16437 35225
rect 16395 35176 16396 35216
rect 16436 35176 16437 35216
rect 16395 35167 16437 35176
rect 16204 35008 16436 35048
rect 15915 34336 15916 34376
rect 15956 34336 16052 34376
rect 16203 34376 16245 34385
rect 16203 34336 16204 34376
rect 16244 34336 16245 34376
rect 15915 34327 15957 34336
rect 16203 34327 16245 34336
rect 15819 34292 15861 34301
rect 15819 34252 15820 34292
rect 15860 34252 15861 34292
rect 15819 34243 15861 34252
rect 15820 32957 15860 34243
rect 15916 34242 15956 34327
rect 16204 34040 16244 34327
rect 16396 34133 16436 35008
rect 16395 34124 16437 34133
rect 16395 34084 16396 34124
rect 16436 34084 16437 34124
rect 16395 34075 16437 34084
rect 16204 34000 16340 34040
rect 15916 33704 15956 33713
rect 15956 33691 16244 33704
rect 15956 33664 16204 33691
rect 15819 32948 15861 32957
rect 15819 32908 15820 32948
rect 15860 32908 15861 32948
rect 15819 32899 15861 32908
rect 15820 32864 15860 32899
rect 15916 32873 15956 33664
rect 16204 33642 16244 33651
rect 16204 33452 16244 33461
rect 16012 33412 16204 33452
rect 15820 32814 15860 32824
rect 15915 32864 15957 32873
rect 15915 32824 15916 32864
rect 15956 32824 15957 32864
rect 15915 32815 15957 32824
rect 15723 32360 15765 32369
rect 15723 32320 15724 32360
rect 15764 32320 15765 32360
rect 15723 32311 15765 32320
rect 15915 32360 15957 32369
rect 15915 32320 15916 32360
rect 15956 32320 15957 32360
rect 15915 32311 15957 32320
rect 15916 32226 15956 32311
rect 15723 32192 15765 32201
rect 15723 32152 15724 32192
rect 15764 32152 15765 32192
rect 15723 32143 15765 32152
rect 15628 32059 15668 32068
rect 15724 32058 15764 32143
rect 15532 32024 15572 32033
rect 15532 31352 15572 31984
rect 15915 31688 15957 31697
rect 15915 31648 15916 31688
rect 15956 31648 15957 31688
rect 15915 31639 15957 31648
rect 15052 30631 15092 30640
rect 15148 31144 15284 31184
rect 15340 31312 15572 31352
rect 14860 30546 14900 30631
rect 15148 30596 15188 31144
rect 15148 30547 15188 30556
rect 15340 30596 15380 31312
rect 15723 31184 15765 31193
rect 15723 31144 15724 31184
rect 15764 31144 15765 31184
rect 15723 31135 15765 31144
rect 15435 30680 15477 30689
rect 15435 30640 15436 30680
rect 15476 30640 15477 30680
rect 15435 30631 15477 30640
rect 15724 30680 15764 31135
rect 15724 30631 15764 30640
rect 15820 30680 15860 30689
rect 15340 30547 15380 30556
rect 15436 30546 15476 30631
rect 14668 30437 14708 30522
rect 15244 30512 15284 30521
rect 14667 30428 14709 30437
rect 14667 30388 14668 30428
rect 14708 30388 14709 30428
rect 14667 30379 14709 30388
rect 15147 30428 15189 30437
rect 15147 30388 15148 30428
rect 15188 30388 15189 30428
rect 15147 30379 15189 30388
rect 14571 30260 14613 30269
rect 14571 30220 14572 30260
rect 14612 30220 14613 30260
rect 14571 30211 14613 30220
rect 14667 30176 14709 30185
rect 14667 30136 14668 30176
rect 14708 30136 14709 30176
rect 15148 30176 15188 30379
rect 15244 30353 15284 30472
rect 15243 30344 15285 30353
rect 15243 30304 15244 30344
rect 15284 30304 15285 30344
rect 15243 30295 15285 30304
rect 15148 30136 15284 30176
rect 14667 30127 14709 30136
rect 14668 29000 14708 30127
rect 14859 29924 14901 29933
rect 14859 29884 14860 29924
rect 14900 29884 14901 29924
rect 14859 29875 14901 29884
rect 14860 29177 14900 29875
rect 14955 29336 14997 29345
rect 14955 29296 14956 29336
rect 14996 29296 14997 29336
rect 14955 29287 14997 29296
rect 14859 29168 14901 29177
rect 14859 29128 14860 29168
rect 14900 29128 14901 29168
rect 14859 29119 14901 29128
rect 14860 29034 14900 29119
rect 14668 28960 14804 29000
rect 14667 28160 14709 28169
rect 14667 28120 14668 28160
rect 14708 28120 14709 28160
rect 14667 28111 14709 28120
rect 14572 27656 14612 27665
rect 14572 27497 14612 27616
rect 14668 27656 14708 28111
rect 14668 27607 14708 27616
rect 14571 27488 14613 27497
rect 14571 27448 14572 27488
rect 14612 27448 14613 27488
rect 14571 27439 14613 27448
rect 14380 26767 14420 26776
rect 14475 26816 14517 26825
rect 14475 26776 14476 26816
rect 14516 26776 14517 26816
rect 14475 26767 14517 26776
rect 14572 26816 14612 26825
rect 14764 26816 14804 28960
rect 14860 27824 14900 27833
rect 14956 27824 14996 29287
rect 15051 29168 15093 29177
rect 15051 29128 15052 29168
rect 15092 29128 15093 29168
rect 15051 29119 15093 29128
rect 14900 27784 14996 27824
rect 15052 28916 15092 29119
rect 14860 27775 14900 27784
rect 14860 27656 14900 27667
rect 15052 27656 15092 28876
rect 15244 28505 15284 30136
rect 15820 30017 15860 30640
rect 15916 30101 15956 31639
rect 16012 30689 16052 33412
rect 16204 33403 16244 33412
rect 16204 32192 16244 32201
rect 16204 31865 16244 32152
rect 16203 31856 16245 31865
rect 16203 31816 16204 31856
rect 16244 31816 16245 31856
rect 16203 31807 16245 31816
rect 16300 30764 16340 34000
rect 16396 33704 16436 33713
rect 16396 33209 16436 33664
rect 16492 33704 16532 36427
rect 16587 35888 16629 35897
rect 16587 35848 16588 35888
rect 16628 35848 16629 35888
rect 16587 35839 16629 35848
rect 16588 35754 16628 35839
rect 16588 35216 16628 35225
rect 16588 34889 16628 35176
rect 16587 34880 16629 34889
rect 16587 34840 16588 34880
rect 16628 34840 16629 34880
rect 16587 34831 16629 34840
rect 16684 34040 16724 37687
rect 16780 37652 16820 38195
rect 16875 38200 16876 38240
rect 16916 38200 16917 38240
rect 16875 38191 16917 38200
rect 16780 37603 16820 37612
rect 16779 36896 16821 36905
rect 16779 36856 16780 36896
rect 16820 36856 16821 36896
rect 16779 36847 16821 36856
rect 16780 36728 16820 36847
rect 16780 36679 16820 36688
rect 16876 36728 16916 38191
rect 16972 37661 17012 39880
rect 17163 39752 17205 39761
rect 17163 39712 17164 39752
rect 17204 39712 17205 39752
rect 17163 39703 17205 39712
rect 17164 39618 17204 39703
rect 17260 38996 17300 40123
rect 18027 40004 18069 40013
rect 18027 39964 18028 40004
rect 18068 39964 18069 40004
rect 18027 39955 18069 39964
rect 17835 39920 17877 39929
rect 17835 39880 17836 39920
rect 17876 39880 17877 39920
rect 17835 39871 17877 39880
rect 18028 39920 18068 39955
rect 17836 39786 17876 39871
rect 18028 39869 18068 39880
rect 17692 39710 17732 39719
rect 17692 39668 17732 39670
rect 18219 39668 18261 39677
rect 17692 39628 17780 39668
rect 17740 39164 17780 39628
rect 18219 39628 18220 39668
rect 18260 39628 18261 39668
rect 18219 39619 18261 39628
rect 18220 39534 18260 39619
rect 17740 39115 17780 39124
rect 17547 39080 17589 39089
rect 17547 39040 17548 39080
rect 17588 39040 17589 39080
rect 17547 39031 17589 39040
rect 17164 38956 17300 38996
rect 17067 38240 17109 38249
rect 17067 38200 17068 38240
rect 17108 38200 17109 38240
rect 17067 38191 17109 38200
rect 17068 38106 17108 38191
rect 17068 37988 17108 37997
rect 16971 37652 17013 37661
rect 16971 37612 16972 37652
rect 17012 37612 17013 37652
rect 16971 37603 17013 37612
rect 16972 37484 17012 37493
rect 16972 37241 17012 37444
rect 17068 37325 17108 37948
rect 17164 37652 17204 38956
rect 17548 38912 17588 39031
rect 17548 38863 17588 38872
rect 17932 38912 17972 38921
rect 17259 38660 17301 38669
rect 17259 38620 17260 38660
rect 17300 38620 17301 38660
rect 17259 38611 17301 38620
rect 17260 38240 17300 38611
rect 17260 37997 17300 38200
rect 17356 38240 17396 38249
rect 17259 37988 17301 37997
rect 17259 37948 17260 37988
rect 17300 37948 17301 37988
rect 17259 37939 17301 37948
rect 17356 37820 17396 38200
rect 17643 38240 17685 38249
rect 17643 38200 17644 38240
rect 17684 38200 17685 38240
rect 17643 38191 17685 38200
rect 17644 38106 17684 38191
rect 17932 37820 17972 38872
rect 17164 37603 17204 37612
rect 17260 37780 17396 37820
rect 17836 37780 17972 37820
rect 18028 38912 18068 38921
rect 17163 37484 17205 37493
rect 17163 37444 17164 37484
rect 17204 37444 17205 37484
rect 17163 37435 17205 37444
rect 17067 37316 17109 37325
rect 17067 37276 17068 37316
rect 17108 37276 17109 37316
rect 17067 37267 17109 37276
rect 16971 37232 17013 37241
rect 16971 37192 16972 37232
rect 17012 37192 17013 37232
rect 16971 37183 17013 37192
rect 17164 37148 17204 37435
rect 17260 37409 17300 37780
rect 17355 37652 17397 37661
rect 17355 37612 17356 37652
rect 17396 37612 17397 37652
rect 17355 37603 17397 37612
rect 17259 37400 17301 37409
rect 17259 37360 17260 37400
rect 17300 37360 17301 37400
rect 17259 37351 17301 37360
rect 17356 37400 17396 37603
rect 17068 37108 17204 37148
rect 16971 36980 17013 36989
rect 16971 36940 16972 36980
rect 17012 36940 17013 36980
rect 16971 36931 17013 36940
rect 16972 36896 17012 36931
rect 16972 36845 17012 36856
rect 16876 36679 16916 36688
rect 17068 36728 17108 37108
rect 17068 36679 17108 36688
rect 17163 36728 17205 36737
rect 17163 36688 17164 36728
rect 17204 36688 17205 36728
rect 17163 36679 17205 36688
rect 16971 36644 17013 36653
rect 16971 36604 16972 36644
rect 17012 36604 17013 36644
rect 16971 36595 17013 36604
rect 16972 36308 17012 36595
rect 17164 36392 17204 36679
rect 17260 36569 17300 37351
rect 17356 37325 17396 37360
rect 17355 37316 17397 37325
rect 17355 37276 17356 37316
rect 17396 37276 17397 37316
rect 17355 37267 17397 37276
rect 17547 37148 17589 37157
rect 17547 37108 17548 37148
rect 17588 37108 17589 37148
rect 17547 37099 17589 37108
rect 17548 36728 17588 37099
rect 17836 36989 17876 37780
rect 18028 36989 18068 38872
rect 18220 38912 18260 38921
rect 18124 38744 18164 38755
rect 18124 38669 18164 38704
rect 18123 38660 18165 38669
rect 18123 38620 18124 38660
rect 18164 38620 18165 38660
rect 18123 38611 18165 38620
rect 18220 38081 18260 38872
rect 18219 38072 18261 38081
rect 18219 38032 18220 38072
rect 18260 38032 18261 38072
rect 18219 38023 18261 38032
rect 18316 37820 18356 40720
rect 18412 40676 18452 42223
rect 18508 42029 18548 42928
rect 18603 42104 18645 42113
rect 18603 42064 18604 42104
rect 18644 42064 18645 42104
rect 18603 42055 18645 42064
rect 18507 42020 18549 42029
rect 18507 41980 18508 42020
rect 18548 41980 18549 42020
rect 18507 41971 18549 41980
rect 18507 41180 18549 41189
rect 18507 41140 18508 41180
rect 18548 41140 18549 41180
rect 18507 41131 18549 41140
rect 18508 41046 18548 41131
rect 18604 40937 18644 42055
rect 18700 41441 18740 42928
rect 18892 42701 18932 42928
rect 18891 42692 18933 42701
rect 18891 42652 18892 42692
rect 18932 42652 18933 42692
rect 18891 42643 18933 42652
rect 18891 42524 18933 42533
rect 18891 42484 18892 42524
rect 18932 42484 18933 42524
rect 18891 42475 18933 42484
rect 18699 41432 18741 41441
rect 18699 41392 18700 41432
rect 18740 41392 18741 41432
rect 18699 41383 18741 41392
rect 18892 41180 18932 42475
rect 19084 41357 19124 42928
rect 19276 42449 19316 42928
rect 19468 42617 19508 42928
rect 19947 42776 19989 42785
rect 19947 42736 19948 42776
rect 19988 42736 19989 42776
rect 19947 42727 19989 42736
rect 19467 42608 19509 42617
rect 19467 42568 19468 42608
rect 19508 42568 19509 42608
rect 19467 42559 19509 42568
rect 19275 42440 19317 42449
rect 19275 42400 19276 42440
rect 19316 42400 19317 42440
rect 19275 42391 19317 42400
rect 19563 42188 19605 42197
rect 19563 42148 19564 42188
rect 19604 42148 19605 42188
rect 19563 42139 19605 42148
rect 19564 41432 19604 42139
rect 19564 41383 19604 41392
rect 19948 41432 19988 42727
rect 20048 41600 20416 41609
rect 20088 41560 20130 41600
rect 20170 41560 20212 41600
rect 20252 41560 20294 41600
rect 20334 41560 20376 41600
rect 20048 41551 20416 41560
rect 19948 41383 19988 41392
rect 19083 41348 19125 41357
rect 19083 41308 19084 41348
rect 19124 41308 19125 41348
rect 19083 41299 19125 41308
rect 18892 41131 18932 41140
rect 19180 41105 19220 41190
rect 19372 41180 19412 41189
rect 19276 41140 19372 41180
rect 19179 41096 19221 41105
rect 19179 41056 19180 41096
rect 19220 41056 19221 41096
rect 19179 41047 19221 41056
rect 18699 41012 18741 41021
rect 18699 40972 18700 41012
rect 18740 40972 18741 41012
rect 18699 40963 18741 40972
rect 18603 40928 18645 40937
rect 18603 40888 18604 40928
rect 18644 40888 18645 40928
rect 18603 40879 18645 40888
rect 18700 40878 18740 40963
rect 18808 40844 19176 40853
rect 18848 40804 18890 40844
rect 18930 40804 18972 40844
rect 19012 40804 19054 40844
rect 19094 40804 19136 40844
rect 18808 40795 19176 40804
rect 18412 40627 18452 40636
rect 18795 40676 18837 40685
rect 18795 40636 18796 40676
rect 18836 40636 18837 40676
rect 18795 40627 18837 40636
rect 18987 40676 19029 40685
rect 18987 40636 18988 40676
rect 19028 40636 19029 40676
rect 18987 40627 19029 40636
rect 18796 40542 18836 40627
rect 18603 40508 18645 40517
rect 18603 40468 18604 40508
rect 18644 40468 18645 40508
rect 18603 40459 18645 40468
rect 18988 40508 19028 40627
rect 18988 40459 19028 40468
rect 19180 40508 19220 40517
rect 18604 40374 18644 40459
rect 19180 40349 19220 40468
rect 19179 40340 19221 40349
rect 19179 40300 19180 40340
rect 19220 40300 19221 40340
rect 19179 40291 19221 40300
rect 18603 40256 18645 40265
rect 18603 40216 18604 40256
rect 18644 40216 18645 40256
rect 18603 40207 18645 40216
rect 18604 39668 18644 40207
rect 19276 39929 19316 41140
rect 19372 41131 19412 41140
rect 19755 41180 19797 41189
rect 19755 41140 19756 41180
rect 19796 41140 19797 41180
rect 19755 41131 19797 41140
rect 20121 41177 20161 41186
rect 19756 41046 19796 41131
rect 20121 40928 20161 41137
rect 19852 40888 20161 40928
rect 19372 40592 19412 40601
rect 19372 40349 19412 40552
rect 19564 40424 19604 40433
rect 19468 40384 19564 40424
rect 19371 40340 19413 40349
rect 19371 40300 19372 40340
rect 19412 40300 19413 40340
rect 19371 40291 19413 40300
rect 19275 39920 19317 39929
rect 19275 39880 19276 39920
rect 19316 39880 19317 39920
rect 19275 39871 19317 39880
rect 18796 39668 18836 39677
rect 18604 39619 18644 39628
rect 18700 39628 18796 39668
rect 18411 39500 18453 39509
rect 18411 39460 18412 39500
rect 18452 39460 18453 39500
rect 18411 39451 18453 39460
rect 18412 39366 18452 39451
rect 18700 39341 18740 39628
rect 18796 39619 18836 39628
rect 19179 39668 19221 39677
rect 19179 39628 19180 39668
rect 19220 39628 19221 39668
rect 19179 39619 19221 39628
rect 18988 39509 19028 39594
rect 19180 39534 19220 39619
rect 18987 39500 19029 39509
rect 19372 39500 19412 39509
rect 18987 39460 18988 39500
rect 19028 39460 19029 39500
rect 18987 39451 19029 39460
rect 19276 39460 19372 39500
rect 18699 39332 18741 39341
rect 18699 39292 18700 39332
rect 18740 39292 18741 39332
rect 18699 39283 18741 39292
rect 18808 39332 19176 39341
rect 18848 39292 18890 39332
rect 18930 39292 18972 39332
rect 19012 39292 19054 39332
rect 19094 39292 19136 39332
rect 18808 39283 19176 39292
rect 18411 39248 18453 39257
rect 18411 39208 18412 39248
rect 18452 39208 18453 39248
rect 18411 39199 18453 39208
rect 18603 39248 18645 39257
rect 18603 39208 18604 39248
rect 18644 39208 18645 39248
rect 18603 39199 18645 39208
rect 18412 38996 18452 39199
rect 18412 38947 18452 38956
rect 18604 38921 18644 39199
rect 18988 38921 19028 39006
rect 19276 39005 19316 39460
rect 19372 39451 19412 39460
rect 19468 39089 19508 40384
rect 19564 40375 19604 40384
rect 19755 40424 19797 40433
rect 19755 40384 19756 40424
rect 19796 40384 19797 40424
rect 19755 40375 19797 40384
rect 19756 40290 19796 40375
rect 19659 40256 19701 40265
rect 19659 40216 19660 40256
rect 19700 40216 19701 40256
rect 19659 40207 19701 40216
rect 19660 40122 19700 40207
rect 19564 39668 19604 39677
rect 19564 39173 19604 39628
rect 19756 39500 19796 39509
rect 19563 39164 19605 39173
rect 19563 39124 19564 39164
rect 19604 39124 19605 39164
rect 19563 39115 19605 39124
rect 19467 39080 19509 39089
rect 19467 39040 19468 39080
rect 19508 39040 19509 39080
rect 19467 39031 19509 39040
rect 19083 38996 19125 39005
rect 19083 38956 19084 38996
rect 19124 38956 19125 38996
rect 19083 38947 19125 38956
rect 19275 38996 19317 39005
rect 19275 38956 19276 38996
rect 19316 38956 19317 38996
rect 19275 38947 19317 38956
rect 19372 38996 19412 39005
rect 18603 38912 18645 38921
rect 18796 38912 18836 38921
rect 18603 38872 18604 38912
rect 18644 38872 18645 38912
rect 18603 38863 18645 38872
rect 18700 38872 18796 38912
rect 18411 38744 18453 38753
rect 18411 38704 18412 38744
rect 18452 38704 18453 38744
rect 18411 38695 18453 38704
rect 18604 38744 18644 38753
rect 18412 38240 18452 38695
rect 18604 38501 18644 38704
rect 18603 38492 18645 38501
rect 18603 38452 18604 38492
rect 18644 38452 18645 38492
rect 18603 38443 18645 38452
rect 18603 38240 18645 38249
rect 18412 38200 18548 38240
rect 18316 37780 18452 37820
rect 18315 37064 18357 37073
rect 18315 37024 18316 37064
rect 18356 37024 18357 37064
rect 18315 37015 18357 37024
rect 17835 36980 17877 36989
rect 17835 36940 17836 36980
rect 17876 36940 17877 36980
rect 17835 36931 17877 36940
rect 18027 36980 18069 36989
rect 18027 36940 18028 36980
rect 18068 36940 18069 36980
rect 18027 36931 18069 36940
rect 17643 36896 17685 36905
rect 17643 36856 17644 36896
rect 17684 36856 17685 36896
rect 17643 36847 17685 36856
rect 17644 36762 17684 36847
rect 17932 36821 17972 36852
rect 17931 36812 17973 36821
rect 17931 36772 17932 36812
rect 17972 36772 17973 36812
rect 17931 36763 17973 36772
rect 18316 36812 18356 37015
rect 18316 36763 18356 36772
rect 17356 36683 17396 36692
rect 17452 36686 17492 36695
rect 17259 36560 17301 36569
rect 17259 36520 17260 36560
rect 17300 36520 17301 36560
rect 17259 36511 17301 36520
rect 17164 36352 17300 36392
rect 16972 36268 17204 36308
rect 17067 35552 17109 35561
rect 17067 35512 17068 35552
rect 17108 35512 17109 35552
rect 17067 35503 17109 35512
rect 16779 35468 16821 35477
rect 16779 35428 16780 35468
rect 16820 35428 16821 35468
rect 16779 35419 16821 35428
rect 16492 33655 16532 33664
rect 16588 34000 16724 34040
rect 16395 33200 16437 33209
rect 16395 33160 16396 33200
rect 16436 33160 16437 33200
rect 16395 33151 16437 33160
rect 16588 33041 16628 34000
rect 16684 33872 16724 33881
rect 16780 33872 16820 35419
rect 17068 35384 17108 35503
rect 17068 35335 17108 35344
rect 17068 35216 17108 35225
rect 16910 35201 16950 35210
rect 16910 35057 16950 35161
rect 16909 35048 16951 35057
rect 16909 35008 16910 35048
rect 16950 35008 16951 35048
rect 16909 34999 16951 35008
rect 17068 34805 17108 35176
rect 17164 35216 17204 36268
rect 17164 35167 17204 35176
rect 17163 35048 17205 35057
rect 17163 35008 17164 35048
rect 17204 35008 17205 35048
rect 17163 34999 17205 35008
rect 17067 34796 17109 34805
rect 17067 34756 17068 34796
rect 17108 34756 17109 34796
rect 17067 34747 17109 34756
rect 17164 34628 17204 34999
rect 16724 33832 16820 33872
rect 17068 34588 17204 34628
rect 16684 33823 16724 33832
rect 16876 33704 16916 33713
rect 16916 33664 17012 33704
rect 16876 33655 16916 33664
rect 16779 33536 16821 33545
rect 16779 33496 16780 33536
rect 16820 33496 16821 33536
rect 16779 33487 16821 33496
rect 16683 33284 16725 33293
rect 16683 33244 16684 33284
rect 16724 33244 16725 33284
rect 16683 33235 16725 33244
rect 16587 33032 16629 33041
rect 16587 32992 16588 33032
rect 16628 32992 16629 33032
rect 16587 32983 16629 32992
rect 16684 32453 16724 33235
rect 16683 32444 16725 32453
rect 16683 32404 16684 32444
rect 16724 32404 16725 32444
rect 16683 32395 16725 32404
rect 16684 31520 16724 31529
rect 16684 31361 16724 31480
rect 16396 31352 16436 31361
rect 16396 31193 16436 31312
rect 16683 31352 16725 31361
rect 16683 31312 16684 31352
rect 16724 31312 16725 31352
rect 16683 31303 16725 31312
rect 16395 31184 16437 31193
rect 16395 31144 16396 31184
rect 16436 31144 16437 31184
rect 16395 31135 16437 31144
rect 16780 30848 16820 33487
rect 16875 32864 16917 32873
rect 16875 32824 16876 32864
rect 16916 32824 16917 32864
rect 16875 32815 16917 32824
rect 16684 30808 16820 30848
rect 16300 30724 16436 30764
rect 16011 30680 16053 30689
rect 16011 30640 16012 30680
rect 16052 30640 16053 30680
rect 16011 30631 16053 30640
rect 16204 30596 16244 30605
rect 15915 30092 15957 30101
rect 15915 30052 15916 30092
rect 15956 30052 15957 30092
rect 15915 30043 15957 30052
rect 15819 30008 15861 30017
rect 15819 29968 15820 30008
rect 15860 29968 15861 30008
rect 15819 29959 15861 29968
rect 15916 29933 15956 30043
rect 15435 29924 15477 29933
rect 15435 29884 15436 29924
rect 15476 29884 15477 29924
rect 15435 29875 15477 29884
rect 15915 29924 15957 29933
rect 15915 29884 15916 29924
rect 15956 29884 15957 29924
rect 15915 29875 15957 29884
rect 15436 29840 15476 29875
rect 15436 29789 15476 29800
rect 15819 29840 15861 29849
rect 15819 29800 15820 29840
rect 15860 29800 15861 29840
rect 15819 29791 15861 29800
rect 15820 29706 15860 29791
rect 15628 29672 15668 29681
rect 15340 29632 15628 29672
rect 15340 29261 15380 29632
rect 15628 29623 15668 29632
rect 15339 29252 15381 29261
rect 15339 29212 15340 29252
rect 15380 29212 15381 29252
rect 15339 29203 15381 29212
rect 15916 29252 15956 29261
rect 16204 29252 16244 30556
rect 15956 29212 16244 29252
rect 16300 30596 16340 30605
rect 15243 28496 15285 28505
rect 15243 28456 15244 28496
rect 15284 28456 15285 28496
rect 15243 28447 15285 28456
rect 15244 28328 15284 28447
rect 15340 28328 15380 29203
rect 15531 29168 15573 29177
rect 15531 29128 15532 29168
rect 15572 29128 15573 29168
rect 15531 29119 15573 29128
rect 15819 29168 15861 29177
rect 15819 29128 15820 29168
rect 15860 29128 15861 29168
rect 15819 29119 15861 29128
rect 15435 29084 15477 29093
rect 15435 29044 15436 29084
rect 15476 29044 15477 29084
rect 15435 29035 15477 29044
rect 15436 28580 15476 29035
rect 15532 29034 15572 29119
rect 15820 29034 15860 29119
rect 15627 29000 15669 29009
rect 15627 28960 15628 29000
rect 15668 28960 15669 29000
rect 15627 28951 15669 28960
rect 15436 28531 15476 28540
rect 15531 28412 15573 28421
rect 15531 28372 15532 28412
rect 15572 28372 15573 28412
rect 15531 28363 15573 28372
rect 15436 28328 15476 28337
rect 15340 28288 15436 28328
rect 15244 28279 15284 28288
rect 15436 28279 15476 28288
rect 15532 28328 15572 28363
rect 15532 28277 15572 28288
rect 15339 27824 15381 27833
rect 15339 27784 15340 27824
rect 15380 27784 15381 27824
rect 15339 27775 15381 27784
rect 15340 27656 15380 27775
rect 15436 27656 15476 27665
rect 15052 27648 15170 27656
rect 15052 27639 15188 27648
rect 15052 27616 15148 27639
rect 14860 27581 14900 27616
rect 15130 27599 15148 27616
rect 15130 27581 15188 27599
rect 15340 27616 15436 27656
rect 14859 27572 14901 27581
rect 14859 27532 14860 27572
rect 14900 27532 14901 27572
rect 15130 27572 15189 27581
rect 15130 27532 15148 27572
rect 15188 27532 15189 27572
rect 14859 27523 14901 27532
rect 15147 27523 15189 27532
rect 15148 27504 15188 27523
rect 15051 27488 15093 27497
rect 15051 27448 15052 27488
rect 15092 27448 15093 27488
rect 15051 27439 15093 27448
rect 14859 27152 14901 27161
rect 14859 27112 14860 27152
rect 14900 27112 14901 27152
rect 14859 27103 14901 27112
rect 14612 26776 14804 26816
rect 14572 26767 14612 26776
rect 14283 26648 14325 26657
rect 14283 26608 14284 26648
rect 14324 26608 14325 26648
rect 14283 26599 14325 26608
rect 13900 24928 14228 24968
rect 13803 23876 13845 23885
rect 13803 23836 13804 23876
rect 13844 23836 13845 23876
rect 13803 23827 13845 23836
rect 13804 23792 13844 23827
rect 13804 23129 13844 23752
rect 13803 23120 13845 23129
rect 13803 23080 13804 23120
rect 13844 23080 13845 23120
rect 13803 23071 13845 23080
rect 13515 22532 13557 22541
rect 13515 22492 13516 22532
rect 13556 22492 13557 22532
rect 13515 22483 13557 22492
rect 13516 22324 13652 22364
rect 13516 22322 13556 22324
rect 13516 22273 13556 22282
rect 13515 22196 13557 22205
rect 13515 22156 13516 22196
rect 13556 22156 13557 22196
rect 13515 22147 13557 22156
rect 13324 21400 13460 21440
rect 13324 20096 13364 21400
rect 13419 20768 13461 20777
rect 13419 20728 13420 20768
rect 13460 20728 13461 20768
rect 13419 20719 13461 20728
rect 13420 20634 13460 20719
rect 13516 20105 13556 22147
rect 13612 22037 13652 22324
rect 13708 22112 13748 22121
rect 13748 22072 13844 22112
rect 13708 22063 13748 22072
rect 13611 22028 13653 22037
rect 13611 21988 13612 22028
rect 13652 21988 13653 22028
rect 13611 21979 13653 21988
rect 13227 19508 13269 19517
rect 13227 19468 13228 19508
rect 13268 19468 13269 19508
rect 13324 19508 13364 20056
rect 13515 20096 13557 20105
rect 13515 20056 13516 20096
rect 13556 20056 13557 20096
rect 13515 20047 13557 20056
rect 13324 19468 13556 19508
rect 13227 19459 13269 19468
rect 13419 19340 13461 19349
rect 13036 19300 13268 19340
rect 13035 19172 13077 19181
rect 13035 19132 13036 19172
rect 13076 19132 13077 19172
rect 13035 19123 13077 19132
rect 13036 19038 13076 19123
rect 13131 17996 13173 18005
rect 13131 17956 13132 17996
rect 13172 17956 13173 17996
rect 13131 17947 13173 17956
rect 12652 17368 12980 17408
rect 13036 17744 13076 17753
rect 12363 15812 12405 15821
rect 12363 15772 12364 15812
rect 12404 15772 12405 15812
rect 12363 15763 12405 15772
rect 12267 15560 12309 15569
rect 12267 15520 12268 15560
rect 12308 15520 12309 15560
rect 12267 15511 12309 15520
rect 12459 15140 12501 15149
rect 12652 15140 12692 17368
rect 13036 17240 13076 17704
rect 13132 17744 13172 17947
rect 13228 17753 13268 19300
rect 13419 19300 13420 19340
rect 13460 19300 13461 19340
rect 13419 19291 13461 19300
rect 13324 19256 13364 19267
rect 13324 19181 13364 19216
rect 13420 19256 13460 19291
rect 13323 19172 13365 19181
rect 13323 19132 13324 19172
rect 13364 19132 13365 19172
rect 13323 19123 13365 19132
rect 13420 18257 13460 19216
rect 13419 18248 13461 18257
rect 13419 18208 13420 18248
rect 13460 18208 13461 18248
rect 13419 18199 13461 18208
rect 13516 17912 13556 19468
rect 13612 18173 13652 21979
rect 13804 21603 13844 22072
rect 13804 21554 13844 21563
rect 13804 20082 13844 20091
rect 13804 19424 13844 20042
rect 13900 19853 13940 24928
rect 13995 24800 14037 24809
rect 13995 24760 13996 24800
rect 14036 24760 14037 24800
rect 13995 24751 14037 24760
rect 13996 22952 14036 24751
rect 14284 24716 14324 26599
rect 14571 25304 14613 25313
rect 14571 25264 14572 25304
rect 14612 25264 14613 25304
rect 14571 25255 14613 25264
rect 14188 24676 14324 24716
rect 14188 24548 14228 24676
rect 14379 24632 14421 24641
rect 14284 24590 14324 24599
rect 14283 24550 14284 24557
rect 14379 24592 14380 24632
rect 14420 24592 14421 24632
rect 14379 24583 14421 24592
rect 14324 24550 14325 24557
rect 14283 24548 14325 24550
rect 14188 24508 14284 24548
rect 14324 24508 14325 24548
rect 14283 24499 14325 24508
rect 14284 24455 14324 24499
rect 14380 23885 14420 24583
rect 14476 24380 14516 24389
rect 14379 23876 14421 23885
rect 14379 23836 14380 23876
rect 14420 23836 14421 23876
rect 14379 23827 14421 23836
rect 14476 23792 14516 24340
rect 14476 23743 14516 23752
rect 14572 23792 14612 25255
rect 14612 23752 14708 23792
rect 14572 23743 14612 23752
rect 14284 23204 14324 23213
rect 14324 23164 14612 23204
rect 14284 23155 14324 23164
rect 14092 23120 14132 23129
rect 14572 23120 14612 23164
rect 14132 23080 14228 23120
rect 14092 23071 14132 23080
rect 13996 22912 14132 22952
rect 13995 21692 14037 21701
rect 13995 21652 13996 21692
rect 14036 21652 14037 21692
rect 13995 21643 14037 21652
rect 13996 21558 14036 21643
rect 13996 20180 14036 20189
rect 13899 19844 13941 19853
rect 13899 19804 13900 19844
rect 13940 19804 13941 19844
rect 13899 19795 13941 19804
rect 13899 19508 13941 19517
rect 13899 19468 13900 19508
rect 13940 19468 13941 19508
rect 13899 19459 13941 19468
rect 13708 19384 13844 19424
rect 13708 18761 13748 19384
rect 13900 19340 13940 19459
rect 13804 19256 13844 19267
rect 13804 19181 13844 19216
rect 13803 19172 13845 19181
rect 13803 19132 13804 19172
rect 13844 19132 13845 19172
rect 13803 19123 13845 19132
rect 13900 19013 13940 19300
rect 13899 19004 13941 19013
rect 13899 18964 13900 19004
rect 13940 18964 13941 19004
rect 13899 18955 13941 18964
rect 13707 18752 13749 18761
rect 13707 18712 13708 18752
rect 13748 18712 13749 18752
rect 13707 18703 13749 18712
rect 13996 18593 14036 20140
rect 14092 19676 14132 22912
rect 14188 22289 14228 23080
rect 14572 23071 14612 23080
rect 14668 23120 14708 23752
rect 14379 23036 14421 23045
rect 14379 22996 14380 23036
rect 14420 22996 14421 23036
rect 14379 22987 14421 22996
rect 14283 22364 14325 22373
rect 14283 22324 14284 22364
rect 14324 22324 14325 22364
rect 14283 22315 14325 22324
rect 14187 22280 14229 22289
rect 14187 22240 14188 22280
rect 14228 22240 14229 22280
rect 14187 22231 14229 22240
rect 14188 20693 14228 22231
rect 14187 20684 14229 20693
rect 14187 20644 14188 20684
rect 14228 20644 14229 20684
rect 14187 20635 14229 20644
rect 14188 19853 14228 19938
rect 14187 19844 14229 19853
rect 14187 19804 14188 19844
rect 14228 19804 14229 19844
rect 14187 19795 14229 19804
rect 14091 19636 14132 19676
rect 14091 19592 14131 19636
rect 14091 19552 14132 19592
rect 14092 18920 14132 19552
rect 14284 19004 14324 22315
rect 14380 20684 14420 22987
rect 14668 22868 14708 23080
rect 14764 23045 14804 26776
rect 14860 24641 14900 27103
rect 15052 26573 15092 27439
rect 15051 26564 15093 26573
rect 15051 26524 15052 26564
rect 15092 26524 15093 26564
rect 15051 26515 15093 26524
rect 15243 26396 15285 26405
rect 15243 26356 15244 26396
rect 15284 26356 15285 26396
rect 15243 26347 15285 26356
rect 15244 26144 15284 26347
rect 15340 26237 15380 27616
rect 15436 27607 15476 27616
rect 15532 27656 15572 27665
rect 15436 26321 15476 26406
rect 15435 26312 15477 26321
rect 15435 26272 15436 26312
rect 15476 26272 15477 26312
rect 15435 26263 15477 26272
rect 15339 26228 15381 26237
rect 15339 26188 15340 26228
rect 15380 26188 15381 26228
rect 15339 26179 15381 26188
rect 15244 25733 15284 26104
rect 15435 26144 15477 26153
rect 15532 26144 15572 27616
rect 15628 27320 15668 28951
rect 15916 28748 15956 29212
rect 16204 28916 16244 28925
rect 15820 28708 15956 28748
rect 16012 28876 16204 28916
rect 15820 28589 15860 28708
rect 15819 28580 15861 28589
rect 16012 28580 16052 28876
rect 16204 28867 16244 28876
rect 15819 28540 15820 28580
rect 15860 28540 15861 28580
rect 15819 28531 15861 28540
rect 15977 28540 16052 28580
rect 15977 28343 16017 28540
rect 16203 28496 16245 28505
rect 16203 28456 16204 28496
rect 16244 28456 16245 28496
rect 16203 28447 16245 28456
rect 15723 28328 15765 28337
rect 15723 28288 15724 28328
rect 15764 28288 15765 28328
rect 15723 28279 15765 28288
rect 15820 28328 15860 28337
rect 15977 28294 16017 28303
rect 16204 28328 16244 28447
rect 15724 28194 15764 28279
rect 15820 27665 15860 28288
rect 16204 28279 16244 28288
rect 16203 28160 16245 28169
rect 16203 28120 16204 28160
rect 16244 28120 16245 28160
rect 16203 28111 16245 28120
rect 15916 27784 16148 27824
rect 15819 27656 15861 27665
rect 15819 27616 15820 27656
rect 15860 27616 15861 27656
rect 15819 27607 15861 27616
rect 15820 27488 15860 27497
rect 15916 27488 15956 27784
rect 15860 27448 15956 27488
rect 16012 27656 16052 27665
rect 15820 27439 15860 27448
rect 15628 27280 15956 27320
rect 15627 27152 15669 27161
rect 15627 27112 15628 27152
rect 15668 27112 15669 27152
rect 15627 27103 15669 27112
rect 15435 26104 15436 26144
rect 15476 26104 15572 26144
rect 15435 26095 15477 26104
rect 15243 25724 15285 25733
rect 15243 25684 15244 25724
rect 15284 25684 15285 25724
rect 15243 25675 15285 25684
rect 15244 25304 15284 25675
rect 15436 25481 15476 26095
rect 15628 25976 15668 27103
rect 15820 26816 15860 26825
rect 15820 26405 15860 26776
rect 15819 26396 15861 26405
rect 15819 26356 15820 26396
rect 15860 26356 15861 26396
rect 15819 26347 15861 26356
rect 15723 26312 15765 26321
rect 15723 26272 15724 26312
rect 15764 26272 15765 26312
rect 15723 26263 15765 26272
rect 15724 26144 15764 26263
rect 15724 26060 15764 26104
rect 15819 26060 15861 26069
rect 15724 26020 15820 26060
rect 15860 26020 15861 26060
rect 15819 26011 15861 26020
rect 15628 25936 15764 25976
rect 15531 25556 15573 25565
rect 15531 25516 15532 25556
rect 15572 25516 15573 25556
rect 15531 25507 15573 25516
rect 15435 25472 15477 25481
rect 15435 25432 15436 25472
rect 15476 25432 15477 25472
rect 15435 25423 15477 25432
rect 15532 25422 15572 25507
rect 15340 25304 15380 25313
rect 15244 25264 15340 25304
rect 15244 25061 15284 25264
rect 15340 25255 15380 25264
rect 15435 25304 15477 25313
rect 15435 25264 15436 25304
rect 15476 25264 15477 25304
rect 15435 25255 15477 25264
rect 15436 25136 15476 25255
rect 15340 25096 15476 25136
rect 15243 25052 15285 25061
rect 15243 25012 15244 25052
rect 15284 25012 15285 25052
rect 15243 25003 15285 25012
rect 14859 24632 14901 24641
rect 14859 24592 14860 24632
rect 14900 24592 14901 24632
rect 14859 24583 14901 24592
rect 14955 24380 14997 24389
rect 14955 24340 14956 24380
rect 14996 24340 14997 24380
rect 14955 24331 14997 24340
rect 14956 23792 14996 24331
rect 14763 23036 14805 23045
rect 14763 22996 14764 23036
rect 14804 22996 14805 23036
rect 14956 23036 14996 23752
rect 15051 23792 15093 23801
rect 15051 23752 15052 23792
rect 15092 23752 15188 23792
rect 15051 23743 15093 23752
rect 15052 23658 15092 23743
rect 15052 23036 15092 23045
rect 14956 22996 15052 23036
rect 14763 22987 14805 22996
rect 14668 22828 14804 22868
rect 14668 21608 14708 21617
rect 14668 21113 14708 21568
rect 14764 21608 14804 22828
rect 14860 22280 14900 22291
rect 14860 22205 14900 22240
rect 14859 22196 14901 22205
rect 14859 22156 14860 22196
rect 14900 22156 14901 22196
rect 14859 22147 14901 22156
rect 14667 21104 14709 21113
rect 14667 21064 14668 21104
rect 14708 21064 14709 21104
rect 14667 21055 14709 21064
rect 14668 20768 14708 20777
rect 14668 20693 14708 20728
rect 14667 20684 14709 20693
rect 14380 20644 14612 20684
rect 14475 20516 14517 20525
rect 14475 20476 14476 20516
rect 14516 20476 14517 20516
rect 14475 20467 14517 20476
rect 14476 20273 14516 20467
rect 14475 20264 14517 20273
rect 14475 20224 14476 20264
rect 14516 20224 14517 20264
rect 14475 20215 14517 20224
rect 14379 20096 14421 20105
rect 14379 20056 14380 20096
rect 14420 20056 14421 20096
rect 14379 20047 14421 20056
rect 14380 19601 14420 20047
rect 14379 19592 14421 19601
rect 14379 19552 14380 19592
rect 14420 19552 14421 19592
rect 14379 19543 14421 19552
rect 14379 19424 14421 19433
rect 14379 19384 14380 19424
rect 14420 19384 14421 19424
rect 14379 19375 14421 19384
rect 14380 19256 14420 19375
rect 14380 19207 14420 19216
rect 14284 18964 14420 19004
rect 14092 18880 14324 18920
rect 14091 18752 14133 18761
rect 14091 18712 14092 18752
rect 14132 18712 14133 18752
rect 14091 18703 14133 18712
rect 14092 18618 14132 18703
rect 13995 18584 14037 18593
rect 13900 18542 13940 18551
rect 13899 18502 13900 18509
rect 13995 18544 13996 18584
rect 14036 18544 14037 18584
rect 13995 18535 14037 18544
rect 13940 18502 13941 18509
rect 13899 18500 13941 18502
rect 13899 18460 13900 18500
rect 13940 18460 13941 18500
rect 13899 18451 13941 18460
rect 14091 18500 14133 18509
rect 14091 18460 14092 18500
rect 14132 18460 14133 18500
rect 14091 18451 14133 18460
rect 13900 18407 13940 18451
rect 13707 18332 13749 18341
rect 14092 18332 14132 18451
rect 13707 18292 13708 18332
rect 13748 18292 13749 18332
rect 13707 18283 13749 18292
rect 13996 18292 14132 18332
rect 13611 18164 13653 18173
rect 13611 18124 13612 18164
rect 13652 18124 13653 18164
rect 13611 18115 13653 18124
rect 13420 17872 13556 17912
rect 13132 17408 13172 17704
rect 13227 17744 13269 17753
rect 13227 17704 13228 17744
rect 13268 17704 13269 17744
rect 13227 17695 13269 17704
rect 13132 17368 13268 17408
rect 13132 17240 13172 17249
rect 13036 17200 13132 17240
rect 13132 17191 13172 17200
rect 12939 17156 12981 17165
rect 12939 17116 12940 17156
rect 12980 17116 12981 17156
rect 12939 17107 12981 17116
rect 12940 17072 12980 17107
rect 12940 17021 12980 17032
rect 12747 16400 12789 16409
rect 12747 16360 12748 16400
rect 12788 16360 12789 16400
rect 12747 16351 12789 16360
rect 12748 15317 12788 16351
rect 13228 15980 13268 17368
rect 12844 15940 13268 15980
rect 13324 17072 13364 17081
rect 12747 15308 12789 15317
rect 12747 15268 12748 15308
rect 12788 15268 12789 15308
rect 12747 15259 12789 15268
rect 12459 15100 12460 15140
rect 12500 15100 12501 15140
rect 12459 15091 12501 15100
rect 12556 15100 12692 15140
rect 12172 15016 12308 15056
rect 12171 14888 12213 14897
rect 12171 14848 12172 14888
rect 12212 14848 12213 14888
rect 12171 14839 12213 14848
rect 12076 14720 12116 14729
rect 11980 14680 12076 14720
rect 11980 14561 12020 14680
rect 12076 14671 12116 14680
rect 12172 14720 12212 14839
rect 12172 14671 12212 14680
rect 11979 14552 12021 14561
rect 11979 14512 11980 14552
rect 12020 14512 12021 14552
rect 11979 14503 12021 14512
rect 11979 14384 12021 14393
rect 11979 14344 11980 14384
rect 12020 14344 12021 14384
rect 11979 14335 12021 14344
rect 11595 14176 11596 14216
rect 11636 14176 11637 14216
rect 11595 14167 11637 14176
rect 11692 14176 11924 14216
rect 11596 13964 11636 14167
rect 11596 13915 11636 13924
rect 11692 13796 11732 14176
rect 11980 14132 12020 14335
rect 11884 14092 12020 14132
rect 11787 13880 11829 13889
rect 11787 13840 11788 13880
rect 11828 13840 11829 13880
rect 11787 13831 11829 13840
rect 11596 13756 11732 13796
rect 11308 13411 11348 13420
rect 11499 13460 11541 13469
rect 11499 13420 11500 13460
rect 11540 13420 11541 13460
rect 11499 13411 11541 13420
rect 11500 13301 11540 13411
rect 11499 13292 11541 13301
rect 11499 13252 11500 13292
rect 11540 13252 11541 13292
rect 11499 13243 11541 13252
rect 11115 13208 11157 13217
rect 11115 13168 11116 13208
rect 11156 13168 11157 13208
rect 11115 13159 11157 13168
rect 11403 13208 11445 13217
rect 11403 13168 11404 13208
rect 11444 13168 11445 13208
rect 11403 13159 11445 13168
rect 11116 13074 11156 13159
rect 11116 12545 11156 12630
rect 11115 12536 11157 12545
rect 11115 12496 11116 12536
rect 11156 12496 11157 12536
rect 11115 12487 11157 12496
rect 11307 12536 11349 12545
rect 11307 12496 11308 12536
rect 11348 12496 11349 12536
rect 11307 12487 11349 12496
rect 11115 12368 11157 12377
rect 11115 12328 11116 12368
rect 11156 12328 11157 12368
rect 11115 12319 11157 12328
rect 11116 11873 11156 12319
rect 11115 11864 11157 11873
rect 11115 11824 11116 11864
rect 11156 11824 11157 11864
rect 11115 11815 11157 11824
rect 10924 11572 11156 11612
rect 11019 11108 11061 11117
rect 11019 11068 11020 11108
rect 11060 11068 11061 11108
rect 11019 11059 11061 11068
rect 11020 10445 11060 11059
rect 11019 10436 11061 10445
rect 11019 10396 11020 10436
rect 11060 10396 11061 10436
rect 11019 10387 11061 10396
rect 10827 10268 10869 10277
rect 10827 10228 10828 10268
rect 10868 10228 10869 10268
rect 10827 10219 10869 10228
rect 11116 9521 11156 11572
rect 11308 11453 11348 12487
rect 11307 11444 11349 11453
rect 11307 11404 11308 11444
rect 11348 11404 11349 11444
rect 11307 11395 11349 11404
rect 11404 11117 11444 13159
rect 11499 13040 11541 13049
rect 11499 13000 11500 13040
rect 11540 13000 11541 13040
rect 11499 12991 11541 13000
rect 11500 12906 11540 12991
rect 11596 11957 11636 13756
rect 11788 13746 11828 13831
rect 11691 13292 11733 13301
rect 11691 13252 11692 13292
rect 11732 13252 11733 13292
rect 11691 13243 11733 13252
rect 11692 13158 11732 13243
rect 11787 13208 11829 13217
rect 11787 13168 11788 13208
rect 11828 13168 11829 13208
rect 11884 13208 11924 14092
rect 11979 13964 12021 13973
rect 11979 13924 11980 13964
rect 12020 13924 12021 13964
rect 11979 13915 12021 13924
rect 11980 13830 12020 13915
rect 12171 13880 12213 13889
rect 12171 13840 12172 13880
rect 12212 13840 12213 13880
rect 12171 13831 12213 13840
rect 12172 13746 12212 13831
rect 12268 13217 12308 15016
rect 12363 13964 12405 13973
rect 12363 13924 12364 13964
rect 12404 13924 12405 13964
rect 12363 13915 12405 13924
rect 12364 13830 12404 13915
rect 11980 13208 12020 13217
rect 11884 13168 11980 13208
rect 11787 13159 11829 13168
rect 11691 12536 11733 12545
rect 11691 12496 11692 12536
rect 11732 12496 11733 12536
rect 11691 12487 11733 12496
rect 11595 11948 11637 11957
rect 11595 11908 11596 11948
rect 11636 11908 11637 11948
rect 11595 11899 11637 11908
rect 11596 11360 11636 11899
rect 11692 11696 11732 12487
rect 11692 11647 11732 11656
rect 11500 11320 11636 11360
rect 11403 11108 11445 11117
rect 11403 11068 11404 11108
rect 11444 11068 11445 11108
rect 11403 11059 11445 11068
rect 11500 11024 11540 11320
rect 11691 11192 11733 11201
rect 11691 11152 11692 11192
rect 11732 11152 11733 11192
rect 11691 11143 11733 11152
rect 11500 10975 11540 10984
rect 11692 11024 11732 11143
rect 11692 10865 11732 10984
rect 11691 10856 11733 10865
rect 11691 10816 11692 10856
rect 11732 10816 11733 10856
rect 11691 10807 11733 10816
rect 11788 10688 11828 13159
rect 11980 12293 12020 13168
rect 12267 13208 12309 13217
rect 12267 13168 12268 13208
rect 12308 13168 12309 13208
rect 12267 13159 12309 13168
rect 12363 12536 12405 12545
rect 12363 12496 12364 12536
rect 12404 12496 12405 12536
rect 12363 12487 12405 12496
rect 12364 12402 12404 12487
rect 11979 12284 12021 12293
rect 11979 12244 11980 12284
rect 12020 12244 12021 12284
rect 11979 12235 12021 12244
rect 12363 12284 12405 12293
rect 12363 12244 12364 12284
rect 12404 12244 12405 12284
rect 12363 12235 12405 12244
rect 12172 11696 12212 11705
rect 11884 11612 11924 11621
rect 12172 11612 12212 11656
rect 12267 11696 12309 11705
rect 12267 11656 12268 11696
rect 12308 11656 12309 11696
rect 12267 11647 12309 11656
rect 11924 11572 12212 11612
rect 11884 11563 11924 11572
rect 12268 11562 12308 11647
rect 12364 11276 12404 12235
rect 12172 11236 12404 11276
rect 11979 10772 12021 10781
rect 11979 10732 11980 10772
rect 12020 10732 12021 10772
rect 11979 10723 12021 10732
rect 11692 10648 11828 10688
rect 11595 10352 11637 10361
rect 11595 10312 11596 10352
rect 11636 10312 11637 10352
rect 11595 10303 11637 10312
rect 11596 10184 11636 10303
rect 11596 10109 11636 10144
rect 11595 10100 11637 10109
rect 11595 10060 11596 10100
rect 11636 10060 11637 10100
rect 11595 10051 11637 10060
rect 11403 10016 11445 10025
rect 11596 10020 11636 10051
rect 11403 9976 11404 10016
rect 11444 9976 11445 10016
rect 11403 9967 11445 9976
rect 11404 9857 11444 9967
rect 11403 9848 11445 9857
rect 11403 9808 11404 9848
rect 11444 9808 11445 9848
rect 11403 9799 11445 9808
rect 11499 9680 11541 9689
rect 11499 9640 11500 9680
rect 11540 9640 11541 9680
rect 11499 9631 11541 9640
rect 10924 9512 10964 9521
rect 10827 8756 10869 8765
rect 10827 8716 10828 8756
rect 10868 8716 10869 8756
rect 10827 8707 10869 8716
rect 10828 8686 10868 8707
rect 10828 8621 10868 8646
rect 10924 8177 10964 9472
rect 11115 9512 11157 9521
rect 11115 9472 11116 9512
rect 11156 9472 11157 9512
rect 11115 9463 11157 9472
rect 11308 9512 11348 9521
rect 11019 9428 11061 9437
rect 11019 9388 11020 9428
rect 11060 9388 11061 9428
rect 11019 9379 11061 9388
rect 11212 9386 11252 9395
rect 11020 9294 11060 9379
rect 11115 9344 11157 9353
rect 11115 9304 11116 9344
rect 11156 9304 11157 9344
rect 11115 9295 11157 9304
rect 11116 9210 11156 9295
rect 11019 9176 11061 9185
rect 11019 9136 11020 9176
rect 11060 9136 11061 9176
rect 11019 9127 11061 9136
rect 11020 8743 11060 9127
rect 11115 8840 11157 8849
rect 11212 8840 11252 9346
rect 11308 9176 11348 9472
rect 11500 9512 11540 9631
rect 11500 9463 11540 9472
rect 11308 9136 11636 9176
rect 11307 9008 11349 9017
rect 11307 8968 11308 9008
rect 11348 8968 11349 9008
rect 11307 8959 11349 8968
rect 11308 8840 11348 8959
rect 11596 8924 11636 9136
rect 11596 8875 11636 8884
rect 11115 8800 11116 8840
rect 11156 8800 11252 8840
rect 11298 8800 11348 8840
rect 11115 8791 11157 8800
rect 11298 8756 11338 8800
rect 11020 8703 11156 8743
rect 11020 8513 11060 8598
rect 11019 8504 11061 8513
rect 11019 8464 11020 8504
rect 11060 8464 11061 8504
rect 11019 8455 11061 8464
rect 10923 8168 10965 8177
rect 10923 8128 10924 8168
rect 10964 8128 10965 8168
rect 10923 8119 10965 8128
rect 10924 8000 10964 8011
rect 10924 7925 10964 7960
rect 10923 7916 10965 7925
rect 10923 7876 10924 7916
rect 10964 7876 10965 7916
rect 10923 7867 10965 7876
rect 11019 7664 11061 7673
rect 11019 7624 11020 7664
rect 11060 7624 11061 7664
rect 11019 7615 11061 7624
rect 10923 7412 10965 7421
rect 10923 7372 10924 7412
rect 10964 7372 10965 7412
rect 10923 7363 10965 7372
rect 10732 7195 10772 7204
rect 10636 5237 10676 7195
rect 10924 6329 10964 7363
rect 10923 6320 10965 6329
rect 10923 6280 10924 6320
rect 10964 6280 10965 6320
rect 10923 6271 10965 6280
rect 10731 5396 10773 5405
rect 10731 5356 10732 5396
rect 10772 5356 10773 5396
rect 10731 5347 10773 5356
rect 10635 5228 10677 5237
rect 10635 5188 10636 5228
rect 10676 5188 10677 5228
rect 10635 5179 10677 5188
rect 10636 4976 10676 5179
rect 10636 4927 10676 4936
rect 10539 4304 10581 4313
rect 10539 4264 10540 4304
rect 10580 4264 10581 4304
rect 10539 4255 10581 4264
rect 10444 4087 10484 4096
rect 10539 4136 10581 4145
rect 10539 4096 10540 4136
rect 10580 4096 10581 4136
rect 10539 4087 10581 4096
rect 10636 4136 10676 4145
rect 10540 4002 10580 4087
rect 10636 3977 10676 4096
rect 10732 4136 10772 5347
rect 10732 4087 10772 4096
rect 10924 4136 10964 4145
rect 10924 3977 10964 4096
rect 10635 3968 10677 3977
rect 10635 3928 10636 3968
rect 10676 3928 10677 3968
rect 10635 3919 10677 3928
rect 10923 3968 10965 3977
rect 10923 3928 10924 3968
rect 10964 3928 10965 3968
rect 10923 3919 10965 3928
rect 10443 3884 10485 3893
rect 10443 3844 10444 3884
rect 10484 3844 10485 3884
rect 10443 3835 10485 3844
rect 10444 3632 10484 3835
rect 11020 3725 11060 7615
rect 11116 5237 11156 8703
rect 11212 8716 11338 8756
rect 11212 7337 11252 8716
rect 11404 8672 11444 8681
rect 11308 8657 11348 8666
rect 11308 8513 11348 8617
rect 11307 8504 11349 8513
rect 11307 8464 11308 8504
rect 11348 8464 11349 8504
rect 11307 8455 11349 8464
rect 11404 8009 11444 8632
rect 11595 8672 11637 8681
rect 11595 8632 11596 8672
rect 11636 8632 11637 8672
rect 11595 8623 11637 8632
rect 11596 8538 11636 8623
rect 11403 8000 11445 8009
rect 11403 7960 11404 8000
rect 11444 7960 11445 8000
rect 11403 7951 11445 7960
rect 11499 7580 11541 7589
rect 11499 7540 11500 7580
rect 11540 7540 11541 7580
rect 11499 7531 11541 7540
rect 11500 7421 11540 7531
rect 11499 7412 11541 7421
rect 11499 7372 11500 7412
rect 11540 7372 11541 7412
rect 11499 7363 11541 7372
rect 11211 7328 11253 7337
rect 11692 7328 11732 10648
rect 11883 10604 11925 10613
rect 11883 10564 11884 10604
rect 11924 10564 11925 10604
rect 11883 10555 11925 10564
rect 11788 10436 11828 10445
rect 11884 10436 11924 10555
rect 11828 10396 11924 10436
rect 11788 10387 11828 10396
rect 11980 10016 12020 10723
rect 12076 10184 12116 10193
rect 12076 10025 12116 10144
rect 12075 10016 12117 10025
rect 11980 9976 12076 10016
rect 12116 9976 12117 10016
rect 11787 9764 11829 9773
rect 11787 9724 11788 9764
rect 11828 9724 11829 9764
rect 11787 9715 11829 9724
rect 11788 7589 11828 9715
rect 11883 8756 11925 8765
rect 11980 8756 12020 9976
rect 12075 9967 12117 9976
rect 12075 9848 12117 9857
rect 12075 9808 12076 9848
rect 12116 9808 12117 9848
rect 12075 9799 12117 9808
rect 11883 8716 11884 8756
rect 11924 8716 12020 8756
rect 11883 8707 11925 8716
rect 11884 8672 11924 8707
rect 11884 8621 11924 8632
rect 11883 8084 11925 8093
rect 11883 8044 11884 8084
rect 11924 8044 11925 8084
rect 11883 8035 11925 8044
rect 11787 7580 11829 7589
rect 11787 7540 11788 7580
rect 11828 7540 11829 7580
rect 11787 7531 11829 7540
rect 11211 7288 11212 7328
rect 11252 7288 11253 7328
rect 11211 7279 11253 7288
rect 11596 7288 11732 7328
rect 11212 7160 11252 7279
rect 11212 7111 11252 7120
rect 11499 6908 11541 6917
rect 11499 6868 11500 6908
rect 11540 6868 11541 6908
rect 11499 6859 11541 6868
rect 11211 5648 11253 5657
rect 11211 5608 11212 5648
rect 11252 5608 11253 5648
rect 11211 5599 11253 5608
rect 11404 5648 11444 5657
rect 11115 5228 11157 5237
rect 11115 5188 11116 5228
rect 11156 5188 11157 5228
rect 11115 5179 11157 5188
rect 11116 4985 11156 5066
rect 11115 4976 11157 4985
rect 11115 4931 11116 4976
rect 11156 4931 11157 4976
rect 11115 4927 11157 4931
rect 11116 4922 11156 4927
rect 11116 4304 11156 4313
rect 11212 4304 11252 5599
rect 11404 5489 11444 5608
rect 11403 5480 11445 5489
rect 11403 5440 11404 5480
rect 11444 5440 11445 5480
rect 11403 5431 11445 5440
rect 11403 5228 11445 5237
rect 11403 5188 11404 5228
rect 11444 5188 11445 5228
rect 11403 5179 11445 5188
rect 11307 5144 11349 5153
rect 11307 5104 11308 5144
rect 11348 5104 11349 5144
rect 11307 5095 11349 5104
rect 11308 5060 11348 5095
rect 11308 5009 11348 5020
rect 11156 4264 11252 4304
rect 11116 4255 11156 4264
rect 11116 4136 11156 4145
rect 11116 3893 11156 4096
rect 11211 4136 11253 4145
rect 11211 4096 11212 4136
rect 11252 4096 11253 4136
rect 11211 4087 11253 4096
rect 11404 4136 11444 5179
rect 11500 5060 11540 6859
rect 11596 6320 11636 7288
rect 11740 7169 11780 7178
rect 11780 7129 11828 7160
rect 11740 7120 11828 7129
rect 11788 6656 11828 7120
rect 11884 7076 11924 8035
rect 12076 7748 12116 9799
rect 12172 9092 12212 11236
rect 12267 11108 12309 11117
rect 12267 11068 12268 11108
rect 12308 11068 12309 11108
rect 12267 11059 12309 11068
rect 12268 9605 12308 11059
rect 12460 10856 12500 15091
rect 12556 14813 12596 15100
rect 12748 15056 12788 15259
rect 12652 15016 12788 15056
rect 12555 14804 12597 14813
rect 12555 14764 12556 14804
rect 12596 14764 12597 14804
rect 12555 14755 12597 14764
rect 12652 14804 12692 15016
rect 12652 14755 12692 14764
rect 12556 14670 12596 14755
rect 12747 14720 12789 14729
rect 12747 14680 12748 14720
rect 12788 14680 12789 14720
rect 12747 14671 12789 14680
rect 12652 14048 12692 14057
rect 12556 14008 12652 14048
rect 12556 12620 12596 14008
rect 12652 13999 12692 14008
rect 12748 14048 12788 14671
rect 12748 13999 12788 14008
rect 12844 13973 12884 15940
rect 13324 15896 13364 17032
rect 13132 15856 13364 15896
rect 13132 15149 13172 15856
rect 13420 15737 13460 17872
rect 13611 17828 13653 17837
rect 13611 17788 13612 17828
rect 13652 17788 13653 17828
rect 13611 17779 13653 17788
rect 13515 17744 13557 17753
rect 13515 17704 13516 17744
rect 13556 17704 13557 17744
rect 13515 17695 13557 17704
rect 13516 16409 13556 17695
rect 13612 17694 13652 17779
rect 13708 17753 13748 18283
rect 13899 18248 13941 18257
rect 13899 18208 13900 18248
rect 13940 18208 13941 18248
rect 13899 18199 13941 18208
rect 13803 18164 13845 18173
rect 13803 18124 13804 18164
rect 13844 18124 13845 18164
rect 13803 18115 13845 18124
rect 13707 17744 13749 17753
rect 13707 17704 13708 17744
rect 13748 17704 13749 17744
rect 13707 17695 13749 17704
rect 13515 16400 13557 16409
rect 13515 16360 13516 16400
rect 13556 16360 13557 16400
rect 13515 16351 13557 16360
rect 13516 16232 13556 16241
rect 13419 15728 13461 15737
rect 13419 15688 13420 15728
rect 13460 15688 13461 15728
rect 13419 15679 13461 15688
rect 13227 15644 13269 15653
rect 13227 15604 13228 15644
rect 13268 15604 13269 15644
rect 13227 15595 13269 15604
rect 13228 15560 13268 15595
rect 13228 15509 13268 15520
rect 13323 15392 13365 15401
rect 13323 15352 13324 15392
rect 13364 15352 13365 15392
rect 13323 15343 13365 15352
rect 13420 15392 13460 15401
rect 13516 15392 13556 16192
rect 13612 16232 13652 16243
rect 13612 16157 13652 16192
rect 13611 16148 13653 16157
rect 13611 16108 13612 16148
rect 13652 16108 13653 16148
rect 13611 16099 13653 16108
rect 13612 15569 13652 16099
rect 13611 15560 13653 15569
rect 13611 15520 13612 15560
rect 13652 15520 13653 15560
rect 13611 15511 13653 15520
rect 13708 15560 13748 17695
rect 13708 15511 13748 15520
rect 13460 15352 13556 15392
rect 13420 15343 13460 15352
rect 13227 15308 13269 15317
rect 13227 15268 13228 15308
rect 13268 15268 13269 15308
rect 13227 15259 13269 15268
rect 13131 15140 13173 15149
rect 13131 15100 13132 15140
rect 13172 15100 13173 15140
rect 13131 15091 13173 15100
rect 12939 14888 12981 14897
rect 12939 14848 12940 14888
rect 12980 14848 12981 14888
rect 12939 14839 12981 14848
rect 12843 13964 12885 13973
rect 12843 13924 12844 13964
rect 12884 13924 12885 13964
rect 12843 13915 12885 13924
rect 12651 13880 12693 13889
rect 12651 13840 12652 13880
rect 12692 13840 12693 13880
rect 12651 13831 12693 13840
rect 12556 12571 12596 12580
rect 12652 12452 12692 13831
rect 12556 12412 12692 12452
rect 12748 12536 12788 12545
rect 12556 11117 12596 12412
rect 12748 12209 12788 12496
rect 12747 12200 12789 12209
rect 12747 12160 12748 12200
rect 12788 12160 12789 12200
rect 12747 12151 12789 12160
rect 12651 11864 12693 11873
rect 12651 11824 12652 11864
rect 12692 11824 12693 11864
rect 12651 11815 12693 11824
rect 12652 11780 12692 11815
rect 12652 11729 12692 11740
rect 12748 11780 12788 11789
rect 12940 11780 12980 14839
rect 13132 14720 13172 14729
rect 13132 14309 13172 14680
rect 13131 14300 13173 14309
rect 13131 14260 13132 14300
rect 13172 14260 13173 14300
rect 13131 14251 13173 14260
rect 13228 14132 13268 15259
rect 13132 14092 13268 14132
rect 13132 14048 13172 14092
rect 13132 13999 13172 14008
rect 13227 13964 13269 13973
rect 13227 13924 13228 13964
rect 13268 13924 13269 13964
rect 13227 13915 13269 13924
rect 13228 13830 13268 13915
rect 13227 13544 13269 13553
rect 13227 13504 13228 13544
rect 13268 13504 13269 13544
rect 13227 13495 13269 13504
rect 13228 13250 13268 13495
rect 13228 13201 13268 13210
rect 13035 12536 13077 12545
rect 13035 12496 13036 12536
rect 13076 12496 13077 12536
rect 13035 12487 13077 12496
rect 12788 11740 12980 11780
rect 12748 11731 12788 11740
rect 12940 11621 12980 11740
rect 12939 11612 12981 11621
rect 12939 11572 12940 11612
rect 12980 11572 12981 11612
rect 12939 11563 12981 11572
rect 12555 11108 12597 11117
rect 12555 11068 12556 11108
rect 12596 11068 12597 11108
rect 12555 11059 12597 11068
rect 12940 11024 12980 11033
rect 13036 11024 13076 12487
rect 13227 11696 13269 11705
rect 13227 11656 13228 11696
rect 13268 11656 13269 11696
rect 13227 11647 13269 11656
rect 13228 11562 13268 11647
rect 13324 11369 13364 15343
rect 13707 15308 13749 15317
rect 13707 15268 13708 15308
rect 13748 15268 13749 15308
rect 13707 15259 13749 15268
rect 13612 14725 13652 14734
rect 13515 14300 13557 14309
rect 13515 14260 13516 14300
rect 13556 14260 13557 14300
rect 13515 14251 13557 14260
rect 13419 13460 13461 13469
rect 13419 13420 13420 13460
rect 13460 13420 13461 13460
rect 13419 13411 13461 13420
rect 13420 13326 13460 13411
rect 13516 12209 13556 14251
rect 13612 13469 13652 14685
rect 13708 14048 13748 15259
rect 13804 14720 13844 18115
rect 13900 16316 13940 18199
rect 13996 17081 14036 18292
rect 14187 18164 14229 18173
rect 14187 18124 14188 18164
rect 14228 18124 14229 18164
rect 14187 18115 14229 18124
rect 14092 17744 14132 17753
rect 14188 17744 14228 18115
rect 14132 17704 14228 17744
rect 14092 17695 14132 17704
rect 13995 17072 14037 17081
rect 13995 17032 13996 17072
rect 14036 17032 14037 17072
rect 13995 17023 14037 17032
rect 13996 16316 14036 16325
rect 13900 16276 13996 16316
rect 13996 16267 14036 16276
rect 14188 16241 14228 17704
rect 14092 16232 14132 16241
rect 13899 16064 13941 16073
rect 13899 16024 13900 16064
rect 13940 16024 13941 16064
rect 13899 16015 13941 16024
rect 13900 15317 13940 16015
rect 13899 15308 13941 15317
rect 13899 15268 13900 15308
rect 13940 15268 13941 15308
rect 13899 15259 13941 15268
rect 13804 14680 13940 14720
rect 13708 13999 13748 14008
rect 13804 14552 13844 14561
rect 13804 13889 13844 14512
rect 13803 13880 13845 13889
rect 13803 13840 13804 13880
rect 13844 13840 13845 13880
rect 13803 13831 13845 13840
rect 13611 13460 13653 13469
rect 13611 13420 13612 13460
rect 13652 13420 13653 13460
rect 13611 13411 13653 13420
rect 13900 13217 13940 14680
rect 13995 14636 14037 14645
rect 13995 14596 13996 14636
rect 14036 14596 14037 14636
rect 13995 14587 14037 14596
rect 13804 13208 13844 13217
rect 13899 13208 13941 13217
rect 13844 13168 13900 13208
rect 13940 13168 13941 13208
rect 13804 13159 13844 13168
rect 13899 13159 13941 13168
rect 13611 13124 13653 13133
rect 13611 13084 13612 13124
rect 13652 13084 13653 13124
rect 13611 13075 13653 13084
rect 13612 12990 13652 13075
rect 13900 12545 13940 13159
rect 13996 12872 14036 14587
rect 14092 13049 14132 16192
rect 14187 16232 14229 16241
rect 14187 16192 14188 16232
rect 14228 16192 14229 16232
rect 14187 16183 14229 16192
rect 14188 15737 14228 16183
rect 14187 15728 14229 15737
rect 14187 15688 14188 15728
rect 14228 15688 14229 15728
rect 14187 15679 14229 15688
rect 14188 14034 14228 14043
rect 14188 13133 14228 13994
rect 14187 13124 14229 13133
rect 14187 13084 14188 13124
rect 14228 13084 14229 13124
rect 14187 13075 14229 13084
rect 14091 13040 14133 13049
rect 14091 13000 14092 13040
rect 14132 13000 14133 13040
rect 14091 12991 14133 13000
rect 13996 12832 14132 12872
rect 14092 12545 14132 12832
rect 13899 12536 13941 12545
rect 13996 12536 14036 12545
rect 13899 12496 13900 12536
rect 13940 12496 13996 12536
rect 13899 12487 13941 12496
rect 13996 12487 14036 12496
rect 14091 12536 14133 12545
rect 14091 12496 14092 12536
rect 14132 12496 14133 12536
rect 14091 12487 14133 12496
rect 13900 12402 13940 12487
rect 13707 12284 13749 12293
rect 13707 12244 13708 12284
rect 13748 12244 13749 12284
rect 13707 12235 13749 12244
rect 13515 12200 13557 12209
rect 13515 12160 13516 12200
rect 13556 12160 13557 12200
rect 13515 12151 13557 12160
rect 13419 12032 13461 12041
rect 13419 11992 13420 12032
rect 13460 11992 13461 12032
rect 13419 11983 13461 11992
rect 13323 11360 13365 11369
rect 13323 11320 13324 11360
rect 13364 11320 13365 11360
rect 13323 11311 13365 11320
rect 13131 11108 13173 11117
rect 13131 11068 13132 11108
rect 13172 11068 13173 11108
rect 13131 11059 13173 11068
rect 13324 11108 13364 11117
rect 12980 10984 13076 11024
rect 12940 10975 12980 10984
rect 12460 10816 12596 10856
rect 12459 10688 12501 10697
rect 12459 10648 12460 10688
rect 12500 10648 12501 10688
rect 12459 10639 12501 10648
rect 12363 10184 12405 10193
rect 12363 10144 12364 10184
rect 12404 10144 12405 10184
rect 12363 10135 12405 10144
rect 12460 10184 12500 10639
rect 12460 10135 12500 10144
rect 12364 10050 12404 10135
rect 12267 9596 12309 9605
rect 12267 9556 12268 9596
rect 12308 9556 12309 9596
rect 12267 9547 12309 9556
rect 12172 9052 12500 9092
rect 12171 8924 12213 8933
rect 12171 8884 12172 8924
rect 12212 8884 12213 8924
rect 12171 8875 12213 8884
rect 12172 8672 12212 8875
rect 12172 8623 12212 8632
rect 12267 8588 12309 8597
rect 12267 8548 12268 8588
rect 12308 8548 12309 8588
rect 12267 8539 12309 8548
rect 12171 8084 12213 8093
rect 12171 8044 12172 8084
rect 12212 8044 12213 8084
rect 12171 8035 12213 8044
rect 12172 8000 12212 8035
rect 12172 7949 12212 7960
rect 12268 7925 12308 8539
rect 12267 7916 12309 7925
rect 12267 7876 12268 7916
rect 12308 7876 12309 7916
rect 12267 7867 12309 7876
rect 12364 7748 12404 7757
rect 12076 7708 12212 7748
rect 11979 7496 12021 7505
rect 11979 7456 11980 7496
rect 12020 7456 12021 7496
rect 11979 7447 12021 7456
rect 11884 7027 11924 7036
rect 11884 6656 11924 6665
rect 11788 6616 11884 6656
rect 11884 6607 11924 6616
rect 11692 6497 11732 6582
rect 11691 6488 11733 6497
rect 11691 6448 11692 6488
rect 11732 6448 11733 6488
rect 11691 6439 11733 6448
rect 11596 6280 11732 6320
rect 11596 5480 11636 5489
rect 11596 5237 11636 5440
rect 11595 5228 11637 5237
rect 11595 5188 11596 5228
rect 11636 5188 11637 5228
rect 11595 5179 11637 5188
rect 11500 5011 11540 5020
rect 11596 4976 11636 4985
rect 11499 4472 11541 4481
rect 11499 4432 11500 4472
rect 11540 4432 11541 4472
rect 11499 4423 11541 4432
rect 11404 4087 11444 4096
rect 11500 4136 11540 4423
rect 11596 4229 11636 4936
rect 11595 4220 11637 4229
rect 11595 4180 11596 4220
rect 11636 4180 11637 4220
rect 11595 4171 11637 4180
rect 11500 4087 11540 4096
rect 11115 3884 11157 3893
rect 11115 3844 11116 3884
rect 11156 3844 11157 3884
rect 11115 3835 11157 3844
rect 10635 3716 10677 3725
rect 10635 3676 10636 3716
rect 10676 3676 10677 3716
rect 10635 3667 10677 3676
rect 11019 3716 11061 3725
rect 11019 3676 11020 3716
rect 11060 3676 11061 3716
rect 11019 3667 11061 3676
rect 10444 3583 10484 3592
rect 10539 3548 10581 3557
rect 10539 3508 10540 3548
rect 10580 3508 10581 3548
rect 10539 3499 10581 3508
rect 10540 3305 10580 3499
rect 10636 3380 10676 3667
rect 11212 3632 11252 4087
rect 11403 3884 11445 3893
rect 11403 3844 11404 3884
rect 11444 3844 11445 3884
rect 11403 3835 11445 3844
rect 11212 3583 11252 3592
rect 11020 3473 11060 3558
rect 11019 3464 11061 3473
rect 11019 3424 11020 3464
rect 11060 3424 11061 3464
rect 11019 3415 11061 3424
rect 11116 3464 11156 3473
rect 10636 3331 10676 3340
rect 10156 2659 10196 2668
rect 10252 3256 10388 3296
rect 10539 3296 10581 3305
rect 10539 3256 10540 3296
rect 10580 3256 10581 3296
rect 10059 2540 10101 2549
rect 10059 2500 10060 2540
rect 10100 2500 10101 2540
rect 10059 2491 10101 2500
rect 10252 2465 10292 3256
rect 10539 3247 10581 3256
rect 11116 3221 11156 3424
rect 11308 3464 11348 3473
rect 11115 3212 11157 3221
rect 11115 3172 11116 3212
rect 11156 3172 11157 3212
rect 11115 3163 11157 3172
rect 11308 3053 11348 3424
rect 11404 3464 11444 3835
rect 11505 3464 11545 3473
rect 11404 3415 11444 3424
rect 11500 3424 11505 3464
rect 11500 3415 11545 3424
rect 11403 3212 11445 3221
rect 11403 3172 11404 3212
rect 11444 3172 11445 3212
rect 11403 3163 11445 3172
rect 11307 3044 11349 3053
rect 11307 3004 11308 3044
rect 11348 3004 11349 3044
rect 11307 2995 11349 3004
rect 10539 2708 10581 2717
rect 10539 2668 10540 2708
rect 10580 2668 10581 2708
rect 10539 2659 10581 2668
rect 11115 2708 11157 2717
rect 11115 2668 11116 2708
rect 11156 2668 11157 2708
rect 11115 2659 11157 2668
rect 11404 2708 11444 3163
rect 10540 2574 10580 2659
rect 10828 2624 10868 2633
rect 10635 2540 10677 2549
rect 10635 2500 10636 2540
rect 10676 2500 10677 2540
rect 10635 2491 10677 2500
rect 10251 2456 10293 2465
rect 10251 2416 10252 2456
rect 10292 2416 10293 2456
rect 10251 2407 10293 2416
rect 10348 2456 10388 2465
rect 9867 2288 9909 2297
rect 9867 2248 9868 2288
rect 9908 2248 9909 2288
rect 9867 2239 9909 2248
rect 9676 1240 9812 1280
rect 9483 1196 9525 1205
rect 9483 1156 9484 1196
rect 9524 1156 9525 1196
rect 9483 1147 9525 1156
rect 9387 1112 9429 1121
rect 9387 1072 9388 1112
rect 9428 1072 9429 1112
rect 9387 1063 9429 1072
rect 9388 944 9428 953
rect 9388 533 9428 904
rect 9387 524 9429 533
rect 9387 484 9388 524
rect 9428 484 9429 524
rect 9387 475 9429 484
rect 9484 80 9524 1147
rect 9579 1112 9621 1121
rect 9579 1072 9580 1112
rect 9620 1072 9621 1112
rect 9579 1063 9621 1072
rect 9580 978 9620 1063
rect 9676 80 9716 1240
rect 9868 80 9908 2239
rect 10252 2045 10292 2407
rect 10251 2036 10293 2045
rect 10251 1996 10252 2036
rect 10292 1996 10293 2036
rect 10251 1987 10293 1996
rect 9964 1952 10004 1961
rect 9964 1037 10004 1912
rect 10060 1952 10100 1963
rect 10060 1877 10100 1912
rect 10059 1868 10101 1877
rect 10059 1828 10060 1868
rect 10100 1828 10101 1868
rect 10059 1819 10101 1828
rect 10348 1280 10388 2416
rect 10539 2456 10581 2465
rect 10539 2416 10540 2456
rect 10580 2416 10581 2456
rect 10539 2407 10581 2416
rect 10540 1952 10580 2407
rect 10540 1903 10580 1912
rect 10444 1868 10484 1877
rect 10444 1784 10484 1828
rect 10444 1744 10580 1784
rect 10443 1616 10485 1625
rect 10443 1576 10444 1616
rect 10484 1576 10485 1616
rect 10443 1567 10485 1576
rect 10060 1240 10388 1280
rect 9963 1028 10005 1037
rect 9963 988 9964 1028
rect 10004 988 10005 1028
rect 9963 979 10005 988
rect 10060 80 10100 1240
rect 10251 860 10293 869
rect 10251 820 10252 860
rect 10292 820 10293 860
rect 10251 811 10293 820
rect 10252 80 10292 811
rect 10444 80 10484 1567
rect 10540 1541 10580 1744
rect 10539 1532 10581 1541
rect 10539 1492 10540 1532
rect 10580 1492 10581 1532
rect 10539 1483 10581 1492
rect 10539 1280 10581 1289
rect 10539 1240 10540 1280
rect 10580 1240 10581 1280
rect 10539 1231 10581 1240
rect 10540 860 10580 1231
rect 10636 944 10676 2491
rect 10828 2213 10868 2584
rect 10923 2624 10965 2633
rect 10923 2584 10924 2624
rect 10964 2584 10965 2624
rect 10923 2575 10965 2584
rect 10827 2204 10869 2213
rect 10827 2164 10828 2204
rect 10868 2164 10869 2204
rect 10827 2155 10869 2164
rect 10924 1877 10964 2575
rect 11019 2540 11061 2549
rect 11019 2500 11020 2540
rect 11060 2500 11061 2540
rect 11019 2491 11061 2500
rect 11020 1952 11060 2491
rect 11020 1903 11060 1912
rect 10923 1868 10965 1877
rect 10923 1828 10924 1868
rect 10964 1828 10965 1868
rect 10923 1819 10965 1828
rect 11020 1280 11060 1289
rect 11116 1280 11156 2659
rect 11308 2624 11348 2633
rect 11308 2213 11348 2584
rect 11404 2465 11444 2668
rect 11403 2456 11445 2465
rect 11403 2416 11404 2456
rect 11444 2416 11445 2456
rect 11403 2407 11445 2416
rect 11500 2381 11540 3415
rect 11595 2456 11637 2465
rect 11595 2416 11596 2456
rect 11636 2416 11637 2456
rect 11595 2407 11637 2416
rect 11499 2372 11541 2381
rect 11499 2332 11500 2372
rect 11540 2332 11541 2372
rect 11499 2323 11541 2332
rect 11307 2204 11349 2213
rect 11307 2164 11308 2204
rect 11348 2164 11349 2204
rect 11307 2155 11349 2164
rect 11500 1938 11540 1947
rect 11211 1868 11253 1877
rect 11211 1828 11212 1868
rect 11252 1828 11253 1868
rect 11211 1819 11253 1828
rect 11212 1289 11252 1819
rect 11060 1240 11156 1280
rect 11211 1280 11253 1289
rect 11211 1240 11212 1280
rect 11252 1240 11253 1280
rect 11020 1231 11060 1240
rect 11211 1231 11253 1240
rect 11500 1205 11540 1898
rect 11499 1196 11541 1205
rect 11499 1156 11500 1196
rect 11540 1156 11541 1196
rect 11499 1147 11541 1156
rect 10828 1112 10868 1121
rect 11211 1112 11253 1121
rect 10868 1072 11156 1112
rect 10828 1063 10868 1072
rect 10636 904 10868 944
rect 10540 820 10676 860
rect 10636 80 10676 820
rect 10828 80 10868 904
rect 11116 869 11156 1072
rect 11211 1072 11212 1112
rect 11252 1072 11348 1112
rect 11211 1063 11253 1072
rect 11212 978 11252 1063
rect 10923 860 10965 869
rect 11115 860 11157 869
rect 10923 820 10924 860
rect 10964 820 11060 860
rect 10923 811 10965 820
rect 11020 80 11060 820
rect 11115 820 11116 860
rect 11156 820 11157 860
rect 11115 811 11157 820
rect 11116 533 11156 811
rect 11211 608 11253 617
rect 11211 568 11212 608
rect 11252 568 11253 608
rect 11211 559 11253 568
rect 11115 524 11157 533
rect 11115 484 11116 524
rect 11156 484 11157 524
rect 11115 475 11157 484
rect 11212 80 11252 559
rect 11308 197 11348 1072
rect 11403 860 11445 869
rect 11403 820 11404 860
rect 11444 820 11445 860
rect 11403 811 11445 820
rect 11307 188 11349 197
rect 11307 148 11308 188
rect 11348 148 11349 188
rect 11307 139 11349 148
rect 11404 80 11444 811
rect 11596 80 11636 2407
rect 11692 2297 11732 6280
rect 11883 6236 11925 6245
rect 11883 6196 11884 6236
rect 11924 6196 11925 6236
rect 11883 6187 11925 6196
rect 11788 5657 11828 5742
rect 11787 5648 11829 5657
rect 11787 5608 11788 5648
rect 11828 5608 11829 5648
rect 11787 5599 11829 5608
rect 11884 5396 11924 6187
rect 11788 5356 11924 5396
rect 11788 5153 11828 5356
rect 11883 5228 11925 5237
rect 11883 5188 11884 5228
rect 11924 5188 11925 5228
rect 11980 5228 12020 7447
rect 12075 6656 12117 6665
rect 12075 6616 12076 6656
rect 12116 6616 12117 6656
rect 12075 6607 12117 6616
rect 12076 6522 12116 6607
rect 11980 5188 12116 5228
rect 11883 5179 11925 5188
rect 11787 5144 11829 5153
rect 11787 5104 11788 5144
rect 11828 5104 11829 5144
rect 11787 5095 11829 5104
rect 11788 4052 11828 5095
rect 11884 4976 11924 5179
rect 11980 4985 12020 5070
rect 11884 4927 11924 4936
rect 11979 4976 12021 4985
rect 11979 4936 11980 4976
rect 12020 4936 12021 4976
rect 11979 4927 12021 4936
rect 12076 4808 12116 5188
rect 11884 4768 12116 4808
rect 11884 4220 11924 4768
rect 11884 4171 11924 4180
rect 11980 4136 12020 4145
rect 11980 4052 12020 4096
rect 11788 4012 12020 4052
rect 12172 3893 12212 7708
rect 12268 7708 12364 7748
rect 12268 7160 12308 7708
rect 12364 7699 12404 7708
rect 12268 7111 12308 7120
rect 12364 7160 12404 7169
rect 12268 6404 12308 6413
rect 12268 5909 12308 6364
rect 12267 5900 12309 5909
rect 12267 5860 12268 5900
rect 12308 5860 12309 5900
rect 12267 5851 12309 5860
rect 12364 5741 12404 7120
rect 12460 6488 12500 9052
rect 12556 9017 12596 10816
rect 13036 10781 13076 10984
rect 13132 10974 13172 11059
rect 13324 10949 13364 11068
rect 13323 10940 13365 10949
rect 13323 10900 13324 10940
rect 13364 10900 13365 10940
rect 13323 10891 13365 10900
rect 13035 10772 13077 10781
rect 13035 10732 13036 10772
rect 13076 10732 13077 10772
rect 13035 10723 13077 10732
rect 12939 10604 12981 10613
rect 12939 10564 12940 10604
rect 12980 10564 12981 10604
rect 12939 10555 12981 10564
rect 12748 10352 12788 10361
rect 12652 10312 12748 10352
rect 12555 9008 12597 9017
rect 12555 8968 12556 9008
rect 12596 8968 12597 9008
rect 12555 8959 12597 8968
rect 12556 8840 12596 8849
rect 12556 8597 12596 8800
rect 12555 8588 12597 8597
rect 12555 8548 12556 8588
rect 12596 8548 12597 8588
rect 12555 8539 12597 8548
rect 12555 8168 12597 8177
rect 12555 8128 12556 8168
rect 12596 8128 12597 8168
rect 12555 8119 12597 8128
rect 12556 8034 12596 8119
rect 12652 8000 12692 10312
rect 12748 10303 12788 10312
rect 12940 10184 12980 10555
rect 12844 10144 12940 10184
rect 12747 10100 12789 10109
rect 12747 10060 12748 10100
rect 12788 10060 12789 10100
rect 12747 10051 12789 10060
rect 12748 9512 12788 10051
rect 12748 9463 12788 9472
rect 12748 8672 12788 8683
rect 12748 8597 12788 8632
rect 12844 8672 12884 10144
rect 12940 10135 12980 10144
rect 13131 10184 13173 10193
rect 13131 10144 13132 10184
rect 13172 10144 13173 10184
rect 13131 10135 13173 10144
rect 13228 10184 13268 10193
rect 13132 10050 13172 10135
rect 13228 10025 13268 10144
rect 13420 10184 13460 11983
rect 13708 11710 13748 12235
rect 13995 12200 14037 12209
rect 13995 12160 13996 12200
rect 14036 12160 14037 12200
rect 13995 12151 14037 12160
rect 13708 11661 13748 11670
rect 13803 11612 13845 11621
rect 13803 11572 13804 11612
rect 13844 11572 13845 11612
rect 13803 11563 13845 11572
rect 13420 10135 13460 10144
rect 13516 11010 13556 11019
rect 13036 10016 13076 10025
rect 12940 9260 12980 9269
rect 12940 8672 12980 9220
rect 13036 9101 13076 9976
rect 13227 10016 13269 10025
rect 13227 9976 13228 10016
rect 13268 9976 13269 10016
rect 13227 9967 13269 9976
rect 13324 9680 13364 9689
rect 13516 9680 13556 10970
rect 13707 10688 13749 10697
rect 13707 10648 13708 10688
rect 13748 10648 13749 10688
rect 13707 10639 13749 10648
rect 13611 10016 13653 10025
rect 13611 9976 13612 10016
rect 13652 9976 13653 10016
rect 13611 9967 13653 9976
rect 13364 9640 13556 9680
rect 13324 9631 13364 9640
rect 13323 9512 13365 9521
rect 13323 9472 13324 9512
rect 13364 9472 13365 9512
rect 13323 9463 13365 9472
rect 13515 9512 13557 9521
rect 13515 9472 13516 9512
rect 13556 9472 13557 9512
rect 13515 9463 13557 9472
rect 13035 9092 13077 9101
rect 13035 9052 13036 9092
rect 13076 9052 13077 9092
rect 13035 9043 13077 9052
rect 13036 8849 13076 8934
rect 13035 8840 13077 8849
rect 13035 8800 13036 8840
rect 13076 8800 13077 8840
rect 13035 8791 13077 8800
rect 13036 8672 13076 8681
rect 12940 8632 13036 8672
rect 12747 8588 12789 8597
rect 12747 8548 12748 8588
rect 12788 8548 12789 8588
rect 12747 8539 12789 8548
rect 12844 8009 12884 8632
rect 12748 8000 12788 8009
rect 12652 7960 12748 8000
rect 12748 7951 12788 7960
rect 12843 8000 12885 8009
rect 12843 7960 12844 8000
rect 12884 7960 12885 8000
rect 12843 7951 12885 7960
rect 13036 8000 13076 8632
rect 13131 8672 13173 8681
rect 13131 8632 13132 8672
rect 13172 8632 13173 8672
rect 13131 8623 13173 8632
rect 13132 8168 13172 8623
rect 13227 8504 13269 8513
rect 13227 8464 13228 8504
rect 13268 8464 13269 8504
rect 13227 8455 13269 8464
rect 13228 8370 13268 8455
rect 13324 8261 13364 9463
rect 13516 9378 13556 9463
rect 13515 9008 13557 9017
rect 13515 8968 13516 9008
rect 13556 8968 13557 9008
rect 13515 8959 13557 8968
rect 13419 8756 13461 8765
rect 13419 8716 13420 8756
rect 13460 8716 13461 8756
rect 13419 8707 13461 8716
rect 13420 8622 13460 8707
rect 13323 8252 13365 8261
rect 13323 8212 13324 8252
rect 13364 8212 13365 8252
rect 13323 8203 13365 8212
rect 13132 8119 13172 8128
rect 13227 8168 13269 8177
rect 13227 8128 13228 8168
rect 13268 8128 13269 8168
rect 13227 8119 13269 8128
rect 13036 7951 13076 7960
rect 12555 7916 12597 7925
rect 12555 7876 12556 7916
rect 12596 7876 12597 7916
rect 12555 7867 12597 7876
rect 12363 5732 12405 5741
rect 12363 5692 12364 5732
rect 12404 5692 12405 5732
rect 12363 5683 12405 5692
rect 12460 5657 12500 6448
rect 12459 5648 12501 5657
rect 12459 5608 12460 5648
rect 12500 5608 12501 5648
rect 12459 5599 12501 5608
rect 12556 5480 12596 7867
rect 12844 7866 12884 7951
rect 12747 7328 12789 7337
rect 12747 7288 12748 7328
rect 12788 7288 12789 7328
rect 12747 7279 12789 7288
rect 12748 7244 12788 7279
rect 12748 7193 12788 7204
rect 12844 7160 12884 7169
rect 13228 7160 13268 8119
rect 13323 8000 13365 8009
rect 13323 7960 13324 8000
rect 13364 7960 13365 8000
rect 13323 7951 13365 7960
rect 13324 7866 13364 7951
rect 13516 7337 13556 8959
rect 13612 8672 13652 9967
rect 13708 9521 13748 10639
rect 13707 9512 13749 9521
rect 13707 9472 13708 9512
rect 13748 9472 13749 9512
rect 13707 9463 13749 9472
rect 13804 9269 13844 11563
rect 13900 11528 13940 11537
rect 13900 11285 13940 11488
rect 13899 11276 13941 11285
rect 13899 11236 13900 11276
rect 13940 11236 13941 11276
rect 13899 11227 13941 11236
rect 13996 11024 14036 12151
rect 14092 12041 14132 12487
rect 14187 12284 14229 12293
rect 14187 12244 14188 12284
rect 14228 12244 14229 12284
rect 14187 12235 14229 12244
rect 14188 12150 14228 12235
rect 14091 12032 14133 12041
rect 14284 12032 14324 18880
rect 14380 18173 14420 18964
rect 14379 18164 14421 18173
rect 14379 18124 14380 18164
rect 14420 18124 14421 18164
rect 14379 18115 14421 18124
rect 14379 17912 14421 17921
rect 14379 17872 14380 17912
rect 14420 17872 14421 17912
rect 14379 17863 14421 17872
rect 14380 16325 14420 17863
rect 14379 16316 14421 16325
rect 14379 16276 14380 16316
rect 14420 16276 14421 16316
rect 14379 16267 14421 16276
rect 14380 14141 14420 14226
rect 14379 14132 14421 14141
rect 14379 14092 14380 14132
rect 14420 14092 14421 14132
rect 14379 14083 14421 14092
rect 14476 14048 14516 20215
rect 14572 17921 14612 20644
rect 14667 20644 14668 20684
rect 14708 20644 14709 20684
rect 14667 20635 14709 20644
rect 14668 18845 14708 20635
rect 14764 20021 14804 21568
rect 15052 21524 15092 22996
rect 15148 23036 15188 23752
rect 15188 22996 15284 23036
rect 15148 22987 15188 22996
rect 15147 21524 15189 21533
rect 15052 21484 15148 21524
rect 15188 21484 15189 21524
rect 15147 21475 15189 21484
rect 15244 21524 15284 22996
rect 15148 21390 15188 21475
rect 14859 21020 14901 21029
rect 14859 20980 14860 21020
rect 14900 20980 14901 21020
rect 14859 20971 14901 20980
rect 14860 20886 14900 20971
rect 14763 20012 14805 20021
rect 14763 19972 14764 20012
rect 14804 19972 14805 20012
rect 14763 19963 14805 19972
rect 15244 19853 15284 21484
rect 14859 19844 14901 19853
rect 14859 19804 14860 19844
rect 14900 19804 14901 19844
rect 14859 19795 14901 19804
rect 15243 19844 15285 19853
rect 15243 19804 15244 19844
rect 15284 19804 15285 19844
rect 15243 19795 15285 19804
rect 14860 19270 14900 19795
rect 14860 19221 14900 19230
rect 15243 19256 15285 19265
rect 15243 19216 15244 19256
rect 15284 19216 15285 19256
rect 15243 19207 15285 19216
rect 15244 19122 15284 19207
rect 14859 19088 14901 19097
rect 14859 19048 14860 19088
rect 14900 19048 14901 19088
rect 14859 19039 14901 19048
rect 15051 19088 15093 19097
rect 15051 19048 15052 19088
rect 15092 19048 15093 19088
rect 15051 19039 15093 19048
rect 14667 18836 14709 18845
rect 14667 18796 14668 18836
rect 14708 18796 14709 18836
rect 14667 18787 14709 18796
rect 14764 18500 14804 18509
rect 14764 18173 14804 18460
rect 14763 18164 14805 18173
rect 14763 18124 14764 18164
rect 14804 18124 14805 18164
rect 14763 18115 14805 18124
rect 14571 17912 14613 17921
rect 14571 17872 14572 17912
rect 14612 17872 14613 17912
rect 14571 17863 14613 17872
rect 14763 17828 14805 17837
rect 14763 17788 14764 17828
rect 14804 17788 14805 17828
rect 14763 17779 14805 17788
rect 14620 17753 14660 17762
rect 14660 17713 14708 17744
rect 14620 17704 14708 17713
rect 14668 17240 14708 17704
rect 14764 17660 14804 17779
rect 14860 17753 14900 19039
rect 15052 18954 15092 19039
rect 14955 18920 14997 18929
rect 14955 18880 14956 18920
rect 14996 18880 14997 18920
rect 14955 18871 14997 18880
rect 15147 18920 15189 18929
rect 15147 18880 15148 18920
rect 15188 18880 15189 18920
rect 15147 18871 15189 18880
rect 14956 18752 14996 18871
rect 14956 18703 14996 18712
rect 15148 18584 15188 18871
rect 15340 18752 15380 25096
rect 15532 23792 15572 23801
rect 15532 23120 15572 23752
rect 15724 23213 15764 25936
rect 15820 25304 15860 26011
rect 15820 25255 15860 25264
rect 15819 25136 15861 25145
rect 15819 25096 15820 25136
rect 15860 25096 15861 25136
rect 15819 25087 15861 25096
rect 15820 23381 15860 25087
rect 15819 23372 15861 23381
rect 15819 23332 15820 23372
rect 15860 23332 15861 23372
rect 15819 23323 15861 23332
rect 15723 23204 15765 23213
rect 15723 23164 15724 23204
rect 15764 23164 15765 23204
rect 15723 23155 15765 23164
rect 15628 23120 15668 23148
rect 15532 23080 15628 23120
rect 15532 22625 15572 23080
rect 15628 23071 15668 23080
rect 15627 22700 15669 22709
rect 15627 22660 15628 22700
rect 15668 22660 15669 22700
rect 15627 22651 15669 22660
rect 15531 22616 15573 22625
rect 15531 22576 15532 22616
rect 15572 22576 15573 22616
rect 15531 22567 15573 22576
rect 15628 21020 15668 22651
rect 15723 22616 15765 22625
rect 15723 22576 15724 22616
rect 15764 22576 15765 22616
rect 15723 22567 15765 22576
rect 15724 21608 15764 22567
rect 15724 21559 15764 21568
rect 15819 21272 15861 21281
rect 15819 21232 15820 21272
rect 15860 21232 15861 21272
rect 15819 21223 15861 21232
rect 15628 20971 15668 20980
rect 15436 20852 15476 20861
rect 15436 20021 15476 20812
rect 15820 20768 15860 21223
rect 15820 20719 15860 20728
rect 15916 20180 15956 27280
rect 16012 27161 16052 27616
rect 16108 27572 16148 27784
rect 16108 27523 16148 27532
rect 16204 27488 16244 28111
rect 16300 27833 16340 30556
rect 16396 30269 16436 30724
rect 16395 30260 16437 30269
rect 16395 30220 16396 30260
rect 16436 30220 16437 30260
rect 16395 30211 16437 30220
rect 16684 29261 16724 30808
rect 16780 30680 16820 30691
rect 16780 30605 16820 30640
rect 16779 30596 16821 30605
rect 16779 30556 16780 30596
rect 16820 30556 16821 30596
rect 16779 30547 16821 30556
rect 16779 29336 16821 29345
rect 16779 29296 16780 29336
rect 16820 29296 16821 29336
rect 16779 29287 16821 29296
rect 16491 29252 16533 29261
rect 16491 29212 16492 29252
rect 16532 29212 16533 29252
rect 16491 29203 16533 29212
rect 16683 29252 16725 29261
rect 16683 29212 16684 29252
rect 16724 29212 16725 29252
rect 16683 29203 16725 29212
rect 16395 29168 16437 29177
rect 16395 29128 16396 29168
rect 16436 29128 16437 29168
rect 16395 29119 16437 29128
rect 16396 29034 16436 29119
rect 16492 29084 16532 29203
rect 16780 29168 16820 29287
rect 16780 29119 16820 29128
rect 16492 29035 16532 29044
rect 16684 29084 16724 29093
rect 16587 29000 16629 29009
rect 16587 28960 16588 29000
rect 16628 28960 16629 29000
rect 16587 28951 16629 28960
rect 16588 28866 16628 28951
rect 16395 28328 16437 28337
rect 16395 28288 16396 28328
rect 16436 28288 16437 28328
rect 16395 28279 16437 28288
rect 16299 27824 16341 27833
rect 16299 27784 16300 27824
rect 16340 27784 16341 27824
rect 16299 27775 16341 27784
rect 16300 27665 16340 27696
rect 16299 27656 16341 27665
rect 16299 27616 16300 27656
rect 16340 27616 16341 27656
rect 16299 27607 16341 27616
rect 16396 27656 16436 28279
rect 16684 28169 16724 29044
rect 16683 28160 16725 28169
rect 16683 28120 16684 28160
rect 16724 28120 16725 28160
rect 16683 28111 16725 28120
rect 16588 27665 16628 27750
rect 16876 27749 16916 32815
rect 16972 32201 17012 33664
rect 17068 33032 17108 34588
rect 17260 33293 17300 36352
rect 17356 35981 17396 36643
rect 17451 36646 17452 36653
rect 17548 36679 17588 36688
rect 17932 36728 17972 36763
rect 17492 36646 17493 36653
rect 17451 36644 17493 36646
rect 17451 36604 17452 36644
rect 17492 36604 17493 36644
rect 17451 36595 17493 36604
rect 17452 36551 17492 36595
rect 17932 36140 17972 36688
rect 18220 36728 18260 36737
rect 18028 36140 18068 36149
rect 17932 36100 18028 36140
rect 18028 36091 18068 36100
rect 18220 36056 18260 36688
rect 18220 36016 18356 36056
rect 17355 35972 17397 35981
rect 17355 35932 17356 35972
rect 17396 35932 17397 35972
rect 17355 35923 17397 35932
rect 17836 35888 17876 35897
rect 18220 35888 18260 35897
rect 17451 35552 17493 35561
rect 17451 35512 17452 35552
rect 17492 35512 17684 35552
rect 17451 35503 17493 35512
rect 17355 35384 17397 35393
rect 17355 35344 17356 35384
rect 17396 35344 17397 35384
rect 17355 35335 17397 35344
rect 17356 35216 17396 35335
rect 17356 35167 17396 35176
rect 17451 35216 17493 35225
rect 17451 35176 17452 35216
rect 17492 35176 17493 35216
rect 17451 35167 17493 35176
rect 17644 35216 17684 35512
rect 17836 35477 17876 35848
rect 18124 35848 18220 35888
rect 18028 35720 18068 35731
rect 18028 35645 18068 35680
rect 18027 35636 18069 35645
rect 18027 35596 18028 35636
rect 18068 35596 18069 35636
rect 18027 35587 18069 35596
rect 17835 35468 17877 35477
rect 17835 35428 17836 35468
rect 17876 35428 17877 35468
rect 17835 35419 17877 35428
rect 18027 35300 18069 35309
rect 17740 35225 17780 35269
rect 17836 35258 17876 35267
rect 17644 35167 17684 35176
rect 17739 35216 17781 35225
rect 17739 35176 17740 35216
rect 17780 35176 17781 35216
rect 17739 35174 17781 35176
rect 17739 35167 17740 35174
rect 17452 35082 17492 35167
rect 17780 35167 17781 35174
rect 18027 35260 18028 35300
rect 18068 35260 18069 35300
rect 18027 35251 18069 35260
rect 17740 35125 17780 35134
rect 17836 35132 17876 35218
rect 18028 35216 18068 35251
rect 18028 35165 18068 35176
rect 17931 35132 17973 35141
rect 17836 35092 17877 35132
rect 17355 34964 17397 34973
rect 17837 34964 17877 35092
rect 17931 35092 17932 35132
rect 17972 35092 17973 35132
rect 17931 35083 17973 35092
rect 17932 34998 17972 35083
rect 17355 34924 17356 34964
rect 17396 34924 17397 34964
rect 17355 34915 17397 34924
rect 17836 34924 17877 34964
rect 17259 33284 17301 33293
rect 17259 33244 17260 33284
rect 17300 33244 17301 33284
rect 17259 33235 17301 33244
rect 17259 33032 17301 33041
rect 17068 32992 17204 33032
rect 17068 32864 17108 32875
rect 17068 32789 17108 32824
rect 17067 32780 17109 32789
rect 17067 32740 17068 32780
rect 17108 32740 17109 32780
rect 17067 32731 17109 32740
rect 16971 32192 17013 32201
rect 16971 32152 16972 32192
rect 17012 32152 17013 32192
rect 16971 32143 17013 32152
rect 17067 31772 17109 31781
rect 17067 31732 17068 31772
rect 17108 31732 17109 31772
rect 17067 31723 17109 31732
rect 17068 31352 17108 31723
rect 17068 31303 17108 31312
rect 16972 31268 17012 31277
rect 16972 29588 17012 31228
rect 17164 31025 17204 32992
rect 17259 32992 17260 33032
rect 17300 32992 17301 33032
rect 17259 32983 17301 32992
rect 17260 32898 17300 32983
rect 17356 31352 17396 34915
rect 17643 34628 17685 34637
rect 17643 34588 17644 34628
rect 17684 34588 17685 34628
rect 17643 34579 17685 34588
rect 17644 34494 17684 34579
rect 17451 34376 17493 34385
rect 17451 34336 17452 34376
rect 17492 34336 17493 34376
rect 17451 34327 17493 34336
rect 17452 32201 17492 34327
rect 17836 34133 17876 34924
rect 17931 34880 17973 34889
rect 17931 34840 17932 34880
rect 17972 34840 17973 34880
rect 17931 34831 17973 34840
rect 17835 34124 17877 34133
rect 17835 34084 17836 34124
rect 17876 34084 17877 34124
rect 17835 34075 17877 34084
rect 17932 33872 17972 34831
rect 18027 34628 18069 34637
rect 18027 34588 18028 34628
rect 18068 34588 18069 34628
rect 18027 34579 18069 34588
rect 18028 34376 18068 34579
rect 18028 34327 18068 34336
rect 18027 34040 18069 34049
rect 18027 34000 18028 34040
rect 18068 34000 18069 34040
rect 18027 33991 18069 34000
rect 17644 33832 17972 33872
rect 17644 32864 17684 33832
rect 17835 33704 17877 33713
rect 17835 33664 17836 33704
rect 17876 33664 17877 33704
rect 17835 33655 17877 33664
rect 17644 32360 17684 32824
rect 17836 32789 17876 33655
rect 17931 33116 17973 33125
rect 17931 33076 17932 33116
rect 17972 33076 17973 33116
rect 17931 33067 17973 33076
rect 17932 32864 17972 33067
rect 18028 32957 18068 33991
rect 18124 33881 18164 35848
rect 18220 35839 18260 35848
rect 18316 35309 18356 36016
rect 18315 35300 18357 35309
rect 18315 35260 18316 35300
rect 18356 35260 18357 35300
rect 18315 35251 18357 35260
rect 18220 35216 18260 35225
rect 18123 33872 18165 33881
rect 18123 33832 18124 33872
rect 18164 33832 18165 33872
rect 18123 33823 18165 33832
rect 18124 33704 18164 33715
rect 18124 33629 18164 33664
rect 18123 33620 18165 33629
rect 18123 33580 18124 33620
rect 18164 33580 18165 33620
rect 18123 33571 18165 33580
rect 18027 32948 18069 32957
rect 18027 32908 18028 32948
rect 18068 32908 18069 32948
rect 18027 32899 18069 32908
rect 17932 32815 17972 32824
rect 18028 32864 18068 32899
rect 18028 32813 18068 32824
rect 17835 32780 17877 32789
rect 17835 32740 17836 32780
rect 17876 32740 17877 32780
rect 17835 32731 17877 32740
rect 18124 32537 18164 33571
rect 18123 32528 18165 32537
rect 18123 32488 18124 32528
rect 18164 32488 18165 32528
rect 18123 32479 18165 32488
rect 18220 32360 18260 35176
rect 18315 34964 18357 34973
rect 18315 34924 18316 34964
rect 18356 34924 18357 34964
rect 18315 34915 18357 34924
rect 18316 34830 18356 34915
rect 18412 34553 18452 37780
rect 18508 35384 18548 38200
rect 18603 38200 18604 38240
rect 18644 38200 18645 38240
rect 18603 38191 18645 38200
rect 18604 37400 18644 38191
rect 18604 36896 18644 37360
rect 18700 37325 18740 38872
rect 18796 38863 18836 38872
rect 18987 38912 19029 38921
rect 18987 38872 18988 38912
rect 19028 38872 19029 38912
rect 18987 38863 19029 38872
rect 19084 38828 19124 38947
rect 19372 38828 19412 38956
rect 19467 38912 19509 38921
rect 19467 38872 19468 38912
rect 19508 38872 19509 38912
rect 19467 38863 19509 38872
rect 19084 38788 19412 38828
rect 18892 38744 18932 38753
rect 18892 38417 18932 38704
rect 19468 38417 19508 38863
rect 19563 38744 19605 38753
rect 19563 38704 19564 38744
rect 19604 38704 19605 38744
rect 19563 38695 19605 38704
rect 19564 38610 19604 38695
rect 19756 38669 19796 39460
rect 19852 39164 19892 40888
rect 19947 40760 19989 40769
rect 19947 40720 19948 40760
rect 19988 40720 19989 40760
rect 19947 40711 19989 40720
rect 19948 40676 19988 40711
rect 19948 40625 19988 40636
rect 20120 40508 20162 40517
rect 20120 40468 20121 40508
rect 20161 40468 20162 40508
rect 20120 40459 20162 40468
rect 20121 40374 20161 40459
rect 20048 40088 20416 40097
rect 20088 40048 20130 40088
rect 20170 40048 20212 40088
rect 20252 40048 20294 40088
rect 20334 40048 20376 40088
rect 20048 40039 20416 40048
rect 19947 39752 19989 39761
rect 19947 39712 19948 39752
rect 19988 39712 19989 39752
rect 19947 39703 19989 39712
rect 20140 39739 20180 39748
rect 19948 39618 19988 39703
rect 20044 39668 20084 39677
rect 19852 39124 19988 39164
rect 19852 38996 19892 39005
rect 19755 38660 19797 38669
rect 19755 38620 19756 38660
rect 19796 38620 19797 38660
rect 19755 38611 19797 38620
rect 19852 38585 19892 38956
rect 19948 38753 19988 39124
rect 20044 39005 20084 39628
rect 20140 39257 20180 39699
rect 20811 39584 20853 39593
rect 20811 39544 20812 39584
rect 20852 39544 20853 39584
rect 20811 39535 20853 39544
rect 20715 39416 20757 39425
rect 20715 39376 20716 39416
rect 20756 39376 20757 39416
rect 20715 39367 20757 39376
rect 20139 39248 20181 39257
rect 20139 39208 20140 39248
rect 20180 39208 20181 39248
rect 20139 39199 20181 39208
rect 20043 38996 20085 39005
rect 20043 38956 20044 38996
rect 20084 38956 20085 38996
rect 20043 38947 20085 38956
rect 20619 38996 20661 39005
rect 20619 38956 20620 38996
rect 20660 38956 20661 38996
rect 20619 38947 20661 38956
rect 20044 38753 20084 38838
rect 19942 38744 19988 38753
rect 19942 38704 19943 38744
rect 19983 38704 19988 38744
rect 20043 38744 20085 38753
rect 20043 38704 20044 38744
rect 20084 38704 20085 38744
rect 19942 38695 19984 38704
rect 20043 38695 20085 38704
rect 19851 38576 19893 38585
rect 19851 38536 19852 38576
rect 19892 38536 19893 38576
rect 19851 38527 19893 38536
rect 20048 38576 20416 38585
rect 20088 38536 20130 38576
rect 20170 38536 20212 38576
rect 20252 38536 20294 38576
rect 20334 38536 20376 38576
rect 20048 38527 20416 38536
rect 18891 38408 18933 38417
rect 18891 38368 18892 38408
rect 18932 38368 18933 38408
rect 18891 38359 18933 38368
rect 19275 38408 19317 38417
rect 19275 38368 19276 38408
rect 19316 38368 19317 38408
rect 19275 38359 19317 38368
rect 19467 38408 19509 38417
rect 19467 38368 19468 38408
rect 19508 38368 19509 38408
rect 19467 38359 19509 38368
rect 20235 38408 20277 38417
rect 20235 38368 20236 38408
rect 20276 38368 20277 38408
rect 20235 38359 20277 38368
rect 19083 38324 19125 38333
rect 19083 38284 19084 38324
rect 19124 38284 19125 38324
rect 19083 38275 19125 38284
rect 18891 38240 18933 38249
rect 18891 38200 18892 38240
rect 18932 38200 18933 38240
rect 18891 38191 18933 38200
rect 18892 38106 18932 38191
rect 19084 38190 19124 38275
rect 19276 37829 19316 38359
rect 20139 38324 20181 38333
rect 20139 38284 20140 38324
rect 20180 38284 20181 38324
rect 20139 38275 20181 38284
rect 20140 38261 20180 38275
rect 20236 38274 20276 38359
rect 20523 38324 20565 38333
rect 20523 38284 20524 38324
rect 20564 38284 20565 38324
rect 20523 38275 20565 38284
rect 19467 38240 19509 38249
rect 19467 38200 19468 38240
rect 19508 38200 19509 38240
rect 19467 38191 19509 38200
rect 19564 38240 19604 38249
rect 19468 38106 19508 38191
rect 19564 37997 19604 38200
rect 19756 38240 19796 38249
rect 19948 38240 19988 38249
rect 19796 38200 19948 38240
rect 19756 38191 19796 38200
rect 19563 37988 19605 37997
rect 19756 37988 19796 37997
rect 19563 37948 19564 37988
rect 19604 37948 19605 37988
rect 19563 37939 19605 37948
rect 19660 37948 19756 37988
rect 18808 37820 19176 37829
rect 18848 37780 18890 37820
rect 18930 37780 18972 37820
rect 19012 37780 19054 37820
rect 19094 37780 19136 37820
rect 18808 37771 19176 37780
rect 19275 37820 19317 37829
rect 19275 37780 19276 37820
rect 19316 37780 19317 37820
rect 19275 37771 19317 37780
rect 18795 37652 18837 37661
rect 18795 37612 18796 37652
rect 18836 37612 18837 37652
rect 18795 37603 18837 37612
rect 18796 37518 18836 37603
rect 18987 37568 19029 37577
rect 19660 37568 19700 37948
rect 19756 37939 19796 37948
rect 19851 37820 19893 37829
rect 19851 37780 19852 37820
rect 19892 37780 19893 37820
rect 19851 37771 19893 37780
rect 18987 37528 18988 37568
rect 19028 37528 19029 37568
rect 18987 37519 19029 37528
rect 19180 37528 19700 37568
rect 19852 37568 19892 37771
rect 19948 37745 19988 38200
rect 20043 38240 20085 38249
rect 20043 38200 20044 38240
rect 20084 38200 20085 38240
rect 20043 38191 20085 38200
rect 20044 38106 20084 38191
rect 20140 38189 20180 38221
rect 19947 37736 19989 37745
rect 19947 37696 19948 37736
rect 19988 37696 19989 37736
rect 19947 37687 19989 37696
rect 19852 37528 19988 37568
rect 18891 37400 18933 37409
rect 18891 37360 18892 37400
rect 18932 37360 18933 37400
rect 18891 37351 18933 37360
rect 18988 37400 19028 37519
rect 18988 37351 19028 37360
rect 19083 37400 19125 37409
rect 19083 37360 19084 37400
rect 19124 37360 19125 37400
rect 19083 37351 19125 37360
rect 19180 37400 19220 37528
rect 19180 37351 19220 37360
rect 19275 37400 19317 37409
rect 19275 37360 19276 37400
rect 19316 37360 19317 37400
rect 19275 37351 19317 37360
rect 19468 37400 19508 37409
rect 18699 37316 18741 37325
rect 18699 37276 18700 37316
rect 18740 37276 18741 37316
rect 18699 37267 18741 37276
rect 18796 37232 18836 37243
rect 18796 37157 18836 37192
rect 18795 37148 18837 37157
rect 18795 37108 18796 37148
rect 18836 37108 18837 37148
rect 18795 37099 18837 37108
rect 18604 36856 18740 36896
rect 18603 36728 18645 36737
rect 18603 36688 18604 36728
rect 18644 36688 18645 36728
rect 18603 36679 18645 36688
rect 18604 36560 18644 36679
rect 18604 36511 18644 36520
rect 18700 35477 18740 36856
rect 18796 36728 18836 36737
rect 18796 36569 18836 36688
rect 18892 36728 18932 37351
rect 19084 37266 19124 37351
rect 19276 37266 19316 37351
rect 18987 37232 19029 37241
rect 18987 37192 18988 37232
rect 19028 37192 19029 37232
rect 18987 37183 19029 37192
rect 18892 36653 18932 36688
rect 18988 36728 19028 37183
rect 19083 36980 19125 36989
rect 19083 36940 19084 36980
rect 19124 36940 19125 36980
rect 19083 36931 19125 36940
rect 19084 36896 19124 36931
rect 19468 36905 19508 37360
rect 19660 37400 19700 37409
rect 19563 37316 19605 37325
rect 19563 37276 19564 37316
rect 19604 37276 19605 37316
rect 19563 37267 19605 37276
rect 19564 37182 19604 37267
rect 19563 36980 19605 36989
rect 19563 36940 19564 36980
rect 19604 36940 19605 36980
rect 19563 36931 19605 36940
rect 19084 36845 19124 36856
rect 19467 36896 19509 36905
rect 19467 36856 19468 36896
rect 19508 36856 19509 36896
rect 19467 36847 19509 36856
rect 19564 36896 19604 36931
rect 19564 36845 19604 36856
rect 19660 36821 19700 37360
rect 19756 37400 19796 37409
rect 19659 36812 19701 36821
rect 19659 36772 19660 36812
rect 19700 36772 19701 36812
rect 19659 36763 19701 36772
rect 18988 36679 19028 36688
rect 19276 36728 19316 36739
rect 19276 36653 19316 36688
rect 19372 36728 19412 36737
rect 18891 36644 18933 36653
rect 18891 36604 18892 36644
rect 18932 36604 18933 36644
rect 18891 36595 18933 36604
rect 19275 36644 19317 36653
rect 19275 36604 19276 36644
rect 19316 36604 19317 36644
rect 19275 36595 19317 36604
rect 18795 36560 18837 36569
rect 18795 36520 18796 36560
rect 18836 36520 18837 36560
rect 18795 36511 18837 36520
rect 19275 36392 19317 36401
rect 19275 36352 19276 36392
rect 19316 36352 19317 36392
rect 19275 36343 19317 36352
rect 18808 36308 19176 36317
rect 18848 36268 18890 36308
rect 18930 36268 18972 36308
rect 19012 36268 19054 36308
rect 19094 36268 19136 36308
rect 18808 36259 19176 36268
rect 19179 35888 19221 35897
rect 19179 35848 19180 35888
rect 19220 35848 19221 35888
rect 19179 35839 19221 35848
rect 19180 35754 19220 35839
rect 18699 35468 18741 35477
rect 18699 35428 18700 35468
rect 18740 35428 18741 35468
rect 18699 35419 18741 35428
rect 18508 35344 18644 35384
rect 18508 35216 18548 35225
rect 18508 34805 18548 35176
rect 18507 34796 18549 34805
rect 18507 34756 18508 34796
rect 18548 34756 18549 34796
rect 18507 34747 18549 34756
rect 18507 34628 18549 34637
rect 18507 34588 18508 34628
rect 18548 34588 18549 34628
rect 18507 34579 18549 34588
rect 18411 34544 18453 34553
rect 18411 34504 18412 34544
rect 18452 34504 18453 34544
rect 18411 34495 18453 34504
rect 18316 34376 18356 34385
rect 18316 34049 18356 34336
rect 18411 34292 18453 34301
rect 18411 34252 18412 34292
rect 18452 34252 18453 34292
rect 18411 34243 18453 34252
rect 18412 34158 18452 34243
rect 18315 34040 18357 34049
rect 18315 34000 18316 34040
rect 18356 34000 18357 34040
rect 18315 33991 18357 34000
rect 18412 33704 18452 33713
rect 18508 33704 18548 34579
rect 18452 33664 18548 33704
rect 18412 33655 18452 33664
rect 18604 33209 18644 35344
rect 18808 34796 19176 34805
rect 18848 34756 18890 34796
rect 18930 34756 18972 34796
rect 19012 34756 19054 34796
rect 19094 34756 19136 34796
rect 18808 34747 19176 34756
rect 18699 34544 18741 34553
rect 18699 34504 18700 34544
rect 18740 34504 18741 34544
rect 18699 34495 18741 34504
rect 18700 34410 18740 34495
rect 19083 34460 19125 34469
rect 19083 34420 19084 34460
rect 19124 34420 19125 34460
rect 19083 34411 19125 34420
rect 18983 34376 19023 34385
rect 19084 34376 19124 34411
rect 19276 34385 19316 36343
rect 19372 36233 19412 36688
rect 19468 36728 19508 36737
rect 19371 36224 19413 36233
rect 19371 36184 19372 36224
rect 19412 36184 19413 36224
rect 19468 36224 19508 36688
rect 19756 36485 19796 37360
rect 19948 37400 19988 37528
rect 20524 37484 20564 38275
rect 20620 37829 20660 38947
rect 20619 37820 20661 37829
rect 20619 37780 20620 37820
rect 20660 37780 20661 37820
rect 20619 37771 20661 37780
rect 20524 37444 20660 37484
rect 19948 37351 19988 37360
rect 20033 37400 20075 37409
rect 20236 37400 20276 37409
rect 20033 37360 20034 37400
rect 20074 37360 20084 37400
rect 20033 37351 20084 37360
rect 20044 37316 20084 37351
rect 20140 37358 20180 37367
rect 20044 37267 20084 37276
rect 20139 37318 20140 37325
rect 20276 37360 20564 37400
rect 20236 37351 20276 37360
rect 20180 37318 20181 37325
rect 20139 37316 20181 37318
rect 20139 37276 20140 37316
rect 20180 37276 20181 37316
rect 20139 37267 20181 37276
rect 20140 37223 20180 37267
rect 19947 37148 19989 37157
rect 19947 37108 19948 37148
rect 19988 37108 19989 37148
rect 19947 37099 19989 37108
rect 19948 36896 19988 37099
rect 20048 37064 20416 37073
rect 20088 37024 20130 37064
rect 20170 37024 20212 37064
rect 20252 37024 20294 37064
rect 20334 37024 20376 37064
rect 20048 37015 20416 37024
rect 20140 36896 20180 36905
rect 20524 36896 20564 37360
rect 19948 36856 20084 36896
rect 19947 36728 19989 36737
rect 19947 36688 19948 36728
rect 19988 36688 19989 36728
rect 19947 36679 19989 36688
rect 20044 36728 20084 36856
rect 20180 36856 20564 36896
rect 20140 36847 20180 36856
rect 20044 36679 20084 36688
rect 20139 36728 20181 36737
rect 20139 36688 20140 36728
rect 20180 36688 20181 36728
rect 20139 36679 20181 36688
rect 20236 36728 20276 36737
rect 20620 36728 20660 37444
rect 20276 36688 20660 36728
rect 20236 36679 20276 36688
rect 19948 36594 19988 36679
rect 20043 36560 20085 36569
rect 20043 36520 20044 36560
rect 20084 36520 20085 36560
rect 20043 36511 20085 36520
rect 19755 36476 19797 36485
rect 19755 36436 19756 36476
rect 19796 36436 19797 36476
rect 19755 36427 19797 36436
rect 19468 36184 19988 36224
rect 19371 36175 19413 36184
rect 19372 34889 19412 36175
rect 19948 36140 19988 36184
rect 19948 36091 19988 36100
rect 19468 35897 19508 35982
rect 20044 35972 20084 36511
rect 20140 36056 20180 36679
rect 20619 36140 20661 36149
rect 20619 36100 20620 36140
rect 20660 36100 20661 36140
rect 20619 36091 20661 36100
rect 20140 36007 20180 36016
rect 19948 35932 20084 35972
rect 19467 35888 19509 35897
rect 19467 35848 19468 35888
rect 19508 35848 19509 35888
rect 19467 35839 19509 35848
rect 19660 35888 19700 35897
rect 19468 35720 19508 35729
rect 19508 35680 19604 35720
rect 19468 35671 19508 35680
rect 19467 34964 19509 34973
rect 19467 34924 19468 34964
rect 19508 34924 19509 34964
rect 19467 34915 19509 34924
rect 19371 34880 19413 34889
rect 19371 34840 19372 34880
rect 19412 34840 19413 34880
rect 19371 34831 19413 34840
rect 19371 34712 19413 34721
rect 19371 34672 19372 34712
rect 19412 34672 19413 34712
rect 19371 34663 19413 34672
rect 19023 34336 19028 34376
rect 18983 34327 19028 34336
rect 18700 33704 18740 33713
rect 18700 33293 18740 33664
rect 18795 33704 18837 33713
rect 18795 33664 18796 33704
rect 18836 33664 18837 33704
rect 18795 33655 18837 33664
rect 18796 33570 18836 33655
rect 18988 33536 19028 34327
rect 19084 34325 19124 34336
rect 19180 34376 19220 34385
rect 19275 34376 19317 34385
rect 19220 34336 19276 34376
rect 19316 34336 19317 34376
rect 19180 34327 19220 34336
rect 19275 34327 19317 34336
rect 19372 34376 19412 34663
rect 19372 34327 19412 34336
rect 19468 34376 19508 34915
rect 19276 34208 19316 34217
rect 19468 34208 19508 34336
rect 19276 33704 19316 34168
rect 19276 33655 19316 33664
rect 19372 34168 19508 34208
rect 19564 34208 19604 35680
rect 19660 35561 19700 35848
rect 19756 35888 19796 35897
rect 19756 35645 19796 35848
rect 19851 35804 19893 35813
rect 19851 35764 19852 35804
rect 19892 35764 19893 35804
rect 19851 35755 19893 35764
rect 19755 35636 19797 35645
rect 19755 35596 19756 35636
rect 19796 35596 19797 35636
rect 19755 35587 19797 35596
rect 19659 35552 19701 35561
rect 19659 35512 19660 35552
rect 19700 35512 19701 35552
rect 19659 35503 19701 35512
rect 19755 35216 19797 35225
rect 19755 35176 19756 35216
rect 19796 35176 19797 35216
rect 19755 35167 19797 35176
rect 19756 35082 19796 35167
rect 19852 34721 19892 35755
rect 19948 35384 19988 35932
rect 20140 35880 20180 35889
rect 20043 35804 20085 35813
rect 20140 35804 20180 35840
rect 20523 35888 20565 35897
rect 20523 35848 20524 35888
rect 20564 35848 20565 35888
rect 20523 35839 20565 35848
rect 20043 35764 20044 35804
rect 20084 35764 20180 35804
rect 20043 35755 20085 35764
rect 20048 35552 20416 35561
rect 20088 35512 20130 35552
rect 20170 35512 20212 35552
rect 20252 35512 20294 35552
rect 20334 35512 20376 35552
rect 20048 35503 20416 35512
rect 19948 35344 20084 35384
rect 19947 34964 19989 34973
rect 19947 34924 19948 34964
rect 19988 34924 19989 34964
rect 19947 34915 19989 34924
rect 19948 34830 19988 34915
rect 19851 34712 19893 34721
rect 19851 34672 19852 34712
rect 19892 34672 19893 34712
rect 19851 34663 19893 34672
rect 19852 34544 19892 34553
rect 19660 34385 19700 34470
rect 19755 34460 19797 34469
rect 19755 34420 19756 34460
rect 19796 34420 19797 34460
rect 19755 34411 19797 34420
rect 19659 34376 19701 34385
rect 19659 34336 19660 34376
rect 19700 34336 19701 34376
rect 19659 34327 19701 34336
rect 19756 34326 19796 34411
rect 19564 34168 19700 34208
rect 19372 33620 19412 34168
rect 19660 33704 19700 34168
rect 19852 33788 19892 34504
rect 19947 34544 19989 34553
rect 19947 34504 19948 34544
rect 19988 34504 19989 34544
rect 19947 34495 19989 34504
rect 19948 34460 19988 34495
rect 19948 34409 19988 34420
rect 20044 34376 20084 35344
rect 20044 34327 20084 34336
rect 20236 35048 20276 35057
rect 20236 34208 20276 35008
rect 19948 34168 20276 34208
rect 19948 33965 19988 34168
rect 20048 34040 20416 34049
rect 20088 34000 20130 34040
rect 20170 34000 20212 34040
rect 20252 34000 20294 34040
rect 20334 34000 20376 34040
rect 20048 33991 20416 34000
rect 19947 33956 19989 33965
rect 19947 33916 19948 33956
rect 19988 33916 19989 33956
rect 19947 33907 19989 33916
rect 20524 33797 20564 35839
rect 20620 34553 20660 36091
rect 20716 35561 20756 39367
rect 20812 35897 20852 39535
rect 21387 39332 21429 39341
rect 21387 39292 21388 39332
rect 21428 39292 21429 39332
rect 21387 39283 21429 39292
rect 21388 39089 21428 39283
rect 21387 39080 21429 39089
rect 21387 39040 21388 39080
rect 21428 39040 21429 39080
rect 21387 39031 21429 39040
rect 20907 37736 20949 37745
rect 20907 37696 20908 37736
rect 20948 37696 20949 37736
rect 20907 37687 20949 37696
rect 20811 35888 20853 35897
rect 20811 35848 20812 35888
rect 20852 35848 20853 35888
rect 20811 35839 20853 35848
rect 20811 35720 20853 35729
rect 20811 35680 20812 35720
rect 20852 35680 20853 35720
rect 20811 35671 20853 35680
rect 20715 35552 20757 35561
rect 20715 35512 20716 35552
rect 20756 35512 20757 35552
rect 20715 35503 20757 35512
rect 20619 34544 20661 34553
rect 20619 34504 20620 34544
rect 20660 34504 20661 34544
rect 20619 34495 20661 34504
rect 20812 34049 20852 35671
rect 20811 34040 20853 34049
rect 20811 34000 20812 34040
rect 20852 34000 20853 34040
rect 20811 33991 20853 34000
rect 19660 33655 19700 33664
rect 19756 33748 19892 33788
rect 20523 33788 20565 33797
rect 20523 33748 20524 33788
rect 20564 33748 20565 33788
rect 19372 33571 19412 33580
rect 19564 33620 19604 33629
rect 19084 33536 19124 33545
rect 18988 33496 19084 33536
rect 19084 33487 19124 33496
rect 19467 33536 19509 33545
rect 19467 33496 19468 33536
rect 19508 33496 19509 33536
rect 19564 33536 19604 33580
rect 19756 33536 19796 33748
rect 20523 33739 20565 33748
rect 19851 33620 19893 33629
rect 19851 33580 19852 33620
rect 19892 33580 19893 33620
rect 19851 33571 19893 33580
rect 19564 33496 19796 33536
rect 19467 33487 19509 33496
rect 19468 33402 19508 33487
rect 19852 33486 19892 33571
rect 20043 33452 20085 33461
rect 20043 33412 20044 33452
rect 20084 33412 20085 33452
rect 20043 33403 20085 33412
rect 20044 33318 20084 33403
rect 18699 33284 18741 33293
rect 18699 33244 18700 33284
rect 18740 33244 18741 33284
rect 18699 33235 18741 33244
rect 18808 33284 19176 33293
rect 18848 33244 18890 33284
rect 18930 33244 18972 33284
rect 19012 33244 19054 33284
rect 19094 33244 19136 33284
rect 18808 33235 19176 33244
rect 18603 33200 18645 33209
rect 18603 33160 18604 33200
rect 18644 33160 18645 33200
rect 18603 33151 18645 33160
rect 20043 33200 20085 33209
rect 20043 33160 20044 33200
rect 20084 33160 20085 33200
rect 20043 33151 20085 33160
rect 19275 33116 19317 33125
rect 19275 33076 19276 33116
rect 19316 33076 19317 33116
rect 19275 33067 19317 33076
rect 18316 33032 18356 33041
rect 18356 32992 18740 33032
rect 18316 32983 18356 32992
rect 18603 32864 18645 32873
rect 18603 32824 18604 32864
rect 18644 32824 18645 32864
rect 18603 32815 18645 32824
rect 18315 32780 18357 32789
rect 18315 32740 18316 32780
rect 18356 32740 18357 32780
rect 18315 32731 18357 32740
rect 17644 32311 17684 32320
rect 17932 32320 18260 32360
rect 17451 32192 17493 32201
rect 17836 32192 17876 32201
rect 17451 32152 17452 32192
rect 17492 32152 17493 32192
rect 17451 32143 17493 32152
rect 17548 32152 17836 32192
rect 17452 32058 17492 32143
rect 17356 31109 17396 31312
rect 17355 31100 17397 31109
rect 17355 31060 17356 31100
rect 17396 31060 17397 31100
rect 17355 31051 17397 31060
rect 17163 31016 17205 31025
rect 17163 30976 17164 31016
rect 17204 30976 17205 31016
rect 17163 30967 17205 30976
rect 17548 30932 17588 32152
rect 17836 32143 17876 32152
rect 17644 31940 17684 31949
rect 17835 31940 17877 31949
rect 17684 31900 17780 31940
rect 17644 31891 17684 31900
rect 17740 31352 17780 31900
rect 17835 31900 17836 31940
rect 17876 31900 17877 31940
rect 17835 31891 17877 31900
rect 17836 31806 17876 31891
rect 17643 31268 17685 31277
rect 17643 31228 17644 31268
rect 17684 31228 17685 31268
rect 17643 31219 17685 31228
rect 17356 30892 17588 30932
rect 17260 30666 17300 30675
rect 17260 30101 17300 30626
rect 17259 30092 17301 30101
rect 17259 30052 17260 30092
rect 17300 30052 17301 30092
rect 17356 30092 17396 30892
rect 17644 30848 17684 31219
rect 17644 30799 17684 30808
rect 17740 30773 17780 31312
rect 17452 30764 17492 30773
rect 17739 30764 17781 30773
rect 17492 30724 17588 30764
rect 17452 30715 17492 30724
rect 17548 30260 17588 30724
rect 17739 30724 17740 30764
rect 17780 30724 17781 30764
rect 17739 30715 17781 30724
rect 17836 30689 17876 30774
rect 17835 30680 17877 30689
rect 17835 30640 17836 30680
rect 17876 30640 17877 30680
rect 17835 30631 17877 30640
rect 17932 30666 17972 32320
rect 18028 32192 18068 32201
rect 18028 31613 18068 32152
rect 18220 32192 18260 32201
rect 18316 32192 18356 32731
rect 18604 32730 18644 32815
rect 18603 32612 18645 32621
rect 18603 32572 18604 32612
rect 18644 32572 18645 32612
rect 18603 32563 18645 32572
rect 18411 32360 18453 32369
rect 18411 32320 18412 32360
rect 18452 32320 18453 32360
rect 18411 32311 18453 32320
rect 18260 32152 18356 32192
rect 18220 32143 18260 32152
rect 18412 31940 18452 32311
rect 18220 31900 18452 31940
rect 18027 31604 18069 31613
rect 18027 31564 18028 31604
rect 18068 31564 18069 31604
rect 18027 31555 18069 31564
rect 18028 31352 18068 31363
rect 18028 31277 18068 31312
rect 18027 31268 18069 31277
rect 18027 31228 18028 31268
rect 18068 31228 18069 31268
rect 18027 31219 18069 31228
rect 18124 31268 18164 31279
rect 18124 31193 18164 31228
rect 18123 31184 18165 31193
rect 18123 31144 18124 31184
rect 18164 31144 18165 31184
rect 18123 31135 18165 31144
rect 18123 30848 18165 30857
rect 18123 30808 18124 30848
rect 18164 30808 18165 30848
rect 18123 30799 18165 30808
rect 18124 30680 18164 30799
rect 17932 30626 17983 30666
rect 18124 30631 18164 30640
rect 17836 30512 17876 30521
rect 17836 30428 17876 30472
rect 17943 30428 17983 30626
rect 18123 30512 18165 30521
rect 18123 30472 18124 30512
rect 18164 30472 18165 30512
rect 18123 30463 18165 30472
rect 17836 30388 17983 30428
rect 17739 30260 17781 30269
rect 17548 30220 17684 30260
rect 17356 30052 17588 30092
rect 17259 30043 17301 30052
rect 17067 29924 17109 29933
rect 17067 29884 17068 29924
rect 17108 29884 17109 29924
rect 17067 29875 17109 29884
rect 17548 29924 17588 30052
rect 17548 29875 17588 29884
rect 17068 29840 17108 29875
rect 17068 29789 17108 29800
rect 17451 29840 17493 29849
rect 17451 29800 17452 29840
rect 17492 29800 17493 29840
rect 17451 29791 17493 29800
rect 17644 29840 17684 30220
rect 17739 30220 17740 30260
rect 17780 30220 17781 30260
rect 17739 30211 17781 30220
rect 17644 29791 17684 29800
rect 17452 29706 17492 29791
rect 17547 29756 17589 29765
rect 17547 29716 17548 29756
rect 17588 29716 17589 29756
rect 17547 29707 17589 29716
rect 16972 29548 17204 29588
rect 17164 29504 17204 29548
rect 17164 29464 17300 29504
rect 16971 29420 17013 29429
rect 16971 29380 16972 29420
rect 17012 29380 17013 29420
rect 16971 29371 17013 29380
rect 16875 27740 16917 27749
rect 16875 27700 16876 27740
rect 16916 27700 16917 27740
rect 16875 27691 16917 27700
rect 16587 27656 16629 27665
rect 16436 27616 16532 27656
rect 16396 27607 16436 27616
rect 16204 27439 16244 27448
rect 16300 27572 16340 27607
rect 16300 27245 16340 27532
rect 16492 27488 16532 27616
rect 16587 27616 16588 27656
rect 16628 27616 16629 27656
rect 16587 27607 16629 27616
rect 16779 27656 16821 27665
rect 16779 27616 16780 27656
rect 16820 27616 16821 27656
rect 16779 27607 16821 27616
rect 16780 27522 16820 27607
rect 16972 27572 17012 29371
rect 17067 29336 17109 29345
rect 17067 29296 17068 29336
rect 17108 29296 17109 29336
rect 17067 29287 17109 29296
rect 17068 29168 17108 29287
rect 17163 29252 17205 29261
rect 17163 29212 17164 29252
rect 17204 29212 17205 29252
rect 17163 29203 17205 29212
rect 17068 29119 17108 29128
rect 16972 27523 17012 27532
rect 16588 27488 16628 27497
rect 16492 27448 16588 27488
rect 16588 27439 16628 27448
rect 17164 27488 17204 29203
rect 17260 28337 17300 29464
rect 17451 29168 17493 29177
rect 17451 29128 17452 29168
rect 17492 29128 17493 29168
rect 17451 29119 17493 29128
rect 17259 28328 17301 28337
rect 17259 28288 17260 28328
rect 17300 28288 17301 28328
rect 17259 28279 17301 28288
rect 17452 28328 17492 29119
rect 17452 28279 17492 28288
rect 17164 27439 17204 27448
rect 16299 27236 16341 27245
rect 16299 27196 16300 27236
rect 16340 27196 16341 27236
rect 16299 27187 16341 27196
rect 17260 27161 17300 28279
rect 17451 27656 17493 27665
rect 17451 27616 17452 27656
rect 17492 27616 17493 27656
rect 17451 27607 17493 27616
rect 17356 27572 17396 27583
rect 17356 27497 17396 27532
rect 17355 27488 17397 27497
rect 17355 27448 17356 27488
rect 17396 27448 17397 27488
rect 17355 27439 17397 27448
rect 16011 27152 16053 27161
rect 16011 27112 16012 27152
rect 16052 27112 16053 27152
rect 16011 27103 16053 27112
rect 17259 27152 17301 27161
rect 17259 27112 17260 27152
rect 17300 27112 17301 27152
rect 17259 27103 17301 27112
rect 17452 27077 17492 27607
rect 17548 27488 17588 29707
rect 17644 28160 17684 28169
rect 17644 27917 17684 28120
rect 17643 27908 17685 27917
rect 17643 27868 17644 27908
rect 17684 27868 17685 27908
rect 17643 27859 17685 27868
rect 17740 27581 17780 30211
rect 17836 30101 17876 30388
rect 17835 30092 17877 30101
rect 17835 30052 17836 30092
rect 17876 30052 17877 30092
rect 17835 30043 17877 30052
rect 17836 29840 17876 29849
rect 17836 29597 17876 29800
rect 18027 29672 18069 29681
rect 18027 29632 18028 29672
rect 18068 29632 18069 29672
rect 18027 29623 18069 29632
rect 17835 29588 17877 29597
rect 17835 29548 17836 29588
rect 17876 29548 17877 29588
rect 17835 29539 17877 29548
rect 17932 28328 17972 28337
rect 17835 27992 17877 28001
rect 17835 27952 17836 27992
rect 17876 27952 17877 27992
rect 17835 27943 17877 27952
rect 17836 27656 17876 27943
rect 17932 27917 17972 28288
rect 18028 28328 18068 29623
rect 17931 27908 17973 27917
rect 17931 27868 17932 27908
rect 17972 27868 17973 27908
rect 17931 27859 17973 27868
rect 17836 27607 17876 27616
rect 17932 27656 17972 27665
rect 17739 27572 17781 27581
rect 17739 27532 17740 27572
rect 17780 27532 17781 27572
rect 17739 27523 17781 27532
rect 17548 27439 17588 27448
rect 17932 27152 17972 27616
rect 17836 27112 17972 27152
rect 16203 27068 16245 27077
rect 16203 27028 16204 27068
rect 16244 27028 16245 27068
rect 16203 27019 16245 27028
rect 17451 27068 17493 27077
rect 17451 27028 17452 27068
rect 17492 27028 17493 27068
rect 17451 27019 17493 27028
rect 17739 27068 17781 27077
rect 17739 27028 17740 27068
rect 17780 27028 17781 27068
rect 17739 27019 17781 27028
rect 16204 26816 16244 27019
rect 16396 26984 16436 26993
rect 17643 26984 17685 26993
rect 16012 26648 16052 26657
rect 16012 26405 16052 26608
rect 16011 26396 16053 26405
rect 16011 26356 16012 26396
rect 16052 26356 16053 26396
rect 16011 26347 16053 26356
rect 16012 26237 16052 26268
rect 16011 26228 16053 26237
rect 16011 26188 16012 26228
rect 16052 26188 16053 26228
rect 16011 26179 16053 26188
rect 16012 26144 16052 26179
rect 16012 24053 16052 26104
rect 16107 26144 16149 26153
rect 16107 26104 16108 26144
rect 16148 26104 16149 26144
rect 16107 26095 16149 26104
rect 16108 26010 16148 26095
rect 16204 25313 16244 26776
rect 16300 26900 16340 26909
rect 16300 25976 16340 26860
rect 16396 26228 16436 26944
rect 16780 26909 16820 26953
rect 17643 26944 17644 26984
rect 17684 26944 17685 26984
rect 17643 26935 17685 26944
rect 16492 26900 16532 26909
rect 16492 26489 16532 26860
rect 16779 26900 16821 26909
rect 16779 26860 16780 26900
rect 16820 26860 16821 26900
rect 16779 26858 16821 26860
rect 16779 26851 16780 26858
rect 16588 26816 16628 26825
rect 16820 26851 16821 26858
rect 16972 26825 17012 26910
rect 17547 26900 17589 26909
rect 17547 26860 17548 26900
rect 17588 26860 17589 26900
rect 17547 26851 17589 26860
rect 16780 26809 16820 26818
rect 16971 26816 17013 26825
rect 16491 26480 16533 26489
rect 16491 26440 16492 26480
rect 16532 26440 16533 26480
rect 16491 26431 16533 26440
rect 16588 26321 16628 26776
rect 16971 26776 16972 26816
rect 17012 26776 17013 26816
rect 16971 26767 17013 26776
rect 17068 26816 17108 26825
rect 17259 26816 17301 26825
rect 17108 26776 17204 26816
rect 17068 26767 17108 26776
rect 16780 26648 16820 26657
rect 16780 26564 16820 26608
rect 17067 26648 17109 26657
rect 17067 26608 17068 26648
rect 17108 26608 17109 26648
rect 17067 26599 17109 26608
rect 16780 26524 16847 26564
rect 16807 26480 16847 26524
rect 16807 26440 17012 26480
rect 16587 26312 16629 26321
rect 16587 26272 16588 26312
rect 16628 26272 16629 26312
rect 16587 26263 16629 26272
rect 16684 26312 16724 26321
rect 16684 26237 16724 26272
rect 16875 26312 16917 26321
rect 16875 26272 16876 26312
rect 16916 26272 16917 26312
rect 16875 26263 16917 26272
rect 16684 26228 16728 26237
rect 16396 26188 16532 26228
rect 16684 26188 16687 26228
rect 16727 26188 16728 26228
rect 16396 25976 16436 25985
rect 16300 25936 16396 25976
rect 16396 25927 16436 25936
rect 16492 25808 16532 26188
rect 16686 26179 16728 26188
rect 16780 26144 16820 26155
rect 16622 26129 16662 26138
rect 16622 25808 16662 26089
rect 16780 26069 16820 26104
rect 16876 26144 16916 26263
rect 16876 26095 16916 26104
rect 16779 26060 16821 26069
rect 16779 26020 16780 26060
rect 16820 26020 16821 26060
rect 16779 26011 16821 26020
rect 16396 25768 16532 25808
rect 16588 25768 16662 25808
rect 16396 25388 16436 25768
rect 16492 25556 16532 25565
rect 16588 25556 16628 25768
rect 16972 25724 17012 26440
rect 17068 26144 17108 26599
rect 17164 26573 17204 26776
rect 17259 26776 17260 26816
rect 17300 26776 17301 26816
rect 17259 26767 17301 26776
rect 17163 26564 17205 26573
rect 17163 26524 17164 26564
rect 17204 26524 17205 26564
rect 17163 26515 17205 26524
rect 17163 26396 17205 26405
rect 17163 26356 17164 26396
rect 17204 26356 17205 26396
rect 17163 26347 17205 26356
rect 17068 26095 17108 26104
rect 17164 26144 17204 26347
rect 17164 25892 17204 26104
rect 16532 25516 16628 25556
rect 16684 25684 17012 25724
rect 17068 25852 17204 25892
rect 16492 25507 16532 25516
rect 16491 25388 16533 25397
rect 16396 25348 16492 25388
rect 16532 25348 16533 25388
rect 16491 25339 16533 25348
rect 16107 25304 16149 25313
rect 16107 25264 16108 25304
rect 16148 25264 16149 25304
rect 16204 25273 16340 25313
rect 16107 25255 16149 25264
rect 16108 25170 16148 25255
rect 16204 25220 16244 25231
rect 16204 25145 16244 25180
rect 16203 25136 16245 25145
rect 16203 25096 16204 25136
rect 16244 25096 16245 25136
rect 16203 25087 16245 25096
rect 16108 24632 16148 24643
rect 16108 24557 16148 24592
rect 16107 24548 16149 24557
rect 16107 24508 16108 24548
rect 16148 24508 16149 24548
rect 16300 24548 16340 25273
rect 16684 25304 16724 25684
rect 17068 25640 17108 25852
rect 17163 25724 17205 25733
rect 17163 25684 17164 25724
rect 17204 25684 17205 25724
rect 17163 25675 17205 25684
rect 16972 25600 17108 25640
rect 16876 25472 16916 25481
rect 16779 25388 16821 25397
rect 16779 25348 16780 25388
rect 16820 25348 16821 25388
rect 16779 25339 16821 25348
rect 16684 25255 16724 25264
rect 16780 25254 16820 25339
rect 16491 25220 16533 25229
rect 16491 25180 16492 25220
rect 16532 25180 16533 25220
rect 16491 25171 16533 25180
rect 16492 24641 16532 25171
rect 16683 25136 16725 25145
rect 16683 25096 16684 25136
rect 16724 25096 16725 25136
rect 16683 25087 16725 25096
rect 16491 24632 16533 24641
rect 16491 24592 16492 24632
rect 16532 24592 16533 24632
rect 16491 24583 16533 24592
rect 16587 24548 16629 24557
rect 16300 24508 16436 24548
rect 16107 24499 16149 24508
rect 16300 24380 16340 24389
rect 16108 24340 16300 24380
rect 16011 24044 16053 24053
rect 16011 24004 16012 24044
rect 16052 24004 16053 24044
rect 16011 23995 16053 24004
rect 16108 23876 16148 24340
rect 16300 24331 16340 24340
rect 16060 23836 16148 23876
rect 16060 23834 16100 23836
rect 16060 23785 16100 23794
rect 16396 23792 16436 24508
rect 16587 24508 16588 24548
rect 16628 24508 16629 24548
rect 16587 24499 16629 24508
rect 16588 23792 16628 24499
rect 16396 23752 16532 23792
rect 16011 23708 16053 23717
rect 16011 23668 16012 23708
rect 16052 23668 16053 23708
rect 16011 23659 16053 23668
rect 16012 22112 16052 23659
rect 16203 23624 16245 23633
rect 16396 23624 16436 23633
rect 16203 23584 16204 23624
rect 16244 23584 16245 23624
rect 16203 23575 16245 23584
rect 16300 23584 16396 23624
rect 16204 23490 16244 23575
rect 16300 23372 16340 23584
rect 16396 23575 16436 23584
rect 16204 23332 16340 23372
rect 16204 23119 16244 23332
rect 16299 23204 16341 23213
rect 16492 23204 16532 23752
rect 16588 23549 16628 23752
rect 16587 23540 16629 23549
rect 16587 23500 16588 23540
rect 16628 23500 16629 23540
rect 16587 23491 16629 23500
rect 16299 23164 16300 23204
rect 16340 23164 16341 23204
rect 16299 23155 16341 23164
rect 16396 23164 16532 23204
rect 16156 23110 16244 23119
rect 16196 23079 16244 23110
rect 16156 23061 16196 23070
rect 16300 22952 16340 23155
rect 16204 22912 16340 22952
rect 16108 22289 16148 22374
rect 16107 22280 16149 22289
rect 16107 22240 16108 22280
rect 16148 22240 16149 22280
rect 16107 22231 16149 22240
rect 16012 22072 16148 22112
rect 16011 21944 16053 21953
rect 16011 21904 16012 21944
rect 16052 21904 16053 21944
rect 16011 21895 16053 21904
rect 15820 20140 15956 20180
rect 15628 20096 15668 20105
rect 15435 20012 15477 20021
rect 15435 19972 15436 20012
rect 15476 19972 15477 20012
rect 15435 19963 15477 19972
rect 15628 19088 15668 20056
rect 15820 20096 15860 20140
rect 15723 19256 15765 19265
rect 15723 19216 15724 19256
rect 15764 19216 15765 19256
rect 15723 19207 15765 19216
rect 15148 18535 15188 18544
rect 15244 18712 15380 18752
rect 15436 19048 15668 19088
rect 15244 18089 15284 18712
rect 15340 18584 15380 18595
rect 15340 18509 15380 18544
rect 15339 18500 15381 18509
rect 15339 18460 15340 18500
rect 15380 18460 15381 18500
rect 15339 18451 15381 18460
rect 15436 18425 15476 19048
rect 15627 18920 15669 18929
rect 15627 18880 15628 18920
rect 15668 18880 15669 18920
rect 15627 18871 15669 18880
rect 15532 18668 15572 18677
rect 15532 18509 15572 18628
rect 15531 18500 15573 18509
rect 15531 18460 15532 18500
rect 15572 18460 15573 18500
rect 15531 18451 15573 18460
rect 15435 18416 15477 18425
rect 15435 18376 15436 18416
rect 15476 18376 15477 18416
rect 15435 18367 15477 18376
rect 15339 18332 15381 18341
rect 15339 18292 15340 18332
rect 15380 18292 15381 18332
rect 15339 18283 15381 18292
rect 15340 18198 15380 18283
rect 15243 18080 15285 18089
rect 15243 18040 15244 18080
rect 15284 18040 15285 18080
rect 15243 18031 15285 18040
rect 14955 17996 14997 18005
rect 14955 17956 14956 17996
rect 14996 17956 14997 17996
rect 14955 17947 14997 17956
rect 15628 17996 15668 18871
rect 15724 18579 15764 19207
rect 15724 18530 15764 18539
rect 15820 18416 15860 20056
rect 15915 19844 15957 19853
rect 15915 19804 15916 19844
rect 15956 19804 15957 19844
rect 15915 19795 15957 19804
rect 15628 17947 15668 17956
rect 15724 18376 15860 18416
rect 14956 17862 14996 17947
rect 15147 17828 15189 17837
rect 15724 17828 15764 18376
rect 15147 17788 15148 17828
rect 15188 17788 15189 17828
rect 15147 17779 15189 17788
rect 15340 17788 15764 17828
rect 15819 17828 15861 17837
rect 15819 17788 15820 17828
rect 15860 17788 15861 17828
rect 14860 17713 14996 17753
rect 14764 17611 14804 17620
rect 14859 17576 14901 17585
rect 14859 17536 14860 17576
rect 14900 17536 14901 17576
rect 14859 17527 14901 17536
rect 14764 17240 14804 17249
rect 14668 17200 14764 17240
rect 14764 17191 14804 17200
rect 14571 17156 14613 17165
rect 14571 17116 14572 17156
rect 14612 17116 14613 17156
rect 14571 17107 14613 17116
rect 14572 17072 14612 17107
rect 14572 17021 14612 17032
rect 14667 17072 14709 17081
rect 14667 17032 14668 17072
rect 14708 17032 14709 17072
rect 14667 17023 14709 17032
rect 14571 16232 14613 16241
rect 14571 16192 14572 16232
rect 14612 16192 14613 16232
rect 14571 16183 14613 16192
rect 14572 16073 14612 16183
rect 14571 16064 14613 16073
rect 14571 16024 14572 16064
rect 14612 16024 14613 16064
rect 14571 16015 14613 16024
rect 14572 14048 14612 14057
rect 14476 14034 14572 14048
rect 14091 11992 14092 12032
rect 14132 11992 14133 12032
rect 14091 11983 14133 11992
rect 14188 11992 14324 12032
rect 14380 14008 14572 14034
rect 14380 13994 14516 14008
rect 14572 13999 14612 14008
rect 14091 11528 14133 11537
rect 14091 11488 14092 11528
rect 14132 11488 14133 11528
rect 14091 11479 14133 11488
rect 14092 11394 14132 11479
rect 13996 10975 14036 10984
rect 14091 10436 14133 10445
rect 14091 10396 14092 10436
rect 14132 10396 14133 10436
rect 14091 10387 14133 10396
rect 14092 9941 14132 10387
rect 14091 9932 14133 9941
rect 14091 9892 14092 9932
rect 14132 9892 14133 9932
rect 14091 9883 14133 9892
rect 13803 9260 13845 9269
rect 13803 9220 13804 9260
rect 13844 9220 13845 9260
rect 13803 9211 13845 9220
rect 13707 9176 13749 9185
rect 13707 9136 13708 9176
rect 13748 9136 13749 9176
rect 13707 9127 13749 9136
rect 13612 8623 13652 8632
rect 13611 7832 13653 7841
rect 13611 7792 13612 7832
rect 13652 7792 13653 7832
rect 13611 7783 13653 7792
rect 13515 7328 13557 7337
rect 13515 7288 13516 7328
rect 13556 7288 13557 7328
rect 13515 7279 13557 7288
rect 13324 7160 13364 7169
rect 13228 7120 13324 7160
rect 12844 6992 12884 7120
rect 13324 7111 13364 7120
rect 12364 5440 12596 5480
rect 12748 6952 12884 6992
rect 12364 4976 12404 5440
rect 12748 4985 12788 6952
rect 12843 6656 12885 6665
rect 12843 6616 12844 6656
rect 12884 6616 12885 6656
rect 12843 6607 12885 6616
rect 12364 4565 12404 4936
rect 12555 4976 12597 4985
rect 12555 4936 12556 4976
rect 12596 4936 12597 4976
rect 12555 4927 12597 4936
rect 12747 4976 12789 4985
rect 12747 4936 12748 4976
rect 12788 4936 12789 4976
rect 12747 4927 12789 4936
rect 12459 4892 12501 4901
rect 12459 4852 12460 4892
rect 12500 4852 12501 4892
rect 12459 4843 12501 4852
rect 12460 4758 12500 4843
rect 12459 4640 12501 4649
rect 12459 4600 12460 4640
rect 12500 4600 12501 4640
rect 12459 4591 12501 4600
rect 12363 4556 12405 4565
rect 12363 4516 12364 4556
rect 12404 4516 12405 4556
rect 12363 4507 12405 4516
rect 12460 4136 12500 4591
rect 12556 4481 12596 4927
rect 12747 4808 12789 4817
rect 12747 4768 12748 4808
rect 12788 4768 12789 4808
rect 12747 4759 12789 4768
rect 12555 4472 12597 4481
rect 12555 4432 12556 4472
rect 12596 4432 12597 4472
rect 12555 4423 12597 4432
rect 12748 4145 12788 4759
rect 12460 4061 12500 4096
rect 12747 4136 12789 4145
rect 12747 4096 12748 4136
rect 12788 4096 12789 4136
rect 12747 4087 12789 4096
rect 12459 4052 12501 4061
rect 12459 4012 12460 4052
rect 12500 4012 12501 4052
rect 12459 4003 12501 4012
rect 12171 3884 12213 3893
rect 12171 3844 12172 3884
rect 12212 3844 12213 3884
rect 12171 3835 12213 3844
rect 12651 3548 12693 3557
rect 12651 3508 12652 3548
rect 12692 3508 12693 3548
rect 12651 3499 12693 3508
rect 11787 3464 11829 3473
rect 11787 3424 11788 3464
rect 11828 3424 11829 3464
rect 11787 3415 11829 3424
rect 11788 3330 11828 3415
rect 11787 3128 11829 3137
rect 11787 3088 11788 3128
rect 11828 3088 11829 3128
rect 11787 3079 11829 3088
rect 11788 2633 11828 3079
rect 11883 2792 11925 2801
rect 11883 2752 11884 2792
rect 11924 2752 11925 2792
rect 11883 2743 11925 2752
rect 11787 2624 11829 2633
rect 11787 2584 11788 2624
rect 11828 2584 11829 2624
rect 11787 2575 11829 2584
rect 11884 2624 11924 2743
rect 11884 2575 11924 2584
rect 12364 2629 12404 2638
rect 12364 2540 12404 2589
rect 11980 2500 12404 2540
rect 12556 2540 12596 2549
rect 12652 2540 12692 3499
rect 12748 2624 12788 4087
rect 12844 3305 12884 6607
rect 12939 5984 12981 5993
rect 12939 5944 12940 5984
rect 12980 5944 12981 5984
rect 13612 5984 13652 7783
rect 13708 7076 13748 9127
rect 14091 7496 14133 7505
rect 14091 7456 14092 7496
rect 14132 7456 14133 7496
rect 14091 7447 14133 7456
rect 13852 7169 13892 7178
rect 13892 7129 13940 7160
rect 13852 7120 13940 7129
rect 13708 7036 13844 7076
rect 13707 6488 13749 6497
rect 13707 6448 13708 6488
rect 13748 6448 13749 6488
rect 13707 6439 13749 6448
rect 13708 6354 13748 6439
rect 13612 5944 13748 5984
rect 12939 5935 12981 5944
rect 12940 4976 12980 5935
rect 13611 5816 13653 5825
rect 13611 5776 13612 5816
rect 13652 5776 13653 5816
rect 13611 5767 13653 5776
rect 13036 5648 13076 5657
rect 13036 5489 13076 5608
rect 13516 5648 13556 5657
rect 13228 5564 13268 5573
rect 13516 5564 13556 5608
rect 13612 5648 13652 5767
rect 13612 5599 13652 5608
rect 13268 5524 13556 5564
rect 13228 5515 13268 5524
rect 13035 5480 13077 5489
rect 13035 5440 13036 5480
rect 13076 5440 13077 5480
rect 13035 5431 13077 5440
rect 13516 4985 13556 5524
rect 13612 5060 13652 5069
rect 13515 4976 13557 4985
rect 13420 4962 13460 4971
rect 12940 4817 12980 4936
rect 13132 4922 13420 4962
rect 13515 4936 13516 4976
rect 13556 4936 13557 4976
rect 13515 4927 13557 4936
rect 12939 4808 12981 4817
rect 12939 4768 12940 4808
rect 12980 4768 12981 4808
rect 12939 4759 12981 4768
rect 12988 4145 13028 4154
rect 13132 4136 13172 4922
rect 13420 4913 13460 4922
rect 13419 4724 13461 4733
rect 13419 4684 13420 4724
rect 13460 4684 13461 4724
rect 13419 4675 13461 4684
rect 13323 4388 13365 4397
rect 13323 4348 13324 4388
rect 13364 4348 13365 4388
rect 13323 4339 13365 4348
rect 13324 4254 13364 4339
rect 13028 4105 13172 4136
rect 12988 4096 13172 4105
rect 13036 3800 13076 4096
rect 13132 3968 13172 3977
rect 13172 3928 13364 3968
rect 13132 3919 13172 3928
rect 13036 3760 13268 3800
rect 13228 3632 13268 3760
rect 13228 3583 13268 3592
rect 13324 3557 13364 3928
rect 13035 3548 13077 3557
rect 13035 3508 13036 3548
rect 13076 3508 13077 3548
rect 13035 3499 13077 3508
rect 13323 3548 13365 3557
rect 13323 3508 13324 3548
rect 13364 3508 13365 3548
rect 13323 3499 13365 3508
rect 13036 3464 13076 3499
rect 12843 3296 12885 3305
rect 12843 3256 12844 3296
rect 12884 3256 12885 3296
rect 12843 3247 12885 3256
rect 13036 2801 13076 3424
rect 13420 2960 13460 4675
rect 13515 4388 13557 4397
rect 13515 4348 13516 4388
rect 13556 4348 13557 4388
rect 13515 4339 13557 4348
rect 13516 4220 13556 4339
rect 13516 4171 13556 4180
rect 13612 4136 13652 5020
rect 13708 4733 13748 5944
rect 13707 4724 13749 4733
rect 13707 4684 13708 4724
rect 13748 4684 13749 4724
rect 13707 4675 13749 4684
rect 13804 4397 13844 7036
rect 13900 6656 13940 7120
rect 13996 7085 14036 7170
rect 13995 7076 14037 7085
rect 13995 7036 13996 7076
rect 14036 7036 14037 7076
rect 13995 7027 14037 7036
rect 14092 7001 14132 7447
rect 14091 6992 14133 7001
rect 14091 6952 14092 6992
rect 14132 6952 14133 6992
rect 14091 6943 14133 6952
rect 14188 6740 14228 11992
rect 14284 11780 14324 11791
rect 14284 11705 14324 11740
rect 14283 11696 14325 11705
rect 14283 11656 14284 11696
rect 14324 11656 14325 11696
rect 14283 11647 14325 11656
rect 14380 11201 14420 13994
rect 14668 12452 14708 17023
rect 14763 16904 14805 16913
rect 14763 16864 14764 16904
rect 14804 16864 14805 16904
rect 14763 16855 14805 16864
rect 14764 14645 14804 16855
rect 14763 14636 14805 14645
rect 14763 14596 14764 14636
rect 14804 14596 14805 14636
rect 14763 14587 14805 14596
rect 14860 12704 14900 17527
rect 14956 17072 14996 17713
rect 15148 17694 15188 17779
rect 14956 16913 14996 17032
rect 14955 16904 14997 16913
rect 14955 16864 14956 16904
rect 14996 16864 14997 16904
rect 14955 16855 14997 16864
rect 14955 16400 14997 16409
rect 14955 16360 14956 16400
rect 14996 16360 14997 16400
rect 14955 16351 14997 16360
rect 14956 15653 14996 16351
rect 15100 16241 15140 16250
rect 15140 16201 15188 16232
rect 15100 16192 15188 16201
rect 15148 15728 15188 16192
rect 15243 16064 15285 16073
rect 15243 16024 15244 16064
rect 15284 16024 15285 16064
rect 15243 16015 15285 16024
rect 15244 15930 15284 16015
rect 15148 15679 15188 15688
rect 14955 15644 14997 15653
rect 14955 15604 14956 15644
rect 14996 15604 14997 15644
rect 14955 15595 14997 15604
rect 14956 15560 14996 15595
rect 14956 15317 14996 15520
rect 14955 15308 14997 15317
rect 14955 15268 14956 15308
rect 14996 15268 14997 15308
rect 14955 15259 14997 15268
rect 15051 15140 15093 15149
rect 15051 15100 15052 15140
rect 15092 15100 15093 15140
rect 15051 15091 15093 15100
rect 15052 13208 15092 15091
rect 15243 14048 15285 14057
rect 15243 14008 15244 14048
rect 15284 14008 15285 14048
rect 15243 13999 15285 14008
rect 15244 13385 15284 13999
rect 15243 13376 15285 13385
rect 15243 13336 15244 13376
rect 15284 13336 15285 13376
rect 15243 13327 15285 13336
rect 15052 13159 15092 13168
rect 15244 13208 15284 13327
rect 15244 13159 15284 13168
rect 14860 12664 14996 12704
rect 14860 12536 14900 12545
rect 14668 12403 14708 12412
rect 14764 12496 14860 12536
rect 14476 12284 14516 12293
rect 14476 12125 14516 12244
rect 14475 12116 14517 12125
rect 14475 12076 14476 12116
rect 14516 12076 14517 12116
rect 14475 12067 14517 12076
rect 14475 11948 14517 11957
rect 14764 11948 14804 12496
rect 14860 12487 14900 12496
rect 14859 12284 14901 12293
rect 14859 12244 14860 12284
rect 14900 12244 14901 12284
rect 14859 12235 14901 12244
rect 14860 12150 14900 12235
rect 14475 11908 14476 11948
rect 14516 11908 14517 11948
rect 14475 11899 14517 11908
rect 14668 11908 14804 11948
rect 14476 11705 14516 11899
rect 14475 11696 14517 11705
rect 14475 11656 14476 11696
rect 14516 11656 14517 11696
rect 14475 11647 14517 11656
rect 14571 11528 14613 11537
rect 14571 11488 14572 11528
rect 14612 11488 14613 11528
rect 14571 11479 14613 11488
rect 14572 11394 14612 11479
rect 14475 11360 14517 11369
rect 14475 11320 14476 11360
rect 14516 11320 14517 11360
rect 14475 11311 14517 11320
rect 14379 11192 14421 11201
rect 14379 11152 14380 11192
rect 14420 11152 14421 11192
rect 14379 11143 14421 11152
rect 14476 11024 14516 11311
rect 14571 11276 14613 11285
rect 14571 11236 14572 11276
rect 14612 11236 14613 11276
rect 14571 11227 14613 11236
rect 14476 10975 14516 10984
rect 14572 11024 14612 11227
rect 14572 10975 14612 10984
rect 14668 10949 14708 11908
rect 14764 11780 14804 11789
rect 14764 11696 14804 11740
rect 14956 11696 14996 12664
rect 15244 12620 15284 12629
rect 15052 12536 15092 12545
rect 15052 11873 15092 12496
rect 15051 11864 15093 11873
rect 15051 11824 15052 11864
rect 15092 11824 15093 11864
rect 15051 11815 15093 11824
rect 14764 11656 14996 11696
rect 15052 11696 15092 11705
rect 14763 11528 14805 11537
rect 14763 11488 14764 11528
rect 14804 11488 14805 11528
rect 14763 11479 14805 11488
rect 14283 10940 14325 10949
rect 14283 10900 14284 10940
rect 14324 10900 14325 10940
rect 14283 10891 14325 10900
rect 14667 10940 14709 10949
rect 14667 10900 14668 10940
rect 14708 10900 14709 10940
rect 14667 10891 14709 10900
rect 14284 7421 14324 10891
rect 14475 10856 14517 10865
rect 14475 10816 14476 10856
rect 14516 10816 14517 10856
rect 14475 10807 14517 10816
rect 14379 10688 14421 10697
rect 14379 10648 14380 10688
rect 14420 10648 14421 10688
rect 14379 10639 14421 10648
rect 14380 9521 14420 10639
rect 14379 9512 14421 9521
rect 14379 9472 14380 9512
rect 14420 9472 14421 9512
rect 14379 9463 14421 9472
rect 14380 7505 14420 9463
rect 14379 7496 14421 7505
rect 14379 7456 14380 7496
rect 14420 7456 14421 7496
rect 14379 7447 14421 7456
rect 14283 7412 14325 7421
rect 14283 7372 14284 7412
rect 14324 7372 14325 7412
rect 14476 7412 14516 10807
rect 14667 10772 14709 10781
rect 14667 10732 14668 10772
rect 14708 10732 14709 10772
rect 14667 10723 14709 10732
rect 14668 10184 14708 10723
rect 14668 10135 14708 10144
rect 14667 10016 14709 10025
rect 14667 9976 14668 10016
rect 14708 9976 14709 10016
rect 14667 9967 14709 9976
rect 14571 8756 14613 8765
rect 14571 8716 14572 8756
rect 14612 8716 14613 8756
rect 14571 8707 14613 8716
rect 14572 8000 14612 8707
rect 14572 7757 14612 7960
rect 14668 7925 14708 9967
rect 14764 9638 14804 11479
rect 15052 11360 15092 11656
rect 14860 11320 15092 11360
rect 15148 11696 15188 11705
rect 14860 10436 14900 11320
rect 15051 11108 15093 11117
rect 15051 11068 15052 11108
rect 15092 11068 15093 11108
rect 15051 11059 15093 11068
rect 14860 10387 14900 10396
rect 14956 11024 14996 11033
rect 14956 10688 14996 10984
rect 15052 11024 15092 11059
rect 15052 10973 15092 10984
rect 15148 10688 15188 11656
rect 15244 11192 15284 12580
rect 15340 12461 15380 17788
rect 15819 17779 15861 17788
rect 15820 17744 15860 17779
rect 15820 17660 15860 17704
rect 15724 17620 15860 17660
rect 15724 16409 15764 17620
rect 15819 17072 15861 17081
rect 15819 17032 15820 17072
rect 15860 17032 15861 17072
rect 15819 17023 15861 17032
rect 15723 16400 15765 16409
rect 15723 16360 15724 16400
rect 15764 16360 15765 16400
rect 15723 16351 15765 16360
rect 15676 16241 15716 16250
rect 15628 16201 15676 16232
rect 15628 16192 15716 16201
rect 15532 16064 15572 16073
rect 15532 15485 15572 16024
rect 15628 15728 15668 16192
rect 15723 15980 15765 15989
rect 15723 15940 15724 15980
rect 15764 15940 15765 15980
rect 15723 15931 15765 15940
rect 15724 15821 15764 15931
rect 15723 15812 15765 15821
rect 15723 15772 15724 15812
rect 15764 15772 15765 15812
rect 15723 15763 15765 15772
rect 15628 15679 15668 15688
rect 15531 15476 15573 15485
rect 15531 15436 15532 15476
rect 15572 15436 15573 15476
rect 15531 15427 15573 15436
rect 15531 15308 15573 15317
rect 15531 15268 15532 15308
rect 15572 15268 15573 15308
rect 15531 15259 15573 15268
rect 15436 14552 15476 14561
rect 15436 13721 15476 14512
rect 15532 14384 15572 15259
rect 15628 14725 15668 14734
rect 15628 14561 15668 14685
rect 15627 14552 15669 14561
rect 15627 14512 15628 14552
rect 15668 14512 15669 14552
rect 15627 14503 15669 14512
rect 15532 14344 15668 14384
rect 15531 13880 15573 13889
rect 15531 13840 15532 13880
rect 15572 13840 15573 13880
rect 15531 13831 15573 13840
rect 15435 13712 15477 13721
rect 15435 13672 15436 13712
rect 15476 13672 15477 13712
rect 15435 13663 15477 13672
rect 15435 12620 15477 12629
rect 15435 12580 15436 12620
rect 15476 12580 15477 12620
rect 15435 12571 15477 12580
rect 15436 12531 15476 12571
rect 15436 12482 15476 12491
rect 15339 12452 15381 12461
rect 15339 12412 15340 12452
rect 15380 12412 15381 12452
rect 15339 12403 15381 12412
rect 15532 12368 15572 13831
rect 15628 13628 15668 14344
rect 15724 13805 15764 15763
rect 15820 15560 15860 17023
rect 15820 14309 15860 15520
rect 15819 14300 15861 14309
rect 15819 14260 15820 14300
rect 15860 14260 15861 14300
rect 15819 14251 15861 14260
rect 15820 14048 15860 14251
rect 15723 13796 15765 13805
rect 15723 13756 15724 13796
rect 15764 13756 15765 13796
rect 15723 13747 15765 13756
rect 15628 13588 15764 13628
rect 15436 12328 15572 12368
rect 15436 11360 15476 12328
rect 15627 11864 15669 11873
rect 15627 11824 15628 11864
rect 15668 11824 15669 11864
rect 15627 11815 15669 11824
rect 15628 11780 15668 11815
rect 15531 11696 15573 11705
rect 15531 11656 15532 11696
rect 15572 11656 15573 11696
rect 15531 11647 15573 11656
rect 15532 11562 15572 11647
rect 15436 11320 15572 11360
rect 15244 11152 15476 11192
rect 15243 11024 15285 11033
rect 15243 10984 15244 11024
rect 15284 10984 15285 11024
rect 15243 10975 15285 10984
rect 15340 11024 15380 11033
rect 14956 10648 15188 10688
rect 14956 9773 14996 10648
rect 15051 10184 15093 10193
rect 15051 10144 15052 10184
rect 15092 10144 15093 10184
rect 15051 10135 15093 10144
rect 15148 10184 15188 10195
rect 15244 10184 15284 10975
rect 15340 10445 15380 10984
rect 15339 10436 15381 10445
rect 15339 10396 15340 10436
rect 15380 10396 15381 10436
rect 15339 10387 15381 10396
rect 15340 10184 15380 10193
rect 15244 10144 15340 10184
rect 15052 10050 15092 10135
rect 15148 10109 15188 10144
rect 15340 10135 15380 10144
rect 15147 10100 15189 10109
rect 15147 10060 15148 10100
rect 15188 10060 15189 10100
rect 15147 10051 15189 10060
rect 15339 10016 15381 10025
rect 15339 9976 15340 10016
rect 15380 9976 15381 10016
rect 15339 9967 15381 9976
rect 15243 9932 15285 9941
rect 15243 9892 15244 9932
rect 15284 9892 15285 9932
rect 15243 9883 15285 9892
rect 14955 9764 14997 9773
rect 14955 9724 14956 9764
rect 14996 9724 14997 9764
rect 14955 9715 14997 9724
rect 14764 9598 14996 9638
rect 14763 9512 14805 9521
rect 14763 9472 14764 9512
rect 14804 9472 14805 9512
rect 14763 9463 14805 9472
rect 14764 9378 14804 9463
rect 14859 8756 14901 8765
rect 14859 8716 14860 8756
rect 14900 8716 14901 8756
rect 14859 8707 14901 8716
rect 14860 8672 14900 8707
rect 14860 8621 14900 8632
rect 14956 8504 14996 9598
rect 15052 9512 15092 9521
rect 15052 9437 15092 9472
rect 15147 9512 15189 9521
rect 15147 9472 15148 9512
rect 15188 9472 15189 9512
rect 15147 9463 15189 9472
rect 15051 9428 15093 9437
rect 15051 9388 15052 9428
rect 15092 9388 15093 9428
rect 15051 9379 15093 9388
rect 15052 8924 15092 9379
rect 15148 9378 15188 9463
rect 15244 9353 15284 9883
rect 15243 9344 15285 9353
rect 15243 9304 15244 9344
rect 15284 9304 15285 9344
rect 15243 9295 15285 9304
rect 15052 8875 15092 8884
rect 15051 8756 15093 8765
rect 15051 8716 15052 8756
rect 15092 8716 15093 8756
rect 15051 8707 15093 8716
rect 14860 8464 14996 8504
rect 14763 8084 14805 8093
rect 14763 8044 14764 8084
rect 14804 8044 14805 8084
rect 14763 8035 14805 8044
rect 14764 7950 14804 8035
rect 14667 7916 14709 7925
rect 14667 7876 14668 7916
rect 14708 7876 14709 7916
rect 14667 7867 14709 7876
rect 14571 7748 14613 7757
rect 14571 7708 14572 7748
rect 14612 7708 14613 7748
rect 14571 7699 14613 7708
rect 14764 7505 14804 7507
rect 14763 7496 14805 7505
rect 14763 7456 14764 7496
rect 14804 7456 14805 7496
rect 14763 7447 14805 7456
rect 14764 7412 14804 7447
rect 14476 7372 14612 7412
rect 14283 7363 14325 7372
rect 14572 7328 14612 7372
rect 14764 7363 14804 7372
rect 14572 7288 14708 7328
rect 14285 7169 14325 7254
rect 14475 7244 14517 7253
rect 14283 7162 14325 7169
rect 14283 7160 14285 7162
rect 14283 7120 14284 7160
rect 14324 7120 14325 7122
rect 14283 7111 14325 7120
rect 14380 7204 14476 7244
rect 14516 7204 14517 7244
rect 14380 7160 14420 7204
rect 14475 7195 14517 7204
rect 14380 7111 14420 7120
rect 14572 7160 14612 7169
rect 14475 6992 14517 7001
rect 14475 6952 14476 6992
rect 14516 6952 14517 6992
rect 14475 6943 14517 6952
rect 14476 6858 14516 6943
rect 13900 6607 13940 6616
rect 13996 6700 14228 6740
rect 13996 5732 14036 6700
rect 14091 6488 14133 6497
rect 14091 6448 14092 6488
rect 14132 6448 14133 6488
rect 14091 6439 14133 6448
rect 14092 6354 14132 6439
rect 14283 6236 14325 6245
rect 14283 6196 14284 6236
rect 14324 6196 14325 6236
rect 14283 6187 14325 6196
rect 14187 5816 14229 5825
rect 14187 5776 14188 5816
rect 14228 5776 14229 5816
rect 14187 5767 14229 5776
rect 13996 5683 14036 5692
rect 14092 5648 14132 5657
rect 14092 5489 14132 5608
rect 14091 5480 14133 5489
rect 14091 5440 14092 5480
rect 14132 5440 14133 5480
rect 14091 5431 14133 5440
rect 13995 5060 14037 5069
rect 13995 5020 13996 5060
rect 14036 5020 14037 5060
rect 13995 5011 14037 5020
rect 13899 4976 13941 4985
rect 13899 4936 13900 4976
rect 13940 4936 13941 4976
rect 13899 4927 13941 4936
rect 13996 4976 14036 5011
rect 13900 4842 13940 4927
rect 13996 4925 14036 4936
rect 13803 4388 13845 4397
rect 13803 4348 13804 4388
rect 13844 4348 13845 4388
rect 13803 4339 13845 4348
rect 14091 4388 14133 4397
rect 14091 4348 14092 4388
rect 14132 4348 14133 4388
rect 14091 4339 14133 4348
rect 13899 4304 13941 4313
rect 13899 4264 13900 4304
rect 13940 4264 13941 4304
rect 13899 4255 13941 4264
rect 13900 4220 13940 4255
rect 13900 4169 13940 4180
rect 14092 4136 14132 4339
rect 14188 4313 14228 5767
rect 14187 4304 14229 4313
rect 14187 4264 14188 4304
rect 14228 4264 14229 4304
rect 14187 4255 14229 4264
rect 13612 4096 13844 4136
rect 13804 4052 13844 4096
rect 14092 4087 14132 4096
rect 13516 4012 13748 4052
rect 13804 4012 13940 4052
rect 13516 3893 13556 4012
rect 13708 3968 13748 4012
rect 13708 3919 13748 3928
rect 13504 3884 13556 3893
rect 13504 3844 13505 3884
rect 13545 3844 13556 3884
rect 13504 3835 13546 3844
rect 13803 3548 13845 3557
rect 13803 3508 13804 3548
rect 13844 3508 13845 3548
rect 13803 3499 13845 3508
rect 13900 3548 13940 4012
rect 14091 3968 14133 3977
rect 14091 3928 14092 3968
rect 14132 3928 14133 3968
rect 14091 3919 14133 3928
rect 13995 3884 14037 3893
rect 13995 3844 13996 3884
rect 14036 3844 14037 3884
rect 13995 3835 14037 3844
rect 13900 3499 13940 3508
rect 13516 3464 13556 3473
rect 13516 3053 13556 3424
rect 13804 3464 13844 3499
rect 13804 3413 13844 3424
rect 13803 3296 13845 3305
rect 13803 3256 13804 3296
rect 13844 3256 13845 3296
rect 13803 3247 13845 3256
rect 13515 3044 13557 3053
rect 13515 3004 13516 3044
rect 13556 3004 13557 3044
rect 13515 2995 13557 3004
rect 13132 2920 13460 2960
rect 13035 2792 13077 2801
rect 13035 2752 13036 2792
rect 13076 2752 13077 2792
rect 13035 2743 13077 2752
rect 12748 2575 12788 2584
rect 12596 2500 12692 2540
rect 11691 2288 11733 2297
rect 11691 2248 11692 2288
rect 11732 2248 11733 2288
rect 11691 2239 11733 2248
rect 11691 2120 11733 2129
rect 11691 2080 11692 2120
rect 11732 2080 11733 2120
rect 11691 2071 11733 2080
rect 11980 2120 12020 2500
rect 12556 2491 12596 2500
rect 11980 2071 12020 2080
rect 11692 1986 11732 2071
rect 12171 2036 12213 2045
rect 12171 1996 12172 2036
rect 12212 1996 12213 2036
rect 12171 1987 12213 1996
rect 12172 1952 12212 1987
rect 12172 1901 12212 1912
rect 12171 1784 12213 1793
rect 12171 1744 12172 1784
rect 12212 1744 12213 1784
rect 12171 1735 12213 1744
rect 11787 1700 11829 1709
rect 11787 1660 11788 1700
rect 11828 1660 11829 1700
rect 11787 1651 11829 1660
rect 11979 1700 12021 1709
rect 11979 1660 11980 1700
rect 12020 1660 12021 1700
rect 11979 1651 12021 1660
rect 11788 80 11828 1651
rect 11980 80 12020 1651
rect 12172 80 12212 1735
rect 12555 1280 12597 1289
rect 12555 1240 12556 1280
rect 12596 1240 12597 1280
rect 12555 1231 12597 1240
rect 12747 1280 12789 1289
rect 12747 1240 12748 1280
rect 12788 1240 12789 1280
rect 12747 1231 12789 1240
rect 12844 1280 12884 1291
rect 12459 1112 12501 1121
rect 12459 1072 12460 1112
rect 12500 1072 12501 1112
rect 12459 1063 12501 1072
rect 12460 978 12500 1063
rect 12363 524 12405 533
rect 12363 484 12364 524
rect 12404 484 12405 524
rect 12363 475 12405 484
rect 12364 80 12404 475
rect 12556 80 12596 1231
rect 12748 80 12788 1231
rect 12844 1205 12884 1240
rect 12939 1280 12981 1289
rect 12939 1240 12940 1280
rect 12980 1240 12981 1280
rect 12939 1231 12981 1240
rect 12843 1196 12885 1205
rect 12843 1156 12844 1196
rect 12884 1156 12885 1196
rect 12843 1147 12885 1156
rect 12940 80 12980 1231
rect 13036 1112 13076 1121
rect 13036 365 13076 1072
rect 13035 356 13077 365
rect 13035 316 13036 356
rect 13076 316 13077 356
rect 13035 307 13077 316
rect 13132 80 13172 2920
rect 13419 2288 13461 2297
rect 13419 2248 13420 2288
rect 13460 2248 13461 2288
rect 13419 2239 13461 2248
rect 13420 1952 13460 2239
rect 13420 1903 13460 1912
rect 13804 1952 13844 3247
rect 13996 2801 14036 3835
rect 13995 2792 14037 2801
rect 13995 2752 13996 2792
rect 14036 2752 14037 2792
rect 13995 2743 14037 2752
rect 13804 1903 13844 1912
rect 13996 2624 14036 2743
rect 13996 1793 14036 2584
rect 13995 1784 14037 1793
rect 13995 1744 13996 1784
rect 14036 1744 14037 1784
rect 13995 1735 14037 1744
rect 13899 1532 13941 1541
rect 13899 1492 13900 1532
rect 13940 1492 13941 1532
rect 13899 1483 13941 1492
rect 13515 1280 13557 1289
rect 13515 1240 13516 1280
rect 13556 1240 13557 1280
rect 13515 1231 13557 1240
rect 13707 1280 13749 1289
rect 13707 1240 13708 1280
rect 13748 1240 13749 1280
rect 13707 1231 13749 1240
rect 13323 1028 13365 1037
rect 13323 988 13324 1028
rect 13364 988 13365 1028
rect 13323 979 13365 988
rect 13324 80 13364 979
rect 13516 80 13556 1231
rect 13708 80 13748 1231
rect 13900 80 13940 1483
rect 14092 80 14132 3919
rect 14187 3296 14229 3305
rect 14187 3256 14188 3296
rect 14228 3256 14229 3296
rect 14187 3247 14229 3256
rect 14188 3162 14228 3247
rect 14187 3044 14229 3053
rect 14187 3004 14188 3044
rect 14228 3004 14229 3044
rect 14187 2995 14229 3004
rect 14188 2876 14228 2995
rect 14188 2827 14228 2836
rect 14284 2540 14324 6187
rect 14572 5909 14612 7120
rect 14571 5900 14613 5909
rect 14571 5860 14572 5900
rect 14612 5860 14613 5900
rect 14571 5851 14613 5860
rect 14572 5657 14612 5742
rect 14571 5648 14613 5657
rect 14571 5608 14572 5648
rect 14612 5608 14613 5648
rect 14571 5599 14613 5608
rect 14380 4892 14420 4901
rect 14380 4565 14420 4852
rect 14475 4892 14517 4901
rect 14475 4852 14476 4892
rect 14516 4852 14517 4892
rect 14475 4843 14517 4852
rect 14476 4758 14516 4843
rect 14379 4556 14421 4565
rect 14379 4516 14380 4556
rect 14420 4516 14421 4556
rect 14379 4507 14421 4516
rect 14475 4388 14517 4397
rect 14475 4348 14476 4388
rect 14516 4348 14517 4388
rect 14475 4339 14517 4348
rect 14379 3380 14421 3389
rect 14379 3340 14380 3380
rect 14420 3340 14421 3380
rect 14379 3331 14421 3340
rect 14380 3246 14420 3331
rect 14379 2876 14421 2885
rect 14379 2836 14380 2876
rect 14420 2836 14421 2876
rect 14379 2827 14421 2836
rect 14380 2742 14420 2827
rect 14188 2500 14324 2540
rect 14188 1037 14228 2500
rect 14283 1196 14325 1205
rect 14283 1156 14284 1196
rect 14324 1156 14325 1196
rect 14283 1147 14325 1156
rect 14284 1112 14324 1147
rect 14284 1061 14324 1072
rect 14187 1028 14229 1037
rect 14187 988 14188 1028
rect 14228 988 14229 1028
rect 14187 979 14229 988
rect 14283 944 14325 953
rect 14283 904 14284 944
rect 14324 904 14325 944
rect 14283 895 14325 904
rect 14284 80 14324 895
rect 14476 80 14516 4339
rect 14668 3977 14708 7288
rect 14667 3968 14709 3977
rect 14667 3928 14668 3968
rect 14708 3928 14709 3968
rect 14667 3919 14709 3928
rect 14572 3212 14612 3221
rect 14764 3212 14804 3221
rect 14612 3172 14708 3212
rect 14572 3163 14612 3172
rect 14571 3044 14613 3053
rect 14571 3004 14572 3044
rect 14612 3004 14613 3044
rect 14571 2995 14613 3004
rect 14572 2708 14612 2995
rect 14572 2659 14612 2668
rect 14571 2372 14613 2381
rect 14571 2332 14572 2372
rect 14612 2332 14613 2372
rect 14571 2323 14613 2332
rect 14572 1280 14612 2323
rect 14668 1448 14708 3172
rect 14860 3212 14900 8464
rect 14956 8168 14996 8177
rect 15052 8168 15092 8707
rect 15244 8672 15284 9295
rect 15244 8623 15284 8632
rect 14996 8128 15092 8168
rect 14956 8119 14996 8128
rect 15148 7986 15188 7995
rect 14955 7748 14997 7757
rect 14955 7708 14956 7748
rect 14996 7708 14997 7748
rect 14955 7699 14997 7708
rect 14956 7160 14996 7699
rect 15051 7580 15093 7589
rect 15051 7540 15052 7580
rect 15092 7540 15093 7580
rect 15051 7531 15093 7540
rect 14956 7111 14996 7120
rect 15052 6404 15092 7531
rect 15148 7505 15188 7946
rect 15340 7841 15380 9967
rect 15436 8597 15476 11152
rect 15532 9689 15572 11320
rect 15531 9680 15573 9689
rect 15531 9640 15532 9680
rect 15572 9640 15573 9680
rect 15531 9631 15573 9640
rect 15532 9428 15572 9437
rect 15532 9269 15572 9388
rect 15628 9428 15668 11740
rect 15724 10445 15764 13588
rect 15820 13553 15860 14008
rect 15819 13544 15861 13553
rect 15819 13504 15820 13544
rect 15860 13504 15861 13544
rect 15819 13495 15861 13504
rect 15820 11201 15860 13495
rect 15916 13250 15956 19795
rect 16012 16409 16052 21895
rect 16108 18845 16148 22072
rect 16204 21953 16244 22912
rect 16300 22112 16340 22121
rect 16203 21944 16245 21953
rect 16203 21904 16204 21944
rect 16244 21904 16245 21944
rect 16203 21895 16245 21904
rect 16300 21608 16340 22072
rect 16252 21598 16340 21608
rect 16292 21568 16340 21598
rect 16396 21776 16436 23164
rect 16588 23120 16628 23129
rect 16252 21549 16292 21558
rect 16396 20516 16436 21736
rect 16492 23080 16588 23120
rect 16492 20777 16532 23080
rect 16588 23071 16628 23080
rect 16684 22448 16724 25087
rect 16779 23540 16821 23549
rect 16779 23500 16780 23540
rect 16820 23500 16821 23540
rect 16779 23491 16821 23500
rect 16588 22408 16724 22448
rect 16588 21776 16628 22408
rect 16780 22289 16820 23491
rect 16876 22448 16916 25432
rect 16972 25388 17012 25600
rect 16972 25339 17012 25348
rect 17068 25304 17108 25313
rect 17164 25304 17204 25675
rect 17260 25565 17300 26767
rect 17548 26766 17588 26851
rect 17356 26648 17396 26657
rect 17356 26489 17396 26608
rect 17355 26480 17397 26489
rect 17355 26440 17356 26480
rect 17396 26440 17397 26480
rect 17355 26431 17397 26440
rect 17356 26144 17396 26431
rect 17451 26312 17493 26321
rect 17451 26272 17452 26312
rect 17492 26272 17493 26312
rect 17451 26263 17493 26272
rect 17452 26178 17492 26263
rect 17548 26153 17588 26238
rect 17356 26069 17396 26104
rect 17547 26144 17589 26153
rect 17547 26104 17548 26144
rect 17588 26104 17589 26144
rect 17547 26095 17589 26104
rect 17355 26060 17397 26069
rect 17355 26020 17356 26060
rect 17396 26020 17397 26060
rect 17355 26011 17397 26020
rect 17356 25980 17396 26011
rect 17644 25976 17684 26935
rect 17740 26934 17780 27019
rect 17836 26732 17876 27112
rect 17932 26909 17972 26994
rect 17931 26900 17973 26909
rect 17931 26860 17932 26900
rect 17972 26860 17973 26900
rect 17931 26851 17973 26860
rect 17836 26692 17972 26732
rect 17835 26564 17877 26573
rect 17835 26524 17836 26564
rect 17876 26524 17877 26564
rect 17835 26515 17877 26524
rect 17740 26144 17780 26153
rect 17740 26069 17780 26104
rect 17739 26060 17781 26069
rect 17739 26020 17740 26060
rect 17780 26020 17781 26060
rect 17739 26011 17781 26020
rect 17452 25936 17684 25976
rect 17259 25556 17301 25565
rect 17259 25516 17260 25556
rect 17300 25516 17301 25556
rect 17259 25507 17301 25516
rect 17452 25472 17492 25936
rect 17740 25901 17780 26011
rect 17739 25892 17781 25901
rect 17739 25852 17740 25892
rect 17780 25852 17781 25892
rect 17739 25843 17781 25852
rect 17547 25808 17589 25817
rect 17547 25768 17548 25808
rect 17588 25768 17589 25808
rect 17547 25759 17589 25768
rect 17548 25481 17588 25759
rect 17108 25264 17204 25304
rect 17356 25432 17492 25472
rect 17547 25472 17589 25481
rect 17547 25432 17548 25472
rect 17588 25432 17589 25472
rect 17068 25255 17108 25264
rect 17260 25220 17300 25229
rect 17356 25220 17396 25432
rect 17547 25423 17589 25432
rect 17451 25304 17493 25313
rect 17451 25264 17452 25304
rect 17492 25264 17493 25304
rect 17451 25255 17493 25264
rect 17300 25180 17396 25220
rect 17260 25171 17300 25180
rect 17452 25061 17492 25255
rect 17451 25052 17493 25061
rect 17451 25012 17452 25052
rect 17492 25012 17493 25052
rect 17451 25003 17493 25012
rect 17259 24632 17301 24641
rect 17259 24592 17260 24632
rect 17300 24592 17301 24632
rect 17259 24583 17301 24592
rect 16876 22408 17012 22448
rect 16684 22280 16724 22289
rect 16684 21953 16724 22240
rect 16779 22280 16821 22289
rect 16779 22240 16780 22280
rect 16820 22240 16821 22280
rect 16779 22231 16821 22240
rect 16876 22280 16916 22289
rect 16780 22112 16820 22121
rect 16683 21944 16725 21953
rect 16683 21904 16684 21944
rect 16724 21904 16725 21944
rect 16683 21895 16725 21904
rect 16588 21736 16724 21776
rect 16587 21608 16629 21617
rect 16587 21568 16588 21608
rect 16628 21568 16629 21608
rect 16587 21559 16629 21568
rect 16588 21474 16628 21559
rect 16491 20768 16533 20777
rect 16491 20728 16492 20768
rect 16532 20728 16533 20768
rect 16491 20719 16533 20728
rect 16396 20476 16532 20516
rect 16395 20348 16437 20357
rect 16395 20308 16396 20348
rect 16436 20308 16437 20348
rect 16395 20299 16437 20308
rect 16107 18836 16149 18845
rect 16107 18796 16108 18836
rect 16148 18796 16149 18836
rect 16107 18787 16149 18796
rect 16108 18509 16148 18787
rect 16204 18584 16244 18593
rect 16107 18500 16149 18509
rect 16107 18460 16108 18500
rect 16148 18460 16149 18500
rect 16107 18451 16149 18460
rect 16204 18257 16244 18544
rect 16203 18248 16245 18257
rect 16203 18208 16204 18248
rect 16244 18208 16245 18248
rect 16203 18199 16245 18208
rect 16396 17081 16436 20299
rect 16492 20189 16532 20476
rect 16491 20180 16533 20189
rect 16684 20180 16724 21736
rect 16780 21449 16820 22072
rect 16876 21533 16916 22240
rect 16875 21524 16917 21533
rect 16875 21484 16876 21524
rect 16916 21484 16917 21524
rect 16875 21475 16917 21484
rect 16779 21440 16821 21449
rect 16779 21400 16780 21440
rect 16820 21400 16821 21440
rect 16779 21391 16821 21400
rect 16972 20264 17012 22408
rect 17068 22280 17108 22289
rect 17068 21029 17108 22240
rect 17163 22280 17205 22289
rect 17163 22240 17164 22280
rect 17204 22240 17205 22280
rect 17163 22231 17205 22240
rect 17164 22146 17204 22231
rect 17260 21281 17300 24583
rect 17451 23624 17493 23633
rect 17451 23584 17452 23624
rect 17492 23584 17493 23624
rect 17451 23575 17493 23584
rect 17355 22112 17397 22121
rect 17355 22072 17356 22112
rect 17396 22072 17397 22112
rect 17355 22063 17397 22072
rect 17356 21978 17396 22063
rect 17452 21860 17492 23575
rect 17356 21820 17492 21860
rect 17259 21272 17301 21281
rect 17259 21232 17260 21272
rect 17300 21232 17301 21272
rect 17259 21223 17301 21232
rect 17163 21104 17205 21113
rect 17163 21064 17164 21104
rect 17204 21064 17205 21104
rect 17163 21055 17205 21064
rect 17067 21020 17109 21029
rect 17067 20980 17068 21020
rect 17108 20980 17109 21020
rect 17067 20971 17109 20980
rect 17068 20768 17108 20777
rect 17164 20768 17204 21055
rect 17259 21020 17301 21029
rect 17259 20980 17260 21020
rect 17300 20980 17301 21020
rect 17259 20971 17301 20980
rect 17260 20886 17300 20971
rect 17108 20728 17204 20768
rect 17068 20719 17108 20728
rect 17356 20357 17396 21820
rect 17548 21785 17588 25423
rect 17739 25220 17781 25229
rect 17739 25180 17740 25220
rect 17780 25180 17781 25220
rect 17739 25171 17781 25180
rect 17740 24632 17780 25171
rect 17644 24592 17740 24632
rect 17644 23213 17684 24592
rect 17740 24583 17780 24592
rect 17836 24557 17876 26515
rect 17932 24884 17972 26692
rect 18028 25229 18068 28288
rect 18124 27068 18164 30463
rect 18220 27152 18260 31900
rect 18411 31520 18453 31529
rect 18411 31480 18412 31520
rect 18452 31480 18453 31520
rect 18411 31471 18453 31480
rect 18412 31386 18452 31471
rect 18604 29177 18644 32563
rect 18700 31688 18740 32992
rect 19276 32982 19316 33067
rect 19948 33032 19988 33041
rect 19852 32948 19892 32957
rect 19755 32864 19797 32873
rect 19755 32824 19756 32864
rect 19796 32824 19797 32864
rect 19755 32815 19797 32824
rect 19275 32780 19317 32789
rect 19468 32780 19508 32789
rect 19275 32740 19276 32780
rect 19316 32740 19317 32780
rect 19275 32731 19317 32740
rect 19372 32740 19468 32780
rect 18808 31772 19176 31781
rect 18848 31732 18890 31772
rect 18930 31732 18972 31772
rect 19012 31732 19054 31772
rect 19094 31732 19136 31772
rect 18808 31723 19176 31732
rect 18700 31648 18774 31688
rect 18734 31367 18774 31648
rect 19276 31604 19316 32731
rect 19084 31564 19316 31604
rect 18734 31318 18774 31327
rect 18892 31352 18932 31361
rect 18892 31109 18932 31312
rect 18988 31352 19028 31361
rect 19084 31352 19124 31564
rect 19276 31361 19316 31446
rect 19028 31312 19124 31352
rect 19180 31352 19220 31361
rect 18988 31303 19028 31312
rect 19083 31184 19125 31193
rect 19083 31144 19084 31184
rect 19124 31144 19125 31184
rect 19083 31135 19125 31144
rect 18891 31100 18933 31109
rect 18891 31060 18892 31100
rect 18932 31060 18933 31100
rect 18891 31051 18933 31060
rect 19084 31050 19124 31135
rect 19180 30857 19220 31312
rect 19275 31352 19317 31361
rect 19275 31312 19276 31352
rect 19316 31312 19317 31352
rect 19275 31303 19317 31312
rect 19372 31184 19412 32740
rect 19468 32731 19508 32740
rect 19756 32730 19796 32815
rect 19852 32360 19892 32908
rect 19564 32320 19892 32360
rect 19468 32201 19508 32286
rect 19467 32192 19509 32201
rect 19467 32152 19468 32192
rect 19508 32152 19509 32192
rect 19467 32143 19509 32152
rect 19564 32024 19604 32320
rect 19948 32276 19988 32992
rect 20044 32948 20084 33151
rect 20908 32957 20948 37687
rect 20044 32873 20084 32908
rect 20139 32948 20181 32957
rect 20139 32908 20140 32948
rect 20180 32908 20181 32948
rect 20139 32906 20181 32908
rect 20139 32899 20140 32906
rect 20043 32864 20085 32873
rect 20043 32824 20044 32864
rect 20084 32824 20085 32864
rect 20043 32815 20085 32824
rect 20180 32899 20181 32906
rect 20907 32948 20949 32957
rect 20907 32908 20908 32948
rect 20948 32908 20949 32948
rect 20907 32899 20949 32908
rect 20140 32789 20180 32866
rect 20619 32864 20661 32873
rect 20619 32824 20620 32864
rect 20660 32824 20661 32864
rect 20619 32815 20661 32824
rect 20139 32780 20181 32789
rect 20139 32740 20140 32780
rect 20180 32740 20181 32780
rect 20139 32731 20181 32740
rect 20048 32528 20416 32537
rect 20088 32488 20130 32528
rect 20170 32488 20212 32528
rect 20252 32488 20294 32528
rect 20334 32488 20376 32528
rect 20048 32479 20416 32488
rect 19468 31984 19604 32024
rect 19756 32236 19988 32276
rect 19468 31529 19508 31984
rect 19660 31940 19700 31949
rect 19564 31900 19660 31940
rect 19467 31520 19509 31529
rect 19467 31480 19468 31520
rect 19508 31480 19509 31520
rect 19467 31471 19509 31480
rect 19564 31436 19604 31900
rect 19660 31891 19700 31900
rect 19564 31361 19604 31396
rect 19660 31520 19700 31529
rect 19468 31352 19508 31361
rect 19468 31193 19508 31312
rect 19563 31352 19605 31361
rect 19563 31312 19564 31352
rect 19604 31312 19605 31352
rect 19563 31303 19605 31312
rect 19564 31272 19604 31303
rect 19276 31144 19412 31184
rect 19467 31184 19509 31193
rect 19467 31144 19468 31184
rect 19508 31144 19509 31184
rect 19179 30848 19221 30857
rect 19179 30808 19180 30848
rect 19220 30808 19221 30848
rect 19179 30799 19221 30808
rect 18808 30260 19176 30269
rect 18848 30220 18890 30260
rect 18930 30220 18972 30260
rect 19012 30220 19054 30260
rect 19094 30220 19136 30260
rect 18808 30211 19176 30220
rect 19276 30092 19316 31144
rect 19467 31135 19509 31144
rect 19564 30764 19604 30775
rect 19564 30689 19604 30724
rect 19371 30680 19413 30689
rect 19371 30640 19372 30680
rect 19412 30640 19413 30680
rect 19371 30631 19413 30640
rect 19563 30680 19605 30689
rect 19563 30640 19564 30680
rect 19604 30640 19605 30680
rect 19563 30631 19605 30640
rect 19372 30546 19412 30631
rect 19180 30052 19316 30092
rect 19084 29840 19124 29849
rect 19084 29177 19124 29800
rect 18315 29168 18357 29177
rect 18315 29128 18316 29168
rect 18356 29128 18357 29168
rect 18315 29119 18357 29128
rect 18603 29168 18645 29177
rect 18603 29128 18604 29168
rect 18644 29128 18645 29168
rect 18603 29119 18645 29128
rect 19083 29168 19125 29177
rect 19083 29128 19084 29168
rect 19124 29128 19125 29168
rect 19083 29119 19125 29128
rect 19180 29168 19220 30052
rect 19564 29840 19604 29849
rect 19276 29756 19316 29765
rect 19564 29756 19604 29800
rect 19316 29716 19604 29756
rect 19276 29707 19316 29716
rect 19660 29588 19700 31480
rect 19756 31436 19796 32236
rect 19851 32108 19893 32117
rect 19851 32068 19852 32108
rect 19892 32068 19893 32108
rect 19851 32059 19893 32068
rect 19852 31974 19892 32059
rect 20043 31940 20085 31949
rect 20043 31900 20044 31940
rect 20084 31900 20085 31940
rect 20043 31891 20085 31900
rect 20044 31806 20084 31891
rect 19756 31387 19796 31396
rect 20043 31436 20085 31445
rect 20043 31396 20044 31436
rect 20084 31396 20085 31436
rect 20043 31387 20085 31396
rect 19852 31352 19892 31361
rect 19755 30932 19797 30941
rect 19755 30892 19756 30932
rect 19796 30892 19797 30932
rect 19755 30883 19797 30892
rect 19756 30680 19796 30883
rect 19852 30848 19892 31312
rect 20044 31302 20084 31387
rect 20236 31184 20276 31193
rect 20276 31144 20564 31184
rect 20236 31135 20276 31144
rect 20048 31016 20416 31025
rect 20088 30976 20130 31016
rect 20170 30976 20212 31016
rect 20252 30976 20294 31016
rect 20334 30976 20376 31016
rect 20048 30967 20416 30976
rect 20044 30848 20084 30857
rect 19852 30808 20044 30848
rect 20044 30799 20084 30808
rect 19756 30631 19796 30640
rect 19851 30680 19893 30689
rect 19851 30640 19852 30680
rect 19892 30640 19893 30680
rect 19851 30631 19893 30640
rect 20044 30680 20084 30691
rect 19852 30546 19892 30631
rect 20044 30605 20084 30640
rect 20043 30596 20085 30605
rect 20043 30556 20044 30596
rect 20084 30556 20085 30596
rect 20043 30547 20085 30556
rect 20235 30008 20277 30017
rect 20235 29968 20236 30008
rect 20276 29968 20277 30008
rect 20235 29959 20277 29968
rect 20236 29874 20276 29959
rect 19852 29840 19892 29849
rect 19180 29119 19220 29128
rect 19276 29548 19700 29588
rect 19756 29800 19852 29840
rect 18316 29034 18356 29119
rect 18700 29084 18740 29093
rect 18508 29000 18548 29009
rect 18548 28960 18644 29000
rect 18508 28951 18548 28960
rect 18412 28328 18452 28337
rect 18412 27824 18452 28288
rect 18507 28328 18549 28337
rect 18507 28288 18508 28328
rect 18548 28288 18549 28328
rect 18507 28279 18549 28288
rect 18508 28194 18548 28279
rect 18604 28001 18644 28960
rect 18700 28673 18740 29044
rect 18891 29000 18933 29009
rect 18891 28960 18892 29000
rect 18932 28960 18933 29000
rect 18891 28951 18933 28960
rect 18892 28866 18932 28951
rect 18808 28748 19176 28757
rect 18848 28708 18890 28748
rect 18930 28708 18972 28748
rect 19012 28708 19054 28748
rect 19094 28708 19136 28748
rect 18808 28699 19176 28708
rect 18699 28664 18741 28673
rect 18699 28624 18700 28664
rect 18740 28624 18741 28664
rect 18699 28615 18741 28624
rect 18988 28328 19028 28337
rect 18603 27992 18645 28001
rect 18603 27952 18604 27992
rect 18644 27952 18645 27992
rect 18603 27943 18645 27952
rect 18412 27784 18740 27824
rect 18316 27572 18356 27581
rect 18316 27329 18356 27532
rect 18412 27572 18452 27583
rect 18412 27497 18452 27532
rect 18603 27572 18645 27581
rect 18603 27532 18604 27572
rect 18644 27532 18645 27572
rect 18603 27523 18645 27532
rect 18411 27488 18453 27497
rect 18411 27448 18412 27488
rect 18452 27448 18453 27488
rect 18411 27439 18453 27448
rect 18315 27320 18357 27329
rect 18315 27280 18316 27320
rect 18356 27280 18357 27320
rect 18315 27271 18357 27280
rect 18220 27112 18356 27152
rect 18124 27019 18164 27028
rect 18316 26911 18356 27112
rect 18316 26862 18356 26871
rect 18412 26816 18452 27439
rect 18316 26776 18452 26816
rect 18508 26984 18548 26993
rect 18219 26564 18261 26573
rect 18219 26524 18220 26564
rect 18260 26524 18261 26564
rect 18219 26515 18261 26524
rect 18220 25481 18260 26515
rect 18219 25472 18261 25481
rect 18219 25432 18220 25472
rect 18260 25432 18261 25472
rect 18219 25423 18261 25432
rect 18027 25220 18069 25229
rect 18027 25180 18028 25220
rect 18068 25180 18069 25220
rect 18027 25171 18069 25180
rect 18316 25061 18356 26776
rect 18411 26648 18453 26657
rect 18508 26648 18548 26944
rect 18411 26608 18412 26648
rect 18452 26608 18548 26648
rect 18604 26648 18644 27523
rect 18700 27077 18740 27784
rect 18891 27656 18933 27665
rect 18891 27616 18892 27656
rect 18932 27616 18933 27656
rect 18891 27607 18933 27616
rect 18892 27522 18932 27607
rect 18988 27404 19028 28288
rect 19276 27749 19316 29548
rect 19756 29000 19796 29800
rect 19852 29791 19892 29800
rect 19948 29756 19988 29765
rect 19564 28960 19796 29000
rect 19851 29000 19893 29009
rect 19851 28960 19852 29000
rect 19892 28960 19893 29000
rect 19371 28916 19413 28925
rect 19371 28876 19372 28916
rect 19412 28876 19413 28916
rect 19371 28867 19413 28876
rect 19372 28085 19412 28867
rect 19468 28333 19508 28342
rect 19371 28076 19413 28085
rect 19371 28036 19372 28076
rect 19412 28036 19413 28076
rect 19371 28027 19413 28036
rect 19468 28001 19508 28293
rect 19467 27992 19509 28001
rect 19467 27952 19468 27992
rect 19508 27952 19509 27992
rect 19467 27943 19509 27952
rect 19371 27908 19413 27917
rect 19371 27868 19372 27908
rect 19412 27868 19413 27908
rect 19371 27859 19413 27868
rect 19275 27740 19317 27749
rect 19275 27700 19276 27740
rect 19316 27700 19317 27740
rect 19275 27691 19317 27700
rect 19372 27651 19412 27859
rect 19564 27740 19604 28960
rect 19851 28951 19893 28960
rect 19852 28866 19892 28951
rect 19852 28421 19892 28506
rect 19851 28412 19893 28421
rect 19851 28372 19852 28412
rect 19892 28372 19893 28412
rect 19851 28363 19893 28372
rect 19660 28244 19700 28253
rect 19948 28244 19988 29716
rect 20048 29504 20416 29513
rect 20088 29464 20130 29504
rect 20170 29464 20212 29504
rect 20252 29464 20294 29504
rect 20334 29464 20376 29504
rect 20048 29455 20416 29464
rect 20524 28505 20564 31144
rect 20620 31109 20660 32815
rect 21003 32276 21045 32285
rect 21003 32236 21004 32276
rect 21044 32236 21045 32276
rect 21003 32227 21045 32236
rect 20619 31100 20661 31109
rect 20619 31060 20620 31100
rect 20660 31060 20661 31100
rect 20619 31051 20661 31060
rect 20523 28496 20565 28505
rect 20523 28456 20524 28496
rect 20564 28456 20565 28496
rect 20523 28447 20565 28456
rect 19700 28204 19988 28244
rect 19660 28195 19700 28204
rect 20044 28160 20084 28169
rect 19564 27691 19604 27700
rect 19948 28120 20044 28160
rect 19372 27602 19412 27611
rect 19948 27581 19988 28120
rect 20044 28111 20084 28120
rect 20048 27992 20416 28001
rect 20088 27952 20130 27992
rect 20170 27952 20212 27992
rect 20252 27952 20294 27992
rect 20334 27952 20376 27992
rect 20048 27943 20416 27952
rect 20127 27643 20167 27652
rect 19755 27572 19797 27581
rect 19755 27532 19756 27572
rect 19796 27532 19797 27572
rect 19755 27523 19797 27532
rect 19947 27572 19989 27581
rect 19947 27532 19948 27572
rect 19988 27532 19989 27572
rect 19947 27523 19989 27532
rect 19756 27438 19796 27523
rect 20127 27413 20167 27603
rect 19948 27404 19988 27413
rect 18988 27364 19316 27404
rect 18808 27236 19176 27245
rect 18848 27196 18890 27236
rect 18930 27196 18972 27236
rect 19012 27196 19054 27236
rect 19094 27196 19136 27236
rect 18808 27187 19176 27196
rect 19276 27161 19316 27364
rect 19275 27152 19317 27161
rect 19275 27112 19276 27152
rect 19316 27112 19317 27152
rect 19275 27103 19317 27112
rect 19948 27077 19988 27364
rect 20126 27404 20168 27413
rect 20126 27364 20127 27404
rect 20167 27364 20168 27404
rect 20126 27355 20168 27364
rect 20235 27404 20277 27413
rect 20235 27364 20236 27404
rect 20276 27364 20277 27404
rect 20235 27355 20277 27364
rect 20236 27270 20276 27355
rect 18699 27068 18741 27077
rect 18699 27028 18700 27068
rect 18740 27028 18741 27068
rect 18699 27019 18741 27028
rect 19947 27068 19989 27077
rect 19947 27028 19948 27068
rect 19988 27028 19989 27068
rect 19947 27019 19989 27028
rect 18795 26984 18837 26993
rect 18795 26944 18796 26984
rect 18836 26944 18837 26984
rect 18795 26935 18837 26944
rect 18699 26900 18741 26909
rect 18699 26860 18700 26900
rect 18740 26860 18741 26900
rect 18699 26851 18741 26860
rect 18700 26816 18740 26851
rect 18700 26765 18740 26776
rect 18796 26816 18836 26935
rect 19564 26900 19604 26911
rect 18988 26816 19028 26825
rect 19180 26816 19220 26825
rect 18796 26767 18836 26776
rect 18892 26776 18988 26816
rect 19028 26776 19180 26816
rect 18604 26608 18740 26648
rect 18411 26599 18453 26608
rect 18411 26480 18453 26489
rect 18411 26440 18412 26480
rect 18452 26440 18453 26480
rect 18411 26431 18453 26440
rect 18315 25052 18357 25061
rect 18315 25012 18316 25052
rect 18356 25012 18357 25052
rect 18315 25003 18357 25012
rect 18027 24884 18069 24893
rect 17932 24844 18028 24884
rect 18068 24844 18069 24884
rect 18027 24835 18069 24844
rect 17932 24716 17972 24727
rect 17932 24641 17972 24676
rect 17931 24632 17973 24641
rect 17931 24592 17932 24632
rect 17972 24592 17973 24632
rect 17931 24583 17973 24592
rect 17835 24548 17877 24557
rect 17835 24508 17836 24548
rect 17876 24508 17877 24548
rect 17835 24499 17877 24508
rect 17931 23960 17973 23969
rect 17931 23920 17932 23960
rect 17972 23920 17973 23960
rect 17931 23911 17973 23920
rect 17739 23876 17781 23885
rect 17739 23836 17740 23876
rect 17780 23836 17781 23876
rect 17739 23827 17781 23836
rect 17643 23204 17685 23213
rect 17643 23164 17644 23204
rect 17684 23164 17685 23204
rect 17643 23155 17685 23164
rect 17643 22616 17685 22625
rect 17643 22576 17644 22616
rect 17684 22576 17685 22616
rect 17643 22567 17685 22576
rect 17644 22280 17684 22567
rect 17644 22231 17684 22240
rect 17740 22280 17780 23827
rect 17835 23792 17877 23801
rect 17835 23752 17836 23792
rect 17876 23752 17877 23792
rect 17835 23743 17877 23752
rect 17836 23658 17876 23743
rect 17835 23204 17877 23213
rect 17835 23164 17836 23204
rect 17876 23164 17877 23204
rect 17835 23155 17877 23164
rect 17836 23120 17876 23155
rect 17836 23069 17876 23080
rect 17932 22448 17972 23911
rect 18028 23801 18068 24835
rect 18219 24716 18261 24725
rect 18202 24676 18220 24716
rect 18260 24676 18261 24716
rect 18202 24667 18261 24676
rect 18202 24647 18242 24667
rect 18202 24598 18242 24607
rect 18027 23792 18069 23801
rect 18027 23752 18028 23792
rect 18068 23752 18069 23792
rect 18027 23743 18069 23752
rect 18124 23792 18164 23801
rect 18028 23288 18068 23297
rect 18124 23288 18164 23752
rect 18316 23633 18356 25003
rect 18412 23969 18452 26431
rect 18507 26396 18549 26405
rect 18507 26356 18508 26396
rect 18548 26356 18549 26396
rect 18507 26347 18549 26356
rect 18508 25649 18548 26347
rect 18507 25640 18549 25649
rect 18507 25600 18508 25640
rect 18548 25600 18549 25640
rect 18507 25591 18549 25600
rect 18508 25136 18548 25591
rect 18700 25565 18740 26608
rect 18892 25901 18932 26776
rect 18988 26767 19028 26776
rect 19180 26767 19220 26776
rect 19372 26816 19412 26827
rect 19564 26825 19604 26860
rect 19948 26900 19988 26909
rect 19372 26741 19412 26776
rect 19563 26816 19605 26825
rect 19563 26776 19564 26816
rect 19604 26776 19605 26816
rect 19563 26767 19605 26776
rect 19371 26732 19413 26741
rect 19371 26692 19372 26732
rect 19412 26692 19413 26732
rect 19371 26683 19413 26692
rect 18988 26648 19028 26657
rect 18988 26321 19028 26608
rect 19276 26648 19316 26657
rect 18987 26312 19029 26321
rect 18987 26272 18988 26312
rect 19028 26272 19029 26312
rect 18987 26263 19029 26272
rect 18987 26144 19029 26153
rect 18987 26104 18988 26144
rect 19028 26104 19029 26144
rect 18987 26095 19029 26104
rect 18988 26010 19028 26095
rect 19180 25901 19220 25986
rect 18891 25892 18933 25901
rect 18891 25852 18892 25892
rect 18932 25852 18933 25892
rect 18891 25843 18933 25852
rect 19179 25892 19221 25901
rect 19179 25852 19180 25892
rect 19220 25852 19221 25892
rect 19179 25843 19221 25852
rect 18808 25724 19176 25733
rect 18848 25684 18890 25724
rect 18930 25684 18972 25724
rect 19012 25684 19054 25724
rect 19094 25684 19136 25724
rect 18808 25675 19176 25684
rect 18699 25556 18741 25565
rect 18699 25516 18700 25556
rect 18740 25516 18741 25556
rect 18699 25507 18741 25516
rect 18987 25556 19029 25565
rect 18987 25516 18988 25556
rect 19028 25516 19029 25556
rect 18987 25507 19029 25516
rect 18891 25472 18933 25481
rect 18891 25432 18892 25472
rect 18932 25432 18933 25472
rect 18891 25423 18933 25432
rect 18700 25304 18740 25313
rect 18892 25304 18932 25423
rect 18740 25264 18932 25304
rect 18988 25304 19028 25507
rect 19276 25481 19316 26608
rect 19756 26648 19796 26657
rect 19796 26608 19892 26648
rect 19756 26599 19796 26608
rect 19755 26312 19797 26321
rect 19755 26272 19756 26312
rect 19796 26272 19797 26312
rect 19755 26263 19797 26272
rect 19372 26144 19412 26153
rect 19275 25472 19317 25481
rect 18700 25255 18740 25264
rect 18508 25096 18740 25136
rect 18603 24716 18645 24725
rect 18603 24676 18604 24716
rect 18644 24676 18645 24716
rect 18603 24667 18645 24676
rect 18508 24632 18548 24641
rect 18411 23960 18453 23969
rect 18411 23920 18412 23960
rect 18452 23920 18453 23960
rect 18411 23911 18453 23920
rect 18508 23885 18548 24592
rect 18604 24582 18644 24667
rect 18507 23876 18549 23885
rect 18507 23836 18508 23876
rect 18548 23836 18549 23876
rect 18507 23827 18549 23836
rect 18411 23792 18453 23801
rect 18411 23752 18412 23792
rect 18452 23752 18453 23792
rect 18411 23743 18453 23752
rect 18412 23658 18452 23743
rect 18507 23708 18549 23717
rect 18507 23668 18508 23708
rect 18548 23668 18549 23708
rect 18507 23659 18549 23668
rect 18315 23624 18357 23633
rect 18315 23584 18316 23624
rect 18356 23584 18357 23624
rect 18315 23575 18357 23584
rect 18508 23574 18548 23659
rect 18068 23248 18164 23288
rect 18028 23239 18068 23248
rect 18411 23120 18453 23129
rect 18411 23080 18412 23120
rect 18452 23080 18453 23120
rect 18411 23071 18453 23080
rect 18412 22986 18452 23071
rect 18219 22952 18261 22961
rect 18219 22912 18220 22952
rect 18260 22912 18261 22952
rect 18219 22903 18261 22912
rect 18028 22868 18068 22877
rect 18028 22625 18068 22828
rect 18027 22616 18069 22625
rect 18027 22576 18028 22616
rect 18068 22576 18069 22616
rect 18027 22567 18069 22576
rect 17932 22408 18068 22448
rect 17932 22280 17972 22289
rect 17740 22240 17932 22280
rect 17547 21776 17589 21785
rect 17547 21736 17548 21776
rect 17588 21736 17589 21776
rect 17547 21727 17589 21736
rect 17451 21608 17493 21617
rect 17451 21568 17452 21608
rect 17492 21568 17493 21608
rect 17451 21559 17493 21568
rect 17452 20768 17492 21559
rect 17740 21197 17780 22240
rect 17932 22231 17972 22240
rect 18028 22280 18068 22408
rect 18220 22280 18260 22903
rect 18316 22457 18356 22542
rect 18315 22448 18357 22457
rect 18315 22408 18316 22448
rect 18356 22408 18357 22448
rect 18315 22399 18357 22408
rect 18507 22280 18549 22289
rect 18220 22240 18452 22280
rect 18028 22231 18068 22240
rect 18315 22112 18357 22121
rect 18315 22072 18316 22112
rect 18356 22072 18357 22112
rect 18315 22063 18357 22072
rect 17835 22028 17877 22037
rect 17835 21988 17836 22028
rect 17876 21988 17877 22028
rect 17835 21979 17877 21988
rect 17836 21608 17876 21979
rect 17836 21559 17876 21568
rect 18220 21608 18260 21617
rect 18028 21449 18068 21480
rect 18220 21449 18260 21568
rect 18316 21608 18356 22063
rect 18412 21776 18452 22240
rect 18507 22240 18508 22280
rect 18548 22240 18549 22280
rect 18507 22231 18549 22240
rect 18508 22146 18548 22231
rect 18508 21776 18548 21785
rect 18412 21736 18508 21776
rect 18508 21727 18548 21736
rect 18316 21559 18356 21568
rect 18411 21608 18453 21617
rect 18411 21568 18412 21608
rect 18452 21568 18453 21608
rect 18411 21559 18453 21568
rect 18700 21608 18740 25096
rect 18988 24641 19028 25264
rect 19180 25432 19276 25472
rect 19316 25432 19317 25472
rect 19180 24800 19220 25432
rect 19275 25423 19317 25432
rect 19372 25388 19412 26104
rect 19756 26144 19796 26263
rect 19756 26095 19796 26104
rect 19468 26060 19508 26069
rect 19468 25901 19508 26020
rect 19660 26060 19700 26069
rect 19564 25976 19604 25985
rect 19467 25892 19509 25901
rect 19467 25852 19468 25892
rect 19508 25852 19509 25892
rect 19467 25843 19509 25852
rect 19468 25556 19508 25843
rect 19564 25733 19604 25936
rect 19660 25808 19700 26020
rect 19852 25985 19892 26608
rect 19948 26573 19988 26860
rect 20140 26648 20180 26657
rect 20180 26608 20564 26648
rect 20140 26599 20180 26608
rect 19947 26564 19989 26573
rect 19947 26524 19948 26564
rect 19988 26524 19989 26564
rect 19947 26515 19989 26524
rect 20048 26480 20416 26489
rect 20088 26440 20130 26480
rect 20170 26440 20212 26480
rect 20252 26440 20294 26480
rect 20334 26440 20376 26480
rect 20048 26431 20416 26440
rect 19947 26060 19989 26069
rect 19947 26020 19948 26060
rect 19988 26020 19989 26060
rect 19947 26011 19989 26020
rect 19851 25976 19893 25985
rect 19851 25936 19852 25976
rect 19892 25936 19893 25976
rect 19851 25927 19893 25936
rect 19948 25926 19988 26011
rect 20524 25985 20564 26608
rect 20523 25976 20565 25985
rect 20523 25936 20524 25976
rect 20564 25936 20565 25976
rect 20523 25927 20565 25936
rect 20140 25892 20180 25901
rect 20180 25852 20372 25892
rect 20140 25843 20180 25852
rect 19660 25768 20084 25808
rect 19563 25724 19605 25733
rect 19563 25684 19564 25724
rect 19604 25684 19605 25724
rect 19563 25675 19605 25684
rect 19660 25565 19700 25650
rect 19659 25556 19701 25565
rect 19468 25516 19604 25556
rect 19564 25388 19604 25516
rect 19659 25516 19660 25556
rect 19700 25516 19701 25556
rect 19659 25507 19701 25516
rect 19851 25472 19893 25481
rect 19851 25432 19852 25472
rect 19892 25432 19893 25472
rect 19851 25423 19893 25432
rect 20044 25472 20084 25768
rect 20129 25556 20171 25565
rect 20129 25516 20130 25556
rect 20170 25516 20171 25556
rect 20129 25507 20171 25516
rect 20044 25423 20084 25432
rect 19372 25348 19508 25388
rect 19564 25348 19700 25388
rect 19275 25304 19317 25313
rect 19275 25264 19276 25304
rect 19316 25264 19317 25304
rect 19275 25255 19317 25264
rect 19276 25170 19316 25255
rect 19372 25220 19412 25231
rect 19372 25145 19412 25180
rect 19371 25136 19413 25145
rect 19371 25096 19372 25136
rect 19412 25096 19413 25136
rect 19371 25087 19413 25096
rect 19468 24800 19508 25348
rect 19563 25220 19605 25229
rect 19563 25180 19564 25220
rect 19604 25180 19605 25220
rect 19563 25171 19605 25180
rect 19180 24760 19412 24800
rect 18987 24632 19029 24641
rect 18987 24592 18988 24632
rect 19028 24592 19029 24632
rect 19275 24632 19317 24641
rect 18987 24583 19029 24592
rect 19118 24617 19158 24626
rect 19275 24592 19276 24632
rect 19316 24592 19317 24632
rect 19275 24583 19317 24592
rect 19372 24632 19412 24760
rect 19468 24751 19508 24760
rect 19372 24583 19412 24592
rect 19564 24632 19604 25171
rect 19564 24583 19604 24592
rect 19660 24632 19700 25348
rect 19852 25304 19892 25423
rect 19947 25388 19989 25397
rect 19947 25348 19948 25388
rect 19988 25348 19989 25388
rect 19947 25339 19989 25348
rect 20130 25388 20170 25507
rect 20130 25339 20170 25348
rect 19852 25255 19892 25264
rect 19948 24641 19988 25339
rect 20236 25313 20276 25398
rect 20235 25304 20277 25313
rect 20235 25264 20236 25304
rect 20276 25264 20277 25304
rect 20235 25255 20277 25264
rect 20332 25145 20372 25852
rect 20331 25136 20373 25145
rect 20331 25096 20332 25136
rect 20372 25096 20373 25136
rect 20331 25087 20373 25096
rect 20048 24968 20416 24977
rect 20088 24928 20130 24968
rect 20170 24928 20212 24968
rect 20252 24928 20294 24968
rect 20334 24928 20376 24968
rect 20048 24919 20416 24928
rect 19660 24583 19700 24592
rect 19947 24632 19989 24641
rect 19947 24592 19948 24632
rect 19988 24592 19989 24632
rect 19947 24583 19989 24592
rect 18892 24464 18932 24473
rect 19118 24464 19158 24577
rect 19276 24498 19316 24583
rect 19851 24548 19893 24557
rect 19851 24508 19852 24548
rect 19892 24508 19893 24548
rect 19851 24499 19893 24508
rect 18932 24424 19158 24464
rect 18892 24415 18932 24424
rect 19852 24414 19892 24499
rect 20043 24464 20085 24473
rect 20043 24424 20044 24464
rect 20084 24424 20085 24464
rect 20043 24415 20085 24424
rect 20044 24330 20084 24415
rect 18808 24212 19176 24221
rect 18848 24172 18890 24212
rect 18930 24172 18972 24212
rect 19012 24172 19054 24212
rect 19094 24172 19136 24212
rect 18808 24163 19176 24172
rect 20620 24044 20660 31051
rect 20811 27740 20853 27749
rect 20811 27700 20812 27740
rect 20852 27700 20853 27740
rect 20811 27691 20853 27700
rect 20715 27404 20757 27413
rect 20715 27364 20716 27404
rect 20756 27364 20757 27404
rect 20715 27355 20757 27364
rect 20236 24004 20660 24044
rect 18796 23960 18836 23969
rect 19467 23960 19509 23969
rect 18836 23920 19062 23960
rect 18796 23911 18836 23920
rect 19022 23807 19062 23920
rect 19467 23920 19468 23960
rect 19508 23920 19509 23960
rect 19467 23911 19509 23920
rect 20139 23960 20181 23969
rect 20139 23920 20140 23960
rect 20180 23920 20181 23960
rect 20139 23911 20181 23920
rect 20236 23960 20276 24004
rect 20236 23911 20276 23920
rect 19022 23758 19062 23767
rect 19180 23792 19220 23801
rect 19180 23129 19220 23752
rect 19275 23792 19317 23801
rect 19275 23752 19276 23792
rect 19316 23752 19317 23792
rect 19275 23743 19317 23752
rect 19468 23792 19508 23911
rect 19755 23876 19797 23885
rect 19755 23836 19756 23876
rect 19796 23836 19797 23876
rect 19755 23827 19797 23836
rect 19468 23743 19508 23752
rect 19564 23792 19604 23801
rect 19276 23658 19316 23743
rect 19372 23624 19412 23633
rect 19179 23120 19221 23129
rect 19179 23080 19180 23120
rect 19220 23080 19221 23120
rect 19179 23071 19221 23080
rect 19372 22952 19412 23584
rect 19276 22912 19412 22952
rect 18808 22700 19176 22709
rect 18848 22660 18890 22700
rect 18930 22660 18972 22700
rect 19012 22660 19054 22700
rect 19094 22660 19136 22700
rect 18808 22651 19176 22660
rect 19083 22532 19125 22541
rect 19083 22492 19084 22532
rect 19124 22492 19125 22532
rect 19083 22483 19125 22492
rect 18795 22448 18837 22457
rect 18795 22408 18796 22448
rect 18836 22408 18837 22448
rect 18795 22399 18837 22408
rect 18412 21474 18452 21559
rect 18027 21440 18069 21449
rect 18027 21400 18028 21440
rect 18068 21400 18069 21440
rect 18027 21391 18069 21400
rect 18219 21440 18261 21449
rect 18219 21400 18220 21440
rect 18260 21400 18261 21440
rect 18219 21391 18261 21400
rect 17835 21356 17877 21365
rect 17835 21316 17836 21356
rect 17876 21316 17877 21356
rect 17835 21307 17877 21316
rect 18028 21356 18068 21391
rect 17739 21188 17781 21197
rect 17739 21148 17740 21188
rect 17780 21148 17781 21188
rect 17739 21139 17781 21148
rect 17547 21020 17589 21029
rect 17547 20980 17548 21020
rect 17588 20980 17589 21020
rect 17547 20971 17589 20980
rect 17452 20719 17492 20728
rect 17548 20768 17588 20971
rect 17548 20719 17588 20728
rect 17643 20768 17685 20777
rect 17643 20728 17644 20768
rect 17684 20728 17685 20768
rect 17643 20719 17685 20728
rect 17740 20768 17780 20777
rect 17644 20634 17684 20719
rect 17740 20609 17780 20728
rect 17739 20600 17781 20609
rect 17739 20560 17740 20600
rect 17780 20560 17781 20600
rect 17739 20551 17781 20560
rect 17355 20348 17397 20357
rect 17355 20308 17356 20348
rect 17396 20308 17397 20348
rect 17355 20299 17397 20308
rect 17643 20348 17685 20357
rect 17643 20308 17644 20348
rect 17684 20308 17685 20348
rect 17643 20299 17685 20308
rect 16972 20224 17204 20264
rect 17164 20180 17204 20224
rect 16491 20140 16492 20180
rect 16532 20140 16628 20180
rect 16684 20140 16916 20180
rect 17164 20140 17396 20180
rect 16491 20131 16533 20140
rect 16491 20012 16533 20021
rect 16491 19972 16492 20012
rect 16532 19972 16533 20012
rect 16491 19963 16533 19972
rect 16492 19256 16532 19963
rect 16492 19207 16532 19216
rect 16491 17996 16533 18005
rect 16491 17956 16492 17996
rect 16532 17956 16533 17996
rect 16491 17947 16533 17956
rect 16203 17072 16245 17081
rect 16203 17032 16204 17072
rect 16244 17032 16245 17072
rect 16203 17023 16245 17032
rect 16395 17072 16437 17081
rect 16395 17032 16396 17072
rect 16436 17032 16437 17072
rect 16395 17023 16437 17032
rect 16204 16938 16244 17023
rect 16299 16820 16341 16829
rect 16396 16820 16436 16829
rect 16299 16780 16300 16820
rect 16340 16780 16396 16820
rect 16299 16771 16341 16780
rect 16396 16771 16436 16780
rect 16011 16400 16053 16409
rect 16011 16360 16012 16400
rect 16052 16360 16053 16400
rect 16011 16351 16053 16360
rect 16203 16232 16245 16241
rect 16203 16192 16204 16232
rect 16244 16192 16245 16232
rect 16203 16183 16245 16192
rect 16011 15728 16053 15737
rect 16011 15688 16012 15728
rect 16052 15688 16053 15728
rect 16011 15679 16053 15688
rect 16012 14552 16052 15679
rect 16204 14981 16244 16183
rect 16299 16064 16341 16073
rect 16299 16024 16300 16064
rect 16340 16024 16341 16064
rect 16299 16015 16341 16024
rect 16203 14972 16245 14981
rect 16203 14932 16204 14972
rect 16244 14932 16245 14972
rect 16203 14923 16245 14932
rect 16107 14804 16149 14813
rect 16107 14764 16108 14804
rect 16148 14764 16149 14804
rect 16107 14755 16149 14764
rect 16108 14720 16148 14755
rect 16108 14669 16148 14680
rect 16203 14552 16245 14561
rect 16012 14512 16148 14552
rect 16011 14132 16053 14141
rect 16011 14092 16012 14132
rect 16052 14092 16053 14132
rect 16011 14083 16053 14092
rect 16012 13998 16052 14083
rect 15916 13210 16052 13250
rect 15916 12536 15956 12545
rect 15916 12209 15956 12496
rect 15915 12200 15957 12209
rect 15915 12160 15916 12200
rect 15956 12160 15957 12200
rect 15915 12151 15957 12160
rect 16012 12032 16052 13210
rect 15916 11992 16052 12032
rect 15819 11192 15861 11201
rect 15819 11152 15820 11192
rect 15860 11152 15861 11192
rect 15819 11143 15861 11152
rect 15916 11033 15956 11992
rect 16108 11696 16148 14512
rect 16203 14512 16204 14552
rect 16244 14512 16245 14552
rect 16203 14503 16245 14512
rect 16204 14216 16244 14503
rect 16204 14167 16244 14176
rect 16203 13796 16245 13805
rect 16203 13756 16204 13796
rect 16244 13756 16245 13796
rect 16203 13747 16245 13756
rect 16108 11360 16148 11656
rect 16012 11320 16148 11360
rect 15915 11024 15957 11033
rect 15915 10984 15916 11024
rect 15956 10984 15957 11024
rect 15915 10975 15957 10984
rect 15723 10436 15765 10445
rect 15723 10396 15724 10436
rect 15764 10396 15765 10436
rect 15723 10387 15765 10396
rect 16012 10277 16052 11320
rect 16107 11108 16149 11117
rect 16107 11068 16108 11108
rect 16148 11068 16149 11108
rect 16107 11059 16149 11068
rect 16011 10268 16053 10277
rect 16011 10228 16012 10268
rect 16052 10228 16053 10268
rect 16011 10219 16053 10228
rect 15819 9848 15861 9857
rect 15819 9808 15820 9848
rect 15860 9808 15861 9848
rect 15819 9799 15861 9808
rect 15531 9260 15573 9269
rect 15531 9220 15532 9260
rect 15572 9220 15573 9260
rect 15531 9211 15573 9220
rect 15628 8849 15668 9388
rect 15723 9260 15765 9269
rect 15723 9220 15724 9260
rect 15764 9220 15765 9260
rect 15723 9211 15765 9220
rect 15627 8840 15669 8849
rect 15627 8800 15628 8840
rect 15668 8800 15669 8840
rect 15627 8791 15669 8800
rect 15435 8588 15477 8597
rect 15435 8548 15436 8588
rect 15476 8548 15477 8588
rect 15435 8539 15477 8548
rect 15627 8420 15669 8429
rect 15627 8380 15628 8420
rect 15668 8380 15669 8420
rect 15627 8371 15669 8380
rect 15628 8000 15668 8371
rect 15628 7951 15668 7960
rect 15339 7832 15381 7841
rect 15339 7792 15340 7832
rect 15380 7792 15381 7832
rect 15339 7783 15381 7792
rect 15147 7496 15189 7505
rect 15147 7456 15148 7496
rect 15188 7456 15189 7496
rect 15147 7447 15189 7456
rect 15340 6488 15380 6497
rect 15052 6364 15188 6404
rect 15051 6236 15093 6245
rect 15051 6196 15052 6236
rect 15092 6196 15093 6236
rect 15051 6187 15093 6196
rect 15052 5662 15092 6187
rect 15052 5069 15092 5622
rect 15051 5060 15093 5069
rect 15051 5020 15052 5060
rect 15092 5020 15093 5060
rect 15051 5011 15093 5020
rect 14956 4976 14996 4985
rect 15148 4962 15188 6364
rect 15243 5648 15285 5657
rect 15243 5608 15244 5648
rect 15284 5608 15285 5648
rect 15243 5599 15285 5608
rect 15244 5564 15284 5599
rect 15244 5513 15284 5524
rect 14956 4313 14996 4936
rect 15052 4922 15188 4962
rect 14955 4304 14997 4313
rect 14955 4264 14956 4304
rect 14996 4264 14997 4304
rect 14955 4255 14997 4264
rect 14955 3800 14997 3809
rect 14955 3760 14956 3800
rect 14996 3760 14997 3800
rect 14955 3751 14997 3760
rect 14956 3380 14996 3751
rect 14956 3331 14996 3340
rect 14860 3172 14996 3212
rect 14764 2969 14804 3172
rect 14859 3044 14901 3053
rect 14859 3004 14860 3044
rect 14900 3004 14901 3044
rect 14859 2995 14901 3004
rect 14763 2960 14805 2969
rect 14763 2920 14764 2960
rect 14804 2920 14805 2960
rect 14763 2911 14805 2920
rect 14860 2792 14900 2995
rect 14764 2752 14900 2792
rect 14764 1961 14804 2752
rect 14956 2708 14996 3172
rect 15052 3053 15092 4922
rect 15340 4136 15380 6448
rect 15724 6488 15764 9211
rect 15820 6656 15860 9799
rect 15915 9680 15957 9689
rect 15915 9640 15916 9680
rect 15956 9640 15957 9680
rect 15915 9631 15957 9640
rect 15916 8765 15956 9631
rect 15915 8756 15957 8765
rect 15915 8716 15916 8756
rect 15956 8716 15957 8756
rect 15915 8707 15957 8716
rect 15915 8504 15957 8513
rect 15915 8464 15916 8504
rect 15956 8464 15957 8504
rect 15915 8455 15957 8464
rect 15820 6607 15860 6616
rect 15724 6439 15764 6448
rect 15819 6488 15861 6497
rect 15819 6448 15820 6488
rect 15860 6448 15861 6488
rect 15819 6439 15861 6448
rect 15916 6488 15956 8455
rect 16012 8429 16052 10219
rect 16108 9773 16148 11059
rect 16107 9764 16149 9773
rect 16107 9724 16108 9764
rect 16148 9724 16149 9764
rect 16107 9715 16149 9724
rect 16108 9512 16148 9715
rect 16108 9463 16148 9472
rect 16107 8756 16149 8765
rect 16107 8716 16108 8756
rect 16148 8716 16149 8756
rect 16107 8707 16149 8716
rect 16011 8420 16053 8429
rect 16011 8380 16012 8420
rect 16052 8380 16053 8420
rect 16011 8371 16053 8380
rect 16011 8252 16053 8261
rect 16011 8212 16012 8252
rect 16052 8212 16053 8252
rect 16011 8203 16053 8212
rect 15916 6439 15956 6448
rect 15531 6236 15573 6245
rect 15531 6196 15532 6236
rect 15572 6196 15573 6236
rect 15531 6187 15573 6196
rect 15532 6102 15572 6187
rect 15820 6152 15860 6439
rect 15820 6112 15956 6152
rect 15436 5825 15476 5910
rect 15435 5816 15477 5825
rect 15435 5776 15436 5816
rect 15476 5776 15477 5816
rect 15435 5767 15477 5776
rect 15819 5648 15861 5657
rect 15819 5608 15820 5648
rect 15860 5608 15861 5648
rect 15819 5599 15861 5608
rect 15724 5564 15764 5573
rect 15531 5396 15573 5405
rect 15531 5356 15532 5396
rect 15572 5356 15573 5396
rect 15531 5347 15573 5356
rect 15435 5060 15477 5069
rect 15435 5020 15436 5060
rect 15476 5020 15477 5060
rect 15435 5011 15477 5020
rect 15436 4971 15476 5011
rect 15436 4922 15476 4931
rect 15532 4388 15572 5347
rect 15628 5144 15668 5153
rect 15724 5144 15764 5524
rect 15820 5514 15860 5599
rect 15668 5104 15764 5144
rect 15628 5095 15668 5104
rect 15820 4808 15860 4817
rect 15532 4339 15572 4348
rect 15628 4768 15820 4808
rect 15340 3893 15380 4096
rect 15339 3884 15381 3893
rect 15339 3844 15340 3884
rect 15380 3844 15381 3884
rect 15339 3835 15381 3844
rect 15339 3716 15381 3725
rect 15339 3676 15340 3716
rect 15380 3676 15381 3716
rect 15339 3667 15381 3676
rect 15244 3464 15284 3473
rect 15051 3044 15093 3053
rect 15051 3004 15052 3044
rect 15092 3004 15093 3044
rect 15051 2995 15093 3004
rect 15052 2717 15092 2738
rect 14860 2668 14996 2708
rect 15051 2708 15093 2717
rect 15051 2668 15052 2708
rect 15092 2668 15093 2708
rect 14763 1952 14805 1961
rect 14763 1912 14764 1952
rect 14804 1912 14805 1952
rect 14763 1903 14805 1912
rect 14860 1877 14900 2668
rect 15051 2659 15093 2668
rect 15052 2643 15092 2659
rect 14956 2604 14996 2613
rect 15052 2594 15092 2603
rect 14956 2540 14996 2564
rect 15244 2540 15284 3424
rect 15340 3464 15380 3667
rect 15340 3415 15380 3424
rect 15435 3212 15477 3221
rect 15435 3172 15436 3212
rect 15476 3172 15477 3212
rect 15435 3163 15477 3172
rect 15436 2708 15476 3163
rect 15531 2960 15573 2969
rect 15531 2920 15532 2960
rect 15572 2920 15573 2960
rect 15531 2911 15573 2920
rect 15436 2659 15476 2668
rect 15532 2708 15572 2911
rect 15532 2659 15572 2668
rect 14956 2500 15284 2540
rect 14955 2372 14997 2381
rect 14955 2332 14956 2372
rect 14996 2332 14997 2372
rect 14955 2323 14997 2332
rect 14859 1868 14901 1877
rect 14859 1828 14860 1868
rect 14900 1828 14901 1868
rect 14859 1819 14901 1828
rect 14668 1408 14900 1448
rect 14572 953 14612 1240
rect 14667 1280 14709 1289
rect 14667 1240 14668 1280
rect 14708 1240 14709 1280
rect 14667 1231 14709 1240
rect 14571 944 14613 953
rect 14571 904 14572 944
rect 14612 904 14613 944
rect 14571 895 14613 904
rect 14668 80 14708 1231
rect 14764 944 14804 953
rect 14764 533 14804 904
rect 14763 524 14805 533
rect 14763 484 14764 524
rect 14804 484 14805 524
rect 14763 475 14805 484
rect 14860 80 14900 1408
rect 14956 1364 14996 2323
rect 15244 2120 15284 2500
rect 15244 2071 15284 2080
rect 15435 2120 15477 2129
rect 15435 2080 15436 2120
rect 15476 2080 15477 2120
rect 15435 2071 15477 2080
rect 15436 1986 15476 2071
rect 15051 1952 15093 1961
rect 15051 1912 15052 1952
rect 15092 1912 15093 1952
rect 15051 1903 15093 1912
rect 15052 1818 15092 1903
rect 15628 1625 15668 4768
rect 15820 4759 15860 4768
rect 15819 4640 15861 4649
rect 15819 4600 15820 4640
rect 15860 4600 15861 4640
rect 15819 4591 15861 4600
rect 15820 3968 15860 4591
rect 15916 4136 15956 6112
rect 15916 4087 15956 4096
rect 16012 4136 16052 8203
rect 16108 8000 16148 8707
rect 16204 8168 16244 13747
rect 16300 8681 16340 16015
rect 16395 15224 16437 15233
rect 16395 15184 16396 15224
rect 16436 15184 16437 15224
rect 16395 15175 16437 15184
rect 16396 14645 16436 15175
rect 16492 14897 16532 17947
rect 16588 15233 16628 20140
rect 16779 19676 16821 19685
rect 16779 19636 16780 19676
rect 16820 19636 16821 19676
rect 16779 19627 16821 19636
rect 16683 19424 16725 19433
rect 16683 19384 16684 19424
rect 16724 19384 16725 19424
rect 16683 19375 16725 19384
rect 16684 19290 16724 19375
rect 16780 18677 16820 19627
rect 16779 18668 16821 18677
rect 16779 18628 16780 18668
rect 16820 18628 16821 18668
rect 16779 18619 16821 18628
rect 16684 18500 16724 18509
rect 16684 18005 16724 18460
rect 16780 18500 16820 18509
rect 16780 18089 16820 18460
rect 16779 18080 16821 18089
rect 16779 18040 16780 18080
rect 16820 18040 16821 18080
rect 16779 18031 16821 18040
rect 16683 17996 16725 18005
rect 16683 17956 16684 17996
rect 16724 17956 16725 17996
rect 16683 17947 16725 17956
rect 16780 17072 16820 17081
rect 16780 16661 16820 17032
rect 16779 16652 16821 16661
rect 16779 16612 16780 16652
rect 16820 16612 16821 16652
rect 16779 16603 16821 16612
rect 16876 16577 16916 20140
rect 16972 20076 17108 20116
rect 16972 20021 17012 20076
rect 17068 20075 17108 20076
rect 17068 20026 17108 20035
rect 16971 20012 17013 20021
rect 16971 19972 16972 20012
rect 17012 19972 17013 20012
rect 16971 19963 17013 19972
rect 17259 19844 17301 19853
rect 17259 19804 17260 19844
rect 17300 19804 17301 19844
rect 17259 19795 17301 19804
rect 17260 19710 17300 19795
rect 17356 19601 17396 20140
rect 17644 20096 17684 20299
rect 17836 20180 17876 21307
rect 17931 21104 17973 21113
rect 17931 21064 17932 21104
rect 17972 21064 17973 21104
rect 17931 21055 17973 21064
rect 17932 20768 17972 21055
rect 18028 20777 18068 21316
rect 18507 20852 18549 20861
rect 18507 20812 18508 20852
rect 18548 20812 18549 20852
rect 18507 20803 18549 20812
rect 17932 20719 17972 20728
rect 18027 20768 18069 20777
rect 18027 20728 18028 20768
rect 18068 20728 18069 20768
rect 18027 20719 18069 20728
rect 18124 20768 18164 20777
rect 18028 20600 18068 20609
rect 18028 20441 18068 20560
rect 18027 20432 18069 20441
rect 18027 20392 18028 20432
rect 18068 20392 18069 20432
rect 18027 20383 18069 20392
rect 18124 20189 18164 20728
rect 18315 20768 18357 20777
rect 18315 20728 18316 20768
rect 18356 20728 18357 20768
rect 18315 20719 18357 20728
rect 18316 20634 18356 20719
rect 18219 20516 18261 20525
rect 18219 20476 18220 20516
rect 18260 20476 18261 20516
rect 18219 20467 18261 20476
rect 18123 20180 18165 20189
rect 17836 20140 17972 20180
rect 17644 19685 17684 20056
rect 17643 19676 17685 19685
rect 17643 19636 17644 19676
rect 17684 19636 17685 19676
rect 17643 19627 17685 19636
rect 17355 19592 17397 19601
rect 17355 19552 17356 19592
rect 17396 19552 17397 19592
rect 17355 19543 17397 19552
rect 17739 19508 17781 19517
rect 17739 19468 17740 19508
rect 17780 19468 17781 19508
rect 17739 19459 17781 19468
rect 17452 19424 17492 19433
rect 17161 19384 17452 19424
rect 17161 19273 17201 19384
rect 17452 19375 17492 19384
rect 17643 19340 17685 19349
rect 17643 19300 17644 19340
rect 17684 19300 17685 19340
rect 17643 19291 17685 19300
rect 17068 19256 17108 19265
rect 17161 19264 17204 19273
rect 17161 19225 17164 19264
rect 16972 19088 17012 19097
rect 16972 17417 17012 19048
rect 17068 18929 17108 19216
rect 17164 19215 17204 19224
rect 17259 19256 17301 19265
rect 17452 19256 17492 19265
rect 17259 19216 17260 19256
rect 17300 19216 17301 19256
rect 17259 19207 17301 19216
rect 17356 19216 17452 19256
rect 17067 18920 17109 18929
rect 17067 18880 17068 18920
rect 17108 18880 17109 18920
rect 17067 18871 17109 18880
rect 17260 18761 17300 19207
rect 17259 18752 17301 18761
rect 17259 18712 17260 18752
rect 17300 18712 17301 18752
rect 17259 18703 17301 18712
rect 17067 18668 17109 18677
rect 17067 18628 17068 18668
rect 17108 18628 17109 18668
rect 17067 18619 17109 18628
rect 17068 17744 17108 18619
rect 17164 18584 17204 18593
rect 17164 18509 17204 18544
rect 17260 18584 17300 18595
rect 17260 18509 17300 18544
rect 17152 18500 17204 18509
rect 17152 18460 17153 18500
rect 17193 18460 17204 18500
rect 17259 18500 17301 18509
rect 17259 18460 17260 18500
rect 17300 18460 17301 18500
rect 17152 18451 17194 18460
rect 17259 18451 17301 18460
rect 17356 17996 17396 19216
rect 17452 19207 17492 19216
rect 17644 19256 17684 19291
rect 17644 18845 17684 19216
rect 17740 19256 17780 19459
rect 17740 19207 17780 19216
rect 17932 18929 17972 20140
rect 18123 20140 18124 20180
rect 18164 20140 18165 20180
rect 18123 20131 18165 20140
rect 18123 19256 18165 19265
rect 18123 19216 18124 19256
rect 18164 19216 18165 19256
rect 18123 19207 18165 19216
rect 18220 19256 18260 20467
rect 18411 20180 18453 20189
rect 18411 20140 18412 20180
rect 18452 20140 18453 20180
rect 18411 20131 18453 20140
rect 18315 19844 18357 19853
rect 18315 19804 18316 19844
rect 18356 19804 18357 19844
rect 18315 19795 18357 19804
rect 18220 19207 18260 19216
rect 17931 18920 17973 18929
rect 17931 18880 17932 18920
rect 17972 18880 17973 18920
rect 17931 18871 17973 18880
rect 17643 18836 17685 18845
rect 17643 18796 17644 18836
rect 17684 18796 17685 18836
rect 17643 18787 17685 18796
rect 17835 18836 17877 18845
rect 17835 18796 17836 18836
rect 17876 18796 17877 18836
rect 17835 18787 17877 18796
rect 17739 18752 17781 18761
rect 17739 18712 17740 18752
rect 17780 18712 17781 18752
rect 17739 18703 17781 18712
rect 17644 18593 17684 18678
rect 17548 18584 17588 18593
rect 17451 18500 17493 18509
rect 17451 18460 17452 18500
rect 17492 18460 17493 18500
rect 17451 18451 17493 18460
rect 17068 17695 17108 17704
rect 17164 17956 17396 17996
rect 16971 17408 17013 17417
rect 16971 17368 16972 17408
rect 17012 17368 17013 17408
rect 16971 17359 17013 17368
rect 17067 17156 17109 17165
rect 17067 17116 17068 17156
rect 17108 17116 17109 17156
rect 17067 17107 17109 17116
rect 16971 17072 17013 17081
rect 16971 17032 16972 17072
rect 17012 17032 17013 17072
rect 16971 17023 17013 17032
rect 17068 17072 17108 17107
rect 16875 16568 16917 16577
rect 16875 16528 16876 16568
rect 16916 16528 16917 16568
rect 16875 16519 16917 16528
rect 16683 16400 16725 16409
rect 16683 16360 16684 16400
rect 16724 16360 16725 16400
rect 16683 16351 16725 16360
rect 16684 16316 16724 16351
rect 16587 15224 16629 15233
rect 16587 15184 16588 15224
rect 16628 15184 16629 15224
rect 16587 15175 16629 15184
rect 16684 15065 16724 16276
rect 16780 16232 16820 16241
rect 16972 16232 17012 17023
rect 17068 17021 17108 17032
rect 17068 16904 17108 16913
rect 17164 16904 17204 17956
rect 17259 17828 17301 17837
rect 17259 17788 17260 17828
rect 17300 17788 17301 17828
rect 17259 17779 17301 17788
rect 17260 17744 17300 17779
rect 17260 17693 17300 17704
rect 17356 17744 17396 17753
rect 17452 17744 17492 18451
rect 17396 17704 17492 17744
rect 17548 17744 17588 18544
rect 17643 18584 17685 18593
rect 17643 18544 17644 18584
rect 17684 18544 17685 18584
rect 17643 18535 17685 18544
rect 17740 18584 17780 18703
rect 17740 18535 17780 18544
rect 17836 18584 17876 18787
rect 17836 18509 17876 18544
rect 17835 18500 17877 18509
rect 17835 18460 17836 18500
rect 17876 18460 17877 18500
rect 17835 18451 17877 18460
rect 18027 18500 18069 18509
rect 18027 18460 18028 18500
rect 18068 18460 18069 18500
rect 18027 18451 18069 18460
rect 17836 18420 17876 18451
rect 17643 18332 17685 18341
rect 17643 18292 17644 18332
rect 17684 18292 17685 18332
rect 17643 18283 17685 18292
rect 17259 17408 17301 17417
rect 17259 17368 17260 17408
rect 17300 17368 17301 17408
rect 17259 17359 17301 17368
rect 17260 17072 17300 17359
rect 17356 17333 17396 17704
rect 17548 17695 17588 17704
rect 17452 17576 17492 17585
rect 17355 17324 17397 17333
rect 17355 17284 17356 17324
rect 17396 17284 17397 17324
rect 17355 17275 17397 17284
rect 17355 17156 17397 17165
rect 17355 17116 17356 17156
rect 17396 17116 17397 17156
rect 17355 17107 17397 17116
rect 17260 17023 17300 17032
rect 17356 17022 17396 17107
rect 17452 17072 17492 17536
rect 17452 17023 17492 17032
rect 17644 17072 17684 18283
rect 18028 18089 18068 18451
rect 18027 18080 18069 18089
rect 18027 18040 18028 18080
rect 18068 18040 18069 18080
rect 18027 18031 18069 18040
rect 17739 17996 17781 18005
rect 17739 17956 17740 17996
rect 17780 17956 17781 17996
rect 17739 17947 17781 17956
rect 17740 17585 17780 17947
rect 17932 17744 17972 17753
rect 17739 17576 17781 17585
rect 17739 17536 17740 17576
rect 17780 17536 17781 17576
rect 17739 17527 17781 17536
rect 17644 17023 17684 17032
rect 17108 16864 17204 16904
rect 17068 16855 17108 16864
rect 17259 16820 17301 16829
rect 17259 16780 17260 16820
rect 17300 16780 17301 16820
rect 17259 16771 17301 16780
rect 17644 16820 17684 16829
rect 17163 16316 17205 16325
rect 17163 16276 17164 16316
rect 17204 16276 17205 16316
rect 17163 16267 17205 16276
rect 16820 16192 17012 16232
rect 17164 16232 17204 16267
rect 16780 15485 16820 16192
rect 17068 15560 17108 15569
rect 16972 15520 17068 15560
rect 16779 15476 16821 15485
rect 16779 15436 16780 15476
rect 16820 15436 16821 15476
rect 16779 15427 16821 15436
rect 16683 15056 16725 15065
rect 16683 15016 16684 15056
rect 16724 15016 16725 15056
rect 16683 15007 16725 15016
rect 16491 14888 16533 14897
rect 16491 14848 16492 14888
rect 16532 14848 16533 14888
rect 16491 14839 16533 14848
rect 16779 14888 16821 14897
rect 16779 14848 16780 14888
rect 16820 14848 16821 14888
rect 16779 14839 16821 14848
rect 16588 14720 16628 14729
rect 16395 14636 16437 14645
rect 16395 14596 16396 14636
rect 16436 14596 16437 14636
rect 16395 14587 16437 14596
rect 16588 14561 16628 14680
rect 16684 14720 16724 14729
rect 16684 14645 16724 14680
rect 16683 14636 16725 14645
rect 16683 14596 16684 14636
rect 16724 14596 16725 14636
rect 16683 14587 16725 14596
rect 16684 14585 16724 14587
rect 16587 14552 16629 14561
rect 16587 14512 16588 14552
rect 16628 14512 16629 14552
rect 16587 14503 16629 14512
rect 16395 14300 16437 14309
rect 16395 14260 16396 14300
rect 16436 14260 16437 14300
rect 16395 14251 16437 14260
rect 16396 14048 16436 14251
rect 16396 13999 16436 14008
rect 16395 13796 16437 13805
rect 16395 13756 16396 13796
rect 16436 13756 16437 13796
rect 16395 13747 16437 13756
rect 16396 12452 16436 13747
rect 16588 13721 16628 14503
rect 16587 13712 16629 13721
rect 16587 13672 16588 13712
rect 16628 13672 16629 13712
rect 16587 13663 16629 13672
rect 16780 13301 16820 14839
rect 16972 14057 17012 15520
rect 17068 15511 17108 15520
rect 17164 15317 17204 16192
rect 17260 16232 17300 16771
rect 17355 16652 17397 16661
rect 17355 16612 17356 16652
rect 17396 16612 17397 16652
rect 17355 16603 17397 16612
rect 17260 16183 17300 16192
rect 17356 16064 17396 16603
rect 17644 16493 17684 16780
rect 17643 16484 17685 16493
rect 17643 16444 17644 16484
rect 17684 16444 17685 16484
rect 17643 16435 17685 16444
rect 17260 16024 17396 16064
rect 17548 16232 17588 16241
rect 17163 15308 17205 15317
rect 17163 15268 17164 15308
rect 17204 15268 17205 15308
rect 17163 15259 17205 15268
rect 17067 15224 17109 15233
rect 17067 15184 17068 15224
rect 17108 15184 17109 15224
rect 17067 15175 17109 15184
rect 17068 14720 17108 15175
rect 16971 14048 17013 14057
rect 16971 14008 16972 14048
rect 17012 14008 17013 14048
rect 16971 13999 17013 14008
rect 17068 13805 17108 14680
rect 17164 14720 17204 14729
rect 17164 14141 17204 14680
rect 17163 14132 17205 14141
rect 17163 14092 17164 14132
rect 17204 14092 17205 14132
rect 17163 14083 17205 14092
rect 17260 13889 17300 16024
rect 17548 15989 17588 16192
rect 17547 15980 17589 15989
rect 17547 15940 17548 15980
rect 17588 15940 17589 15980
rect 17547 15931 17589 15940
rect 17355 15560 17397 15569
rect 17355 15520 17356 15560
rect 17396 15520 17397 15560
rect 17355 15511 17397 15520
rect 17452 15560 17492 15569
rect 17356 15426 17396 15511
rect 17452 15149 17492 15520
rect 17548 15560 17588 15569
rect 17451 15140 17493 15149
rect 17451 15100 17452 15140
rect 17492 15100 17493 15140
rect 17451 15091 17493 15100
rect 17355 15056 17397 15065
rect 17355 15016 17356 15056
rect 17396 15016 17397 15056
rect 17355 15007 17397 15016
rect 17259 13880 17301 13889
rect 17259 13840 17260 13880
rect 17300 13840 17301 13880
rect 17259 13831 17301 13840
rect 17067 13796 17109 13805
rect 17067 13756 17068 13796
rect 17108 13756 17109 13796
rect 17067 13747 17109 13756
rect 16779 13292 16821 13301
rect 16779 13252 16780 13292
rect 16820 13252 16821 13292
rect 16779 13243 16821 13252
rect 16491 13208 16533 13217
rect 16491 13168 16492 13208
rect 16532 13168 16533 13208
rect 16491 13159 16533 13168
rect 17164 13208 17204 13217
rect 16492 13074 16532 13159
rect 16684 13040 16724 13049
rect 16587 12536 16629 12545
rect 16396 12284 16436 12412
rect 16492 12496 16588 12536
rect 16628 12496 16629 12536
rect 16492 12452 16532 12496
rect 16587 12487 16629 12496
rect 16492 12403 16532 12412
rect 16396 12244 16532 12284
rect 16395 11192 16437 11201
rect 16395 11152 16396 11192
rect 16436 11152 16437 11192
rect 16395 11143 16437 11152
rect 16299 8672 16341 8681
rect 16299 8632 16300 8672
rect 16340 8632 16341 8672
rect 16299 8623 16341 8632
rect 16204 8128 16340 8168
rect 16108 7421 16148 7960
rect 16203 8000 16245 8009
rect 16203 7960 16204 8000
rect 16244 7960 16245 8000
rect 16203 7951 16245 7960
rect 16204 7866 16244 7951
rect 16107 7412 16149 7421
rect 16107 7372 16108 7412
rect 16148 7372 16149 7412
rect 16107 7363 16149 7372
rect 16107 7244 16149 7253
rect 16107 7204 16108 7244
rect 16148 7204 16149 7244
rect 16107 7195 16149 7204
rect 16108 6833 16148 7195
rect 16204 7160 16244 7169
rect 16300 7160 16340 8128
rect 16244 7120 16340 7160
rect 16107 6824 16149 6833
rect 16107 6784 16108 6824
rect 16148 6784 16149 6824
rect 16107 6775 16149 6784
rect 16108 6497 16148 6775
rect 16204 6665 16244 7120
rect 16299 6992 16341 7001
rect 16299 6952 16300 6992
rect 16340 6952 16341 6992
rect 16299 6943 16341 6952
rect 16203 6656 16245 6665
rect 16203 6616 16204 6656
rect 16244 6616 16245 6656
rect 16203 6607 16245 6616
rect 16107 6488 16149 6497
rect 16107 6448 16108 6488
rect 16148 6448 16149 6488
rect 16107 6439 16149 6448
rect 16300 6488 16340 6943
rect 16396 6656 16436 11143
rect 16492 11117 16532 12244
rect 16684 11780 16724 13000
rect 17164 12713 17204 13168
rect 17163 12704 17205 12713
rect 17163 12664 17164 12704
rect 17204 12664 17205 12704
rect 17163 12655 17205 12664
rect 17259 12620 17301 12629
rect 17259 12580 17260 12620
rect 17300 12580 17301 12620
rect 17259 12571 17301 12580
rect 16876 12536 16916 12545
rect 16636 11740 16724 11780
rect 16780 12496 16876 12536
rect 16636 11738 16676 11740
rect 16780 11705 16820 12496
rect 16876 12487 16916 12496
rect 16972 12536 17012 12545
rect 16972 11948 17012 12496
rect 17260 12486 17300 12571
rect 17356 12461 17396 15007
rect 17451 13964 17493 13973
rect 17451 13924 17452 13964
rect 17492 13924 17493 13964
rect 17451 13915 17493 13924
rect 17452 12713 17492 13915
rect 17451 12704 17493 12713
rect 17451 12664 17452 12704
rect 17492 12664 17493 12704
rect 17451 12655 17493 12664
rect 17452 12536 17492 12545
rect 17163 12452 17205 12461
rect 17163 12412 17164 12452
rect 17204 12412 17205 12452
rect 17163 12403 17205 12412
rect 17355 12452 17397 12461
rect 17355 12412 17356 12452
rect 17396 12412 17397 12452
rect 17355 12403 17397 12412
rect 17164 12284 17204 12403
rect 17164 12244 17396 12284
rect 16876 11908 17012 11948
rect 16636 11689 16676 11698
rect 16779 11696 16821 11705
rect 16779 11656 16780 11696
rect 16820 11656 16821 11696
rect 16779 11647 16821 11656
rect 16779 11528 16821 11537
rect 16779 11488 16780 11528
rect 16820 11488 16821 11528
rect 16779 11479 16821 11488
rect 16780 11394 16820 11479
rect 16780 11192 16820 11201
rect 16876 11192 16916 11908
rect 17164 11780 17204 11789
rect 16972 11537 17012 11622
rect 16971 11528 17013 11537
rect 16971 11488 16972 11528
rect 17012 11488 17013 11528
rect 16971 11479 17013 11488
rect 16971 11360 17013 11369
rect 16971 11320 16972 11360
rect 17012 11320 17013 11360
rect 16971 11311 17013 11320
rect 16820 11152 16916 11192
rect 16780 11143 16820 11152
rect 16491 11108 16533 11117
rect 16972 11108 17012 11311
rect 17067 11192 17109 11201
rect 17067 11152 17068 11192
rect 17108 11152 17109 11192
rect 17067 11143 17109 11152
rect 16491 11068 16492 11108
rect 16532 11068 16533 11108
rect 16491 11059 16533 11068
rect 16876 11068 17012 11108
rect 16588 11024 16628 11033
rect 16588 10781 16628 10984
rect 16876 10949 16916 11068
rect 16972 10982 17012 10991
rect 16875 10940 16917 10949
rect 16875 10900 16876 10940
rect 16916 10900 16917 10940
rect 16875 10891 16917 10900
rect 16587 10772 16629 10781
rect 16587 10732 16588 10772
rect 16628 10732 16629 10772
rect 16587 10723 16629 10732
rect 16972 10529 17012 10942
rect 16971 10520 17013 10529
rect 16971 10480 16972 10520
rect 17012 10480 17013 10520
rect 16971 10471 17013 10480
rect 16587 10436 16629 10445
rect 16587 10396 16588 10436
rect 16628 10396 16629 10436
rect 16587 10387 16629 10396
rect 16588 10184 16628 10387
rect 17068 10352 17108 11143
rect 17164 10613 17204 11740
rect 17356 11696 17396 12244
rect 17356 11647 17396 11656
rect 17452 10781 17492 12496
rect 17451 10772 17493 10781
rect 17451 10732 17452 10772
rect 17492 10732 17493 10772
rect 17451 10723 17493 10732
rect 17163 10604 17205 10613
rect 17163 10564 17164 10604
rect 17204 10564 17205 10604
rect 17163 10555 17205 10564
rect 17259 10436 17301 10445
rect 17259 10396 17260 10436
rect 17300 10396 17301 10436
rect 17259 10387 17301 10396
rect 16491 10100 16533 10109
rect 16491 10060 16492 10100
rect 16532 10060 16533 10100
rect 16491 10051 16533 10060
rect 16492 8840 16532 10051
rect 16588 9689 16628 10144
rect 16972 10312 17108 10352
rect 16972 10184 17012 10312
rect 16972 10135 17012 10144
rect 17067 10184 17109 10193
rect 17067 10144 17068 10184
rect 17108 10144 17109 10184
rect 17067 10135 17109 10144
rect 17260 10184 17300 10387
rect 17260 10135 17300 10144
rect 17452 10184 17492 10193
rect 17068 10050 17108 10135
rect 17452 10025 17492 10144
rect 16780 10016 16820 10025
rect 16684 9976 16780 10016
rect 16587 9680 16629 9689
rect 16587 9640 16588 9680
rect 16628 9640 16629 9680
rect 16587 9631 16629 9640
rect 16684 9521 16724 9976
rect 16780 9967 16820 9976
rect 17164 10016 17204 10025
rect 17164 9764 17204 9976
rect 17451 10016 17493 10025
rect 17451 9976 17452 10016
rect 17492 9976 17493 10016
rect 17451 9967 17493 9976
rect 17164 9724 17396 9764
rect 16779 9680 16821 9689
rect 16779 9640 16780 9680
rect 16820 9640 16821 9680
rect 16779 9631 16821 9640
rect 16780 9546 16820 9631
rect 16683 9512 16725 9521
rect 16588 9498 16628 9507
rect 16683 9472 16684 9512
rect 16724 9472 16725 9512
rect 16683 9463 16725 9472
rect 16972 9512 17012 9523
rect 16588 8924 16628 9458
rect 16972 9437 17012 9472
rect 17068 9512 17108 9521
rect 16971 9428 17013 9437
rect 16971 9388 16972 9428
rect 17012 9388 17013 9428
rect 16971 9379 17013 9388
rect 16684 8924 16724 8933
rect 16588 8884 16684 8924
rect 16724 8884 16916 8924
rect 16684 8875 16724 8884
rect 16492 8800 16628 8840
rect 16492 8672 16532 8683
rect 16492 8597 16532 8632
rect 16491 8588 16533 8597
rect 16491 8548 16492 8588
rect 16532 8548 16533 8588
rect 16491 8539 16533 8548
rect 16491 8336 16533 8345
rect 16491 8296 16492 8336
rect 16532 8296 16533 8336
rect 16491 8287 16533 8296
rect 16492 7589 16532 8287
rect 16588 8252 16628 8800
rect 16876 8681 16916 8884
rect 16972 8743 17012 9379
rect 17068 8849 17108 9472
rect 17163 9512 17205 9521
rect 17163 9472 17164 9512
rect 17204 9472 17205 9512
rect 17163 9463 17205 9472
rect 17260 9512 17300 9521
rect 17164 9378 17204 9463
rect 17260 8849 17300 9472
rect 17356 8924 17396 9724
rect 17548 9689 17588 15520
rect 17644 15560 17684 15569
rect 17644 14561 17684 15520
rect 17740 15317 17780 17527
rect 17835 17156 17877 17165
rect 17835 17116 17836 17156
rect 17876 17116 17877 17156
rect 17835 17107 17877 17116
rect 17836 17072 17876 17107
rect 17836 17021 17876 17032
rect 17932 15653 17972 17704
rect 17931 15644 17973 15653
rect 17931 15604 17932 15644
rect 17972 15604 17973 15644
rect 17931 15595 17973 15604
rect 17835 15560 17877 15569
rect 17835 15520 17836 15560
rect 17876 15520 17877 15560
rect 17835 15511 17877 15520
rect 17836 15426 17876 15511
rect 17739 15308 17781 15317
rect 17739 15268 17740 15308
rect 17780 15268 17781 15308
rect 17739 15259 17781 15268
rect 17739 15140 17781 15149
rect 17739 15100 17740 15140
rect 17780 15100 17781 15140
rect 17739 15091 17781 15100
rect 17740 14720 17780 15091
rect 17835 14972 17877 14981
rect 17835 14932 17836 14972
rect 17876 14932 17877 14972
rect 17835 14923 17877 14932
rect 17643 14552 17685 14561
rect 17643 14512 17644 14552
rect 17684 14512 17685 14552
rect 17643 14503 17685 14512
rect 17643 14384 17685 14393
rect 17643 14344 17644 14384
rect 17684 14344 17685 14384
rect 17643 14335 17685 14344
rect 17644 14048 17684 14335
rect 17644 10697 17684 14008
rect 17740 13469 17780 14680
rect 17836 14720 17876 14923
rect 18028 14888 18068 18031
rect 18124 17828 18164 19207
rect 18124 17779 18164 17788
rect 18316 18584 18356 19795
rect 18412 18929 18452 20131
rect 18411 18920 18453 18929
rect 18411 18880 18412 18920
rect 18452 18880 18453 18920
rect 18411 18871 18453 18880
rect 18220 17744 18260 17753
rect 18316 17744 18356 18544
rect 18412 18584 18452 18593
rect 18508 18584 18548 20803
rect 18452 18544 18548 18584
rect 18412 18535 18452 18544
rect 18260 17704 18356 17744
rect 18411 17744 18453 17753
rect 18411 17704 18412 17744
rect 18452 17704 18453 17744
rect 18220 17695 18260 17704
rect 18411 17695 18453 17704
rect 18412 17610 18452 17695
rect 18700 17669 18740 21568
rect 18796 21524 18836 22399
rect 18987 22112 19029 22121
rect 18987 22072 18988 22112
rect 19028 22072 19029 22112
rect 18987 22063 19029 22072
rect 18891 21608 18933 21617
rect 18891 21568 18892 21608
rect 18932 21568 18933 21608
rect 18891 21559 18933 21568
rect 18796 21475 18836 21484
rect 18892 21440 18932 21559
rect 18988 21524 19028 22063
rect 19084 21608 19124 22483
rect 19084 21559 19124 21568
rect 19276 21608 19316 22912
rect 19564 22868 19604 23752
rect 19756 23742 19796 23827
rect 20140 23805 20180 23911
rect 20140 23756 20180 23765
rect 19947 23624 19989 23633
rect 19947 23584 19948 23624
rect 19988 23584 19989 23624
rect 19947 23575 19989 23584
rect 19948 23490 19988 23575
rect 20048 23456 20416 23465
rect 20088 23416 20130 23456
rect 20170 23416 20212 23456
rect 20252 23416 20294 23456
rect 20334 23416 20376 23456
rect 20048 23407 20416 23416
rect 19659 23204 19701 23213
rect 19659 23164 19660 23204
rect 19700 23164 19701 23204
rect 19659 23155 19701 23164
rect 19468 22828 19604 22868
rect 19660 23120 19700 23155
rect 20236 23129 20276 23214
rect 19371 22784 19413 22793
rect 19468 22784 19508 22828
rect 19371 22744 19372 22784
rect 19412 22744 19508 22784
rect 19371 22735 19413 22744
rect 19276 21559 19316 21568
rect 18988 21475 19028 21484
rect 19372 21524 19412 22735
rect 19563 22700 19605 22709
rect 19563 22660 19564 22700
rect 19604 22660 19605 22700
rect 19563 22651 19605 22660
rect 19564 22373 19604 22651
rect 19563 22364 19605 22373
rect 19563 22324 19564 22364
rect 19604 22324 19605 22364
rect 19563 22315 19605 22324
rect 19564 21776 19604 22315
rect 19660 22280 19700 23080
rect 19947 23120 19989 23129
rect 19947 23080 19948 23120
rect 19988 23080 19989 23120
rect 19947 23071 19989 23080
rect 20044 23120 20084 23129
rect 19852 22952 19892 22961
rect 19756 22912 19852 22952
rect 19756 22793 19796 22912
rect 19852 22903 19892 22912
rect 19755 22784 19797 22793
rect 19755 22744 19756 22784
rect 19796 22744 19797 22784
rect 19755 22735 19797 22744
rect 19851 22700 19893 22709
rect 19851 22660 19852 22700
rect 19892 22660 19893 22700
rect 19851 22651 19893 22660
rect 19756 22280 19796 22289
rect 19660 22240 19756 22280
rect 19756 22231 19796 22240
rect 19852 21785 19892 22651
rect 19948 22532 19988 23071
rect 20044 22709 20084 23080
rect 20235 23120 20277 23129
rect 20235 23080 20236 23120
rect 20276 23080 20277 23120
rect 20235 23071 20277 23080
rect 20139 23036 20181 23045
rect 20139 22996 20140 23036
rect 20180 22996 20181 23036
rect 20139 22987 20181 22996
rect 20140 22902 20180 22987
rect 20043 22700 20085 22709
rect 20043 22660 20044 22700
rect 20084 22660 20085 22700
rect 20043 22651 20085 22660
rect 20236 22532 20276 22541
rect 19948 22492 20236 22532
rect 20236 22483 20276 22492
rect 20127 22269 20167 22278
rect 19948 22196 19988 22205
rect 20127 22196 20167 22229
rect 19988 22156 20167 22196
rect 19851 21776 19893 21785
rect 19564 21736 19796 21776
rect 19563 21608 19605 21617
rect 19563 21568 19564 21608
rect 19604 21568 19605 21608
rect 19563 21559 19605 21568
rect 19660 21608 19700 21617
rect 19756 21608 19796 21736
rect 19851 21736 19852 21776
rect 19892 21736 19893 21776
rect 19851 21727 19893 21736
rect 19852 21608 19892 21617
rect 19756 21568 19852 21608
rect 19372 21475 19412 21484
rect 19564 21524 19604 21559
rect 19564 21473 19604 21484
rect 18892 21391 18932 21400
rect 19275 21440 19317 21449
rect 19275 21400 19276 21440
rect 19316 21400 19317 21440
rect 19275 21391 19317 21400
rect 19467 21440 19509 21449
rect 19467 21400 19468 21440
rect 19508 21400 19509 21440
rect 19660 21440 19700 21568
rect 19852 21559 19892 21568
rect 19948 21608 19988 22156
rect 20236 22121 20276 22206
rect 20235 22112 20277 22121
rect 20235 22072 20236 22112
rect 20276 22072 20277 22112
rect 20235 22063 20277 22072
rect 20048 21944 20416 21953
rect 20088 21904 20130 21944
rect 20170 21904 20212 21944
rect 20252 21904 20294 21944
rect 20334 21904 20376 21944
rect 20048 21895 20416 21904
rect 20139 21776 20181 21785
rect 20139 21736 20140 21776
rect 20180 21736 20181 21776
rect 20139 21727 20181 21736
rect 20043 21692 20085 21701
rect 20043 21652 20044 21692
rect 20084 21652 20085 21692
rect 20043 21643 20085 21652
rect 19948 21559 19988 21568
rect 19948 21440 19988 21449
rect 19660 21400 19948 21440
rect 19467 21391 19509 21400
rect 19948 21391 19988 21400
rect 18808 21188 19176 21197
rect 18848 21148 18890 21188
rect 18930 21148 18972 21188
rect 19012 21148 19054 21188
rect 19094 21148 19136 21188
rect 18808 21139 19176 21148
rect 19276 21020 19316 21391
rect 19468 21306 19508 21391
rect 20044 21104 20084 21643
rect 20140 21622 20180 21727
rect 20140 21573 20180 21582
rect 20044 21064 20180 21104
rect 19180 20980 19316 21020
rect 18891 20768 18933 20777
rect 18891 20728 18892 20768
rect 18932 20728 18933 20768
rect 18891 20719 18933 20728
rect 18892 20096 18932 20719
rect 18987 20600 19029 20609
rect 18987 20560 18988 20600
rect 19028 20560 19029 20600
rect 18987 20551 19029 20560
rect 18892 20021 18932 20056
rect 18891 20012 18933 20021
rect 18891 19972 18892 20012
rect 18932 19972 18933 20012
rect 18891 19963 18933 19972
rect 18988 19937 19028 20551
rect 19083 20096 19125 20105
rect 19083 20056 19084 20096
rect 19124 20056 19125 20096
rect 19083 20047 19125 20056
rect 18987 19928 19029 19937
rect 18987 19888 18988 19928
rect 19028 19888 19029 19928
rect 18987 19879 19029 19888
rect 19084 19853 19124 20047
rect 19083 19844 19125 19853
rect 19083 19804 19084 19844
rect 19124 19804 19125 19844
rect 19180 19844 19220 20980
rect 20140 20810 20180 21064
rect 19563 20768 19605 20777
rect 19563 20728 19564 20768
rect 19604 20728 19605 20768
rect 19563 20719 19605 20728
rect 19948 20768 19988 20777
rect 19564 20634 19604 20719
rect 19756 20684 19796 20693
rect 19948 20684 19988 20728
rect 19660 20644 19756 20684
rect 19796 20644 19988 20684
rect 20044 20768 20084 20777
rect 19660 20264 19700 20644
rect 19756 20635 19796 20644
rect 20044 20600 20084 20728
rect 20140 20609 20180 20770
rect 19948 20560 20084 20600
rect 20139 20600 20181 20609
rect 20139 20560 20140 20600
rect 20180 20560 20181 20600
rect 19468 20224 19700 20264
rect 19275 20096 19317 20105
rect 19275 20056 19276 20096
rect 19316 20056 19317 20096
rect 19275 20047 19317 20056
rect 19372 20096 19412 20105
rect 19276 19962 19316 20047
rect 19180 19804 19316 19844
rect 19083 19795 19125 19804
rect 18808 19676 19176 19685
rect 18848 19636 18890 19676
rect 18930 19636 18972 19676
rect 19012 19636 19054 19676
rect 19094 19636 19136 19676
rect 18808 19627 19176 19636
rect 19276 18761 19316 19804
rect 19372 19088 19412 20056
rect 19468 20096 19508 20224
rect 19468 20047 19508 20056
rect 19564 20096 19604 20105
rect 19467 19676 19509 19685
rect 19467 19636 19468 19676
rect 19508 19636 19509 19676
rect 19467 19627 19509 19636
rect 19468 19256 19508 19627
rect 19564 19349 19604 20056
rect 19660 19844 19700 20224
rect 19755 20264 19797 20273
rect 19755 20224 19756 20264
rect 19796 20224 19797 20264
rect 19755 20215 19797 20224
rect 19948 20264 19988 20560
rect 20139 20551 20181 20560
rect 20236 20600 20276 20609
rect 20276 20560 20564 20600
rect 20236 20551 20276 20560
rect 20048 20432 20416 20441
rect 20088 20392 20130 20432
rect 20170 20392 20212 20432
rect 20252 20392 20294 20432
rect 20334 20392 20376 20432
rect 20048 20383 20416 20392
rect 19948 20215 19988 20224
rect 19756 20111 19796 20215
rect 19756 20045 19796 20071
rect 19852 20096 19892 20105
rect 19852 19853 19892 20056
rect 20044 20096 20084 20105
rect 19851 19844 19893 19853
rect 19660 19804 19768 19844
rect 19728 19760 19768 19804
rect 19851 19804 19852 19844
rect 19892 19804 19988 19844
rect 19851 19795 19893 19804
rect 19728 19720 19796 19760
rect 19659 19676 19701 19685
rect 19659 19636 19660 19676
rect 19700 19636 19701 19676
rect 19659 19627 19701 19636
rect 19660 19508 19700 19627
rect 19660 19459 19700 19468
rect 19563 19340 19605 19349
rect 19563 19300 19564 19340
rect 19604 19300 19605 19340
rect 19563 19291 19605 19300
rect 19468 19207 19508 19216
rect 19756 19088 19796 19720
rect 19851 19424 19893 19433
rect 19851 19384 19852 19424
rect 19892 19384 19893 19424
rect 19851 19375 19893 19384
rect 19852 19256 19892 19375
rect 19852 19207 19892 19216
rect 19948 19256 19988 19804
rect 20044 19265 20084 20056
rect 20139 19424 20181 19433
rect 20139 19384 20140 19424
rect 20180 19384 20181 19424
rect 20139 19375 20181 19384
rect 20140 19267 20180 19375
rect 19948 19207 19988 19216
rect 20043 19256 20085 19265
rect 20043 19216 20044 19256
rect 20084 19216 20085 19256
rect 20140 19218 20180 19227
rect 20043 19207 20085 19216
rect 20044 19088 20084 19097
rect 19372 19048 19508 19088
rect 19756 19048 19892 19088
rect 19468 18845 19508 19048
rect 19467 18836 19509 18845
rect 19467 18796 19468 18836
rect 19508 18796 19509 18836
rect 19467 18787 19509 18796
rect 19275 18752 19317 18761
rect 19275 18712 19276 18752
rect 19316 18712 19317 18752
rect 19275 18703 19317 18712
rect 19372 18584 19412 18593
rect 19276 18544 19372 18584
rect 18795 18500 18837 18509
rect 18795 18460 18796 18500
rect 18836 18460 18837 18500
rect 18795 18451 18837 18460
rect 18892 18500 18932 18509
rect 18796 18366 18836 18451
rect 18892 18341 18932 18460
rect 18891 18332 18933 18341
rect 18891 18292 18892 18332
rect 18932 18292 18933 18332
rect 18891 18283 18933 18292
rect 19276 18257 19316 18544
rect 19372 18535 19412 18544
rect 19371 18332 19413 18341
rect 19371 18292 19372 18332
rect 19412 18292 19413 18332
rect 19371 18283 19413 18292
rect 19275 18248 19317 18257
rect 19275 18208 19276 18248
rect 19316 18208 19317 18248
rect 19275 18199 19317 18208
rect 18808 18164 19176 18173
rect 18848 18124 18890 18164
rect 18930 18124 18972 18164
rect 19012 18124 19054 18164
rect 19094 18124 19136 18164
rect 18808 18115 19176 18124
rect 19179 17996 19221 18005
rect 19179 17956 19180 17996
rect 19220 17956 19221 17996
rect 19179 17947 19221 17956
rect 18699 17660 18741 17669
rect 18699 17620 18700 17660
rect 18740 17620 18741 17660
rect 18699 17611 18741 17620
rect 18124 17072 18164 17083
rect 19180 17081 19220 17947
rect 18124 16997 18164 17032
rect 18699 17072 18741 17081
rect 18699 17032 18700 17072
rect 18740 17032 18741 17072
rect 18699 17023 18741 17032
rect 19179 17072 19221 17081
rect 19179 17032 19180 17072
rect 19220 17032 19221 17072
rect 19179 17023 19221 17032
rect 18123 16988 18165 16997
rect 18123 16948 18124 16988
rect 18164 16948 18165 16988
rect 18123 16939 18165 16948
rect 18700 16232 18740 17023
rect 18808 16652 19176 16661
rect 18848 16612 18890 16652
rect 18930 16612 18972 16652
rect 19012 16612 19054 16652
rect 19094 16612 19136 16652
rect 18808 16603 19176 16612
rect 19083 16484 19125 16493
rect 19083 16444 19084 16484
rect 19124 16444 19125 16484
rect 19276 16484 19316 18199
rect 19372 17240 19412 18283
rect 19468 18005 19508 18787
rect 19852 18579 19892 19048
rect 19852 18530 19892 18539
rect 19948 19048 20044 19088
rect 19659 18080 19701 18089
rect 19659 18040 19660 18080
rect 19700 18040 19701 18080
rect 19659 18031 19701 18040
rect 19467 17996 19509 18005
rect 19467 17956 19468 17996
rect 19508 17956 19509 17996
rect 19467 17947 19509 17956
rect 19660 17744 19700 18031
rect 19948 17744 19988 19048
rect 20044 19039 20084 19048
rect 20048 18920 20416 18929
rect 20088 18880 20130 18920
rect 20170 18880 20212 18920
rect 20252 18880 20294 18920
rect 20334 18880 20376 18920
rect 20048 18871 20416 18880
rect 20043 18752 20085 18761
rect 20043 18712 20044 18752
rect 20084 18712 20085 18752
rect 20043 18703 20085 18712
rect 20235 18752 20277 18761
rect 20235 18712 20236 18752
rect 20276 18712 20277 18752
rect 20235 18703 20277 18712
rect 20044 18618 20084 18703
rect 20236 17996 20276 18703
rect 20236 17947 20276 17956
rect 20044 17744 20084 17753
rect 19948 17704 20044 17744
rect 19660 17695 19700 17704
rect 20044 17695 20084 17704
rect 20236 17744 20276 17753
rect 20524 17744 20564 20560
rect 20716 20180 20756 27355
rect 20812 21953 20852 27691
rect 21004 23969 21044 32227
rect 21291 28916 21333 28925
rect 21291 28876 21292 28916
rect 21332 28876 21333 28916
rect 21291 28867 21333 28876
rect 21099 25724 21141 25733
rect 21099 25684 21100 25724
rect 21140 25684 21141 25724
rect 21099 25675 21141 25684
rect 21003 23960 21045 23969
rect 21003 23920 21004 23960
rect 21044 23920 21045 23960
rect 21003 23911 21045 23920
rect 20811 21944 20853 21953
rect 20811 21904 20812 21944
rect 20852 21904 20853 21944
rect 20811 21895 20853 21904
rect 20276 17704 20564 17744
rect 20620 20140 20756 20180
rect 20236 17695 20276 17704
rect 19852 17576 19892 17585
rect 19892 17536 19988 17576
rect 19852 17527 19892 17536
rect 19372 17200 19508 17240
rect 19371 17072 19413 17081
rect 19371 17032 19372 17072
rect 19412 17032 19413 17072
rect 19371 17023 19413 17032
rect 19372 16938 19412 17023
rect 19276 16444 19412 16484
rect 19083 16435 19125 16444
rect 18796 16232 18836 16241
rect 18700 16192 18796 16232
rect 18700 15905 18740 16192
rect 18796 16183 18836 16192
rect 18987 16232 19029 16241
rect 18987 16192 18988 16232
rect 19028 16192 19029 16232
rect 18987 16183 19029 16192
rect 19084 16232 19124 16435
rect 19179 16400 19221 16409
rect 19179 16360 19180 16400
rect 19220 16360 19313 16400
rect 19179 16351 19221 16360
rect 19273 16316 19313 16360
rect 19273 16276 19316 16316
rect 19180 16232 19220 16241
rect 19084 16192 19180 16232
rect 18988 16064 19028 16183
rect 18699 15896 18741 15905
rect 18699 15856 18700 15896
rect 18740 15856 18741 15896
rect 18699 15847 18741 15856
rect 18411 15728 18453 15737
rect 18411 15688 18412 15728
rect 18452 15688 18453 15728
rect 18411 15679 18453 15688
rect 18699 15728 18741 15737
rect 18699 15688 18700 15728
rect 18740 15688 18741 15728
rect 18699 15679 18741 15688
rect 18796 15732 18836 15741
rect 18124 15560 18164 15571
rect 18124 15485 18164 15520
rect 18123 15476 18165 15485
rect 18123 15436 18124 15476
rect 18164 15436 18165 15476
rect 18123 15427 18165 15436
rect 18316 15317 18356 15402
rect 18124 15308 18164 15317
rect 18124 15065 18164 15268
rect 18315 15308 18357 15317
rect 18315 15268 18316 15308
rect 18356 15268 18357 15308
rect 18315 15259 18357 15268
rect 18412 15140 18452 15679
rect 18316 15100 18452 15140
rect 18604 15560 18644 15569
rect 18123 15056 18165 15065
rect 18123 15016 18124 15056
rect 18164 15016 18165 15056
rect 18123 15007 18165 15016
rect 18028 14848 18164 14888
rect 17836 14671 17876 14680
rect 17932 14720 17972 14729
rect 17835 14048 17877 14057
rect 17835 14008 17836 14048
rect 17876 14008 17877 14048
rect 17835 13999 17877 14008
rect 17836 13914 17876 13999
rect 17932 13889 17972 14680
rect 18028 14552 18068 14561
rect 17931 13880 17973 13889
rect 17931 13840 17932 13880
rect 17972 13840 17973 13880
rect 17931 13831 17973 13840
rect 17739 13460 17781 13469
rect 17739 13420 17740 13460
rect 17780 13420 17781 13460
rect 17739 13411 17781 13420
rect 17739 13292 17781 13301
rect 17739 13252 17740 13292
rect 17780 13252 17781 13292
rect 17739 13243 17781 13252
rect 17740 13049 17780 13243
rect 17739 13040 17781 13049
rect 17739 13000 17740 13040
rect 17780 13000 17781 13040
rect 17739 12991 17781 13000
rect 17740 11537 17780 12991
rect 17739 11528 17781 11537
rect 17739 11488 17740 11528
rect 17780 11488 17781 11528
rect 17739 11479 17781 11488
rect 17643 10688 17685 10697
rect 17643 10648 17644 10688
rect 17684 10648 17685 10688
rect 17643 10639 17685 10648
rect 17446 9680 17488 9689
rect 17547 9680 17589 9689
rect 17446 9640 17447 9680
rect 17487 9640 17492 9680
rect 17446 9631 17492 9640
rect 17547 9640 17548 9680
rect 17588 9640 17589 9680
rect 17547 9631 17589 9640
rect 17452 9512 17492 9631
rect 17452 9463 17492 9472
rect 17643 9512 17685 9521
rect 17643 9472 17644 9512
rect 17684 9472 17685 9512
rect 17643 9463 17685 9472
rect 17644 9378 17684 9463
rect 17451 9260 17493 9269
rect 17451 9220 17452 9260
rect 17492 9220 17493 9260
rect 17451 9211 17493 9220
rect 17452 9126 17492 9211
rect 17356 8884 17492 8924
rect 17067 8840 17109 8849
rect 17067 8800 17068 8840
rect 17108 8800 17109 8840
rect 17067 8791 17109 8800
rect 17259 8840 17301 8849
rect 17259 8800 17260 8840
rect 17300 8800 17301 8840
rect 17259 8791 17301 8800
rect 16972 8703 17097 8743
rect 17057 8686 17097 8703
rect 16875 8672 16917 8681
rect 16875 8632 16876 8672
rect 16916 8632 16917 8672
rect 17057 8672 17108 8686
rect 17356 8681 17396 8766
rect 17452 8765 17492 8884
rect 17451 8756 17493 8765
rect 17451 8716 17452 8756
rect 17492 8716 17493 8756
rect 17451 8707 17493 8716
rect 16875 8623 16917 8632
rect 16972 8651 17012 8660
rect 16588 8212 16820 8252
rect 16683 8084 16725 8093
rect 16683 8044 16684 8084
rect 16724 8044 16725 8084
rect 16683 8035 16725 8044
rect 16588 8000 16628 8009
rect 16588 7832 16628 7960
rect 16684 8000 16724 8035
rect 16684 7949 16724 7960
rect 16588 7792 16724 7832
rect 16491 7580 16533 7589
rect 16491 7540 16492 7580
rect 16532 7540 16533 7580
rect 16491 7531 16533 7540
rect 16684 7505 16724 7792
rect 16780 7748 16820 8212
rect 16876 8009 16916 8623
rect 17057 8646 17068 8672
rect 17068 8623 17108 8632
rect 17355 8672 17397 8681
rect 17355 8632 17356 8672
rect 17396 8632 17397 8672
rect 17355 8623 17397 8632
rect 17644 8672 17684 8681
rect 17740 8672 17780 11479
rect 17932 11360 17972 13831
rect 18028 12629 18068 14512
rect 18124 14468 18164 14848
rect 18219 14720 18261 14729
rect 18219 14680 18220 14720
rect 18260 14680 18261 14720
rect 18219 14671 18261 14680
rect 18316 14720 18356 15100
rect 18507 15056 18549 15065
rect 18507 15016 18508 15056
rect 18548 15016 18549 15056
rect 18507 15007 18549 15016
rect 18508 14813 18548 15007
rect 18507 14804 18549 14813
rect 18507 14764 18508 14804
rect 18548 14764 18549 14804
rect 18507 14755 18549 14764
rect 18316 14671 18356 14680
rect 18412 14720 18452 14731
rect 18604 14729 18644 15520
rect 18700 15560 18740 15679
rect 18700 15511 18740 15520
rect 18796 15485 18836 15692
rect 18988 15569 19028 16024
rect 19084 15737 19124 16192
rect 19180 16183 19220 16192
rect 19276 16232 19316 16276
rect 19276 16183 19316 16192
rect 19275 16064 19317 16073
rect 19275 16024 19276 16064
rect 19316 16024 19317 16064
rect 19275 16015 19317 16024
rect 19083 15728 19125 15737
rect 19083 15688 19084 15728
rect 19124 15688 19125 15728
rect 19083 15679 19125 15688
rect 18987 15560 19029 15569
rect 18987 15520 18988 15560
rect 19028 15520 19029 15560
rect 18987 15511 19029 15520
rect 19084 15560 19124 15679
rect 18795 15476 18837 15485
rect 18795 15436 18796 15476
rect 18836 15436 18837 15476
rect 18795 15427 18837 15436
rect 19084 15317 19124 15520
rect 18699 15308 18741 15317
rect 18699 15268 18700 15308
rect 18740 15268 18741 15308
rect 18699 15259 18741 15268
rect 19083 15308 19125 15317
rect 19083 15268 19084 15308
rect 19124 15268 19125 15308
rect 19083 15259 19125 15268
rect 18220 14586 18260 14671
rect 18412 14645 18452 14680
rect 18603 14720 18645 14729
rect 18603 14680 18604 14720
rect 18644 14680 18645 14720
rect 18603 14671 18645 14680
rect 18700 14720 18740 15259
rect 18808 15140 19176 15149
rect 18848 15100 18890 15140
rect 18930 15100 18972 15140
rect 19012 15100 19054 15140
rect 19094 15100 19136 15140
rect 18808 15091 19176 15100
rect 19276 14972 19316 16015
rect 19372 15560 19412 16444
rect 19468 16325 19508 17200
rect 19756 17081 19796 17166
rect 19755 17072 19797 17081
rect 19755 17032 19756 17072
rect 19796 17032 19797 17072
rect 19755 17023 19797 17032
rect 19564 16820 19604 16829
rect 19564 16400 19604 16780
rect 19755 16820 19797 16829
rect 19755 16780 19756 16820
rect 19796 16780 19797 16820
rect 19755 16771 19797 16780
rect 19756 16686 19796 16771
rect 19948 16493 19988 17536
rect 20048 17408 20416 17417
rect 20088 17368 20130 17408
rect 20170 17368 20212 17408
rect 20252 17368 20294 17408
rect 20334 17368 20376 17408
rect 20048 17359 20416 17368
rect 20044 17072 20084 17081
rect 19947 16484 19989 16493
rect 19947 16444 19948 16484
rect 19988 16444 19989 16484
rect 19947 16435 19989 16444
rect 19564 16360 19892 16400
rect 19467 16316 19509 16325
rect 19467 16276 19468 16316
rect 19508 16276 19509 16316
rect 19467 16267 19509 16276
rect 19468 16064 19508 16073
rect 19468 15737 19508 16024
rect 19467 15728 19509 15737
rect 19467 15688 19468 15728
rect 19508 15688 19509 15728
rect 19467 15679 19509 15688
rect 19372 15233 19412 15520
rect 19467 15560 19509 15569
rect 19467 15520 19468 15560
rect 19508 15520 19509 15560
rect 19467 15511 19509 15520
rect 19468 15426 19508 15511
rect 19467 15308 19509 15317
rect 19467 15268 19468 15308
rect 19508 15268 19509 15308
rect 19467 15259 19509 15268
rect 19371 15224 19413 15233
rect 19371 15184 19372 15224
rect 19412 15184 19413 15224
rect 19371 15175 19413 15184
rect 19468 15140 19508 15259
rect 19564 15224 19604 16360
rect 19659 16232 19701 16241
rect 19659 16192 19660 16232
rect 19700 16192 19701 16232
rect 19659 16183 19701 16192
rect 19852 16232 19892 16360
rect 19852 16183 19892 16192
rect 19948 16232 19988 16241
rect 19660 16098 19700 16183
rect 19755 16064 19797 16073
rect 19755 16024 19756 16064
rect 19796 16024 19797 16064
rect 19755 16015 19797 16024
rect 19756 15930 19796 16015
rect 19948 15812 19988 16192
rect 20044 16073 20084 17032
rect 20043 16064 20085 16073
rect 20043 16024 20044 16064
rect 20084 16024 20085 16064
rect 20043 16015 20085 16024
rect 20620 15989 20660 20140
rect 20715 17996 20757 18005
rect 20715 17956 20716 17996
rect 20756 17956 20757 17996
rect 20715 17947 20757 17956
rect 20619 15980 20661 15989
rect 20619 15940 20620 15980
rect 20660 15940 20661 15980
rect 20619 15931 20661 15940
rect 20048 15896 20416 15905
rect 20088 15856 20130 15896
rect 20170 15856 20212 15896
rect 20252 15856 20294 15896
rect 20334 15856 20376 15896
rect 20048 15847 20416 15856
rect 19756 15772 19988 15812
rect 19756 15392 19796 15772
rect 20043 15728 20085 15737
rect 20043 15688 20044 15728
rect 20084 15688 20180 15728
rect 20043 15679 20085 15688
rect 20140 15602 20180 15688
rect 19948 15560 19988 15569
rect 19756 15343 19796 15352
rect 19852 15520 19948 15560
rect 20140 15553 20180 15562
rect 20236 15560 20276 15569
rect 19852 15233 19892 15520
rect 19948 15511 19988 15520
rect 19947 15308 19989 15317
rect 19947 15268 19948 15308
rect 19988 15268 19989 15308
rect 19947 15259 19989 15268
rect 19659 15224 19701 15233
rect 19564 15184 19660 15224
rect 19700 15184 19701 15224
rect 19659 15175 19701 15184
rect 19851 15224 19893 15233
rect 19851 15184 19852 15224
rect 19892 15184 19893 15224
rect 19851 15175 19893 15184
rect 19948 15174 19988 15259
rect 19468 15100 19604 15140
rect 19371 15056 19413 15065
rect 19371 15016 19372 15056
rect 19412 15016 19413 15056
rect 19371 15007 19413 15016
rect 18988 14932 19316 14972
rect 18891 14888 18933 14897
rect 18891 14848 18892 14888
rect 18932 14848 18933 14888
rect 18891 14839 18933 14848
rect 18700 14671 18740 14680
rect 18796 14804 18836 14813
rect 18411 14636 18453 14645
rect 18411 14596 18412 14636
rect 18452 14596 18453 14636
rect 18411 14587 18453 14596
rect 18508 14552 18548 14561
rect 18796 14552 18836 14764
rect 18892 14754 18932 14839
rect 18988 14804 19028 14932
rect 18988 14755 19028 14764
rect 19083 14804 19125 14813
rect 19083 14764 19084 14804
rect 19124 14764 19125 14804
rect 19083 14755 19125 14764
rect 19084 14720 19124 14755
rect 19084 14669 19124 14680
rect 19275 14720 19317 14729
rect 19275 14680 19276 14720
rect 19316 14680 19317 14720
rect 19275 14671 19317 14680
rect 19372 14720 19412 15007
rect 19467 14972 19509 14981
rect 19467 14932 19468 14972
rect 19508 14932 19509 14972
rect 19467 14923 19509 14932
rect 19372 14671 19412 14680
rect 19468 14720 19508 14923
rect 19564 14897 19604 15100
rect 20236 15065 20276 15520
rect 19659 15056 19701 15065
rect 19659 15016 19660 15056
rect 19700 15016 19701 15056
rect 19659 15007 19701 15016
rect 20235 15056 20277 15065
rect 20235 15016 20236 15056
rect 20276 15016 20277 15056
rect 20235 15007 20277 15016
rect 19563 14888 19605 14897
rect 19563 14848 19564 14888
rect 19604 14848 19605 14888
rect 19563 14839 19605 14848
rect 19468 14671 19508 14680
rect 19564 14720 19604 14839
rect 19564 14671 19604 14680
rect 19276 14586 19316 14671
rect 18548 14512 18836 14552
rect 19563 14552 19605 14561
rect 19563 14512 19564 14552
rect 19604 14512 19605 14552
rect 18508 14503 18548 14512
rect 19563 14503 19605 14512
rect 18411 14468 18453 14477
rect 18124 14428 18260 14468
rect 18123 13460 18165 13469
rect 18123 13420 18124 13460
rect 18164 13420 18165 13460
rect 18123 13411 18165 13420
rect 18027 12620 18069 12629
rect 18027 12580 18028 12620
rect 18068 12580 18069 12620
rect 18027 12571 18069 12580
rect 17836 11320 17972 11360
rect 17836 9512 17876 11320
rect 18027 10772 18069 10781
rect 18027 10732 18028 10772
rect 18068 10732 18069 10772
rect 18027 10723 18069 10732
rect 18028 10193 18068 10723
rect 18027 10184 18069 10193
rect 18027 10144 18028 10184
rect 18068 10144 18069 10184
rect 18027 10135 18069 10144
rect 17931 9680 17973 9689
rect 17931 9640 17932 9680
rect 17972 9640 17973 9680
rect 17931 9631 17973 9640
rect 17932 9546 17972 9631
rect 17836 9176 17876 9472
rect 18028 9512 18068 10135
rect 18028 9463 18068 9472
rect 18124 9512 18164 13411
rect 18220 13217 18260 14428
rect 18411 14428 18412 14468
rect 18452 14428 18453 14468
rect 18411 14419 18453 14428
rect 19083 14468 19125 14477
rect 19083 14428 19084 14468
rect 19124 14428 19125 14468
rect 19083 14419 19125 14428
rect 18219 13208 18261 13217
rect 18219 13168 18220 13208
rect 18260 13168 18261 13208
rect 18219 13159 18261 13168
rect 18412 13208 18452 14419
rect 19084 14048 19124 14419
rect 19468 14048 19508 14057
rect 19084 13999 19124 14008
rect 19372 14008 19468 14048
rect 19275 13880 19317 13889
rect 19275 13840 19276 13880
rect 19316 13840 19317 13880
rect 19275 13831 19317 13840
rect 19276 13746 19316 13831
rect 18808 13628 19176 13637
rect 18848 13588 18890 13628
rect 18930 13588 18972 13628
rect 19012 13588 19054 13628
rect 19094 13588 19136 13628
rect 18808 13579 19176 13588
rect 18603 13460 18645 13469
rect 18603 13420 18604 13460
rect 18644 13420 18645 13460
rect 18603 13411 18645 13420
rect 18891 13460 18933 13469
rect 18891 13420 18892 13460
rect 18932 13420 18933 13460
rect 18891 13411 18933 13420
rect 18604 13326 18644 13411
rect 18452 13168 18644 13208
rect 18412 13159 18452 13168
rect 18604 11696 18644 13168
rect 18892 12762 18932 13411
rect 18987 13376 19029 13385
rect 18987 13336 18988 13376
rect 19028 13336 19029 13376
rect 18987 13327 19029 13336
rect 19179 13376 19221 13385
rect 19179 13336 19180 13376
rect 19220 13336 19221 13376
rect 19179 13327 19221 13336
rect 18892 12713 18932 12722
rect 18988 12713 19028 13327
rect 19180 13208 19220 13327
rect 19180 13159 19220 13168
rect 18987 12704 19029 12713
rect 18987 12664 18988 12704
rect 19028 12664 19029 12704
rect 18987 12655 19029 12664
rect 18700 12536 18740 12545
rect 18700 12041 18740 12496
rect 18988 12536 19028 12655
rect 19083 12620 19125 12629
rect 19083 12580 19084 12620
rect 19124 12580 19125 12620
rect 19083 12571 19125 12580
rect 18988 12487 19028 12496
rect 19084 12536 19124 12571
rect 19084 12485 19124 12496
rect 19275 12536 19317 12545
rect 19275 12496 19276 12536
rect 19316 12496 19317 12536
rect 19275 12487 19317 12496
rect 19276 12293 19316 12487
rect 19372 12368 19412 14008
rect 19468 13999 19508 14008
rect 19564 13964 19604 14503
rect 19660 14141 19700 15007
rect 19756 14888 19796 14897
rect 20043 14888 20085 14897
rect 19796 14848 19891 14888
rect 19756 14839 19796 14848
rect 19851 14813 19891 14848
rect 20043 14848 20044 14888
rect 20084 14848 20085 14888
rect 20043 14839 20085 14848
rect 19851 14804 19893 14813
rect 19851 14764 19852 14804
rect 19892 14764 19893 14804
rect 19851 14755 19893 14764
rect 19756 14678 19796 14731
rect 19755 14638 19756 14645
rect 19947 14720 19989 14729
rect 19947 14680 19948 14720
rect 19988 14680 19989 14720
rect 19947 14671 19989 14680
rect 20044 14720 20084 14839
rect 19796 14638 19797 14645
rect 19755 14636 19797 14638
rect 19755 14596 19756 14636
rect 19796 14596 19797 14636
rect 19755 14587 19797 14596
rect 19948 14586 19988 14671
rect 20044 14645 20084 14680
rect 20043 14636 20085 14645
rect 20043 14596 20044 14636
rect 20084 14596 20085 14636
rect 20043 14587 20085 14596
rect 19947 14468 19989 14477
rect 19947 14428 19948 14468
rect 19988 14428 19989 14468
rect 19947 14419 19989 14428
rect 19659 14132 19701 14141
rect 19659 14092 19660 14132
rect 19700 14092 19701 14132
rect 19659 14083 19701 14092
rect 19851 14048 19893 14057
rect 19851 14008 19852 14048
rect 19892 14008 19893 14048
rect 19948 14048 19988 14419
rect 20048 14384 20416 14393
rect 20088 14344 20130 14384
rect 20170 14344 20212 14384
rect 20252 14344 20294 14384
rect 20334 14344 20376 14384
rect 20048 14335 20416 14344
rect 20139 14132 20181 14141
rect 20139 14092 20140 14132
rect 20180 14092 20181 14132
rect 20139 14083 20181 14092
rect 20044 14048 20084 14057
rect 19948 14008 20044 14048
rect 19851 13999 19893 14008
rect 20044 13999 20084 14008
rect 19564 13915 19604 13924
rect 19756 13964 19796 13973
rect 19467 13880 19509 13889
rect 19467 13840 19468 13880
rect 19508 13840 19509 13880
rect 19467 13831 19509 13840
rect 19660 13880 19700 13889
rect 19468 13712 19508 13831
rect 19468 13672 19604 13712
rect 19467 13208 19509 13217
rect 19467 13168 19468 13208
rect 19508 13168 19509 13208
rect 19467 13159 19509 13168
rect 19564 13208 19604 13672
rect 19564 13159 19604 13168
rect 19468 13074 19508 13159
rect 19660 12872 19700 13840
rect 19372 12319 19412 12328
rect 19468 12832 19700 12872
rect 19275 12284 19317 12293
rect 19275 12244 19276 12284
rect 19316 12244 19317 12284
rect 19275 12235 19317 12244
rect 18808 12116 19176 12125
rect 18848 12076 18890 12116
rect 18930 12076 18972 12116
rect 19012 12076 19054 12116
rect 19094 12076 19136 12116
rect 18808 12067 19176 12076
rect 18699 12032 18741 12041
rect 18699 11992 18700 12032
rect 18740 11992 18741 12032
rect 18699 11983 18741 11992
rect 19468 11957 19508 12832
rect 19564 12704 19604 12713
rect 19756 12704 19796 13924
rect 19852 13914 19892 13999
rect 20140 13998 20180 14083
rect 20236 14048 20276 14057
rect 20716 14048 20756 17947
rect 21100 17417 21140 25675
rect 21195 24800 21237 24809
rect 21195 24760 21196 24800
rect 21236 24760 21237 24800
rect 21195 24751 21237 24760
rect 21196 22457 21236 24751
rect 21195 22448 21237 22457
rect 21195 22408 21196 22448
rect 21236 22408 21237 22448
rect 21195 22399 21237 22408
rect 21292 20180 21332 28867
rect 21387 26648 21429 26657
rect 21387 26608 21388 26648
rect 21428 26608 21429 26648
rect 21387 26599 21429 26608
rect 21388 26489 21428 26599
rect 21387 26480 21429 26489
rect 21387 26440 21388 26480
rect 21428 26440 21429 26480
rect 21387 26431 21429 26440
rect 21387 25808 21429 25817
rect 21387 25768 21388 25808
rect 21428 25768 21429 25808
rect 21387 25759 21429 25768
rect 21388 25481 21428 25759
rect 21387 25472 21429 25481
rect 21387 25432 21388 25472
rect 21428 25432 21429 25472
rect 21387 25423 21429 25432
rect 21387 25136 21429 25145
rect 21387 25096 21388 25136
rect 21428 25096 21429 25136
rect 21387 25087 21429 25096
rect 21388 24977 21428 25087
rect 21387 24968 21429 24977
rect 21387 24928 21388 24968
rect 21428 24928 21429 24968
rect 21387 24919 21429 24928
rect 21196 20140 21332 20180
rect 21099 17408 21141 17417
rect 21099 17368 21100 17408
rect 21140 17368 21141 17408
rect 21099 17359 21141 17368
rect 21196 15401 21236 20140
rect 21387 19760 21429 19769
rect 21387 19720 21388 19760
rect 21428 19720 21429 19760
rect 21387 19711 21429 19720
rect 21388 18929 21428 19711
rect 21387 18920 21429 18929
rect 21387 18880 21388 18920
rect 21428 18880 21429 18920
rect 21387 18871 21429 18880
rect 21195 15392 21237 15401
rect 21195 15352 21196 15392
rect 21236 15352 21237 15392
rect 21195 15343 21237 15352
rect 21195 14384 21237 14393
rect 21195 14344 21196 14384
rect 21236 14344 21237 14384
rect 21195 14335 21237 14344
rect 20276 14008 20756 14048
rect 19947 13880 19989 13889
rect 19947 13840 19948 13880
rect 19988 13840 19989 13880
rect 19947 13831 19989 13840
rect 19851 13376 19893 13385
rect 19851 13336 19852 13376
rect 19892 13336 19893 13376
rect 19851 13327 19893 13336
rect 19852 13242 19892 13327
rect 19851 13040 19893 13049
rect 19851 13000 19852 13040
rect 19892 13000 19893 13040
rect 19851 12991 19893 13000
rect 19852 12713 19892 12991
rect 19467 11948 19509 11957
rect 19467 11908 19468 11948
rect 19508 11908 19509 11948
rect 19467 11899 19509 11908
rect 19083 11864 19125 11873
rect 19083 11824 19084 11864
rect 19124 11824 19125 11864
rect 19083 11815 19125 11824
rect 19084 11730 19124 11815
rect 18604 11360 18644 11656
rect 19467 11696 19509 11705
rect 19467 11656 19468 11696
rect 19508 11656 19509 11696
rect 19467 11647 19509 11656
rect 18795 11612 18837 11621
rect 18795 11572 18796 11612
rect 18836 11572 18837 11612
rect 18795 11563 18837 11572
rect 19372 11612 19412 11623
rect 18796 11478 18836 11563
rect 19372 11537 19412 11572
rect 19468 11562 19508 11647
rect 19371 11528 19413 11537
rect 19371 11488 19372 11528
rect 19412 11488 19413 11528
rect 19371 11479 19413 11488
rect 19564 11360 19604 12664
rect 18220 11320 18836 11360
rect 18220 11024 18260 11320
rect 18411 11192 18453 11201
rect 18411 11152 18412 11192
rect 18452 11152 18453 11192
rect 18411 11143 18453 11152
rect 18699 11192 18741 11201
rect 18699 11152 18700 11192
rect 18740 11152 18741 11192
rect 18699 11143 18741 11152
rect 18412 11058 18452 11143
rect 18220 10975 18260 10984
rect 18507 11024 18549 11033
rect 18507 10984 18508 11024
rect 18548 10984 18549 11024
rect 18507 10975 18549 10984
rect 18700 11024 18740 11143
rect 18700 10975 18740 10984
rect 18219 10100 18261 10109
rect 18219 10060 18220 10100
rect 18260 10060 18261 10100
rect 18219 10051 18261 10060
rect 18124 9463 18164 9472
rect 18220 9260 18260 10051
rect 18315 9512 18357 9521
rect 18315 9472 18316 9512
rect 18356 9472 18357 9512
rect 18315 9463 18357 9472
rect 18316 9378 18356 9463
rect 18220 9220 18356 9260
rect 17836 9136 18068 9176
rect 18028 8849 18068 9136
rect 17835 8840 17877 8849
rect 17835 8800 17836 8840
rect 17876 8800 17877 8840
rect 17835 8791 17877 8800
rect 18027 8840 18069 8849
rect 18027 8800 18028 8840
rect 18068 8800 18069 8840
rect 18027 8791 18069 8800
rect 18220 8840 18260 8849
rect 17684 8632 17780 8672
rect 17836 8672 17876 8791
rect 16972 8597 17012 8611
rect 16971 8588 17013 8597
rect 16971 8548 16972 8588
rect 17012 8548 17013 8588
rect 16971 8539 17013 8548
rect 17164 8588 17204 8597
rect 17204 8548 17300 8588
rect 17164 8539 17204 8548
rect 16972 8516 17012 8539
rect 17260 8345 17300 8548
rect 17452 8504 17492 8513
rect 17356 8464 17452 8504
rect 17259 8336 17301 8345
rect 17259 8296 17260 8336
rect 17300 8296 17301 8336
rect 17259 8287 17301 8296
rect 17163 8168 17205 8177
rect 17163 8128 17164 8168
rect 17204 8128 17205 8168
rect 17163 8119 17205 8128
rect 16971 8084 17013 8093
rect 16971 8044 16972 8084
rect 17012 8044 17013 8084
rect 16971 8035 17013 8044
rect 16875 8000 16917 8009
rect 16875 7960 16876 8000
rect 16916 7960 16917 8000
rect 16875 7951 16917 7960
rect 16972 8000 17012 8035
rect 17164 8034 17204 8119
rect 16972 7949 17012 7960
rect 17067 8000 17109 8009
rect 17067 7960 17068 8000
rect 17108 7960 17109 8000
rect 17067 7951 17109 7960
rect 17260 8000 17300 8009
rect 17356 8000 17396 8464
rect 17452 8455 17492 8464
rect 17644 8345 17684 8632
rect 17836 8623 17876 8632
rect 18028 8672 18068 8681
rect 17931 8504 17973 8513
rect 17931 8464 17932 8504
rect 17972 8464 17973 8504
rect 17931 8455 17973 8464
rect 17835 8420 17877 8429
rect 17835 8380 17836 8420
rect 17876 8380 17877 8420
rect 17835 8371 17877 8380
rect 17451 8336 17493 8345
rect 17451 8296 17452 8336
rect 17492 8296 17493 8336
rect 17451 8287 17493 8296
rect 17643 8336 17685 8345
rect 17643 8296 17644 8336
rect 17684 8296 17685 8336
rect 17643 8287 17685 8296
rect 17300 7960 17396 8000
rect 17452 8000 17492 8287
rect 17547 8168 17589 8177
rect 17547 8128 17548 8168
rect 17588 8128 17589 8168
rect 17547 8119 17589 8128
rect 17548 8034 17588 8119
rect 17260 7951 17300 7960
rect 17452 7951 17492 7960
rect 17643 8000 17685 8009
rect 17643 7960 17644 8000
rect 17684 7960 17685 8000
rect 17643 7951 17685 7960
rect 17740 8000 17780 8009
rect 17836 8000 17876 8371
rect 17932 8370 17972 8455
rect 18028 8177 18068 8632
rect 18220 8261 18260 8800
rect 18316 8681 18356 9220
rect 18508 8756 18548 10975
rect 18603 10940 18645 10949
rect 18603 10900 18604 10940
rect 18644 10900 18645 10940
rect 18603 10891 18645 10900
rect 18604 8840 18644 10891
rect 18796 10856 18836 11320
rect 19276 11320 19604 11360
rect 19660 12664 19796 12704
rect 19851 12704 19893 12713
rect 19851 12664 19852 12704
rect 19892 12664 19893 12704
rect 18987 11276 19029 11285
rect 18987 11236 18988 11276
rect 19028 11236 19029 11276
rect 18987 11227 19029 11236
rect 19179 11276 19221 11285
rect 19179 11236 19180 11276
rect 19220 11236 19221 11276
rect 19179 11227 19221 11236
rect 18988 11024 19028 11227
rect 19180 11117 19220 11227
rect 19179 11108 19221 11117
rect 19179 11068 19180 11108
rect 19220 11068 19221 11108
rect 19179 11059 19221 11068
rect 18988 10975 19028 10984
rect 19084 11024 19124 11033
rect 19084 10865 19124 10984
rect 18700 10816 18836 10856
rect 19083 10856 19125 10865
rect 19083 10816 19084 10856
rect 19124 10816 19125 10856
rect 18700 10184 18740 10816
rect 19083 10807 19125 10816
rect 18808 10604 19176 10613
rect 18848 10564 18890 10604
rect 18930 10564 18972 10604
rect 19012 10564 19054 10604
rect 19094 10564 19136 10604
rect 18808 10555 19176 10564
rect 18795 10436 18837 10445
rect 18892 10436 18932 10445
rect 18795 10396 18796 10436
rect 18836 10396 18892 10436
rect 18795 10387 18837 10396
rect 18892 10387 18932 10396
rect 18700 9521 18740 10144
rect 18699 9512 18741 9521
rect 18699 9472 18700 9512
rect 18740 9472 18741 9512
rect 18699 9463 18741 9472
rect 18796 9260 18836 10387
rect 19084 10352 19124 10361
rect 19084 10193 19124 10312
rect 19083 10184 19125 10193
rect 19083 10144 19084 10184
rect 19124 10144 19125 10184
rect 19083 10135 19125 10144
rect 18700 9220 18836 9260
rect 18700 8924 18740 9220
rect 18808 9092 19176 9101
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 18808 9043 19176 9052
rect 18700 8884 18836 8924
rect 18604 8800 18740 8840
rect 18412 8716 18548 8756
rect 18315 8672 18357 8681
rect 18315 8632 18316 8672
rect 18356 8632 18357 8672
rect 18315 8623 18357 8632
rect 18219 8252 18261 8261
rect 18219 8212 18220 8252
rect 18260 8212 18261 8252
rect 18219 8203 18261 8212
rect 18027 8168 18069 8177
rect 18027 8128 18028 8168
rect 18068 8128 18069 8168
rect 18027 8119 18069 8128
rect 17931 8000 17973 8009
rect 17836 7960 17932 8000
rect 17972 7960 17973 8000
rect 17068 7866 17108 7951
rect 17644 7866 17684 7951
rect 17643 7748 17685 7757
rect 16780 7708 17204 7748
rect 17067 7580 17109 7589
rect 17067 7540 17068 7580
rect 17108 7540 17109 7580
rect 17067 7531 17109 7540
rect 16683 7496 16725 7505
rect 16683 7456 16684 7496
rect 16724 7456 16725 7496
rect 16683 7447 16725 7456
rect 16587 7412 16629 7421
rect 16587 7372 16588 7412
rect 16628 7372 16629 7412
rect 16587 7363 16629 7372
rect 16492 7160 16532 7169
rect 16492 6740 16532 7120
rect 16588 7160 16628 7363
rect 17068 7244 17108 7531
rect 17068 7195 17108 7204
rect 16588 7111 16628 7120
rect 16972 7160 17012 7169
rect 16972 7001 17012 7120
rect 16971 6992 17013 7001
rect 16971 6952 16972 6992
rect 17012 6952 17013 6992
rect 16971 6943 17013 6952
rect 16492 6700 16628 6740
rect 16396 6616 16532 6656
rect 16300 6439 16340 6448
rect 16396 6488 16436 6499
rect 16108 6354 16148 6439
rect 16396 6413 16436 6448
rect 16395 6404 16437 6413
rect 16395 6364 16396 6404
rect 16436 6364 16437 6404
rect 16395 6355 16437 6364
rect 16108 6236 16148 6245
rect 16108 5825 16148 6196
rect 16203 6236 16245 6245
rect 16203 6196 16204 6236
rect 16244 6196 16245 6236
rect 16203 6187 16245 6196
rect 16107 5816 16149 5825
rect 16107 5776 16108 5816
rect 16148 5776 16149 5816
rect 16107 5767 16149 5776
rect 16108 5648 16148 5657
rect 16108 5405 16148 5608
rect 16107 5396 16149 5405
rect 16107 5356 16108 5396
rect 16148 5356 16149 5396
rect 16107 5347 16149 5356
rect 16012 4087 16052 4096
rect 16108 4976 16148 4985
rect 15820 3928 15956 3968
rect 15723 3884 15765 3893
rect 15723 3844 15724 3884
rect 15764 3844 15765 3884
rect 15723 3835 15765 3844
rect 15724 3464 15764 3835
rect 15819 3548 15861 3557
rect 15819 3508 15820 3548
rect 15860 3508 15861 3548
rect 15819 3499 15861 3508
rect 15724 3415 15764 3424
rect 15820 3464 15860 3499
rect 15820 2717 15860 3424
rect 15916 2969 15956 3928
rect 16108 3473 16148 4936
rect 16204 3968 16244 6187
rect 16395 6152 16437 6161
rect 16395 6112 16396 6152
rect 16436 6112 16437 6152
rect 16395 6103 16437 6112
rect 16299 5816 16341 5825
rect 16299 5776 16300 5816
rect 16340 5776 16341 5816
rect 16299 5767 16341 5776
rect 16204 3919 16244 3928
rect 16300 3632 16340 5767
rect 16396 5648 16436 6103
rect 16396 5599 16436 5608
rect 16396 4145 16436 4230
rect 16395 4136 16437 4145
rect 16395 4096 16396 4136
rect 16436 4096 16437 4136
rect 16395 4087 16437 4096
rect 16492 3968 16532 6616
rect 16588 6581 16628 6700
rect 16587 6572 16629 6581
rect 16587 6532 16588 6572
rect 16628 6532 16629 6572
rect 16587 6523 16629 6532
rect 16683 6488 16725 6497
rect 16683 6448 16684 6488
rect 16724 6448 16725 6488
rect 16683 6439 16725 6448
rect 16972 6488 17012 6497
rect 17012 6448 17108 6488
rect 16972 6439 17012 6448
rect 16587 6320 16629 6329
rect 16587 6280 16588 6320
rect 16628 6280 16629 6320
rect 16587 6271 16629 6280
rect 16588 6186 16628 6271
rect 16587 5480 16629 5489
rect 16587 5440 16588 5480
rect 16628 5440 16629 5480
rect 16587 5431 16629 5440
rect 16204 3592 16340 3632
rect 16396 3928 16532 3968
rect 16107 3464 16149 3473
rect 16107 3424 16108 3464
rect 16148 3424 16149 3464
rect 16107 3415 16149 3424
rect 15915 2960 15957 2969
rect 15915 2920 15916 2960
rect 15956 2920 15957 2960
rect 15915 2911 15957 2920
rect 16204 2801 16244 3592
rect 16299 3464 16341 3473
rect 16299 3424 16300 3464
rect 16340 3424 16341 3464
rect 16299 3415 16341 3424
rect 16300 3330 16340 3415
rect 16203 2792 16245 2801
rect 16203 2752 16204 2792
rect 16244 2752 16245 2792
rect 16203 2743 16245 2752
rect 15819 2708 15861 2717
rect 15819 2668 15820 2708
rect 15860 2668 15861 2708
rect 15819 2659 15861 2668
rect 16012 2633 16052 2718
rect 16011 2624 16053 2633
rect 16011 2584 16012 2624
rect 16052 2584 16053 2624
rect 16011 2575 16053 2584
rect 15723 2204 15765 2213
rect 15723 2164 15724 2204
rect 15764 2164 15765 2204
rect 15723 2155 15765 2164
rect 15724 1952 15764 2155
rect 16011 2036 16053 2045
rect 16011 1996 16012 2036
rect 16052 1996 16053 2036
rect 16011 1987 16053 1996
rect 15724 1903 15764 1912
rect 15627 1616 15669 1625
rect 15627 1576 15628 1616
rect 15668 1576 15669 1616
rect 15627 1567 15669 1576
rect 14956 1324 15092 1364
rect 14956 1196 14996 1205
rect 14956 953 14996 1156
rect 14955 944 14997 953
rect 14955 904 14956 944
rect 14996 904 14997 944
rect 14955 895 14997 904
rect 15052 80 15092 1324
rect 15435 1280 15477 1289
rect 15435 1240 15436 1280
rect 15476 1240 15477 1280
rect 15435 1231 15477 1240
rect 15627 1280 15669 1289
rect 15627 1240 15628 1280
rect 15668 1240 15669 1280
rect 15627 1231 15669 1240
rect 15243 1112 15285 1121
rect 15243 1072 15244 1112
rect 15284 1072 15285 1112
rect 15243 1063 15285 1072
rect 15244 978 15284 1063
rect 15243 608 15285 617
rect 15243 568 15244 608
rect 15284 568 15285 608
rect 15243 559 15285 568
rect 15244 80 15284 559
rect 15436 80 15476 1231
rect 15628 80 15668 1231
rect 15819 356 15861 365
rect 15819 316 15820 356
rect 15860 316 15861 356
rect 15819 307 15861 316
rect 15820 80 15860 307
rect 16012 80 16052 1987
rect 16107 272 16149 281
rect 16107 232 16108 272
rect 16148 232 16244 272
rect 16107 223 16149 232
rect 16204 80 16244 232
rect 16396 80 16436 3928
rect 16588 2885 16628 5431
rect 16587 2876 16629 2885
rect 16587 2836 16588 2876
rect 16628 2836 16629 2876
rect 16587 2827 16629 2836
rect 16540 2666 16580 2675
rect 16580 2626 16628 2643
rect 16540 2603 16628 2626
rect 16588 2372 16628 2603
rect 16684 2540 16724 6439
rect 16971 5144 17013 5153
rect 16971 5104 16972 5144
rect 17012 5104 17013 5144
rect 16971 5095 17013 5104
rect 16972 3632 17012 5095
rect 16972 3583 17012 3592
rect 16684 2491 16724 2500
rect 16780 3450 16820 3459
rect 16780 2372 16820 3410
rect 17068 3380 17108 6448
rect 17164 6320 17204 7708
rect 17643 7708 17644 7748
rect 17684 7708 17685 7748
rect 17740 7748 17780 7960
rect 17931 7951 17973 7960
rect 18220 8000 18260 8009
rect 17932 7866 17972 7951
rect 18028 7748 18068 7757
rect 17740 7708 18028 7748
rect 17643 7699 17685 7708
rect 17547 7244 17589 7253
rect 17547 7204 17548 7244
rect 17588 7204 17589 7244
rect 17547 7195 17589 7204
rect 17548 7160 17588 7195
rect 17548 6749 17588 7120
rect 17547 6740 17589 6749
rect 17547 6700 17548 6740
rect 17588 6700 17589 6740
rect 17547 6691 17589 6700
rect 17260 6497 17300 6582
rect 17547 6572 17589 6581
rect 17547 6532 17548 6572
rect 17588 6532 17589 6572
rect 17547 6523 17589 6532
rect 17259 6488 17301 6497
rect 17259 6448 17260 6488
rect 17300 6448 17301 6488
rect 17259 6439 17301 6448
rect 17356 6488 17396 6497
rect 17164 6280 17300 6320
rect 17163 6068 17205 6077
rect 17163 6028 17164 6068
rect 17204 6028 17205 6068
rect 17163 6019 17205 6028
rect 17164 4985 17204 6019
rect 17163 4976 17205 4985
rect 17163 4936 17164 4976
rect 17204 4936 17205 4976
rect 17163 4927 17205 4936
rect 17164 3893 17204 4927
rect 17163 3884 17205 3893
rect 17163 3844 17164 3884
rect 17204 3844 17205 3884
rect 17163 3835 17205 3844
rect 17164 3464 17204 3835
rect 17260 3464 17300 6280
rect 17356 5153 17396 6448
rect 17451 6488 17493 6497
rect 17451 6448 17452 6488
rect 17492 6448 17493 6488
rect 17451 6439 17493 6448
rect 17355 5144 17397 5153
rect 17355 5104 17356 5144
rect 17396 5104 17397 5144
rect 17355 5095 17397 5104
rect 17356 4976 17396 4985
rect 17356 3809 17396 4936
rect 17355 3800 17397 3809
rect 17355 3760 17356 3800
rect 17396 3760 17397 3800
rect 17355 3751 17397 3760
rect 17356 3632 17396 3641
rect 17452 3632 17492 6439
rect 17396 3592 17492 3632
rect 17548 5060 17588 6523
rect 17644 6320 17684 7699
rect 18028 7412 18068 7708
rect 18220 7673 18260 7960
rect 18219 7664 18261 7673
rect 18219 7624 18220 7664
rect 18260 7624 18261 7664
rect 18219 7615 18261 7624
rect 18028 7372 18356 7412
rect 17931 7328 17973 7337
rect 17931 7288 17932 7328
rect 17972 7288 18164 7328
rect 17931 7279 17973 7288
rect 18028 7165 18068 7174
rect 18028 6740 18068 7125
rect 17644 6271 17684 6280
rect 17740 6700 18068 6740
rect 17643 6152 17685 6161
rect 17643 6112 17644 6152
rect 17684 6112 17685 6152
rect 17643 6103 17685 6112
rect 17356 3583 17396 3592
rect 17452 3464 17492 3473
rect 17548 3464 17588 5020
rect 17644 5648 17684 6103
rect 17644 4136 17684 5608
rect 17740 5144 17780 6700
rect 18027 6572 18069 6581
rect 18027 6532 18028 6572
rect 18068 6532 18069 6572
rect 18027 6523 18069 6532
rect 17835 6488 17877 6497
rect 17835 6448 17836 6488
rect 17876 6448 17877 6488
rect 17835 6439 17877 6448
rect 18028 6488 18068 6523
rect 17836 6354 17876 6439
rect 17836 6236 17876 6245
rect 17836 5741 17876 6196
rect 18028 6161 18068 6448
rect 18124 6488 18164 7288
rect 18124 6439 18164 6448
rect 18220 6992 18260 7001
rect 18027 6152 18069 6161
rect 18027 6112 18028 6152
rect 18068 6112 18069 6152
rect 18027 6103 18069 6112
rect 17931 5816 17973 5825
rect 17931 5776 17932 5816
rect 17972 5776 17973 5816
rect 17931 5767 17973 5776
rect 17835 5732 17877 5741
rect 17835 5692 17836 5732
rect 17876 5692 17877 5732
rect 17835 5683 17877 5692
rect 17835 5480 17877 5489
rect 17835 5440 17836 5480
rect 17876 5440 17877 5480
rect 17835 5431 17877 5440
rect 17836 5346 17876 5431
rect 17835 5144 17877 5153
rect 17740 5104 17836 5144
rect 17876 5104 17877 5144
rect 17835 5095 17877 5104
rect 17739 4976 17781 4985
rect 17739 4936 17740 4976
rect 17780 4936 17781 4976
rect 17739 4927 17781 4936
rect 17740 4842 17780 4927
rect 17836 4388 17876 5095
rect 17836 4339 17876 4348
rect 17739 4220 17781 4229
rect 17739 4180 17740 4220
rect 17780 4180 17781 4220
rect 17739 4171 17781 4180
rect 17644 3809 17684 4096
rect 17740 3893 17780 4171
rect 17836 3968 17876 3977
rect 17739 3884 17781 3893
rect 17739 3844 17740 3884
rect 17780 3844 17781 3884
rect 17739 3835 17781 3844
rect 17836 3809 17876 3928
rect 17643 3800 17685 3809
rect 17643 3760 17644 3800
rect 17684 3760 17685 3800
rect 17643 3751 17685 3760
rect 17835 3800 17877 3809
rect 17835 3760 17836 3800
rect 17876 3760 17877 3800
rect 17835 3751 17877 3760
rect 17643 3632 17685 3641
rect 17643 3592 17644 3632
rect 17684 3592 17685 3632
rect 17643 3583 17685 3592
rect 17260 3424 17396 3464
rect 17164 3415 17204 3424
rect 16972 3340 17108 3380
rect 16875 2456 16917 2465
rect 16875 2416 16876 2456
rect 16916 2416 16917 2456
rect 16875 2407 16917 2416
rect 16588 2332 16820 2372
rect 16588 2129 16628 2332
rect 16876 2322 16916 2407
rect 16587 2120 16629 2129
rect 16972 2120 17012 3340
rect 17067 3212 17109 3221
rect 17067 3172 17068 3212
rect 17108 3172 17109 3212
rect 17067 3163 17109 3172
rect 17068 2708 17108 3163
rect 17068 2659 17108 2668
rect 17260 2456 17300 2465
rect 17164 2129 17204 2214
rect 16587 2080 16588 2120
rect 16628 2080 16629 2120
rect 16587 2071 16629 2080
rect 16684 2080 17012 2120
rect 17163 2120 17205 2129
rect 17163 2080 17164 2120
rect 17204 2080 17205 2120
rect 16491 1784 16533 1793
rect 16491 1744 16492 1784
rect 16532 1744 16533 1784
rect 16491 1735 16533 1744
rect 16492 1112 16532 1735
rect 16684 1280 16724 2080
rect 17163 2071 17205 2080
rect 16971 1952 17013 1961
rect 17260 1952 17300 2416
rect 16971 1912 16972 1952
rect 17012 1912 17013 1952
rect 16971 1903 17013 1912
rect 17164 1912 17300 1952
rect 16684 1231 16724 1240
rect 16492 953 16532 1072
rect 16491 944 16533 953
rect 16491 904 16492 944
rect 16532 904 16533 944
rect 16491 895 16533 904
rect 16779 944 16821 953
rect 16779 904 16780 944
rect 16820 904 16821 944
rect 16779 895 16821 904
rect 16876 944 16916 953
rect 16780 524 16820 895
rect 16876 701 16916 904
rect 16972 860 17012 1903
rect 17164 1457 17204 1912
rect 17356 1868 17396 3424
rect 17492 3424 17588 3464
rect 17452 3415 17492 3424
rect 17644 2792 17684 3583
rect 17835 3548 17877 3557
rect 17835 3508 17836 3548
rect 17876 3508 17877 3548
rect 17835 3499 17877 3508
rect 17451 2708 17493 2717
rect 17451 2668 17452 2708
rect 17492 2668 17493 2708
rect 17451 2659 17493 2668
rect 17452 2574 17492 2659
rect 17644 2540 17684 2752
rect 17260 1828 17396 1868
rect 17548 2500 17684 2540
rect 17740 3464 17780 3473
rect 17740 2624 17780 3424
rect 17836 3464 17876 3499
rect 17836 3413 17876 3424
rect 17932 2969 17972 5767
rect 18028 5648 18068 6103
rect 18220 5825 18260 6952
rect 18316 6488 18356 7372
rect 18412 6749 18452 8716
rect 18603 8672 18645 8681
rect 18603 8632 18604 8672
rect 18644 8632 18645 8672
rect 18603 8623 18645 8632
rect 18507 8588 18549 8597
rect 18507 8548 18508 8588
rect 18548 8548 18549 8588
rect 18507 8539 18549 8548
rect 18508 8454 18548 8539
rect 18604 8538 18644 8623
rect 18603 8000 18645 8009
rect 18603 7960 18604 8000
rect 18644 7960 18645 8000
rect 18603 7951 18645 7960
rect 18604 7589 18644 7951
rect 18603 7580 18645 7589
rect 18603 7540 18604 7580
rect 18644 7540 18645 7580
rect 18603 7531 18645 7540
rect 18604 7328 18644 7337
rect 18604 7169 18644 7288
rect 18603 7160 18645 7169
rect 18603 7120 18604 7160
rect 18644 7120 18645 7160
rect 18603 7111 18645 7120
rect 18411 6740 18453 6749
rect 18411 6700 18412 6740
rect 18452 6700 18453 6740
rect 18411 6691 18453 6700
rect 18508 6665 18548 6750
rect 18507 6656 18549 6665
rect 18507 6616 18508 6656
rect 18548 6616 18549 6656
rect 18507 6607 18549 6616
rect 18316 6439 18356 6448
rect 18412 6488 18452 6497
rect 18412 6161 18452 6448
rect 18508 6477 18644 6488
rect 18508 6448 18604 6477
rect 18411 6152 18453 6161
rect 18411 6112 18412 6152
rect 18452 6112 18453 6152
rect 18411 6103 18453 6112
rect 18508 5984 18548 6448
rect 18604 6428 18644 6437
rect 18316 5944 18548 5984
rect 18219 5816 18261 5825
rect 18219 5776 18220 5816
rect 18260 5776 18261 5816
rect 18219 5767 18261 5776
rect 18028 5599 18068 5608
rect 18123 5648 18165 5657
rect 18123 5608 18124 5648
rect 18164 5608 18165 5648
rect 18123 5599 18165 5608
rect 18220 5648 18260 5657
rect 18124 5514 18164 5599
rect 18123 5396 18165 5405
rect 18123 5356 18124 5396
rect 18164 5356 18165 5396
rect 18123 5347 18165 5356
rect 18027 4976 18069 4985
rect 18027 4936 18028 4976
rect 18068 4936 18069 4976
rect 18027 4927 18069 4936
rect 18124 4976 18164 5347
rect 18220 5153 18260 5608
rect 18316 5648 18356 5944
rect 18316 5599 18356 5608
rect 18508 5648 18548 5657
rect 18508 5237 18548 5608
rect 18507 5228 18549 5237
rect 18507 5188 18508 5228
rect 18548 5188 18549 5228
rect 18507 5179 18549 5188
rect 18219 5144 18261 5153
rect 18219 5104 18220 5144
rect 18260 5104 18261 5144
rect 18219 5095 18261 5104
rect 18411 5144 18453 5153
rect 18411 5104 18412 5144
rect 18452 5104 18453 5144
rect 18411 5095 18453 5104
rect 18028 4842 18068 4927
rect 18027 4556 18069 4565
rect 18027 4516 18028 4556
rect 18068 4516 18069 4556
rect 18027 4507 18069 4516
rect 18028 4136 18068 4507
rect 18028 4087 18068 4096
rect 18124 4136 18164 4936
rect 18219 4976 18261 4985
rect 18219 4936 18220 4976
rect 18260 4936 18261 4976
rect 18219 4927 18261 4936
rect 18316 4976 18356 4985
rect 18412 4976 18452 5095
rect 18356 4936 18452 4976
rect 18508 4976 18548 4985
rect 18603 4976 18645 4985
rect 18548 4936 18604 4976
rect 18644 4936 18645 4976
rect 18316 4927 18356 4936
rect 18508 4927 18548 4936
rect 18603 4927 18645 4936
rect 18124 4087 18164 4096
rect 18220 4052 18260 4927
rect 18700 4817 18740 8800
rect 18796 8093 18836 8884
rect 19179 8840 19221 8849
rect 19179 8800 19180 8840
rect 19220 8800 19221 8840
rect 19179 8791 19221 8800
rect 18892 8672 18932 8681
rect 18892 8177 18932 8632
rect 19180 8672 19220 8791
rect 19276 8672 19316 11320
rect 19660 11117 19700 12664
rect 19851 12655 19893 12664
rect 19756 12536 19796 12547
rect 19756 12461 19796 12496
rect 19852 12536 19892 12655
rect 19852 12487 19892 12496
rect 19755 12452 19797 12461
rect 19755 12412 19756 12452
rect 19796 12412 19797 12452
rect 19755 12403 19797 12412
rect 19851 12284 19893 12293
rect 19851 12244 19852 12284
rect 19892 12244 19893 12284
rect 19851 12235 19893 12244
rect 19756 11696 19796 11705
rect 19756 11285 19796 11656
rect 19755 11276 19797 11285
rect 19755 11236 19756 11276
rect 19796 11236 19797 11276
rect 19755 11227 19797 11236
rect 19659 11108 19701 11117
rect 19852 11108 19892 12235
rect 19948 11957 19988 13831
rect 20044 13208 20084 13217
rect 20044 13049 20084 13168
rect 20140 13133 20180 13218
rect 20236 13208 20276 14008
rect 20236 13159 20276 13168
rect 20139 13124 20181 13133
rect 20139 13084 20140 13124
rect 20180 13084 20181 13124
rect 20139 13075 20181 13084
rect 20043 13040 20085 13049
rect 20043 13000 20044 13040
rect 20084 13000 20085 13040
rect 20043 12991 20085 13000
rect 20048 12872 20416 12881
rect 20088 12832 20130 12872
rect 20170 12832 20212 12872
rect 20252 12832 20294 12872
rect 20334 12832 20376 12872
rect 20048 12823 20416 12832
rect 20236 12452 20276 12461
rect 20276 12412 20372 12452
rect 20236 12403 20276 12412
rect 20043 12284 20085 12293
rect 20043 12244 20044 12284
rect 20084 12244 20085 12284
rect 20043 12235 20085 12244
rect 20044 12150 20084 12235
rect 20332 12032 20372 12412
rect 20524 12209 20564 14008
rect 20523 12200 20565 12209
rect 20523 12160 20524 12200
rect 20564 12160 20565 12200
rect 20523 12151 20565 12160
rect 20620 12076 20948 12116
rect 20620 12032 20660 12076
rect 20332 11992 20660 12032
rect 19947 11948 19989 11957
rect 19947 11908 19948 11948
rect 19988 11908 19989 11948
rect 19947 11899 19989 11908
rect 20715 11948 20757 11957
rect 20715 11908 20716 11948
rect 20756 11908 20757 11948
rect 20715 11899 20757 11908
rect 19948 11621 19988 11899
rect 20236 11780 20276 11789
rect 20276 11740 20660 11780
rect 20236 11731 20276 11740
rect 19947 11612 19989 11621
rect 19947 11572 19948 11612
rect 19988 11572 19989 11612
rect 19947 11563 19989 11572
rect 20044 11537 20084 11622
rect 20043 11528 20085 11537
rect 20043 11488 20044 11528
rect 20084 11488 20085 11528
rect 20043 11479 20085 11488
rect 20048 11360 20416 11369
rect 20620 11360 20660 11740
rect 20088 11320 20130 11360
rect 20170 11320 20212 11360
rect 20252 11320 20294 11360
rect 20334 11320 20376 11360
rect 20048 11311 20416 11320
rect 20524 11320 20660 11360
rect 20043 11192 20085 11201
rect 20043 11152 20044 11192
rect 20084 11152 20085 11192
rect 20043 11143 20085 11152
rect 20235 11192 20277 11201
rect 20235 11152 20236 11192
rect 20276 11152 20277 11192
rect 20235 11143 20277 11152
rect 19659 11068 19660 11108
rect 19700 11068 19701 11108
rect 19659 11059 19701 11068
rect 19756 11068 19892 11108
rect 19563 11024 19605 11033
rect 19563 10984 19564 11024
rect 19604 10984 19605 11024
rect 19563 10975 19605 10984
rect 19564 10890 19604 10975
rect 19659 10940 19701 10949
rect 19659 10900 19660 10940
rect 19700 10900 19701 10940
rect 19659 10891 19701 10900
rect 19660 10806 19700 10891
rect 19756 10856 19796 11068
rect 19948 11024 19988 11033
rect 19756 10807 19796 10816
rect 19852 10940 19892 10949
rect 19372 10772 19412 10781
rect 19412 10732 19604 10772
rect 19372 10723 19412 10732
rect 19371 10436 19413 10445
rect 19371 10396 19372 10436
rect 19412 10396 19413 10436
rect 19371 10387 19413 10396
rect 19372 10184 19412 10387
rect 19467 10268 19509 10277
rect 19467 10228 19468 10268
rect 19508 10228 19509 10268
rect 19467 10219 19509 10228
rect 19372 10135 19412 10144
rect 19468 10184 19508 10219
rect 19468 10133 19508 10144
rect 19564 9638 19604 10732
rect 19755 10520 19797 10529
rect 19755 10480 19756 10520
rect 19796 10480 19797 10520
rect 19755 10471 19797 10480
rect 19756 10184 19796 10471
rect 19564 9598 19700 9638
rect 19563 9512 19605 9521
rect 19563 9472 19564 9512
rect 19604 9472 19605 9512
rect 19563 9463 19605 9472
rect 19564 9378 19604 9463
rect 19467 9176 19509 9185
rect 19467 9136 19468 9176
rect 19508 9136 19509 9176
rect 19467 9127 19509 9136
rect 19468 8849 19508 9127
rect 19467 8840 19509 8849
rect 19660 8840 19700 9598
rect 19756 9437 19796 10144
rect 19755 9428 19797 9437
rect 19755 9388 19756 9428
rect 19796 9388 19797 9428
rect 19755 9379 19797 9388
rect 19756 9260 19796 9269
rect 19852 9260 19892 10900
rect 19948 9689 19988 10984
rect 20044 10529 20084 11143
rect 20236 11024 20276 11143
rect 20236 10975 20276 10984
rect 20139 10772 20181 10781
rect 20139 10732 20140 10772
rect 20180 10732 20181 10772
rect 20139 10723 20181 10732
rect 20140 10638 20180 10723
rect 20043 10520 20085 10529
rect 20043 10480 20044 10520
rect 20084 10480 20085 10520
rect 20043 10471 20085 10480
rect 20044 10352 20084 10361
rect 20044 10109 20084 10312
rect 20235 10268 20277 10277
rect 20235 10228 20236 10268
rect 20276 10228 20277 10268
rect 20235 10219 20277 10228
rect 20236 10134 20276 10219
rect 20043 10100 20085 10109
rect 20043 10060 20044 10100
rect 20084 10060 20085 10100
rect 20043 10051 20085 10060
rect 20048 9848 20416 9857
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20048 9799 20416 9808
rect 19947 9680 19989 9689
rect 19947 9640 19948 9680
rect 19988 9640 19989 9680
rect 19947 9631 19989 9640
rect 20236 9521 20276 9606
rect 19947 9512 19989 9521
rect 19947 9472 19948 9512
rect 19988 9472 19989 9512
rect 19947 9463 19989 9472
rect 20044 9512 20084 9521
rect 19948 9378 19988 9463
rect 20044 9260 20084 9472
rect 20235 9512 20277 9521
rect 20235 9472 20236 9512
rect 20276 9472 20277 9512
rect 20235 9463 20277 9472
rect 20140 9260 20180 9297
rect 19852 9220 19988 9260
rect 20044 9220 20180 9260
rect 19756 9017 19796 9220
rect 19755 9008 19797 9017
rect 19755 8968 19756 9008
rect 19796 8968 19797 9008
rect 19755 8959 19797 8968
rect 19467 8800 19468 8840
rect 19508 8800 19509 8840
rect 19467 8791 19509 8800
rect 19564 8800 19700 8840
rect 19755 8840 19797 8849
rect 19755 8800 19756 8840
rect 19796 8800 19797 8840
rect 19372 8672 19412 8681
rect 19276 8632 19372 8672
rect 19180 8623 19220 8632
rect 19372 8623 19412 8632
rect 19467 8672 19509 8681
rect 19467 8632 19468 8672
rect 19508 8632 19509 8672
rect 19467 8623 19509 8632
rect 19468 8538 19508 8623
rect 19276 8504 19316 8513
rect 19276 8345 19316 8464
rect 19371 8504 19413 8513
rect 19371 8464 19372 8504
rect 19412 8464 19413 8504
rect 19371 8455 19413 8464
rect 19275 8336 19317 8345
rect 19275 8296 19276 8336
rect 19316 8296 19317 8336
rect 19275 8287 19317 8296
rect 18891 8168 18933 8177
rect 18891 8128 18892 8168
rect 18932 8128 18933 8168
rect 18891 8119 18933 8128
rect 19275 8168 19317 8177
rect 19275 8128 19276 8168
rect 19316 8128 19317 8168
rect 19275 8119 19317 8128
rect 18795 8084 18837 8093
rect 18795 8044 18796 8084
rect 18836 8044 18837 8084
rect 18795 8035 18837 8044
rect 18808 7580 19176 7589
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 18808 7531 19176 7540
rect 18891 7328 18933 7337
rect 18891 7288 18892 7328
rect 18932 7288 18933 7328
rect 18891 7279 18933 7288
rect 18892 7160 18932 7279
rect 18987 7244 19029 7253
rect 18987 7204 18988 7244
rect 19028 7204 19029 7244
rect 18987 7195 19029 7204
rect 18892 7111 18932 7120
rect 18988 7160 19028 7195
rect 18988 7109 19028 7120
rect 19083 7160 19125 7169
rect 19083 7120 19084 7160
rect 19124 7120 19125 7160
rect 19083 7111 19125 7120
rect 19276 7160 19316 8119
rect 19084 6245 19124 7111
rect 19276 6572 19316 7120
rect 19188 6532 19316 6572
rect 19188 6488 19228 6532
rect 19188 6329 19228 6448
rect 19179 6320 19228 6329
rect 19179 6280 19180 6320
rect 19220 6280 19316 6320
rect 19179 6271 19228 6280
rect 19083 6236 19125 6245
rect 19083 6196 19084 6236
rect 19124 6196 19125 6236
rect 19083 6187 19125 6196
rect 19188 6164 19228 6271
rect 18808 6068 19176 6077
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 18808 6019 19176 6028
rect 18315 4808 18357 4817
rect 18315 4768 18316 4808
rect 18356 4768 18357 4808
rect 18315 4759 18357 4768
rect 18699 4808 18741 4817
rect 18699 4768 18700 4808
rect 18740 4768 18741 4808
rect 18699 4759 18741 4768
rect 18316 4674 18356 4759
rect 18699 4640 18741 4649
rect 18604 4600 18700 4640
rect 18740 4600 18741 4640
rect 18604 4472 18644 4600
rect 18699 4591 18741 4600
rect 18808 4556 19176 4565
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 18808 4507 19176 4516
rect 18316 4432 18644 4472
rect 19276 4472 19316 6280
rect 19372 5237 19412 8455
rect 19564 8168 19604 8800
rect 19755 8791 19797 8800
rect 19659 8672 19701 8681
rect 19659 8632 19660 8672
rect 19700 8632 19701 8672
rect 19659 8623 19701 8632
rect 19756 8651 19796 8791
rect 19851 8756 19893 8765
rect 19851 8716 19852 8756
rect 19892 8716 19893 8756
rect 19851 8707 19893 8716
rect 19660 8538 19700 8623
rect 19852 8672 19892 8707
rect 19852 8621 19892 8632
rect 19948 8672 19988 9220
rect 20137 9185 20180 9220
rect 20235 9260 20277 9269
rect 20235 9220 20236 9260
rect 20276 9220 20277 9260
rect 20235 9211 20277 9220
rect 20137 9176 20181 9185
rect 20137 9136 20140 9176
rect 20180 9136 20181 9176
rect 20139 9127 20181 9136
rect 20236 9126 20276 9211
rect 20126 9008 20168 9017
rect 20126 8968 20127 9008
rect 20167 8968 20168 9008
rect 20126 8959 20168 8968
rect 19948 8623 19988 8632
rect 20127 8661 20167 8959
rect 19756 8602 19796 8611
rect 20127 8513 20167 8621
rect 20236 8513 20276 8598
rect 20126 8504 20168 8513
rect 20126 8464 20127 8504
rect 20167 8464 20168 8504
rect 20126 8455 20168 8464
rect 20235 8504 20277 8513
rect 20235 8464 20236 8504
rect 20276 8464 20277 8504
rect 20235 8455 20277 8464
rect 20048 8336 20416 8345
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20048 8287 20416 8296
rect 19756 8212 19988 8252
rect 19756 8168 19796 8212
rect 19564 8128 19796 8168
rect 19851 8084 19893 8093
rect 19851 8044 19852 8084
rect 19892 8044 19893 8084
rect 19851 8035 19893 8044
rect 19467 8000 19509 8009
rect 19467 7960 19468 8000
rect 19508 7960 19509 8000
rect 19467 7951 19509 7960
rect 19852 8000 19892 8035
rect 19468 7866 19508 7951
rect 19852 7949 19892 7960
rect 19948 8000 19988 8212
rect 20139 8168 20181 8177
rect 20139 8128 20140 8168
rect 20180 8128 20181 8168
rect 20139 8119 20181 8128
rect 20140 8034 20180 8119
rect 19948 7951 19988 7960
rect 19660 7748 19700 7757
rect 19660 7589 19700 7708
rect 19659 7580 19701 7589
rect 19659 7540 19660 7580
rect 19700 7540 19701 7580
rect 19659 7531 19701 7540
rect 19467 7496 19509 7505
rect 19467 7456 19468 7496
rect 19508 7456 19509 7496
rect 19467 7447 19509 7456
rect 19468 6917 19508 7447
rect 19659 7412 19701 7421
rect 20139 7412 20181 7421
rect 19659 7372 19660 7412
rect 19700 7372 19796 7412
rect 19659 7363 19701 7372
rect 19756 7328 19796 7372
rect 20139 7372 20140 7412
rect 20180 7372 20181 7412
rect 20139 7363 20181 7372
rect 19756 7279 19796 7288
rect 20140 7278 20180 7363
rect 19660 7244 19700 7253
rect 19564 7160 19604 7171
rect 19564 7085 19604 7120
rect 19563 7076 19605 7085
rect 19563 7036 19564 7076
rect 19604 7036 19605 7076
rect 19563 7027 19605 7036
rect 19660 6917 19700 7204
rect 19852 7244 19892 7253
rect 19467 6908 19509 6917
rect 19467 6868 19468 6908
rect 19508 6868 19509 6908
rect 19467 6859 19509 6868
rect 19659 6908 19701 6917
rect 19659 6868 19660 6908
rect 19700 6868 19701 6908
rect 19659 6859 19701 6868
rect 19467 6572 19509 6581
rect 19467 6532 19468 6572
rect 19508 6532 19509 6572
rect 19467 6523 19509 6532
rect 19468 6488 19508 6523
rect 19564 6497 19604 6582
rect 19468 6437 19508 6448
rect 19563 6488 19605 6497
rect 19563 6448 19564 6488
rect 19604 6448 19605 6488
rect 19852 6477 19892 7204
rect 19947 7160 19989 7169
rect 19947 7120 19948 7160
rect 19988 7120 19989 7160
rect 19947 7111 19989 7120
rect 20235 7160 20277 7169
rect 20235 7120 20236 7160
rect 20276 7120 20277 7160
rect 20235 7111 20277 7120
rect 19948 7026 19988 7111
rect 20236 7026 20276 7111
rect 20048 6824 20416 6833
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20048 6775 20416 6784
rect 20235 6656 20277 6665
rect 20235 6616 20236 6656
rect 20276 6616 20277 6656
rect 20235 6607 20277 6616
rect 20044 6488 20084 6497
rect 19563 6439 19605 6448
rect 19660 6437 19892 6477
rect 19948 6448 20044 6488
rect 19371 5228 19413 5237
rect 19371 5188 19372 5228
rect 19412 5188 19413 5228
rect 19371 5179 19413 5188
rect 19371 4472 19413 4481
rect 19276 4432 19372 4472
rect 19412 4432 19413 4472
rect 18316 4136 18356 4432
rect 19371 4423 19413 4432
rect 18699 4388 18741 4397
rect 18699 4348 18700 4388
rect 18740 4348 18741 4388
rect 18699 4339 18741 4348
rect 18411 4304 18453 4313
rect 18411 4264 18412 4304
rect 18452 4264 18453 4304
rect 18411 4255 18453 4264
rect 18316 4087 18356 4096
rect 18220 4003 18260 4012
rect 18315 3884 18357 3893
rect 18315 3844 18316 3884
rect 18356 3844 18357 3884
rect 18315 3835 18357 3844
rect 18027 3800 18069 3809
rect 18027 3760 18028 3800
rect 18068 3760 18069 3800
rect 18027 3751 18069 3760
rect 18028 3305 18068 3751
rect 18123 3716 18165 3725
rect 18123 3676 18124 3716
rect 18164 3676 18165 3716
rect 18123 3667 18165 3676
rect 18027 3296 18069 3305
rect 18027 3256 18028 3296
rect 18068 3256 18069 3296
rect 18027 3247 18069 3256
rect 17931 2960 17973 2969
rect 17931 2920 17932 2960
rect 17972 2920 17973 2960
rect 17931 2911 17973 2920
rect 18124 2717 18164 3667
rect 18219 3464 18261 3473
rect 18219 3424 18220 3464
rect 18260 3424 18261 3464
rect 18219 3415 18261 3424
rect 18316 3464 18356 3835
rect 18316 3415 18356 3424
rect 18220 3330 18260 3415
rect 18123 2708 18165 2717
rect 18123 2668 18124 2708
rect 18164 2668 18165 2708
rect 18123 2659 18165 2668
rect 18028 2624 18068 2633
rect 17740 2584 18028 2624
rect 17548 1868 17588 2500
rect 17163 1448 17205 1457
rect 17163 1408 17164 1448
rect 17204 1408 17205 1448
rect 17163 1399 17205 1408
rect 17068 1196 17108 1205
rect 17068 1037 17108 1156
rect 17067 1028 17109 1037
rect 17067 988 17068 1028
rect 17108 988 17109 1028
rect 17067 979 17109 988
rect 16972 820 17204 860
rect 16875 692 16917 701
rect 16875 652 16876 692
rect 16916 652 16917 692
rect 16875 643 16917 652
rect 16780 484 17012 524
rect 16587 188 16629 197
rect 16587 148 16588 188
rect 16628 148 16629 188
rect 16587 139 16629 148
rect 16588 80 16628 139
rect 16779 104 16821 113
rect 16779 80 16780 104
rect 6068 64 6088 80
rect 6008 0 6088 64
rect 6200 0 6280 80
rect 6392 0 6472 80
rect 6584 0 6664 80
rect 6776 0 6856 80
rect 6968 0 7048 80
rect 7160 0 7240 80
rect 7352 0 7432 80
rect 7544 0 7624 80
rect 7736 0 7816 80
rect 7928 0 8008 80
rect 8120 0 8200 80
rect 8312 0 8392 80
rect 8504 0 8584 80
rect 8696 0 8776 80
rect 8888 0 8968 80
rect 9080 0 9160 80
rect 9272 0 9352 80
rect 9464 0 9544 80
rect 9656 0 9736 80
rect 9848 0 9928 80
rect 10040 0 10120 80
rect 10232 0 10312 80
rect 10424 0 10504 80
rect 10616 0 10696 80
rect 10808 0 10888 80
rect 11000 0 11080 80
rect 11192 0 11272 80
rect 11384 0 11464 80
rect 11576 0 11656 80
rect 11768 0 11848 80
rect 11960 0 12040 80
rect 12152 0 12232 80
rect 12344 0 12424 80
rect 12536 0 12616 80
rect 12728 0 12808 80
rect 12920 0 13000 80
rect 13112 0 13192 80
rect 13304 0 13384 80
rect 13496 0 13576 80
rect 13688 0 13768 80
rect 13880 0 13960 80
rect 14072 0 14152 80
rect 14264 0 14344 80
rect 14456 0 14536 80
rect 14648 0 14728 80
rect 14840 0 14920 80
rect 15032 0 15112 80
rect 15224 0 15304 80
rect 15416 0 15496 80
rect 15608 0 15688 80
rect 15800 0 15880 80
rect 15992 0 16072 80
rect 16184 0 16264 80
rect 16376 0 16456 80
rect 16568 0 16648 80
rect 16760 64 16780 80
rect 16820 80 16821 104
rect 16972 80 17012 484
rect 17164 80 17204 820
rect 17260 776 17300 1828
rect 17548 1819 17588 1828
rect 17355 1700 17397 1709
rect 17740 1700 17780 2584
rect 18028 2575 18068 2584
rect 18124 2624 18164 2659
rect 18124 2574 18164 2584
rect 18412 2540 18452 4255
rect 18507 4136 18549 4145
rect 18507 4096 18508 4136
rect 18548 4096 18549 4136
rect 18507 4087 18549 4096
rect 18508 4002 18548 4087
rect 18700 3212 18740 4339
rect 19179 4136 19221 4145
rect 19179 4096 19180 4136
rect 19220 4096 19221 4136
rect 19179 4087 19221 4096
rect 18795 3464 18837 3473
rect 18795 3424 18796 3464
rect 18836 3424 18837 3464
rect 18795 3415 18837 3424
rect 18796 3330 18836 3415
rect 19180 3296 19220 4087
rect 19371 3968 19413 3977
rect 19371 3928 19372 3968
rect 19412 3928 19413 3968
rect 19371 3919 19413 3928
rect 19372 3716 19412 3919
rect 19372 3676 19604 3716
rect 19372 3464 19412 3676
rect 19324 3454 19412 3464
rect 19364 3424 19412 3454
rect 19468 3548 19508 3557
rect 19324 3405 19364 3414
rect 19180 3256 19316 3296
rect 18508 3172 18740 3212
rect 18508 2708 18548 3172
rect 18808 3044 19176 3053
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 18808 2995 19176 3004
rect 18508 2659 18548 2668
rect 19084 2633 19124 2718
rect 18604 2624 18644 2633
rect 18604 2540 18644 2584
rect 19083 2624 19125 2633
rect 19083 2584 19084 2624
rect 19124 2584 19125 2624
rect 19083 2575 19125 2584
rect 18412 2500 18644 2540
rect 17931 1952 17973 1961
rect 17931 1912 17932 1952
rect 17972 1912 17973 1952
rect 17931 1903 17973 1912
rect 19180 1952 19220 1961
rect 19276 1952 19316 3256
rect 19220 1912 19316 1952
rect 19180 1903 19220 1912
rect 17932 1818 17972 1903
rect 17355 1660 17356 1700
rect 17396 1660 17397 1700
rect 17355 1651 17397 1660
rect 17644 1660 17780 1700
rect 17356 1566 17396 1651
rect 17451 1616 17493 1625
rect 17451 1576 17452 1616
rect 17492 1576 17493 1616
rect 17451 1567 17493 1576
rect 17452 1280 17492 1567
rect 17452 1231 17492 1240
rect 17547 1280 17589 1289
rect 17547 1240 17548 1280
rect 17588 1240 17589 1280
rect 17547 1231 17589 1240
rect 17644 1280 17684 1660
rect 18808 1532 19176 1541
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 18808 1483 19176 1492
rect 17644 1231 17684 1240
rect 17739 1280 17781 1289
rect 17739 1240 17740 1280
rect 17780 1240 17781 1280
rect 17739 1231 17781 1240
rect 18315 1280 18357 1289
rect 18315 1240 18316 1280
rect 18356 1240 18357 1280
rect 18315 1231 18357 1240
rect 18987 1280 19029 1289
rect 18987 1240 18988 1280
rect 19028 1240 19029 1280
rect 18987 1231 19029 1240
rect 17260 736 17396 776
rect 17356 80 17396 736
rect 17548 80 17588 1231
rect 17740 80 17780 1231
rect 17836 1112 17876 1123
rect 17836 1037 17876 1072
rect 17835 1028 17877 1037
rect 17835 988 17836 1028
rect 17876 988 17877 1028
rect 17835 979 17877 988
rect 17931 440 17973 449
rect 17931 400 17932 440
rect 17972 400 17973 440
rect 17931 391 17973 400
rect 17932 80 17972 391
rect 18123 272 18165 281
rect 18123 232 18124 272
rect 18164 232 18165 272
rect 18123 223 18165 232
rect 18124 80 18164 223
rect 18316 80 18356 1231
rect 18507 1196 18549 1205
rect 18507 1156 18508 1196
rect 18548 1156 18549 1196
rect 18507 1147 18549 1156
rect 18508 80 18548 1147
rect 18699 860 18741 869
rect 18699 820 18700 860
rect 18740 820 18741 860
rect 18699 811 18741 820
rect 18891 860 18933 869
rect 18891 820 18892 860
rect 18932 820 18933 860
rect 18988 860 19028 1231
rect 19083 1112 19125 1121
rect 19083 1072 19084 1112
rect 19124 1072 19125 1112
rect 19083 1063 19125 1072
rect 19084 978 19124 1063
rect 19276 1037 19316 1912
rect 19372 1700 19412 1709
rect 19372 1112 19412 1660
rect 19468 1112 19508 3508
rect 19564 2638 19604 3676
rect 19660 3641 19700 6437
rect 19851 6320 19893 6329
rect 19851 6280 19852 6320
rect 19892 6280 19893 6320
rect 19851 6271 19893 6280
rect 19852 6186 19892 6271
rect 19948 5732 19988 6448
rect 20044 6439 20084 6448
rect 20236 6488 20276 6607
rect 20236 6439 20276 6448
rect 20043 6236 20085 6245
rect 20043 6196 20044 6236
rect 20084 6196 20085 6236
rect 20043 6187 20085 6196
rect 20044 6102 20084 6187
rect 20139 5900 20181 5909
rect 20139 5860 20140 5900
rect 20180 5860 20181 5900
rect 20139 5851 20181 5860
rect 20140 5766 20180 5851
rect 19852 5692 19988 5732
rect 19755 5648 19797 5657
rect 19755 5608 19756 5648
rect 19796 5608 19797 5648
rect 19755 5599 19797 5608
rect 19756 4976 19796 5599
rect 19756 4145 19796 4936
rect 19755 4136 19797 4145
rect 19755 4096 19756 4136
rect 19796 4096 19797 4136
rect 19755 4087 19797 4096
rect 19659 3632 19701 3641
rect 19659 3592 19660 3632
rect 19700 3592 19701 3632
rect 19852 3632 19892 5692
rect 20236 5648 20276 5659
rect 20236 5573 20276 5608
rect 19947 5564 19989 5573
rect 19947 5524 19948 5564
rect 19988 5524 19989 5564
rect 19947 5515 19989 5524
rect 20235 5564 20277 5573
rect 20235 5524 20236 5564
rect 20276 5524 20277 5564
rect 20235 5515 20277 5524
rect 19948 5430 19988 5515
rect 20048 5312 20416 5321
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20048 5263 20416 5272
rect 20427 4808 20469 4817
rect 20427 4768 20428 4808
rect 20468 4768 20469 4808
rect 20427 4759 20469 4768
rect 19948 4724 19988 4733
rect 19948 4481 19988 4684
rect 19947 4472 19989 4481
rect 19947 4432 19948 4472
rect 19988 4432 19989 4472
rect 19947 4423 19989 4432
rect 20428 4061 20468 4759
rect 20427 4052 20469 4061
rect 20427 4012 20428 4052
rect 20468 4012 20469 4052
rect 20427 4003 20469 4012
rect 19947 3968 19989 3977
rect 19947 3928 19948 3968
rect 19988 3928 19989 3968
rect 19947 3919 19989 3928
rect 19948 3834 19988 3919
rect 20048 3800 20416 3809
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20048 3751 20416 3760
rect 19948 3632 19988 3641
rect 19852 3592 19948 3632
rect 19659 3583 19701 3592
rect 19948 3583 19988 3592
rect 20043 3632 20085 3641
rect 20043 3592 20044 3632
rect 20084 3592 20085 3632
rect 20043 3583 20085 3592
rect 19755 3548 19797 3557
rect 19755 3508 19756 3548
rect 19796 3508 19797 3548
rect 19755 3499 19797 3508
rect 19660 3464 19700 3473
rect 19660 3305 19700 3424
rect 19756 3464 19796 3499
rect 19756 3413 19796 3424
rect 19852 3464 19892 3475
rect 20044 3464 20084 3583
rect 19852 3389 19892 3424
rect 19948 3424 20084 3464
rect 19851 3380 19893 3389
rect 19851 3340 19852 3380
rect 19892 3340 19893 3380
rect 19851 3331 19893 3340
rect 19659 3296 19701 3305
rect 19659 3256 19660 3296
rect 19700 3256 19701 3296
rect 19659 3247 19701 3256
rect 19659 2960 19701 2969
rect 19659 2920 19660 2960
rect 19700 2920 19701 2960
rect 19659 2911 19701 2920
rect 19564 2589 19604 2598
rect 19660 2540 19700 2911
rect 19948 2624 19988 3424
rect 20139 3380 20181 3389
rect 20139 3340 20140 3380
rect 20180 3340 20181 3380
rect 20139 3331 20181 3340
rect 20140 3246 20180 3331
rect 20235 2876 20277 2885
rect 20235 2836 20236 2876
rect 20276 2836 20277 2876
rect 20235 2827 20277 2836
rect 20043 2792 20085 2801
rect 20043 2752 20044 2792
rect 20084 2752 20085 2792
rect 20043 2743 20085 2752
rect 19948 2575 19988 2584
rect 20044 2624 20084 2743
rect 20044 2575 20084 2584
rect 20139 2624 20181 2633
rect 20139 2584 20140 2624
rect 20180 2584 20181 2624
rect 20139 2575 20181 2584
rect 20236 2624 20276 2827
rect 20236 2575 20276 2584
rect 19557 2500 19700 2540
rect 19557 2456 19597 2500
rect 20140 2490 20180 2575
rect 19756 2456 19796 2465
rect 19557 2416 19604 2456
rect 19564 1952 19604 2416
rect 19659 2120 19701 2129
rect 19659 2080 19660 2120
rect 19700 2080 19701 2120
rect 19756 2120 19796 2416
rect 20524 2381 20564 11320
rect 20619 11108 20661 11117
rect 20619 11068 20620 11108
rect 20660 11068 20661 11108
rect 20619 11059 20661 11068
rect 20620 9269 20660 11059
rect 20716 9521 20756 11899
rect 20811 9596 20853 9605
rect 20811 9556 20812 9596
rect 20852 9556 20853 9596
rect 20811 9547 20853 9556
rect 20715 9512 20757 9521
rect 20715 9472 20716 9512
rect 20756 9472 20757 9512
rect 20715 9463 20757 9472
rect 20619 9260 20661 9269
rect 20619 9220 20620 9260
rect 20660 9220 20661 9260
rect 20619 9211 20661 9220
rect 20715 8504 20757 8513
rect 20715 8464 20716 8504
rect 20756 8464 20757 8504
rect 20715 8455 20757 8464
rect 20619 5564 20661 5573
rect 20619 5524 20620 5564
rect 20660 5524 20661 5564
rect 20619 5515 20661 5524
rect 20523 2372 20565 2381
rect 20523 2332 20524 2372
rect 20564 2332 20565 2372
rect 20523 2323 20565 2332
rect 20048 2288 20416 2297
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20048 2239 20416 2248
rect 20043 2120 20085 2129
rect 19756 2080 19892 2120
rect 19659 2071 19701 2080
rect 19660 1986 19700 2071
rect 19564 1903 19604 1912
rect 19755 1952 19797 1961
rect 19755 1912 19756 1952
rect 19796 1912 19797 1952
rect 19755 1903 19797 1912
rect 19756 1818 19796 1903
rect 19660 1112 19700 1121
rect 19468 1072 19660 1112
rect 19372 1063 19412 1072
rect 19660 1063 19700 1072
rect 19756 1112 19796 1121
rect 19852 1112 19892 2080
rect 20043 2080 20044 2120
rect 20084 2080 20085 2120
rect 20043 2071 20085 2080
rect 19947 1952 19989 1961
rect 19947 1912 19948 1952
rect 19988 1912 19989 1952
rect 19947 1903 19989 1912
rect 20044 1952 20084 2071
rect 20044 1903 20084 1912
rect 20236 1952 20276 1961
rect 20620 1952 20660 5515
rect 20716 4649 20756 8455
rect 20812 7169 20852 9547
rect 20908 7757 20948 12076
rect 21003 11780 21045 11789
rect 21003 11740 21004 11780
rect 21044 11740 21045 11780
rect 21003 11731 21045 11740
rect 21004 8345 21044 11731
rect 21099 10856 21141 10865
rect 21099 10816 21100 10856
rect 21140 10816 21141 10856
rect 21099 10807 21141 10816
rect 21003 8336 21045 8345
rect 21003 8296 21004 8336
rect 21044 8296 21045 8336
rect 21003 8287 21045 8296
rect 20907 7748 20949 7757
rect 20907 7708 20908 7748
rect 20948 7708 20949 7748
rect 20907 7699 20949 7708
rect 20811 7160 20853 7169
rect 20811 7120 20812 7160
rect 20852 7120 20853 7160
rect 20811 7111 20853 7120
rect 20812 5825 20852 7111
rect 20907 6908 20949 6917
rect 20907 6868 20908 6908
rect 20948 6868 20949 6908
rect 20907 6859 20949 6868
rect 20811 5816 20853 5825
rect 20811 5776 20812 5816
rect 20852 5776 20853 5816
rect 20811 5767 20853 5776
rect 20811 5228 20853 5237
rect 20811 5188 20812 5228
rect 20852 5188 20853 5228
rect 20811 5179 20853 5188
rect 20715 4640 20757 4649
rect 20715 4600 20716 4640
rect 20756 4600 20757 4640
rect 20715 4591 20757 4600
rect 20812 4472 20852 5179
rect 20716 4432 20852 4472
rect 20716 2885 20756 4432
rect 20811 4304 20853 4313
rect 20811 4264 20812 4304
rect 20852 4264 20853 4304
rect 20811 4255 20853 4264
rect 20812 3893 20852 4255
rect 20811 3884 20853 3893
rect 20811 3844 20812 3884
rect 20852 3844 20853 3884
rect 20811 3835 20853 3844
rect 20715 2876 20757 2885
rect 20715 2836 20716 2876
rect 20756 2836 20757 2876
rect 20715 2827 20757 2836
rect 20908 2540 20948 6859
rect 21003 5816 21045 5825
rect 21003 5776 21004 5816
rect 21044 5776 21045 5816
rect 21003 5767 21045 5776
rect 21004 3473 21044 5767
rect 21003 3464 21045 3473
rect 21003 3424 21004 3464
rect 21044 3424 21045 3464
rect 21003 3415 21045 3424
rect 21100 2717 21140 10807
rect 21196 4901 21236 14335
rect 21195 4892 21237 4901
rect 21195 4852 21196 4892
rect 21236 4852 21237 4892
rect 21195 4843 21237 4852
rect 21387 4136 21429 4145
rect 21387 4096 21388 4136
rect 21428 4096 21429 4136
rect 21387 4087 21429 4096
rect 21388 3809 21428 4087
rect 21387 3800 21429 3809
rect 21387 3760 21388 3800
rect 21428 3760 21429 3800
rect 21387 3751 21429 3760
rect 21099 2708 21141 2717
rect 21099 2668 21100 2708
rect 21140 2668 21141 2708
rect 21099 2659 21141 2668
rect 20276 1912 20660 1952
rect 20716 2500 20948 2540
rect 20236 1903 20276 1912
rect 19948 1818 19988 1903
rect 20716 1868 20756 2500
rect 20332 1828 20756 1868
rect 20043 1784 20085 1793
rect 20043 1744 20044 1784
rect 20084 1744 20085 1784
rect 20043 1735 20085 1744
rect 20236 1784 20276 1793
rect 20332 1784 20372 1828
rect 20276 1744 20372 1784
rect 20236 1735 20276 1744
rect 20044 1364 20084 1735
rect 20044 1315 20084 1324
rect 19796 1072 19892 1112
rect 19756 1063 19796 1072
rect 19275 1028 19317 1037
rect 19275 988 19276 1028
rect 19316 988 19317 1028
rect 19275 979 19317 988
rect 18988 820 19124 860
rect 18891 811 18933 820
rect 18700 80 18740 811
rect 18892 80 18932 811
rect 19084 80 19124 820
rect 20048 776 20416 785
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20048 727 20416 736
rect 19275 692 19317 701
rect 19275 652 19276 692
rect 19316 652 19317 692
rect 19275 643 19317 652
rect 19276 80 19316 643
rect 19467 524 19509 533
rect 19467 484 19468 524
rect 19508 484 19509 524
rect 19467 475 19509 484
rect 19468 80 19508 475
rect 16820 64 16840 80
rect 16760 0 16840 64
rect 16952 0 17032 80
rect 17144 0 17224 80
rect 17336 0 17416 80
rect 17528 0 17608 80
rect 17720 0 17800 80
rect 17912 0 17992 80
rect 18104 0 18184 80
rect 18296 0 18376 80
rect 18488 0 18568 80
rect 18680 0 18760 80
rect 18872 0 18952 80
rect 19064 0 19144 80
rect 19256 0 19336 80
rect 19448 0 19528 80
<< via2 >>
rect 76 42736 116 42776
rect 1612 42568 1652 42608
rect 748 42400 788 42440
rect 268 42064 308 42104
rect 172 39628 212 39668
rect 364 40384 404 40424
rect 268 33580 308 33620
rect 364 31900 404 31940
rect 1420 41728 1460 41768
rect 1324 41140 1364 41180
rect 1516 41560 1556 41600
rect 1516 41140 1556 41180
rect 1420 40468 1460 40508
rect 1228 39460 1268 39500
rect 1900 42400 1940 42440
rect 1804 42232 1844 42272
rect 1612 39376 1652 39416
rect 1708 39208 1748 39248
rect 1900 40300 1940 40340
rect 2188 42904 2228 42944
rect 2188 41980 2228 42020
rect 2092 40552 2132 40592
rect 2092 40300 2132 40340
rect 1996 40132 2036 40172
rect 1516 38872 1556 38912
rect 1708 38872 1748 38912
rect 1708 38620 1748 38660
rect 1612 38452 1652 38492
rect 2092 39712 2132 39752
rect 2092 39460 2132 39500
rect 1996 38956 2036 38996
rect 1804 38536 1844 38576
rect 1804 38368 1844 38408
rect 1228 37780 1268 37820
rect 1228 37612 1268 37652
rect 1516 38116 1556 38156
rect 1324 37444 1364 37484
rect 1324 37192 1364 37232
rect 1420 37024 1460 37064
rect 1900 37696 1940 37736
rect 1708 37192 1748 37232
rect 1900 37024 1940 37064
rect 1612 36520 1652 36560
rect 1900 36520 1940 36560
rect 940 35932 980 35972
rect 1708 36100 1748 36140
rect 844 30976 884 31016
rect 748 29884 788 29924
rect 460 29548 500 29588
rect 172 28960 212 29000
rect 76 28792 116 28832
rect 652 26692 692 26732
rect 1324 35596 1364 35636
rect 1324 34756 1364 34796
rect 1036 34420 1076 34460
rect 940 29044 980 29084
rect 1132 33580 1172 33620
rect 1228 33160 1268 33200
rect 1420 34420 1460 34460
rect 1612 34588 1652 34628
rect 1612 34336 1652 34376
rect 1516 34252 1556 34292
rect 1420 33832 1460 33872
rect 2284 40384 2324 40424
rect 2476 42484 2516 42524
rect 2380 38956 2420 38996
rect 2284 38620 2324 38660
rect 2188 38116 2228 38156
rect 2380 38116 2420 38156
rect 2092 37528 2132 37568
rect 2092 36604 2132 36644
rect 1996 36100 2036 36140
rect 1900 35512 1940 35552
rect 1804 35260 1844 35300
rect 1804 34840 1844 34880
rect 1804 34084 1844 34124
rect 2764 42484 2804 42524
rect 2668 39964 2708 40004
rect 2668 39628 2708 39668
rect 2668 39376 2708 39416
rect 2764 39124 2804 39164
rect 2572 38284 2612 38324
rect 2572 38116 2612 38156
rect 2572 37276 2612 37316
rect 2476 36604 2516 36644
rect 2380 36100 2420 36140
rect 2572 35596 2612 35636
rect 2380 35260 2420 35300
rect 2188 35176 2228 35216
rect 3340 41224 3380 41264
rect 3148 40972 3188 41012
rect 3148 40720 3188 40760
rect 2956 39124 2996 39164
rect 2956 38704 2996 38744
rect 2956 38536 2996 38576
rect 2764 38116 2804 38156
rect 2956 37864 2996 37904
rect 2764 37780 2804 37820
rect 2668 35008 2708 35048
rect 2188 34672 2228 34712
rect 2380 34341 2420 34376
rect 2380 34336 2420 34341
rect 2188 34252 2228 34292
rect 2284 34084 2324 34124
rect 2188 33916 2228 33956
rect 1324 32572 1364 32612
rect 1516 32068 1556 32108
rect 1420 31984 1460 32024
rect 1708 32404 1748 32444
rect 2092 32152 2132 32192
rect 1708 31984 1748 32024
rect 1228 31732 1268 31772
rect 1420 31480 1460 31520
rect 1132 31396 1172 31436
rect 1324 31144 1364 31184
rect 1324 30892 1364 30932
rect 1324 30388 1364 30428
rect 1132 30304 1172 30344
rect 1228 29884 1268 29924
rect 1228 29632 1268 29672
rect 1132 28960 1172 29000
rect 1612 31228 1652 31268
rect 1516 30388 1556 30428
rect 3148 39040 3188 39080
rect 3148 38788 3188 38828
rect 3148 38368 3188 38408
rect 3148 37948 3188 37988
rect 2860 36856 2900 36896
rect 2860 35932 2900 35972
rect 3148 37360 3188 37400
rect 3052 36520 3092 36560
rect 3148 36184 3188 36224
rect 3148 35512 3188 35552
rect 2956 35428 2996 35468
rect 3148 35176 3188 35216
rect 3340 40636 3380 40676
rect 3724 42316 3764 42356
rect 4108 42400 4148 42440
rect 3916 41140 3956 41180
rect 3688 40804 3728 40844
rect 3770 40804 3810 40844
rect 3852 40804 3892 40844
rect 3934 40804 3974 40844
rect 4016 40804 4056 40844
rect 3532 40636 3572 40676
rect 4108 40636 4148 40676
rect 3532 40468 3572 40508
rect 3436 40384 3476 40424
rect 3916 40300 3956 40340
rect 3340 38872 3380 38912
rect 3340 38704 3380 38744
rect 3916 40132 3956 40172
rect 3532 39796 3572 39836
rect 3724 39628 3764 39668
rect 4396 41728 4436 41768
rect 3688 39292 3728 39332
rect 3770 39292 3810 39332
rect 3852 39292 3892 39332
rect 3934 39292 3974 39332
rect 4016 39292 4056 39332
rect 4012 39124 4052 39164
rect 3628 39040 3668 39080
rect 3532 38956 3572 38996
rect 4300 40048 4340 40088
rect 4204 39124 4244 39164
rect 4108 39040 4148 39080
rect 4108 38872 4148 38912
rect 3820 38788 3860 38828
rect 3628 38452 3668 38492
rect 3724 38116 3764 38156
rect 3628 38032 3668 38072
rect 4012 38620 4052 38660
rect 3820 37948 3860 37988
rect 3688 37780 3728 37820
rect 3770 37780 3810 37820
rect 3852 37780 3892 37820
rect 3934 37780 3974 37820
rect 4016 37780 4056 37820
rect 3532 37108 3572 37148
rect 3532 36856 3572 36896
rect 3820 37360 3860 37400
rect 3820 37192 3860 37232
rect 4108 37444 4148 37484
rect 4492 41560 4532 41600
rect 4588 41476 4628 41516
rect 4492 40720 4532 40760
rect 5068 42568 5108 42608
rect 5452 42820 5492 42860
rect 4876 41728 4916 41768
rect 5452 41644 5492 41684
rect 4928 41560 4968 41600
rect 5010 41560 5050 41600
rect 5092 41560 5132 41600
rect 5174 41560 5214 41600
rect 5256 41560 5296 41600
rect 5356 41476 5396 41516
rect 4492 40216 4532 40256
rect 4492 39628 4532 39668
rect 4684 40216 4724 40256
rect 4684 39628 4724 39668
rect 4588 39124 4628 39164
rect 4492 38872 4532 38912
rect 4396 38620 4436 38660
rect 4396 38452 4436 38492
rect 4300 37612 4340 37652
rect 4588 37948 4628 37988
rect 4588 37696 4628 37736
rect 4492 37444 4532 37484
rect 4492 37108 4532 37148
rect 4972 40720 5012 40760
rect 5068 40552 5108 40592
rect 5356 40300 5396 40340
rect 4928 40048 4968 40088
rect 5010 40048 5050 40088
rect 5092 40048 5132 40088
rect 5174 40048 5214 40088
rect 5256 40048 5296 40088
rect 6028 41812 6068 41852
rect 5644 41728 5684 41768
rect 5932 41728 5972 41768
rect 5836 41560 5876 41600
rect 5740 41392 5780 41432
rect 5548 40804 5588 40844
rect 5068 39712 5108 39752
rect 4876 39628 4916 39668
rect 5260 39460 5300 39500
rect 5356 39124 5396 39164
rect 5644 40468 5684 40508
rect 4928 38536 4968 38576
rect 5010 38536 5050 38576
rect 5092 38536 5132 38576
rect 5174 38536 5214 38576
rect 5256 38536 5296 38576
rect 5068 38200 5108 38240
rect 4876 38032 4916 38072
rect 5740 39712 5780 39752
rect 6316 41728 6356 41768
rect 6028 41308 6068 41348
rect 6220 41392 6260 41432
rect 6700 42484 6740 42524
rect 6604 41392 6644 41432
rect 6604 41224 6644 41264
rect 6412 40384 6452 40424
rect 6220 39796 6260 39836
rect 6124 39628 6164 39668
rect 5836 39208 5876 39248
rect 5740 37948 5780 37988
rect 5260 37696 5300 37736
rect 5260 37528 5300 37568
rect 5452 37528 5492 37568
rect 3340 36520 3380 36560
rect 2764 34588 2804 34628
rect 2668 34336 2708 34376
rect 2572 33916 2612 33956
rect 2284 33832 2324 33872
rect 2860 34252 2900 34292
rect 3052 35092 3092 35132
rect 3340 34924 3380 34964
rect 3244 34588 3284 34628
rect 3688 36268 3728 36308
rect 3770 36268 3810 36308
rect 3852 36268 3892 36308
rect 3934 36268 3974 36308
rect 4016 36268 4056 36308
rect 4928 37024 4968 37064
rect 5010 37024 5050 37064
rect 5092 37024 5132 37064
rect 5174 37024 5214 37064
rect 5256 37024 5296 37064
rect 3820 36016 3860 36056
rect 4300 36520 4340 36560
rect 4204 35848 4244 35888
rect 4396 35848 4436 35888
rect 3820 35764 3860 35804
rect 4300 35596 4340 35636
rect 3628 35512 3668 35552
rect 3532 35428 3572 35468
rect 3820 35344 3860 35384
rect 3724 35092 3764 35132
rect 3827 35092 3867 35132
rect 4204 35176 4244 35216
rect 4060 35008 4100 35048
rect 3532 34924 3572 34964
rect 3916 34924 3956 34964
rect 3688 34756 3728 34796
rect 3770 34756 3810 34796
rect 3852 34756 3892 34796
rect 3934 34756 3974 34796
rect 4016 34756 4056 34796
rect 3148 34420 3188 34460
rect 3436 34336 3476 34376
rect 2956 33748 2996 33788
rect 2284 32656 2324 32696
rect 2188 31480 2228 31520
rect 3148 34000 3188 34040
rect 2860 33244 2900 33284
rect 2572 32320 2612 32360
rect 2188 31060 2228 31100
rect 2092 30808 2132 30848
rect 1804 30724 1844 30764
rect 1708 30220 1748 30260
rect 1804 30136 1844 30176
rect 1708 30052 1748 30092
rect 1612 29128 1652 29168
rect 1516 29044 1556 29084
rect 2092 29968 2132 30008
rect 1036 28204 1076 28244
rect 940 25600 980 25640
rect 844 24004 884 24044
rect 652 23920 692 23960
rect 460 23584 500 23624
rect 556 22828 596 22868
rect 172 21316 212 21356
rect 268 14092 308 14132
rect 172 12496 212 12536
rect 172 10144 212 10184
rect 460 13840 500 13880
rect 364 12580 404 12620
rect 364 10312 404 10352
rect 1036 22996 1076 23036
rect 940 18628 980 18668
rect 940 13168 980 13208
rect 748 13000 788 13040
rect 652 12748 692 12788
rect 556 11824 596 11864
rect 460 8800 500 8840
rect 556 7540 596 7580
rect 268 5776 308 5816
rect 1036 11572 1076 11612
rect 940 11152 980 11192
rect 844 9472 884 9512
rect 748 7456 788 7496
rect 1324 28120 1364 28160
rect 1324 27700 1364 27740
rect 1324 27364 1364 27404
rect 1228 26776 1268 26816
rect 1996 28960 2036 29000
rect 1708 28876 1748 28916
rect 1900 28456 1940 28496
rect 1708 28288 1748 28328
rect 1612 28120 1652 28160
rect 1420 26440 1460 26480
rect 1228 26020 1268 26060
rect 1324 25348 1364 25388
rect 1420 24592 1460 24632
rect 1804 27784 1844 27824
rect 1804 26860 1844 26900
rect 1708 25096 1748 25136
rect 1612 23836 1652 23876
rect 1708 23332 1748 23372
rect 1516 23164 1556 23204
rect 1516 22828 1556 22868
rect 1420 22660 1460 22700
rect 1324 22492 1364 22532
rect 1708 22996 1748 23036
rect 2092 28792 2132 28832
rect 2572 31816 2612 31856
rect 2572 31564 2612 31604
rect 2572 31144 2612 31184
rect 2764 32656 2804 32696
rect 3052 33244 3092 33284
rect 2956 32992 2996 33032
rect 2956 32656 2996 32696
rect 3052 32404 3092 32444
rect 3916 34336 3956 34376
rect 4396 35428 4436 35468
rect 4588 35848 4628 35888
rect 4492 35344 4532 35384
rect 5452 36604 5492 36644
rect 5260 36520 5300 36560
rect 5068 36436 5108 36476
rect 5356 36436 5396 36476
rect 4876 36100 4916 36140
rect 4780 35680 4820 35720
rect 4928 35512 4968 35552
rect 5010 35512 5050 35552
rect 5092 35512 5132 35552
rect 5174 35512 5214 35552
rect 5256 35512 5296 35552
rect 4492 35092 4532 35132
rect 4396 34924 4436 34964
rect 4204 34168 4244 34208
rect 3628 33916 3668 33956
rect 3820 33916 3860 33956
rect 4108 33832 4148 33872
rect 3532 33496 3572 33536
rect 3820 33580 3860 33620
rect 3436 33244 3476 33284
rect 3244 32992 3284 33032
rect 3436 32824 3476 32864
rect 3244 32404 3284 32444
rect 2956 32320 2996 32360
rect 3148 32320 3188 32360
rect 2764 32152 2804 32192
rect 2476 30808 2516 30848
rect 2668 30724 2708 30764
rect 2476 30556 2516 30596
rect 2572 30556 2612 30596
rect 2284 30472 2324 30512
rect 2668 30472 2708 30512
rect 2572 30388 2612 30428
rect 2380 30220 2420 30260
rect 2284 29716 2324 29756
rect 2188 26776 2228 26816
rect 2092 26356 2132 26396
rect 1996 24592 2036 24632
rect 1900 23752 1940 23792
rect 1804 22576 1844 22616
rect 1708 22240 1748 22280
rect 1420 21652 1460 21692
rect 1612 21568 1652 21608
rect 1228 21316 1268 21356
rect 1324 20728 1364 20768
rect 1516 20308 1556 20348
rect 1324 19720 1364 19760
rect 1900 20644 1940 20684
rect 1228 18460 1268 18500
rect 1228 18208 1268 18248
rect 1228 17788 1268 17828
rect 1516 18460 1556 18500
rect 1516 17704 1556 17744
rect 1324 17284 1364 17324
rect 1708 19132 1748 19172
rect 2476 29128 2516 29168
rect 2380 28456 2420 28496
rect 3688 33244 3728 33284
rect 3770 33244 3810 33284
rect 3852 33244 3892 33284
rect 3934 33244 3974 33284
rect 4016 33244 4056 33284
rect 4684 35008 4724 35048
rect 4684 34756 4724 34796
rect 4588 34336 4628 34376
rect 4492 34168 4532 34208
rect 4396 33328 4436 33368
rect 4684 34084 4724 34124
rect 4972 35176 5012 35216
rect 4876 34756 4916 34796
rect 5356 34672 5396 34712
rect 4972 34168 5012 34208
rect 4780 34000 4820 34040
rect 4928 34000 4968 34040
rect 5010 34000 5050 34040
rect 5092 34000 5132 34040
rect 5174 34000 5214 34040
rect 5256 34000 5296 34040
rect 4684 33916 4724 33956
rect 3820 33076 3860 33116
rect 4300 33076 4340 33116
rect 4108 32908 4148 32948
rect 4300 32908 4340 32948
rect 4588 32824 4628 32864
rect 4492 32740 4532 32780
rect 3628 32656 3668 32696
rect 4204 32656 4244 32696
rect 4396 32656 4436 32696
rect 3724 32320 3764 32360
rect 4012 32320 4052 32360
rect 3052 31816 3092 31856
rect 2956 31732 2996 31772
rect 2860 30724 2900 30764
rect 2860 30220 2900 30260
rect 2668 30136 2708 30176
rect 2764 30052 2804 30092
rect 2668 28960 2708 29000
rect 3148 31228 3188 31268
rect 3052 30808 3092 30848
rect 3052 30304 3092 30344
rect 3340 30724 3380 30764
rect 3340 30472 3380 30512
rect 2956 29380 2996 29420
rect 2860 29212 2900 29252
rect 2764 27868 2804 27908
rect 2476 27784 2516 27824
rect 2860 27784 2900 27824
rect 2572 27700 2612 27740
rect 2764 27616 2804 27656
rect 2668 27448 2708 27488
rect 2764 27364 2804 27404
rect 2865 27364 2900 27404
rect 2900 27364 2905 27404
rect 2860 27196 2900 27236
rect 2572 26608 2612 26648
rect 2476 26104 2516 26144
rect 2764 26104 2804 26144
rect 3244 29716 3284 29756
rect 3148 29464 3188 29504
rect 3052 28960 3092 29000
rect 3244 29296 3284 29336
rect 3148 28372 3188 28412
rect 3052 28120 3092 28160
rect 3244 27952 3284 27992
rect 3244 27784 3284 27824
rect 3148 27700 3188 27740
rect 3148 27448 3188 27488
rect 3052 27364 3092 27404
rect 3244 27196 3284 27236
rect 3244 26944 3284 26984
rect 3916 32152 3956 32192
rect 3688 31732 3728 31772
rect 3770 31732 3810 31772
rect 3852 31732 3892 31772
rect 3934 31732 3974 31772
rect 4016 31732 4056 31772
rect 3628 31480 3668 31520
rect 3820 31228 3860 31268
rect 3724 30640 3764 30680
rect 4012 31144 4052 31184
rect 3628 30472 3668 30512
rect 3820 30472 3860 30512
rect 4012 30388 4052 30428
rect 4204 31228 4244 31268
rect 4204 30892 4244 30932
rect 4300 30808 4340 30848
rect 4396 30388 4436 30428
rect 4204 30304 4244 30344
rect 3532 30220 3572 30260
rect 3688 30220 3728 30260
rect 3770 30220 3810 30260
rect 3852 30220 3892 30260
rect 3934 30220 3974 30260
rect 4016 30220 4056 30260
rect 4108 29044 4148 29084
rect 3820 28960 3860 29000
rect 3436 28708 3476 28748
rect 3688 28708 3728 28748
rect 3770 28708 3810 28748
rect 3852 28708 3892 28748
rect 3934 28708 3974 28748
rect 4016 28708 4056 28748
rect 3916 28540 3956 28580
rect 4492 30136 4532 30176
rect 4300 29884 4340 29924
rect 5644 36856 5684 36896
rect 5932 37696 5972 37736
rect 6028 37612 6068 37652
rect 5932 37276 5972 37316
rect 6028 37108 6068 37148
rect 5932 36772 5972 36812
rect 5836 36688 5876 36728
rect 6220 39208 6260 39248
rect 6316 37948 6356 37988
rect 6796 41644 6836 41684
rect 6988 40468 7028 40508
rect 7276 41476 7316 41516
rect 7276 41224 7316 41264
rect 7372 40972 7412 41012
rect 7756 41980 7796 42020
rect 7660 41392 7700 41432
rect 7564 40636 7604 40676
rect 7852 41224 7892 41264
rect 7756 40468 7796 40508
rect 6988 40300 7028 40340
rect 7276 40300 7316 40340
rect 6988 39712 7028 39752
rect 6796 39124 6836 39164
rect 6220 37696 6260 37736
rect 6220 36772 6260 36812
rect 6412 37360 6452 37400
rect 6508 37024 6548 37064
rect 6316 36604 6356 36644
rect 6508 36520 6548 36560
rect 6220 35596 6260 35636
rect 5452 34000 5492 34040
rect 6028 35260 6068 35300
rect 6124 35176 6164 35216
rect 6412 35680 6452 35720
rect 6412 35512 6452 35552
rect 6316 35344 6356 35384
rect 5260 33664 5300 33704
rect 4876 33580 4916 33620
rect 4780 33328 4820 33368
rect 4780 32740 4820 32780
rect 5356 33580 5396 33620
rect 4876 32656 4916 32696
rect 4928 32488 4968 32528
rect 5010 32488 5050 32528
rect 5092 32488 5132 32528
rect 5174 32488 5214 32528
rect 5256 32488 5296 32528
rect 4780 32320 4820 32360
rect 5356 32236 5396 32276
rect 4780 31900 4820 31940
rect 4684 31480 4724 31520
rect 4928 30976 4968 31016
rect 5010 30976 5050 31016
rect 5092 30976 5132 31016
rect 5174 30976 5214 31016
rect 5256 30976 5296 31016
rect 5068 30808 5108 30848
rect 4780 30220 4820 30260
rect 5452 31480 5492 31520
rect 5452 30976 5492 31016
rect 5452 30808 5492 30848
rect 5452 30472 5492 30512
rect 5356 30220 5396 30260
rect 5068 29716 5108 29756
rect 4928 29464 4968 29504
rect 5010 29464 5050 29504
rect 5092 29464 5132 29504
rect 5174 29464 5214 29504
rect 5256 29464 5296 29504
rect 5452 29716 5492 29756
rect 5356 29380 5396 29420
rect 5068 29296 5108 29336
rect 4684 28960 4724 29000
rect 4492 28792 4532 28832
rect 4204 28540 4244 28580
rect 4012 28372 4052 28412
rect 4204 28372 4244 28412
rect 4300 28288 4340 28328
rect 3724 28204 3764 28244
rect 4492 28120 4532 28160
rect 4300 27784 4340 27824
rect 3532 27532 3572 27572
rect 3916 27616 3956 27656
rect 4108 27616 4148 27656
rect 3820 27448 3860 27488
rect 3688 27196 3728 27236
rect 3770 27196 3810 27236
rect 3852 27196 3892 27236
rect 3934 27196 3974 27236
rect 4016 27196 4056 27236
rect 3436 27028 3476 27068
rect 3532 26692 3572 26732
rect 4204 26944 4244 26984
rect 4012 26692 4052 26732
rect 4396 26860 4436 26900
rect 4204 26524 4244 26564
rect 3436 26440 3476 26480
rect 3628 26272 3668 26312
rect 2956 26104 2996 26144
rect 2476 25012 2516 25052
rect 2668 25096 2708 25136
rect 2668 24760 2708 24800
rect 2476 24592 2516 24632
rect 2284 24172 2324 24212
rect 2668 24424 2708 24464
rect 2572 23752 2612 23792
rect 2188 23584 2228 23624
rect 2188 23332 2228 23372
rect 2476 22576 2516 22616
rect 2380 22324 2420 22364
rect 2188 22240 2228 22280
rect 2092 21988 2132 22028
rect 2284 21484 2324 21524
rect 2284 19804 2324 19844
rect 2284 19636 2324 19676
rect 2092 18880 2132 18920
rect 2092 18628 2132 18668
rect 1324 17116 1364 17156
rect 1612 17116 1652 17156
rect 1900 17704 1940 17744
rect 1804 17032 1844 17072
rect 1420 16444 1460 16484
rect 1804 16108 1844 16148
rect 2284 17788 2324 17828
rect 2284 17284 2324 17324
rect 2188 16444 2228 16484
rect 3241 26188 3281 26228
rect 4012 26272 4052 26312
rect 3340 25852 3380 25892
rect 3244 25432 3284 25472
rect 4108 26104 4148 26144
rect 3628 26020 3668 26060
rect 4204 25936 4244 25976
rect 3628 25852 3668 25892
rect 3436 25768 3476 25808
rect 3688 25684 3728 25724
rect 3770 25684 3810 25724
rect 3852 25684 3892 25724
rect 3934 25684 3974 25724
rect 4016 25684 4056 25724
rect 3628 25516 3668 25556
rect 5260 28372 5300 28412
rect 5644 33664 5684 33704
rect 5740 33496 5780 33536
rect 6220 34341 6260 34376
rect 6220 34336 6260 34341
rect 6508 35176 6548 35216
rect 6508 34336 6548 34376
rect 6220 34084 6260 34124
rect 6412 34084 6452 34124
rect 6316 33916 6356 33956
rect 6508 33832 6548 33872
rect 6412 33580 6452 33620
rect 6220 33328 6260 33368
rect 6316 33160 6356 33200
rect 5932 32992 5972 33032
rect 5740 32824 5780 32864
rect 6316 32824 6356 32864
rect 6220 32404 6260 32444
rect 7372 40216 7412 40256
rect 7276 40048 7316 40088
rect 7180 39747 7220 39752
rect 7180 39712 7220 39747
rect 7180 39040 7220 39080
rect 7180 38536 7220 38576
rect 7660 39796 7700 39836
rect 7468 38872 7508 38912
rect 7852 40048 7892 40088
rect 7852 39880 7892 39920
rect 7564 38704 7604 38744
rect 7564 38032 7604 38072
rect 7564 37780 7604 37820
rect 7084 37444 7124 37484
rect 6892 37192 6932 37232
rect 6796 37024 6836 37064
rect 6700 36856 6740 36896
rect 6892 36520 6932 36560
rect 6892 35848 6932 35888
rect 6892 35596 6932 35636
rect 6796 35260 6836 35300
rect 6700 35092 6740 35132
rect 6988 35260 7028 35300
rect 6892 34672 6932 34712
rect 6988 34504 7028 34544
rect 6700 34420 6740 34460
rect 6892 34252 6932 34292
rect 6796 33580 6836 33620
rect 6700 33496 6740 33536
rect 6604 33076 6644 33116
rect 6700 32320 6740 32360
rect 6412 32236 6452 32276
rect 5740 31648 5780 31688
rect 5644 31396 5684 31436
rect 5836 31480 5876 31520
rect 6124 31648 6164 31688
rect 6988 33412 7028 33452
rect 6412 31480 6452 31520
rect 6796 31396 6836 31436
rect 5932 30724 5972 30764
rect 5644 30220 5684 30260
rect 5740 29884 5780 29924
rect 5836 29800 5876 29840
rect 5452 28288 5492 28328
rect 4928 27952 4968 27992
rect 5010 27952 5050 27992
rect 5092 27952 5132 27992
rect 5174 27952 5214 27992
rect 5256 27952 5296 27992
rect 5356 27952 5396 27992
rect 4780 27616 4820 27656
rect 4684 26188 4724 26228
rect 5644 29128 5684 29168
rect 5836 29380 5876 29420
rect 5644 28120 5684 28160
rect 5548 27868 5588 27908
rect 5452 27784 5492 27824
rect 6028 30472 6068 30512
rect 6316 31144 6356 31184
rect 6604 31060 6644 31100
rect 6316 30640 6356 30680
rect 6700 30052 6740 30092
rect 6700 29296 6740 29336
rect 7180 36940 7220 36980
rect 7180 36520 7220 36560
rect 7372 37612 7412 37652
rect 7852 38704 7892 38744
rect 7852 38452 7892 38492
rect 7756 38032 7796 38072
rect 7852 37864 7892 37904
rect 7660 37612 7700 37652
rect 7372 37276 7412 37316
rect 7564 37024 7604 37064
rect 7372 36016 7412 36056
rect 7372 34756 7412 34796
rect 7180 34588 7220 34628
rect 7180 34336 7220 34376
rect 7276 34000 7316 34040
rect 7276 33496 7316 33536
rect 8332 42736 8372 42776
rect 8524 41896 8564 41936
rect 8716 41812 8756 41852
rect 8140 41560 8180 41600
rect 8236 41224 8276 41264
rect 8140 40636 8180 40676
rect 8044 40552 8084 40592
rect 8332 40468 8372 40508
rect 8236 39544 8276 39584
rect 8140 39292 8180 39332
rect 8044 39040 8084 39080
rect 8236 38956 8276 38996
rect 8140 38872 8180 38912
rect 8524 39880 8564 39920
rect 8428 39376 8468 39416
rect 8044 38452 8084 38492
rect 8140 38368 8180 38408
rect 8044 38284 8084 38324
rect 7756 36268 7796 36308
rect 7948 36520 7988 36560
rect 7852 36016 7892 36056
rect 7756 35932 7796 35972
rect 7852 35848 7892 35888
rect 7756 35176 7796 35216
rect 7948 35092 7988 35132
rect 7852 35008 7892 35048
rect 7756 34840 7796 34880
rect 7660 34336 7700 34376
rect 7756 34084 7796 34124
rect 7564 33832 7604 33872
rect 7756 33832 7796 33872
rect 7756 33076 7796 33116
rect 7372 32908 7412 32948
rect 6988 30052 7028 30092
rect 6988 29800 7028 29840
rect 7084 29716 7124 29756
rect 7276 30808 7316 30848
rect 7564 32824 7604 32864
rect 7564 32404 7604 32444
rect 7468 31480 7508 31520
rect 7468 30976 7508 31016
rect 7948 34840 7988 34880
rect 7948 34000 7988 34040
rect 8140 37612 8180 37652
rect 8140 37024 8180 37064
rect 8140 36856 8180 36896
rect 8140 36268 8180 36308
rect 8716 39040 8756 39080
rect 8620 38872 8660 38912
rect 8428 38452 8468 38492
rect 8332 38284 8372 38324
rect 8428 37864 8468 37904
rect 8332 36352 8372 36392
rect 8332 35848 8372 35888
rect 8236 35428 8276 35468
rect 8140 35008 8180 35048
rect 8332 35176 8372 35216
rect 8236 34840 8276 34880
rect 8620 36688 8660 36728
rect 8428 34672 8468 34712
rect 8140 34504 8180 34544
rect 8332 34504 8372 34544
rect 8236 34336 8276 34376
rect 9100 42232 9140 42272
rect 9196 42064 9236 42104
rect 9100 41056 9140 41096
rect 9100 40300 9140 40340
rect 9100 39712 9140 39752
rect 9100 39292 9140 39332
rect 9004 38872 9044 38912
rect 9004 37948 9044 37988
rect 9676 42652 9716 42692
rect 9484 42148 9524 42188
rect 10060 42148 10100 42188
rect 11020 41728 11060 41768
rect 10444 41476 10484 41516
rect 10252 41392 10292 41432
rect 9484 41140 9524 41180
rect 9676 40972 9716 41012
rect 9292 40300 9332 40340
rect 9292 39880 9332 39920
rect 9292 39628 9332 39668
rect 9292 38200 9332 38240
rect 9580 40552 9620 40592
rect 9484 40300 9524 40340
rect 9484 39880 9524 39920
rect 9676 40132 9716 40172
rect 9676 39880 9716 39920
rect 9676 39460 9716 39500
rect 9484 38956 9524 38996
rect 10156 41140 10196 41180
rect 10156 40720 10196 40760
rect 9964 40384 10004 40424
rect 10060 40132 10100 40172
rect 10156 39880 10196 39920
rect 9964 39796 10004 39836
rect 9868 39460 9908 39500
rect 9868 39292 9908 39332
rect 10060 39712 10100 39752
rect 10636 41224 10676 41264
rect 10540 41140 10580 41180
rect 10828 41476 10868 41516
rect 10732 40468 10772 40508
rect 10443 40398 10483 40438
rect 10732 40300 10772 40340
rect 10348 40048 10388 40088
rect 10348 39880 10388 39920
rect 10540 39880 10580 39920
rect 10348 39460 10388 39500
rect 11020 41140 11060 41180
rect 11020 40132 11060 40172
rect 10060 38704 10100 38744
rect 9580 38452 9620 38492
rect 9580 38032 9620 38072
rect 9484 37780 9524 37820
rect 9004 37612 9044 37652
rect 9004 37360 9044 37400
rect 9196 37612 9236 37652
rect 9484 37612 9524 37652
rect 8812 36940 8852 36980
rect 9004 36856 9044 36896
rect 9100 36688 9140 36728
rect 8908 36604 8948 36644
rect 8812 36520 8852 36560
rect 9196 36520 9236 36560
rect 9388 37444 9428 37484
rect 9868 38200 9908 38240
rect 10060 38200 10100 38240
rect 9772 37948 9812 37988
rect 9772 37612 9812 37652
rect 9772 36940 9812 36980
rect 9004 35764 9044 35804
rect 8812 35680 8852 35720
rect 8908 35092 8948 35132
rect 8332 33916 8372 33956
rect 7948 33076 7988 33116
rect 8236 33412 8276 33452
rect 7852 32068 7892 32108
rect 7660 31648 7700 31688
rect 7660 31480 7700 31520
rect 7852 31228 7892 31268
rect 8140 32068 8180 32108
rect 8044 31984 8084 32024
rect 8140 31396 8180 31436
rect 8428 33748 8468 33788
rect 8332 33076 8372 33116
rect 8428 32656 8468 32696
rect 8332 32152 8372 32192
rect 8812 34252 8852 34292
rect 8716 34168 8756 34208
rect 8620 33916 8660 33956
rect 8620 33160 8660 33200
rect 8524 32572 8564 32612
rect 8620 32488 8660 32528
rect 8524 32152 8564 32192
rect 8620 31984 8660 32024
rect 7756 30640 7796 30680
rect 6892 29464 6932 29504
rect 6316 28540 6356 28580
rect 5932 28372 5972 28412
rect 6028 28288 6068 28328
rect 5836 27868 5876 27908
rect 5740 27700 5780 27740
rect 5740 27112 5780 27152
rect 5644 27028 5684 27068
rect 5452 26524 5492 26564
rect 4928 26440 4968 26480
rect 5010 26440 5050 26480
rect 5092 26440 5132 26480
rect 5174 26440 5214 26480
rect 5256 26440 5296 26480
rect 4876 26188 4916 26228
rect 4588 26020 4628 26060
rect 4588 25852 4628 25892
rect 4300 25432 4340 25472
rect 3244 25096 3284 25136
rect 3532 25096 3572 25136
rect 3148 24676 3188 24716
rect 2860 24424 2900 24464
rect 3052 24424 3092 24464
rect 2860 23080 2900 23120
rect 3052 23752 3092 23792
rect 3436 24424 3476 24464
rect 3436 24004 3476 24044
rect 3340 23920 3380 23960
rect 4012 25180 4052 25220
rect 3628 24844 3668 24884
rect 3820 24592 3860 24632
rect 3628 24340 3668 24380
rect 4396 24676 4436 24716
rect 4108 24592 4148 24632
rect 3688 24172 3728 24212
rect 3770 24172 3810 24212
rect 3852 24172 3892 24212
rect 3934 24172 3974 24212
rect 4016 24172 4056 24212
rect 4012 24004 4052 24044
rect 3340 23752 3380 23792
rect 4204 23920 4244 23960
rect 4396 24340 4436 24380
rect 3244 23080 3284 23120
rect 2956 22996 2996 23036
rect 2956 22828 2996 22868
rect 2860 22660 2900 22700
rect 3436 22660 3476 22700
rect 3340 22576 3380 22616
rect 3820 22828 3860 22868
rect 5356 26104 5396 26144
rect 5068 26020 5108 26060
rect 4876 25348 4916 25388
rect 5164 25264 5204 25304
rect 5644 26440 5684 26480
rect 5932 26692 5972 26732
rect 6220 28288 6260 28328
rect 6124 27784 6164 27824
rect 6124 27364 6164 27404
rect 6220 27112 6260 27152
rect 6604 28456 6644 28496
rect 6508 28372 6548 28412
rect 6412 28036 6452 28076
rect 6604 27784 6644 27824
rect 6412 27112 6452 27152
rect 6508 26944 6548 26984
rect 6124 26776 6164 26816
rect 6412 26692 6452 26732
rect 6513 26692 6553 26732
rect 5932 26020 5972 26060
rect 5068 25180 5108 25220
rect 5260 25180 5300 25220
rect 5356 25096 5396 25136
rect 5548 25264 5588 25304
rect 5932 25264 5972 25304
rect 6508 26440 6548 26480
rect 6316 26356 6356 26396
rect 6412 26272 6452 26312
rect 5644 25096 5684 25136
rect 5836 25096 5876 25136
rect 4928 24928 4968 24968
rect 5010 24928 5050 24968
rect 5092 24928 5132 24968
rect 5174 24928 5214 24968
rect 5256 24928 5296 24968
rect 4780 24676 4820 24716
rect 4492 23752 4532 23792
rect 4588 23668 4628 23708
rect 4876 24088 4916 24128
rect 4780 23836 4820 23876
rect 5548 24592 5588 24632
rect 5356 24508 5396 24548
rect 6220 25096 6260 25136
rect 5644 24004 5684 24044
rect 4972 23920 5012 23960
rect 4780 23416 4820 23456
rect 4928 23416 4968 23456
rect 5010 23416 5050 23456
rect 5092 23416 5132 23456
rect 5174 23416 5214 23456
rect 5256 23416 5296 23456
rect 4108 22996 4148 23036
rect 4492 22996 4532 23036
rect 5356 22996 5396 23036
rect 3688 22660 3728 22700
rect 3770 22660 3810 22700
rect 3852 22660 3892 22700
rect 3934 22660 3974 22700
rect 4016 22660 4056 22700
rect 4300 22576 4340 22616
rect 3148 22408 3188 22448
rect 2668 22072 2708 22112
rect 2860 22072 2900 22112
rect 2572 21904 2612 21944
rect 2668 21568 2708 21608
rect 2476 21484 2516 21524
rect 2860 21484 2900 21524
rect 2572 21148 2612 21188
rect 3436 21904 3476 21944
rect 3340 21820 3380 21860
rect 3052 21568 3092 21608
rect 2956 20980 2996 21020
rect 2860 20896 2900 20936
rect 2668 20644 2708 20684
rect 3340 21484 3380 21524
rect 3148 21400 3188 21440
rect 2572 20392 2612 20432
rect 3052 20392 3092 20432
rect 2956 20224 2996 20264
rect 2476 20056 2516 20096
rect 2956 20056 2996 20096
rect 2668 19468 2708 19508
rect 2476 19216 2516 19256
rect 2764 19384 2804 19424
rect 2476 17788 2516 17828
rect 2476 17620 2516 17660
rect 1996 15940 2036 15980
rect 1516 15856 1556 15896
rect 1516 15520 1556 15560
rect 1228 14932 1268 14972
rect 1228 14680 1268 14720
rect 1228 14512 1268 14552
rect 1228 14008 1268 14048
rect 1708 15436 1748 15476
rect 2668 18544 2708 18584
rect 2668 17704 2708 17744
rect 2956 19468 2996 19508
rect 2956 19216 2996 19256
rect 2860 19132 2900 19172
rect 3244 20812 3284 20852
rect 3148 19636 3188 19676
rect 3148 19132 3188 19172
rect 3340 20392 3380 20432
rect 3724 21820 3764 21860
rect 4492 22408 4532 22448
rect 4396 22324 4436 22364
rect 3916 21736 3956 21776
rect 3916 21484 3956 21524
rect 3820 21400 3860 21440
rect 4300 21820 4340 21860
rect 4396 21736 4436 21776
rect 4684 22240 4724 22280
rect 4204 21568 4244 21608
rect 4588 21568 4628 21608
rect 4396 21400 4436 21440
rect 3688 21148 3728 21188
rect 3770 21148 3810 21188
rect 3852 21148 3892 21188
rect 3934 21148 3974 21188
rect 4016 21148 4056 21188
rect 4012 20896 4052 20936
rect 3532 20812 3572 20852
rect 3820 20560 3860 20600
rect 3436 20224 3476 20264
rect 3628 20224 3668 20264
rect 3532 20056 3572 20096
rect 3436 19720 3476 19760
rect 3436 19384 3476 19424
rect 3436 19216 3476 19256
rect 3340 19048 3380 19088
rect 3340 18628 3380 18668
rect 3244 18292 3284 18332
rect 2956 17032 2996 17072
rect 3244 17704 3284 17744
rect 2764 16780 2804 16820
rect 2572 16024 2612 16064
rect 1996 14848 2036 14888
rect 1900 14512 1940 14552
rect 1708 14260 1748 14300
rect 1420 13924 1460 13964
rect 1420 13672 1460 13712
rect 1324 11992 1364 12032
rect 1324 11656 1364 11696
rect 1324 10984 1364 11024
rect 1132 10816 1172 10856
rect 1804 14008 1844 14048
rect 2476 14932 2516 14972
rect 2476 14680 2516 14720
rect 2380 14344 2420 14384
rect 3244 16780 3284 16820
rect 3244 15604 3284 15644
rect 2764 15520 2804 15560
rect 3052 15520 3092 15560
rect 2668 15352 2708 15392
rect 2668 14932 2708 14972
rect 3052 14764 3092 14804
rect 2956 14680 2996 14720
rect 2284 14176 2324 14216
rect 2092 14008 2132 14048
rect 1708 13168 1748 13208
rect 1708 12580 1748 12620
rect 1612 11068 1652 11108
rect 2188 13840 2228 13880
rect 2860 14092 2900 14132
rect 2572 13924 2612 13964
rect 2764 13840 2804 13880
rect 2380 13588 2420 13628
rect 2284 12244 2324 12284
rect 2092 12160 2132 12200
rect 1900 11488 1940 11528
rect 1804 11068 1844 11108
rect 1228 9472 1268 9512
rect 1420 10144 1460 10184
rect 1612 9724 1652 9764
rect 1612 9304 1652 9344
rect 1420 9220 1460 9260
rect 1228 8800 1268 8840
rect 1331 8800 1371 8840
rect 844 6952 884 6992
rect 652 6448 692 6488
rect 652 6196 692 6236
rect 556 2500 596 2540
rect 268 904 308 944
rect 748 2500 788 2540
rect 748 2080 788 2120
rect 1036 5356 1076 5396
rect 844 1828 884 1868
rect 652 400 692 440
rect 1420 8716 1460 8756
rect 1996 10900 2036 10940
rect 1996 9808 2036 9848
rect 1900 9304 1940 9344
rect 1804 9052 1844 9092
rect 2188 10396 2228 10436
rect 2188 10228 2228 10268
rect 1804 8716 1844 8756
rect 1516 8464 1556 8504
rect 1420 7456 1460 7496
rect 1324 7120 1364 7160
rect 1324 6952 1364 6992
rect 1228 5608 1268 5648
rect 1612 7960 1652 8000
rect 2284 9892 2324 9932
rect 2476 12412 2516 12452
rect 2476 11404 2516 11444
rect 2476 10984 2516 11024
rect 2380 9808 2420 9848
rect 2380 9472 2420 9512
rect 2668 13336 2708 13376
rect 2860 13336 2900 13376
rect 3148 14512 3188 14552
rect 3052 14176 3092 14216
rect 2956 13084 2996 13124
rect 2860 12580 2900 12620
rect 3244 13756 3284 13796
rect 3244 13588 3284 13628
rect 3436 17956 3476 17996
rect 4204 20728 4244 20768
rect 4108 20392 4148 20432
rect 4396 20896 4436 20936
rect 4396 20644 4436 20684
rect 4406 20392 4446 20432
rect 4684 20728 4724 20768
rect 4876 22828 4916 22868
rect 5356 22744 5396 22784
rect 4876 22576 4916 22616
rect 5452 22324 5492 22364
rect 4928 21904 4968 21944
rect 5010 21904 5050 21944
rect 5092 21904 5132 21944
rect 5174 21904 5214 21944
rect 5256 21904 5296 21944
rect 5356 21400 5396 21440
rect 4876 21064 4916 21104
rect 4780 20644 4820 20684
rect 5356 20728 5396 20768
rect 4684 20560 4724 20600
rect 4876 20560 4916 20600
rect 3916 19888 3956 19928
rect 4396 19972 4436 20012
rect 4108 19888 4148 19928
rect 3628 19804 3668 19844
rect 3688 19636 3728 19676
rect 3770 19636 3810 19676
rect 3852 19636 3892 19676
rect 3934 19636 3974 19676
rect 4016 19636 4056 19676
rect 4012 19468 4052 19508
rect 3628 19384 3668 19424
rect 3820 19216 3860 19256
rect 3916 18712 3956 18752
rect 3628 18544 3668 18584
rect 3820 18544 3860 18584
rect 3628 18376 3668 18416
rect 4204 19804 4244 19844
rect 4928 20392 4968 20432
rect 5010 20392 5050 20432
rect 5092 20392 5132 20432
rect 5174 20392 5214 20432
rect 5256 20392 5296 20432
rect 4492 19468 4532 19508
rect 5260 19468 5300 19508
rect 5548 20224 5588 20264
rect 5740 22156 5780 22196
rect 5836 22072 5876 22112
rect 6796 28288 6836 28328
rect 6892 28204 6932 28244
rect 7276 28372 7316 28412
rect 7660 29800 7700 29840
rect 7564 28876 7604 28916
rect 7372 27700 7412 27740
rect 7564 27700 7604 27740
rect 7468 27616 7508 27656
rect 7084 27112 7124 27152
rect 6796 26776 6836 26816
rect 6604 26356 6644 26396
rect 6892 26272 6932 26312
rect 7180 27028 7220 27068
rect 7276 26860 7316 26900
rect 6604 26104 6644 26144
rect 7180 26692 7220 26732
rect 6508 25768 6548 25808
rect 7372 26524 7412 26564
rect 7276 26440 7316 26480
rect 6988 25768 7028 25808
rect 7180 25768 7220 25808
rect 6604 25264 6644 25304
rect 6316 24592 6356 24632
rect 6508 24760 6548 24800
rect 6508 24424 6548 24464
rect 6412 23836 6452 23876
rect 6124 23080 6164 23120
rect 6220 22744 6260 22784
rect 6124 21904 6164 21944
rect 6028 21736 6068 21776
rect 6124 21568 6164 21608
rect 5836 20728 5876 20768
rect 5836 20392 5876 20432
rect 5740 19888 5780 19928
rect 4396 19048 4436 19088
rect 4204 18796 4244 18836
rect 4108 18376 4148 18416
rect 4012 18292 4052 18332
rect 3688 18124 3728 18164
rect 3770 18124 3810 18164
rect 3852 18124 3892 18164
rect 3934 18124 3974 18164
rect 4016 18124 4056 18164
rect 4928 18880 4968 18920
rect 5010 18880 5050 18920
rect 5092 18880 5132 18920
rect 5174 18880 5214 18920
rect 5256 18880 5296 18920
rect 5260 18628 5300 18668
rect 3532 17536 3572 17576
rect 3916 17116 3956 17156
rect 4108 16948 4148 16988
rect 3628 16780 3668 16820
rect 4108 16780 4148 16820
rect 3688 16612 3728 16652
rect 3770 16612 3810 16652
rect 3852 16612 3892 16652
rect 3934 16612 3974 16652
rect 4016 16612 4056 16652
rect 3436 16360 3476 16400
rect 3916 16360 3956 16400
rect 3820 16276 3860 16316
rect 3724 16192 3764 16232
rect 3724 15772 3764 15812
rect 4204 16360 4244 16400
rect 4204 16192 4244 16232
rect 4012 15520 4052 15560
rect 3688 15100 3728 15140
rect 3770 15100 3810 15140
rect 3852 15100 3892 15140
rect 3934 15100 3974 15140
rect 4016 15100 4056 15140
rect 3340 13420 3380 13460
rect 3340 13000 3380 13040
rect 2956 11740 2996 11780
rect 2860 11656 2900 11696
rect 2764 11572 2804 11612
rect 2668 11404 2708 11444
rect 2572 10144 2612 10184
rect 2860 11236 2900 11276
rect 2764 11068 2804 11108
rect 2668 9472 2708 9512
rect 2284 8800 2324 8840
rect 1996 8128 2036 8168
rect 1900 6952 1940 6992
rect 1804 6868 1844 6908
rect 1516 6448 1556 6488
rect 1324 4096 1364 4136
rect 1516 4180 1556 4220
rect 1516 3340 1556 3380
rect 1516 1996 1556 2036
rect 1228 1828 1268 1868
rect 1420 1660 1460 1700
rect 1900 6784 1940 6824
rect 1708 6280 1748 6320
rect 2188 7876 2228 7916
rect 2092 7120 2132 7160
rect 1996 6700 2036 6740
rect 2092 6616 2132 6656
rect 2188 6280 2228 6320
rect 2092 4852 2132 4892
rect 2380 6448 2420 6488
rect 2380 6280 2420 6320
rect 2572 8548 2612 8588
rect 2572 6952 2612 6992
rect 2572 6280 2612 6320
rect 3148 11908 3188 11948
rect 3244 10816 3284 10856
rect 3052 9808 3092 9848
rect 3532 14680 3572 14720
rect 3916 14848 3956 14888
rect 4012 14764 4052 14804
rect 4396 15268 4436 15308
rect 4300 14932 4340 14972
rect 5740 19216 5780 19256
rect 5644 18964 5684 19004
rect 6316 21568 6356 21608
rect 6604 23332 6644 23372
rect 6700 23080 6740 23120
rect 6892 24508 6932 24548
rect 6892 23752 6932 23792
rect 6604 21988 6644 22028
rect 6508 21736 6548 21776
rect 6412 20896 6452 20936
rect 6316 20728 6356 20768
rect 5452 18544 5492 18584
rect 5836 18544 5876 18584
rect 6028 19804 6068 19844
rect 6028 19216 6068 19256
rect 6412 19720 6452 19760
rect 6316 19468 6356 19508
rect 5452 18292 5492 18332
rect 5932 18292 5972 18332
rect 4588 17452 4628 17492
rect 4928 17368 4968 17408
rect 5010 17368 5050 17408
rect 5092 17368 5132 17408
rect 5174 17368 5214 17408
rect 5256 17368 5296 17408
rect 4972 16948 5012 16988
rect 4684 16864 4724 16904
rect 5164 17032 5204 17072
rect 5932 17704 5972 17744
rect 6220 19132 6260 19172
rect 6124 18712 6164 18752
rect 6124 18544 6164 18584
rect 5489 17116 5529 17156
rect 5740 17452 5780 17492
rect 5836 17200 5876 17240
rect 6316 18124 6356 18164
rect 6412 17956 6452 17996
rect 6796 22660 6836 22700
rect 7180 24592 7220 24632
rect 6988 22660 7028 22700
rect 6988 22492 7028 22532
rect 7084 22324 7124 22364
rect 7372 26272 7412 26312
rect 7564 26776 7604 26816
rect 7564 25852 7604 25892
rect 7468 25264 7508 25304
rect 7180 22240 7220 22280
rect 6892 21736 6932 21776
rect 6796 21568 6836 21608
rect 6892 21316 6932 21356
rect 6892 20980 6932 21020
rect 6604 19216 6644 19256
rect 6892 19888 6932 19928
rect 6700 18880 6740 18920
rect 7084 21568 7124 21608
rect 7084 19804 7124 19844
rect 6988 18796 7028 18836
rect 6604 18628 6644 18668
rect 7372 21568 7412 21608
rect 7372 19972 7412 20012
rect 7948 30472 7988 30512
rect 7948 30136 7988 30176
rect 8428 31060 8468 31100
rect 8428 30892 8468 30932
rect 7852 29632 7892 29672
rect 8332 29800 8372 29840
rect 8524 29800 8564 29840
rect 8428 29296 8468 29336
rect 9004 34000 9044 34040
rect 8812 33916 8852 33956
rect 8812 33748 8852 33788
rect 9004 33244 9044 33284
rect 9004 33076 9044 33116
rect 9388 36016 9428 36056
rect 9196 35092 9236 35132
rect 9196 34336 9236 34376
rect 9580 35848 9620 35888
rect 9388 35596 9428 35636
rect 9388 34756 9428 34796
rect 9292 34000 9332 34040
rect 9196 32824 9236 32864
rect 9388 32824 9428 32864
rect 9388 32152 9428 32192
rect 9100 31480 9140 31520
rect 9196 31228 9236 31268
rect 8908 30556 8948 30596
rect 8812 29800 8852 29840
rect 9388 30640 9428 30680
rect 9100 30304 9140 30344
rect 9580 35176 9620 35216
rect 9580 34588 9620 34628
rect 9580 33664 9620 33704
rect 9964 37948 10004 37988
rect 10060 37864 10100 37904
rect 10444 38956 10484 38996
rect 10252 38872 10292 38912
rect 10252 38536 10292 38576
rect 10252 36940 10292 36980
rect 10252 36772 10292 36812
rect 10156 35428 10196 35468
rect 10060 35344 10100 35384
rect 9964 35092 10004 35132
rect 10156 35260 10196 35300
rect 9868 33748 9908 33788
rect 9868 33496 9908 33536
rect 9676 33244 9716 33284
rect 9676 32824 9716 32864
rect 10060 33832 10100 33872
rect 10060 33412 10100 33452
rect 10540 37780 10580 37820
rect 10444 36688 10484 36728
rect 10348 36016 10388 36056
rect 10252 33832 10292 33872
rect 10444 35092 10484 35132
rect 10444 34252 10484 34292
rect 10444 34084 10484 34124
rect 10636 35512 10676 35552
rect 10924 39208 10964 39248
rect 10924 39040 10964 39080
rect 11308 41560 11348 41600
rect 11212 40048 11252 40088
rect 11500 40972 11540 41012
rect 11500 40216 11540 40256
rect 11404 39880 11444 39920
rect 11116 39376 11156 39416
rect 11020 38536 11060 38576
rect 10924 37444 10964 37484
rect 10828 37108 10868 37148
rect 10828 36772 10868 36812
rect 11404 39712 11444 39752
rect 11212 39208 11252 39248
rect 11212 39040 11252 39080
rect 11692 42148 11732 42188
rect 11692 40384 11732 40424
rect 11980 42064 12020 42104
rect 11884 41308 11924 41348
rect 12364 42484 12404 42524
rect 12556 41560 12596 41600
rect 12652 41392 12692 41432
rect 12556 41308 12596 41348
rect 12460 41224 12500 41264
rect 12172 41140 12212 41180
rect 11596 38620 11636 38660
rect 11308 38116 11348 38156
rect 11596 38116 11636 38156
rect 11212 37864 11252 37904
rect 11596 37864 11636 37904
rect 11116 37780 11156 37820
rect 11020 37024 11060 37064
rect 10828 36520 10868 36560
rect 10732 35260 10772 35300
rect 11692 37528 11732 37568
rect 11596 37360 11636 37400
rect 12268 40972 12308 41012
rect 11980 39544 12020 39584
rect 11884 38872 11924 38912
rect 11980 38788 12020 38828
rect 11884 38620 11924 38660
rect 11212 36856 11252 36896
rect 11212 35932 11252 35972
rect 11596 36016 11636 36056
rect 11116 35512 11156 35552
rect 11020 35344 11060 35384
rect 10924 35092 10964 35132
rect 10924 34504 10964 34544
rect 10252 33076 10292 33116
rect 10348 32908 10388 32948
rect 9580 32488 9620 32528
rect 9580 31984 9620 32024
rect 9676 31228 9716 31268
rect 9676 30640 9716 30680
rect 10060 32656 10100 32696
rect 9868 32488 9908 32528
rect 10060 31816 10100 31856
rect 10540 33664 10580 33704
rect 10828 34168 10868 34208
rect 10540 32824 10580 32864
rect 10444 32656 10484 32696
rect 10732 32488 10772 32528
rect 10636 32320 10676 32360
rect 10636 32068 10676 32108
rect 10636 31732 10676 31772
rect 10156 31396 10196 31436
rect 9964 31228 10004 31268
rect 10444 31228 10484 31268
rect 9868 30808 9908 30848
rect 9484 30136 9524 30176
rect 10444 30472 10484 30512
rect 10156 30388 10196 30428
rect 9100 30052 9140 30092
rect 9964 30052 10004 30092
rect 8716 29632 8756 29672
rect 9004 29632 9044 29672
rect 8716 29296 8756 29336
rect 9196 29632 9236 29672
rect 8236 29128 8276 29168
rect 8524 29128 8564 29168
rect 8908 29128 8948 29168
rect 8140 27952 8180 27992
rect 8044 27784 8084 27824
rect 8044 27616 8084 27656
rect 7756 27448 7796 27488
rect 8812 28708 8852 28748
rect 8716 28624 8756 28664
rect 8428 28372 8468 28412
rect 8620 28288 8660 28328
rect 8908 28288 8948 28328
rect 8524 28204 8564 28244
rect 8428 27952 8468 27992
rect 8332 27784 8372 27824
rect 8812 27784 8852 27824
rect 9484 29800 9524 29840
rect 10252 30220 10292 30260
rect 10060 29632 10100 29672
rect 9196 29212 9236 29252
rect 9388 29044 9428 29084
rect 9580 29044 9620 29084
rect 9964 29212 10004 29252
rect 9772 28960 9812 29000
rect 9484 28708 9524 28748
rect 9676 28708 9716 28748
rect 9868 28624 9908 28664
rect 9388 28372 9428 28412
rect 9100 28288 9140 28328
rect 9484 28288 9524 28328
rect 9868 28288 9908 28328
rect 10156 28960 10196 29000
rect 7852 26272 7892 26312
rect 7660 25180 7700 25220
rect 7852 26104 7892 26144
rect 7756 24004 7796 24044
rect 7852 23500 7892 23540
rect 8524 27616 8564 27656
rect 8908 27700 8948 27740
rect 8428 27532 8468 27572
rect 9004 27532 9044 27572
rect 8524 27448 8564 27488
rect 8620 27196 8660 27236
rect 8428 26272 8468 26312
rect 8428 26104 8468 26144
rect 8236 25768 8276 25808
rect 8236 24928 8276 24968
rect 8140 24340 8180 24380
rect 8140 24172 8180 24212
rect 8140 23500 8180 23540
rect 7660 22408 7700 22448
rect 7564 22240 7604 22280
rect 7564 22072 7604 22112
rect 8044 23080 8084 23120
rect 8332 24592 8372 24632
rect 8332 23836 8372 23876
rect 8332 22996 8372 23036
rect 8812 27028 8852 27068
rect 9388 27700 9428 27740
rect 9484 27448 9524 27488
rect 9100 27028 9140 27068
rect 8716 26776 8756 26816
rect 11212 35176 11252 35216
rect 11596 35344 11636 35384
rect 11596 35176 11636 35216
rect 11020 34420 11060 34460
rect 11020 33748 11060 33788
rect 11212 33580 11252 33620
rect 11116 33412 11156 33452
rect 11020 32740 11060 32780
rect 11116 31144 11156 31184
rect 11020 30136 11060 30176
rect 10444 29808 10484 29840
rect 10444 29800 10484 29808
rect 10444 29632 10484 29672
rect 10348 29296 10388 29336
rect 10636 29800 10676 29840
rect 10540 29212 10580 29252
rect 10060 28120 10100 28160
rect 10060 27700 10100 27740
rect 9868 27448 9908 27488
rect 8812 25936 8852 25976
rect 8812 25516 8852 25556
rect 9004 25768 9044 25808
rect 9580 26608 9620 26648
rect 9964 26776 10004 26816
rect 9868 26524 9908 26564
rect 10636 29128 10676 29168
rect 11020 29632 11060 29672
rect 11308 32404 11348 32444
rect 11308 32236 11348 32276
rect 11596 33832 11636 33872
rect 11788 36604 11828 36644
rect 11980 38452 12020 38492
rect 11980 38116 12020 38156
rect 13132 41644 13172 41684
rect 13324 41560 13364 41600
rect 13708 41896 13748 41936
rect 13516 41476 13556 41516
rect 14380 42400 14420 42440
rect 14284 42316 14324 42356
rect 14092 41728 14132 41768
rect 13900 41392 13940 41432
rect 13708 41224 13748 41264
rect 14188 41056 14228 41096
rect 13900 40972 13940 41012
rect 13036 40636 13076 40676
rect 12652 40300 12692 40340
rect 12556 39544 12596 39584
rect 12172 38872 12212 38912
rect 12172 38452 12212 38492
rect 12076 37696 12116 37736
rect 12076 37528 12116 37568
rect 11884 35848 11924 35888
rect 11788 34504 11828 34544
rect 11692 33664 11732 33704
rect 11596 33496 11636 33536
rect 11596 33328 11636 33368
rect 11500 32152 11540 32192
rect 11596 31732 11636 31772
rect 11308 31648 11348 31688
rect 11692 31648 11732 31688
rect 11596 31480 11636 31520
rect 11308 31396 11348 31436
rect 11404 30472 11444 30512
rect 11308 30304 11348 30344
rect 11692 31312 11732 31352
rect 11692 31060 11732 31100
rect 11596 30472 11636 30512
rect 11692 29968 11732 30008
rect 11308 29212 11348 29252
rect 11212 29128 11252 29168
rect 10540 28540 10580 28580
rect 10444 28288 10484 28328
rect 10828 28960 10868 29000
rect 10828 28792 10868 28832
rect 10732 28708 10772 28748
rect 10924 28456 10964 28496
rect 9868 26104 9908 26144
rect 10060 26104 10100 26144
rect 9676 25936 9716 25976
rect 9868 25936 9908 25976
rect 8620 25180 8660 25220
rect 8620 24928 8660 24968
rect 8524 24760 8564 24800
rect 8524 24592 8564 24632
rect 8524 23080 8564 23120
rect 8716 24760 8756 24800
rect 9004 24592 9044 24632
rect 8908 24256 8948 24296
rect 8716 24172 8756 24212
rect 8716 23920 8756 23960
rect 8716 23752 8756 23792
rect 8716 23584 8756 23624
rect 8812 22996 8852 23036
rect 8332 22828 8372 22868
rect 8236 22324 8276 22364
rect 7948 22156 7988 22196
rect 8236 22072 8276 22112
rect 8044 21484 8084 21524
rect 7660 19720 7700 19760
rect 7276 19048 7316 19088
rect 7372 18712 7412 18752
rect 6988 18628 7028 18668
rect 6508 17704 6548 17744
rect 6316 17620 6356 17660
rect 4684 16024 4724 16064
rect 4588 15100 4628 15140
rect 4108 14596 4148 14636
rect 4108 14260 4148 14300
rect 3820 14008 3860 14048
rect 3532 13588 3572 13628
rect 3688 13588 3728 13628
rect 3770 13588 3810 13628
rect 3852 13588 3892 13628
rect 3934 13588 3974 13628
rect 4016 13588 4056 13628
rect 3628 13336 3668 13376
rect 3724 12748 3764 12788
rect 3532 12496 3572 12536
rect 4012 12580 4052 12620
rect 4204 14008 4244 14048
rect 4300 13840 4340 13880
rect 4300 13588 4340 13628
rect 4972 16024 5012 16064
rect 5260 16108 5300 16148
rect 5164 16024 5204 16064
rect 4928 15856 4968 15896
rect 5010 15856 5050 15896
rect 5092 15856 5132 15896
rect 5174 15856 5214 15896
rect 5256 15856 5296 15896
rect 4780 15688 4820 15728
rect 5164 15688 5204 15728
rect 4972 14512 5012 14552
rect 4780 14428 4820 14468
rect 4588 13420 4628 13460
rect 4588 13168 4628 13208
rect 3916 12244 3956 12284
rect 3688 12076 3728 12116
rect 3770 12076 3810 12116
rect 3852 12076 3892 12116
rect 3934 12076 3974 12116
rect 4016 12076 4056 12116
rect 3436 11404 3476 11444
rect 3436 11068 3476 11108
rect 3820 10984 3860 11024
rect 2956 9556 2996 9596
rect 2860 9304 2900 9344
rect 3340 9556 3380 9596
rect 3688 10564 3728 10604
rect 3770 10564 3810 10604
rect 3852 10564 3892 10604
rect 3934 10564 3974 10604
rect 4016 10564 4056 10604
rect 3532 10312 3572 10352
rect 3436 9220 3476 9260
rect 3340 8968 3380 9008
rect 3244 8884 3284 8924
rect 2956 8464 2996 8504
rect 3148 8632 3188 8672
rect 2860 8296 2900 8336
rect 3052 8296 3092 8336
rect 2764 8128 2804 8168
rect 3052 8128 3092 8168
rect 2956 7960 2996 8000
rect 2764 7876 2804 7916
rect 2860 6952 2900 6992
rect 2764 6616 2804 6656
rect 2860 6448 2900 6488
rect 2476 5608 2516 5648
rect 2284 4684 2324 4724
rect 2668 5524 2708 5564
rect 2572 5020 2612 5060
rect 2380 4600 2420 4640
rect 2284 4348 2324 4388
rect 1996 3592 2036 3632
rect 1804 2836 1844 2876
rect 2188 3459 2228 3464
rect 2188 3424 2228 3459
rect 2092 2668 2132 2708
rect 1900 2164 1940 2204
rect 1612 1408 1652 1448
rect 1804 1324 1844 1364
rect 1996 1828 2036 1868
rect 2188 1660 2228 1700
rect 2860 5776 2900 5816
rect 2860 5188 2900 5228
rect 3244 8548 3284 8588
rect 3148 5860 3188 5900
rect 4204 12244 4244 12284
rect 4012 9388 4052 9428
rect 4108 9304 4148 9344
rect 3916 9220 3956 9260
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 3532 8380 3572 8420
rect 3820 8716 3860 8756
rect 4396 12832 4436 12872
rect 4588 12496 4628 12536
rect 4928 14344 4968 14384
rect 5010 14344 5050 14384
rect 5092 14344 5132 14384
rect 5174 14344 5214 14384
rect 5256 14344 5296 14384
rect 5740 16612 5780 16652
rect 5644 16360 5684 16400
rect 5452 15100 5492 15140
rect 5932 16276 5972 16316
rect 5836 15688 5876 15728
rect 6028 15772 6068 15812
rect 5932 15604 5972 15644
rect 5836 15352 5876 15392
rect 5644 14764 5684 14804
rect 5356 14260 5396 14300
rect 4972 14176 5012 14216
rect 5452 14176 5492 14216
rect 5260 13168 5300 13208
rect 5740 14428 5780 14468
rect 5740 14176 5780 14216
rect 5644 13420 5684 13460
rect 6028 14932 6068 14972
rect 5932 14680 5972 14720
rect 6028 14092 6068 14132
rect 6028 13924 6068 13964
rect 5548 13168 5588 13208
rect 4928 12832 4968 12872
rect 5010 12832 5050 12872
rect 5092 12832 5132 12872
rect 5174 12832 5214 12872
rect 5256 12832 5296 12872
rect 4972 12496 5012 12536
rect 5164 12496 5204 12536
rect 4780 12328 4820 12368
rect 4684 12076 4724 12116
rect 4684 11824 4724 11864
rect 6028 13168 6068 13208
rect 5932 12748 5972 12788
rect 5932 12412 5972 12452
rect 5068 12076 5108 12116
rect 5356 12244 5396 12284
rect 5644 12244 5684 12284
rect 5164 11908 5204 11948
rect 4972 11572 5012 11612
rect 4492 11488 4532 11528
rect 4396 11236 4436 11276
rect 4300 10732 4340 10772
rect 4300 10480 4340 10520
rect 4492 10816 4532 10856
rect 4588 10732 4628 10772
rect 4492 10060 4532 10100
rect 4396 9388 4436 9428
rect 4492 9052 4532 9092
rect 4684 10312 4724 10352
rect 4684 10144 4724 10184
rect 4928 11320 4968 11360
rect 5010 11320 5050 11360
rect 5092 11320 5132 11360
rect 5174 11320 5214 11360
rect 5256 11320 5296 11360
rect 5548 11320 5588 11360
rect 5452 11236 5492 11276
rect 5068 11068 5108 11108
rect 5836 11992 5876 12032
rect 5932 11740 5972 11780
rect 5836 11656 5876 11696
rect 5932 11488 5972 11528
rect 6892 18292 6932 18332
rect 6892 17620 6932 17660
rect 6220 16276 6260 16316
rect 6316 16192 6356 16232
rect 6220 14680 6260 14720
rect 6316 13924 6356 13964
rect 6220 12496 6260 12536
rect 8044 20056 8084 20096
rect 7852 19384 7892 19424
rect 7564 19132 7604 19172
rect 8428 22072 8468 22112
rect 7756 18544 7796 18584
rect 7756 17872 7796 17912
rect 7276 17200 7316 17240
rect 7180 17032 7220 17072
rect 7084 16612 7124 16652
rect 6508 16192 6548 16232
rect 6508 14512 6548 14552
rect 6412 12412 6452 12452
rect 6316 12328 6356 12368
rect 6124 11908 6164 11948
rect 7180 16360 7220 16400
rect 6892 16192 6932 16232
rect 7084 16197 7124 16232
rect 7084 16192 7124 16197
rect 6892 16024 6932 16064
rect 7276 15856 7316 15896
rect 7180 14680 7220 14720
rect 6796 14008 6836 14048
rect 6988 14008 7028 14048
rect 6700 13924 6740 13964
rect 6796 13504 6836 13544
rect 6700 12580 6740 12620
rect 6796 12496 6836 12536
rect 6700 12160 6740 12200
rect 6892 11992 6932 12032
rect 6316 11740 6356 11780
rect 6508 11740 6548 11780
rect 5452 10816 5492 10856
rect 6220 11236 6260 11276
rect 6028 11152 6068 11192
rect 5836 10564 5876 10604
rect 5260 10228 5300 10268
rect 5452 10144 5492 10184
rect 5644 9976 5684 10016
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 4780 9556 4820 9596
rect 4780 8800 4820 8840
rect 4972 9472 5012 9512
rect 3916 8128 3956 8168
rect 4012 7876 4052 7916
rect 3532 7624 3572 7664
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 4300 8296 4340 8336
rect 4204 8128 4244 8168
rect 4108 7372 4148 7412
rect 3532 7204 3572 7244
rect 3436 6280 3476 6320
rect 3052 5608 3092 5648
rect 3340 5608 3380 5648
rect 4204 6616 4244 6656
rect 4396 6532 4436 6572
rect 4012 6448 4052 6488
rect 4300 6448 4340 6488
rect 4204 6112 4244 6152
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 3148 5272 3188 5312
rect 2668 3928 2708 3968
rect 2668 3508 2708 3548
rect 2668 3256 2708 3296
rect 2764 3172 2804 3212
rect 2380 2332 2420 2372
rect 2668 1912 2708 1952
rect 1036 316 1076 356
rect 1996 988 2036 1028
rect 2572 1240 2612 1280
rect 2380 400 2420 440
rect 3148 4600 3188 4640
rect 3532 5608 3572 5648
rect 3532 5440 3572 5480
rect 3436 5104 3476 5144
rect 3052 4180 3092 4220
rect 3340 4180 3380 4220
rect 2956 3760 2996 3800
rect 2956 3592 2996 3632
rect 2860 2584 2900 2624
rect 3244 3844 3284 3884
rect 3148 3172 3188 3212
rect 3436 3760 3476 3800
rect 3340 3088 3380 3128
rect 3244 2752 3284 2792
rect 3148 2668 3188 2708
rect 3628 5356 3668 5396
rect 3820 5776 3860 5816
rect 3916 5608 3956 5648
rect 3724 5188 3764 5228
rect 3628 4936 3668 4976
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 5068 8632 5108 8672
rect 5356 8632 5396 8672
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 5260 8128 5300 8168
rect 5068 7960 5108 8000
rect 5164 7372 5204 7412
rect 5164 7204 5204 7244
rect 4972 7120 5012 7160
rect 4588 6616 4628 6656
rect 5548 9472 5588 9512
rect 5452 8212 5492 8252
rect 6028 10816 6068 10856
rect 6028 10396 6068 10436
rect 5548 8128 5588 8168
rect 5452 7960 5492 8000
rect 5356 7120 5396 7160
rect 5452 6952 5492 6992
rect 5740 8212 5780 8252
rect 5644 7036 5684 7076
rect 4780 6784 4820 6824
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 5548 6784 5588 6824
rect 5644 6700 5684 6740
rect 5068 6616 5108 6656
rect 4684 6532 4724 6572
rect 5548 6448 5588 6488
rect 4492 5944 4532 5984
rect 4396 5860 4436 5900
rect 4300 4936 4340 4976
rect 4204 4180 4244 4220
rect 4492 5608 4532 5648
rect 5932 9472 5972 9512
rect 6220 10312 6260 10352
rect 6220 10060 6260 10100
rect 6124 8632 6164 8672
rect 5836 7876 5876 7916
rect 6124 7708 6164 7748
rect 5836 7540 5876 7580
rect 5932 7120 5972 7160
rect 6028 7036 6068 7076
rect 5836 6616 5876 6656
rect 6028 6448 6068 6488
rect 5836 6364 5876 6404
rect 5740 6280 5780 6320
rect 5644 6196 5684 6236
rect 5260 6112 5300 6152
rect 4684 5608 4724 5648
rect 5068 5608 5108 5648
rect 4588 5356 4628 5396
rect 4492 5104 4532 5144
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 4396 4432 4436 4472
rect 4396 4012 4436 4052
rect 4108 3844 4148 3884
rect 3916 3760 3956 3800
rect 3724 3508 3764 3548
rect 3628 3340 3668 3380
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 4396 3676 4436 3716
rect 4300 3004 4340 3044
rect 3532 2752 3572 2792
rect 3820 2752 3860 2792
rect 3628 2668 3668 2708
rect 3148 1240 3188 1280
rect 3052 148 3092 188
rect 4012 2416 4052 2456
rect 4108 2248 4148 2288
rect 3628 1912 3668 1952
rect 4012 1912 4052 1952
rect 4396 2920 4436 2960
rect 4396 2164 4436 2204
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 4396 1660 4436 1700
rect 3724 1240 3764 1280
rect 4108 1240 4148 1280
rect 4684 4180 4724 4220
rect 4588 4096 4628 4136
rect 5356 4012 5396 4052
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 4588 3508 4628 3548
rect 5356 3340 5396 3380
rect 4780 3256 4820 3296
rect 4684 2836 4724 2876
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 4684 2164 4724 2204
rect 5068 1828 5108 1868
rect 4876 1744 4916 1784
rect 3532 1156 3572 1196
rect 4108 1072 4148 1112
rect 3916 568 3956 608
rect 4300 904 4340 944
rect 5260 1072 5300 1112
rect 6124 6196 6164 6236
rect 5548 5440 5588 5480
rect 6412 9388 6452 9428
rect 6796 11740 6836 11780
rect 6796 11572 6836 11612
rect 6700 11068 6740 11108
rect 6604 10060 6644 10100
rect 6316 9304 6356 9344
rect 6412 9220 6452 9260
rect 6316 9052 6356 9092
rect 6604 9388 6644 9428
rect 7276 14176 7316 14216
rect 7468 17704 7508 17744
rect 7564 17620 7604 17660
rect 8140 18460 8180 18500
rect 8044 17872 8084 17912
rect 7852 17200 7892 17240
rect 7564 16276 7604 16316
rect 7564 16108 7604 16148
rect 7756 16024 7796 16064
rect 8332 19216 8372 19256
rect 8428 19132 8468 19172
rect 8332 17872 8372 17912
rect 8332 17704 8372 17744
rect 8236 17200 8276 17240
rect 7948 16360 7988 16400
rect 8236 16612 8276 16652
rect 7852 15856 7892 15896
rect 7564 15604 7604 15644
rect 7468 14680 7508 14720
rect 7660 15100 7700 15140
rect 7660 14428 7700 14468
rect 7756 14176 7796 14216
rect 7756 13588 7796 13628
rect 7564 13420 7604 13460
rect 8044 15352 8084 15392
rect 8236 15520 8276 15560
rect 8716 22912 8756 22952
rect 8620 22828 8660 22868
rect 9196 25012 9236 25052
rect 9388 24928 9428 24968
rect 9292 24592 9332 24632
rect 9196 24256 9236 24296
rect 9292 24172 9332 24212
rect 9388 24004 9428 24044
rect 9100 23080 9140 23120
rect 8716 22660 8756 22700
rect 9004 22660 9044 22700
rect 8716 22072 8756 22112
rect 8620 18964 8660 19004
rect 8524 16612 8564 16652
rect 8524 15940 8564 15980
rect 8620 15688 8660 15728
rect 8620 15520 8660 15560
rect 8140 14932 8180 14972
rect 7852 13336 7892 13376
rect 7276 11824 7316 11864
rect 7468 12412 7508 12452
rect 7660 13000 7700 13040
rect 7756 12580 7796 12620
rect 7852 12496 7892 12536
rect 7468 11992 7508 12032
rect 6988 11068 7028 11108
rect 6892 10228 6932 10268
rect 6604 9052 6644 9092
rect 6508 8968 6548 9008
rect 6796 8968 6836 9008
rect 6700 8632 6740 8672
rect 6604 8128 6644 8168
rect 6508 7288 6548 7328
rect 6316 7036 6356 7076
rect 6316 6700 6356 6740
rect 6508 6784 6548 6824
rect 6412 6616 6452 6656
rect 6700 7876 6740 7916
rect 8140 13756 8180 13796
rect 8140 13084 8180 13124
rect 8236 12580 8276 12620
rect 7660 11908 7700 11948
rect 7564 11404 7604 11444
rect 7180 11320 7220 11360
rect 7372 10984 7412 11024
rect 7084 10480 7124 10520
rect 7180 10312 7220 10352
rect 7468 10228 7508 10268
rect 7276 10060 7316 10100
rect 7084 9472 7124 9512
rect 6988 9220 7028 9260
rect 6892 7876 6932 7916
rect 7180 8632 7220 8672
rect 7948 11404 7988 11444
rect 7852 11236 7892 11276
rect 7852 10564 7892 10604
rect 8236 11992 8276 12032
rect 8140 11236 8180 11276
rect 8140 10732 8180 10772
rect 8140 10480 8180 10520
rect 7468 8968 7508 9008
rect 7948 10144 7988 10184
rect 8524 14596 8564 14636
rect 8428 14512 8468 14552
rect 8524 14344 8564 14384
rect 8428 14008 8468 14048
rect 8428 13084 8468 13124
rect 8332 10312 8372 10352
rect 8332 9892 8372 9932
rect 7660 9388 7700 9428
rect 7180 7960 7220 8000
rect 8044 9724 8084 9764
rect 8044 9472 8084 9512
rect 6796 7456 6836 7496
rect 6700 7288 6740 7328
rect 6700 7120 6740 7160
rect 5836 5692 5876 5732
rect 5740 5356 5780 5396
rect 5644 4432 5684 4472
rect 5932 5440 5972 5480
rect 5836 4348 5876 4388
rect 5836 4180 5876 4220
rect 7180 7792 7220 7832
rect 7276 7456 7316 7496
rect 6892 6532 6932 6572
rect 7852 7204 7892 7244
rect 7468 7120 7508 7160
rect 7372 7036 7412 7076
rect 7084 6784 7124 6824
rect 7468 6784 7508 6824
rect 7660 7120 7700 7160
rect 7372 6700 7412 6740
rect 7564 6700 7604 6740
rect 7276 6616 7316 6656
rect 6508 5944 6548 5984
rect 6700 6112 6740 6152
rect 7468 6532 7508 6572
rect 7468 6364 7508 6404
rect 7948 6532 7988 6572
rect 7372 6280 7412 6320
rect 6892 6112 6932 6152
rect 6796 6028 6836 6068
rect 6412 5440 6452 5480
rect 6700 5440 6740 5480
rect 6124 5020 6164 5060
rect 6316 4768 6356 4808
rect 6316 4180 6356 4220
rect 6220 4096 6260 4136
rect 6604 5188 6644 5228
rect 6508 4348 6548 4388
rect 5740 3760 5780 3800
rect 5644 3340 5684 3380
rect 5548 2584 5588 2624
rect 6028 3760 6068 3800
rect 5932 3340 5972 3380
rect 5644 2248 5684 2288
rect 6124 2584 6164 2624
rect 6028 2332 6068 2372
rect 5932 1912 5972 1952
rect 5740 1492 5780 1532
rect 5644 1156 5684 1196
rect 4876 988 4916 1028
rect 5068 988 5108 1028
rect 5452 904 5492 944
rect 4684 736 4724 776
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 5356 736 5396 776
rect 4396 652 4436 692
rect 4492 232 4532 272
rect 5068 568 5108 608
rect 4876 316 4916 356
rect 5836 1240 5876 1280
rect 6124 1156 6164 1196
rect 5548 484 5588 524
rect 5452 232 5492 272
rect 5260 148 5300 188
rect 5836 820 5876 860
rect 6028 64 6068 104
rect 6796 5188 6836 5228
rect 7276 5944 7316 5984
rect 7180 5524 7220 5564
rect 6892 4852 6932 4892
rect 6796 4348 6836 4388
rect 7084 4768 7124 4808
rect 6988 4600 7028 4640
rect 6508 3340 6548 3380
rect 6700 3340 6740 3380
rect 6604 3088 6644 3128
rect 6604 2589 6644 2624
rect 6604 2584 6644 2589
rect 6796 2500 6836 2540
rect 7084 3256 7124 3296
rect 6988 2668 7028 2708
rect 7180 2416 7220 2456
rect 7564 6280 7604 6320
rect 7852 6280 7892 6320
rect 7660 6112 7700 6152
rect 7468 5944 7508 5984
rect 7372 3928 7412 3968
rect 8524 11656 8564 11696
rect 8812 21568 8852 21608
rect 9100 22576 9140 22616
rect 9292 23332 9332 23372
rect 9292 22408 9332 22448
rect 9196 21904 9236 21944
rect 8908 21484 8948 21524
rect 10060 25012 10100 25052
rect 9868 24844 9908 24884
rect 9868 24592 9908 24632
rect 9772 24424 9812 24464
rect 9868 24088 9908 24128
rect 9676 23920 9716 23960
rect 9841 23920 9881 23960
rect 9964 23920 10004 23960
rect 9484 23584 9524 23624
rect 9772 23752 9812 23792
rect 10540 26188 10580 26228
rect 10444 24592 10484 24632
rect 10348 24508 10388 24548
rect 10060 23836 10100 23876
rect 9676 22240 9716 22280
rect 9580 21904 9620 21944
rect 9484 21568 9524 21608
rect 9868 23584 9908 23624
rect 9772 21988 9812 22028
rect 9100 20896 9140 20936
rect 9388 20812 9428 20852
rect 9004 20728 9044 20768
rect 9388 20644 9428 20684
rect 9100 19216 9140 19256
rect 9196 19132 9236 19172
rect 9100 18964 9140 19004
rect 9388 19132 9428 19172
rect 9388 18712 9428 18752
rect 8812 17872 8852 17912
rect 8908 17620 8948 17660
rect 8812 17536 8852 17576
rect 8908 16024 8948 16064
rect 8812 14512 8852 14552
rect 8716 12580 8756 12620
rect 8620 10564 8660 10604
rect 8716 10396 8756 10436
rect 8524 9304 8564 9344
rect 8812 10060 8852 10100
rect 9004 14680 9044 14720
rect 9004 13924 9044 13964
rect 9388 18376 9428 18416
rect 9292 17872 9332 17912
rect 9388 17704 9428 17744
rect 9964 23332 10004 23372
rect 10156 23416 10196 23456
rect 10156 22828 10196 22868
rect 10156 22324 10196 22364
rect 10444 24088 10484 24128
rect 11116 27784 11156 27824
rect 11020 27616 11060 27656
rect 11020 26776 11060 26816
rect 11404 28960 11444 29000
rect 11404 28204 11444 28244
rect 11404 27700 11444 27740
rect 11404 26944 11444 26984
rect 11212 26776 11252 26816
rect 10924 24592 10964 24632
rect 10732 24256 10772 24296
rect 11884 32824 11924 32864
rect 11884 32656 11924 32696
rect 12556 38620 12596 38660
rect 12556 38452 12596 38492
rect 12940 39712 12980 39752
rect 12940 39460 12980 39500
rect 12844 39208 12884 39248
rect 13036 39292 13076 39332
rect 13036 38956 13076 38996
rect 12940 38788 12980 38828
rect 12748 38704 12788 38744
rect 14284 40636 14324 40676
rect 13612 40384 13652 40424
rect 13900 40384 13940 40424
rect 13516 40300 13556 40340
rect 13324 39628 13364 39668
rect 13132 38872 13172 38912
rect 12748 37528 12788 37568
rect 12460 37276 12500 37316
rect 12172 36268 12212 36308
rect 12076 34504 12116 34544
rect 12076 34252 12116 34292
rect 12076 34084 12116 34124
rect 12364 35260 12404 35300
rect 12652 37360 12692 37400
rect 12460 34336 12500 34376
rect 12748 37276 12788 37316
rect 12940 37864 12980 37904
rect 12844 35932 12884 35972
rect 12652 34084 12692 34124
rect 12460 32740 12500 32780
rect 12460 32320 12500 32360
rect 12268 32236 12308 32276
rect 12364 32152 12404 32192
rect 12460 31648 12500 31688
rect 12364 31564 12404 31604
rect 12172 31312 12212 31352
rect 11980 30808 12020 30848
rect 11884 30724 11924 30764
rect 11884 27616 11924 27656
rect 11692 26692 11732 26732
rect 11116 26272 11156 26312
rect 11500 26272 11540 26312
rect 11020 24172 11060 24212
rect 10540 23920 10580 23960
rect 10540 23668 10580 23708
rect 10348 23164 10388 23204
rect 10348 22324 10388 22364
rect 10252 22240 10292 22280
rect 10156 22156 10196 22196
rect 10252 21988 10292 22028
rect 10924 23920 10964 23960
rect 11596 25348 11636 25388
rect 11308 24508 11348 24548
rect 11212 24088 11252 24128
rect 11404 24004 11444 24044
rect 11116 23836 11156 23876
rect 11020 23752 11060 23792
rect 10732 23416 10772 23456
rect 10540 23332 10580 23372
rect 10540 22324 10580 22364
rect 10060 21484 10100 21524
rect 10348 21904 10388 21944
rect 11116 23164 11156 23204
rect 10828 22996 10868 23036
rect 11308 22996 11348 23036
rect 11308 22828 11348 22868
rect 11116 22660 11156 22700
rect 11020 22576 11060 22616
rect 11020 22240 11060 22280
rect 11500 23332 11540 23372
rect 11884 26272 11924 26312
rect 11788 24844 11828 24884
rect 12172 30724 12212 30764
rect 12364 31144 12404 31184
rect 12268 30556 12308 30596
rect 12076 30052 12116 30092
rect 12172 29884 12212 29924
rect 12652 33160 12692 33200
rect 12844 33916 12884 33956
rect 12844 33748 12884 33788
rect 12844 33412 12884 33452
rect 12748 32404 12788 32444
rect 12748 30892 12788 30932
rect 12748 30556 12788 30596
rect 12460 29884 12500 29924
rect 12076 29632 12116 29672
rect 12172 27868 12212 27908
rect 12076 26944 12116 26984
rect 12076 26188 12116 26228
rect 12460 29212 12500 29252
rect 13036 37780 13076 37820
rect 13228 38452 13268 38492
rect 13420 39544 13460 39584
rect 13804 40216 13844 40256
rect 13708 39712 13748 39752
rect 13420 38116 13460 38156
rect 13036 37024 13076 37064
rect 13228 37276 13268 37316
rect 13420 37360 13460 37400
rect 13420 37024 13460 37064
rect 13324 36772 13364 36812
rect 13612 38704 13652 38744
rect 13708 38620 13748 38660
rect 14092 40300 14132 40340
rect 14284 40216 14324 40256
rect 14572 42568 14612 42608
rect 14476 41644 14516 41684
rect 14668 41980 14708 42020
rect 14764 41812 14804 41852
rect 14572 40720 14612 40760
rect 14572 40552 14612 40592
rect 13996 39880 14036 39920
rect 14188 39544 14228 39584
rect 14092 39460 14132 39500
rect 13708 38116 13748 38156
rect 13516 36520 13556 36560
rect 13324 35848 13364 35888
rect 13228 35764 13268 35804
rect 13324 35596 13364 35636
rect 13132 34336 13172 34376
rect 12940 31648 12980 31688
rect 12940 31312 12980 31352
rect 13132 31312 13172 31352
rect 12940 31144 12980 31184
rect 12844 29464 12884 29504
rect 12844 29128 12884 29168
rect 12652 28876 12692 28916
rect 12844 28540 12884 28580
rect 12652 28456 12692 28496
rect 12844 28288 12884 28328
rect 12652 27784 12692 27824
rect 12844 27364 12884 27404
rect 12844 27196 12884 27236
rect 12748 26776 12788 26816
rect 12364 25768 12404 25808
rect 12268 25600 12308 25640
rect 12364 25348 12404 25388
rect 12268 25264 12308 25304
rect 11692 23248 11732 23288
rect 11596 23164 11636 23204
rect 11692 22996 11732 23036
rect 11980 24508 12020 24548
rect 11884 24088 11924 24128
rect 12748 25348 12788 25388
rect 12652 24340 12692 24380
rect 12556 23752 12596 23792
rect 13036 30976 13076 31016
rect 13420 35176 13460 35216
rect 13324 35092 13364 35132
rect 13708 35428 13748 35468
rect 13228 30976 13268 31016
rect 13228 30724 13268 30764
rect 13996 37696 14036 37736
rect 13900 35848 13940 35888
rect 13900 35512 13940 35552
rect 13804 35260 13844 35300
rect 13708 34504 13748 34544
rect 13612 34168 13652 34208
rect 13996 35176 14036 35216
rect 14188 37780 14228 37820
rect 14380 39712 14420 39752
rect 14380 39292 14420 39332
rect 14956 42820 14996 42860
rect 14860 41140 14900 41180
rect 15244 42484 15284 42524
rect 15052 42064 15092 42104
rect 14956 41056 14996 41096
rect 14956 40384 14996 40424
rect 14572 40216 14612 40256
rect 14764 40216 14804 40256
rect 14860 39712 14900 39752
rect 14764 39460 14804 39500
rect 14572 39040 14612 39080
rect 14476 38368 14516 38408
rect 14668 38200 14708 38240
rect 14284 35596 14324 35636
rect 13708 34084 13748 34124
rect 13900 34000 13940 34040
rect 13804 33916 13844 33956
rect 14188 34084 14228 34124
rect 14668 37444 14708 37484
rect 14860 38032 14900 38072
rect 14860 37360 14900 37400
rect 14860 36940 14900 36980
rect 14860 36520 14900 36560
rect 14572 35932 14612 35972
rect 14764 36352 14804 36392
rect 15340 41224 15380 41264
rect 15244 40216 15284 40256
rect 15148 40048 15188 40088
rect 15052 39712 15092 39752
rect 15340 39880 15380 39920
rect 15052 38872 15092 38912
rect 15052 38200 15092 38240
rect 15244 37780 15284 37820
rect 15628 40384 15668 40424
rect 16012 42148 16052 42188
rect 15820 40636 15860 40676
rect 16588 41560 16628 41600
rect 15532 39460 15572 39500
rect 15724 39628 15764 39668
rect 16396 40048 16436 40088
rect 16300 39964 16340 40004
rect 16204 39712 16244 39752
rect 16300 39292 16340 39332
rect 16012 39040 16052 39080
rect 15628 38872 15668 38912
rect 16300 38788 16340 38828
rect 16012 38368 16052 38408
rect 15916 38200 15956 38240
rect 15532 38032 15572 38072
rect 15628 37864 15668 37904
rect 15052 37612 15092 37652
rect 15436 37612 15476 37652
rect 15532 37528 15572 37568
rect 15148 37360 15188 37400
rect 15436 37360 15476 37400
rect 15532 37192 15572 37232
rect 15052 36688 15092 36728
rect 15156 36688 15196 36728
rect 15628 37108 15668 37148
rect 15052 36520 15092 36560
rect 14764 35596 14804 35636
rect 14668 35260 14708 35300
rect 14476 35176 14516 35216
rect 14572 35092 14612 35132
rect 14956 35260 14996 35300
rect 15436 36520 15476 36560
rect 15916 37948 15956 37988
rect 15916 37360 15956 37400
rect 16396 38032 16436 38072
rect 16876 41644 16916 41684
rect 16780 41560 16820 41600
rect 16780 41308 16820 41348
rect 16684 40720 16724 40760
rect 16972 41560 17012 41600
rect 17836 42316 17876 42356
rect 17548 42232 17588 42272
rect 17740 42232 17780 42272
rect 17740 41896 17780 41936
rect 17356 41812 17396 41852
rect 17260 41728 17300 41768
rect 17164 41308 17204 41348
rect 17164 40972 17204 41012
rect 16972 40804 17012 40844
rect 17164 40552 17204 40592
rect 17356 41476 17396 41516
rect 17644 41308 17684 41348
rect 17548 40972 17588 41012
rect 17548 40552 17588 40592
rect 18412 42232 18452 42272
rect 18316 41728 18356 41768
rect 18124 41560 18164 41600
rect 17932 41476 17972 41516
rect 18220 41476 18260 41516
rect 17932 40972 17972 41012
rect 18124 40888 18164 40928
rect 17932 40552 17972 40592
rect 18316 40972 18356 41012
rect 16684 40300 16724 40340
rect 17164 40300 17204 40340
rect 17260 40132 17300 40172
rect 16780 39880 16820 39920
rect 16588 39628 16628 39668
rect 16684 38452 16724 38492
rect 16588 38368 16628 38408
rect 16108 37780 16148 37820
rect 16492 37780 16532 37820
rect 16684 37696 16724 37736
rect 16588 37612 16628 37652
rect 16204 37444 16244 37484
rect 16108 37360 16148 37400
rect 16108 36940 16148 36980
rect 15820 36856 15860 36896
rect 15724 36688 15764 36728
rect 15820 36520 15860 36560
rect 15340 36436 15380 36476
rect 15340 35596 15380 35636
rect 14764 34924 14804 34964
rect 14668 34756 14708 34796
rect 14572 34672 14612 34712
rect 14476 34336 14516 34376
rect 13804 33412 13844 33452
rect 13804 32908 13844 32948
rect 14284 33664 14324 33704
rect 14188 33580 14228 33620
rect 14380 33580 14420 33620
rect 14188 33244 14228 33284
rect 13996 32824 14036 32864
rect 13804 32236 13844 32276
rect 14380 33412 14420 33452
rect 14956 34084 14996 34124
rect 14668 34000 14708 34040
rect 14572 33496 14612 33536
rect 14476 33076 14516 33116
rect 14476 32152 14516 32192
rect 14668 32992 14708 33032
rect 14668 32656 14708 32696
rect 14860 33832 14900 33872
rect 15244 35092 15284 35132
rect 15148 34840 15188 34880
rect 15532 36436 15572 36476
rect 15532 36184 15572 36224
rect 15340 34084 15380 34124
rect 15628 35260 15668 35300
rect 15532 35008 15572 35048
rect 15436 34000 15476 34040
rect 15532 33664 15572 33704
rect 16492 37276 16532 37316
rect 16396 36940 16436 36980
rect 16300 36688 16340 36728
rect 15916 36436 15956 36476
rect 16012 36352 16052 36392
rect 15724 35008 15764 35048
rect 15724 34672 15764 34712
rect 15148 33580 15188 33620
rect 15052 32824 15092 32864
rect 14764 32320 14804 32360
rect 14284 31648 14324 31688
rect 13612 31480 13652 31520
rect 13804 31480 13844 31520
rect 14188 31480 14228 31520
rect 13516 31396 13556 31436
rect 13420 31312 13460 31352
rect 13324 30052 13364 30092
rect 13228 29884 13268 29924
rect 13708 31060 13748 31100
rect 13612 30724 13652 30764
rect 13996 31396 14036 31436
rect 14188 31312 14228 31352
rect 14092 31144 14132 31184
rect 13900 30724 13940 30764
rect 14188 30976 14228 31016
rect 13708 30472 13748 30512
rect 13996 30472 14036 30512
rect 13612 30052 13652 30092
rect 13612 29884 13652 29924
rect 13420 29800 13460 29840
rect 13996 30304 14036 30344
rect 14188 29884 14228 29924
rect 13900 29800 13940 29840
rect 13324 29716 13364 29756
rect 13804 29716 13844 29756
rect 13612 29464 13652 29504
rect 13324 29380 13364 29420
rect 13324 29128 13364 29168
rect 13804 29380 13844 29420
rect 13996 29128 14036 29168
rect 13228 28876 13268 28916
rect 13132 28540 13172 28580
rect 13324 28288 13364 28328
rect 13521 28540 13561 28580
rect 13036 28120 13076 28160
rect 13132 27616 13172 27656
rect 13708 28288 13748 28328
rect 14380 31480 14420 31520
rect 14380 30892 14420 30932
rect 14380 29800 14420 29840
rect 14284 29548 14324 29588
rect 14284 29212 14324 29252
rect 14188 29044 14228 29084
rect 13612 28120 13652 28160
rect 13804 28120 13844 28160
rect 13708 27784 13748 27824
rect 13612 27700 13652 27740
rect 13804 27532 13844 27572
rect 13516 27448 13556 27488
rect 13420 27364 13460 27404
rect 13420 26776 13460 26816
rect 13228 26608 13268 26648
rect 13420 26608 13460 26648
rect 13036 24592 13076 24632
rect 12844 24172 12884 24212
rect 12844 24004 12884 24044
rect 12748 23752 12788 23792
rect 12460 23248 12500 23288
rect 11884 22660 11924 22700
rect 11404 22156 11444 22196
rect 10732 21988 10772 22028
rect 10636 21904 10676 21944
rect 11500 21904 11540 21944
rect 11020 21820 11060 21860
rect 10540 21568 10580 21608
rect 9868 21400 9908 21440
rect 10444 21232 10484 21272
rect 10252 21148 10292 21188
rect 10156 20896 10196 20936
rect 9868 19972 9908 20012
rect 9676 19216 9716 19256
rect 9772 18460 9812 18500
rect 9676 17620 9716 17660
rect 9580 17536 9620 17576
rect 9772 17368 9812 17408
rect 9676 17200 9716 17240
rect 10156 20056 10196 20096
rect 10156 17704 10196 17744
rect 9964 17284 10004 17324
rect 9484 17032 9524 17072
rect 9388 16360 9428 16400
rect 9292 16024 9332 16064
rect 9196 14176 9236 14216
rect 9100 12580 9140 12620
rect 9004 12244 9044 12284
rect 9100 11656 9140 11696
rect 9004 10060 9044 10100
rect 8908 9724 8948 9764
rect 9484 15520 9524 15560
rect 9484 14260 9524 14300
rect 10060 16864 10100 16904
rect 10060 16360 10100 16400
rect 9868 16192 9908 16232
rect 9964 15100 10004 15140
rect 10348 20644 10388 20684
rect 10348 20224 10388 20264
rect 10348 20056 10388 20096
rect 11116 21736 11156 21776
rect 10636 20728 10676 20768
rect 11020 20644 11060 20684
rect 11308 21568 11348 21608
rect 10828 19300 10868 19340
rect 10636 18712 10676 18752
rect 10636 18460 10676 18500
rect 11020 18292 11060 18332
rect 10252 16276 10292 16316
rect 10252 15520 10292 15560
rect 10540 16276 10580 16316
rect 10444 16192 10484 16232
rect 10540 15940 10580 15980
rect 10444 15856 10484 15896
rect 10444 15520 10484 15560
rect 9964 14680 10004 14720
rect 10156 14680 10196 14720
rect 9676 14344 9716 14384
rect 9580 14176 9620 14216
rect 9868 14176 9908 14216
rect 9580 14008 9620 14048
rect 10060 14008 10100 14048
rect 9388 13084 9428 13124
rect 9388 12832 9428 12872
rect 9772 13336 9812 13376
rect 9868 13168 9908 13208
rect 9772 12832 9812 12872
rect 9292 12412 9332 12452
rect 9484 12496 9524 12536
rect 9388 12328 9428 12368
rect 9292 12244 9332 12284
rect 9388 11656 9428 11696
rect 9580 11656 9620 11696
rect 9868 12160 9908 12200
rect 9772 11908 9812 11948
rect 9676 11488 9716 11528
rect 9388 11236 9428 11276
rect 9868 11824 9908 11864
rect 10348 14680 10388 14720
rect 10252 13084 10292 13124
rect 10060 12496 10100 12536
rect 10924 18208 10964 18248
rect 10828 17200 10868 17240
rect 11212 20140 11252 20180
rect 11116 16612 11156 16652
rect 11116 16276 11156 16316
rect 11020 16192 11060 16232
rect 11116 15856 11156 15896
rect 11404 20476 11444 20516
rect 11980 22576 12020 22616
rect 12076 22240 12116 22280
rect 11692 22156 11732 22196
rect 11596 19384 11636 19424
rect 11404 18880 11444 18920
rect 11308 18292 11348 18332
rect 11308 18040 11348 18080
rect 11596 18796 11636 18836
rect 11596 17620 11636 17660
rect 11788 21988 11828 22028
rect 12076 21484 12116 21524
rect 12364 21484 12404 21524
rect 11788 21400 11828 21440
rect 11404 16528 11444 16568
rect 11692 16612 11732 16652
rect 11980 21232 12020 21272
rect 11884 19384 11924 19424
rect 11788 16528 11828 16568
rect 11404 16108 11444 16148
rect 11692 16024 11732 16064
rect 10924 15604 10964 15644
rect 11212 15604 11252 15644
rect 10828 14848 10868 14888
rect 10732 14596 10772 14636
rect 10636 14008 10676 14048
rect 10540 13924 10580 13964
rect 10828 13000 10868 13040
rect 10348 12496 10388 12536
rect 10156 12244 10196 12284
rect 9964 11488 10004 11528
rect 9868 11320 9908 11360
rect 9676 10648 9716 10688
rect 9004 9388 9044 9428
rect 8908 9052 8948 9092
rect 8716 8968 8756 9008
rect 8428 8128 8468 8168
rect 8140 7372 8180 7412
rect 8428 6952 8468 6992
rect 8140 6700 8180 6740
rect 8332 6700 8372 6740
rect 8236 6616 8276 6656
rect 8332 6448 8372 6488
rect 8812 8651 8852 8657
rect 8812 8617 8852 8651
rect 9196 9472 9236 9512
rect 9388 9472 9428 9512
rect 9292 8968 9332 9008
rect 8716 8548 8756 8588
rect 10060 10732 10100 10772
rect 9868 10228 9908 10268
rect 10060 10228 10100 10268
rect 9772 10144 9812 10184
rect 9964 10144 10004 10184
rect 9676 9304 9716 9344
rect 9580 8968 9620 9008
rect 7660 5356 7700 5396
rect 7564 4852 7604 4892
rect 7660 3928 7700 3968
rect 7660 3676 7700 3716
rect 7948 4684 7988 4724
rect 7852 4180 7892 4220
rect 7948 3592 7988 3632
rect 7756 3424 7796 3464
rect 7468 3172 7508 3212
rect 7372 3088 7412 3128
rect 7372 2920 7412 2960
rect 7756 2668 7796 2708
rect 8140 5524 8180 5564
rect 8140 5188 8180 5228
rect 8140 3928 8180 3968
rect 8044 2500 8084 2540
rect 7468 2416 7508 2456
rect 7276 2248 7316 2288
rect 6412 1240 6452 1280
rect 6796 1240 6836 1280
rect 6988 1240 7028 1280
rect 7180 1240 7220 1280
rect 6604 316 6644 356
rect 7372 904 7412 944
rect 7276 652 7316 692
rect 7276 232 7316 272
rect 7564 2080 7604 2120
rect 7660 1912 7700 1952
rect 7564 1072 7604 1112
rect 7468 820 7508 860
rect 7756 1240 7796 1280
rect 8140 1240 8180 1280
rect 7756 904 7796 944
rect 8044 904 8084 944
rect 7660 568 7700 608
rect 7948 652 7988 692
rect 9100 7960 9140 8000
rect 9004 7708 9044 7748
rect 8812 7540 8852 7580
rect 8716 7372 8756 7412
rect 8716 7120 8756 7160
rect 9196 7876 9236 7916
rect 9484 7876 9524 7916
rect 9676 8212 9716 8252
rect 9868 8632 9908 8672
rect 10444 12244 10484 12284
rect 10444 11824 10484 11864
rect 10348 11320 10388 11360
rect 10636 11992 10676 12032
rect 10732 11908 10772 11948
rect 10732 11740 10772 11780
rect 10252 10564 10292 10604
rect 10540 11152 10580 11192
rect 10348 10396 10388 10436
rect 10252 10312 10292 10352
rect 10252 10144 10292 10184
rect 10348 9892 10388 9932
rect 10444 9472 10484 9512
rect 10348 8800 10388 8840
rect 10252 8464 10292 8504
rect 9964 8128 10004 8168
rect 9772 7708 9812 7748
rect 8716 6952 8756 6992
rect 9004 6952 9044 6992
rect 9292 7036 9332 7076
rect 9676 7204 9716 7244
rect 9100 6868 9140 6908
rect 9004 6784 9044 6824
rect 8812 6532 8852 6572
rect 8716 6448 8756 6488
rect 8332 6112 8372 6152
rect 8332 5944 8372 5984
rect 8332 5188 8372 5228
rect 9100 6532 9140 6572
rect 8716 6112 8756 6152
rect 8620 5860 8660 5900
rect 8812 5860 8852 5900
rect 8524 5524 8564 5564
rect 8428 4600 8468 4640
rect 8812 4936 8852 4976
rect 8812 4768 8852 4808
rect 8716 4348 8756 4388
rect 8716 4180 8756 4220
rect 9004 5524 9044 5564
rect 9388 6952 9428 6992
rect 9580 7036 9620 7076
rect 9292 6616 9332 6656
rect 10156 7708 10196 7748
rect 10636 8716 10676 8756
rect 10540 8548 10580 8588
rect 10444 7960 10484 8000
rect 10348 7204 10388 7244
rect 10348 6700 10388 6740
rect 9580 6280 9620 6320
rect 10060 6364 10100 6404
rect 9676 5608 9716 5648
rect 10252 6280 10292 6320
rect 9004 4684 9044 4724
rect 8908 3760 8948 3800
rect 9196 5020 9236 5060
rect 9100 4096 9140 4136
rect 9004 3340 9044 3380
rect 8716 2752 8756 2792
rect 8428 1912 8468 1952
rect 8332 1240 8372 1280
rect 8524 1240 8564 1280
rect 8236 904 8276 944
rect 8812 2416 8852 2456
rect 9676 4936 9716 4976
rect 10444 6280 10484 6320
rect 10348 6028 10388 6068
rect 10348 5776 10388 5816
rect 10156 4936 10196 4976
rect 10252 4852 10292 4892
rect 10060 4180 10100 4220
rect 10348 4180 10388 4220
rect 9676 3424 9716 3464
rect 9484 3172 9524 3212
rect 9388 2668 9428 2708
rect 9100 2500 9140 2540
rect 9004 2416 9044 2456
rect 9004 2164 9044 2204
rect 8908 2080 8948 2120
rect 9004 1912 9044 1952
rect 9292 2080 9332 2120
rect 9964 2836 10004 2876
rect 9772 2668 9812 2708
rect 9484 2332 9524 2372
rect 9676 2248 9716 2288
rect 9484 2080 9524 2120
rect 9388 1912 9428 1952
rect 9676 1828 9716 1868
rect 9388 1660 9428 1700
rect 9676 1660 9716 1700
rect 9388 1324 9428 1364
rect 8908 652 8948 692
rect 9100 1072 9140 1112
rect 9004 316 9044 356
rect 9196 988 9236 1028
rect 10156 3760 10196 3800
rect 10252 3508 10292 3548
rect 10636 7708 10676 7748
rect 10636 7204 10676 7244
rect 11500 15520 11540 15560
rect 12268 21400 12308 21440
rect 12652 22828 12692 22868
rect 12748 22576 12788 22616
rect 12556 22156 12596 22196
rect 12844 21568 12884 21608
rect 12460 21232 12500 21272
rect 12652 21148 12692 21188
rect 12652 20980 12692 21020
rect 12076 19636 12116 19676
rect 11980 16948 12020 16988
rect 11884 16024 11924 16064
rect 11884 15856 11924 15896
rect 11212 14344 11252 14384
rect 11308 14176 11348 14216
rect 11788 14512 11828 14552
rect 11692 14344 11732 14384
rect 12076 15856 12116 15896
rect 12364 20056 12404 20096
rect 12652 20056 12692 20096
rect 12748 19972 12788 20012
rect 12844 19888 12884 19928
rect 12844 19552 12884 19592
rect 12268 18544 12308 18584
rect 12556 18544 12596 18584
rect 12652 18460 12692 18500
rect 12652 17704 12692 17744
rect 12364 17536 12404 17576
rect 12652 17536 12692 17576
rect 12268 17032 12308 17072
rect 13420 24256 13460 24296
rect 13324 24172 13364 24212
rect 13228 22576 13268 22616
rect 13132 21568 13172 21608
rect 14092 27028 14132 27068
rect 13996 26944 14036 26984
rect 13804 26776 13844 26816
rect 13996 26104 14036 26144
rect 13900 25600 13940 25640
rect 13996 25516 14036 25556
rect 14092 25180 14132 25220
rect 13996 25096 14036 25136
rect 14380 27112 14420 27152
rect 14380 26944 14420 26984
rect 14284 26860 14324 26900
rect 14572 31648 14612 31688
rect 15340 33244 15380 33284
rect 15244 32824 15284 32864
rect 15436 33076 15476 33116
rect 14956 31984 14996 32024
rect 14668 31480 14708 31520
rect 14860 31480 14900 31520
rect 14956 31144 14996 31184
rect 14668 30808 14708 30848
rect 14860 30640 14900 30680
rect 15148 31984 15188 32024
rect 15148 31648 15188 31688
rect 15628 32656 15668 32696
rect 16588 36520 16628 36560
rect 16492 36436 16532 36476
rect 16396 36184 16436 36224
rect 16204 35932 16244 35972
rect 16204 35596 16244 35636
rect 16300 35344 16340 35384
rect 16108 35260 16148 35300
rect 16396 35176 16436 35216
rect 15916 34336 15956 34376
rect 16204 34336 16244 34376
rect 15820 34252 15860 34292
rect 16396 34084 16436 34124
rect 15820 32908 15860 32948
rect 15916 32824 15956 32864
rect 15724 32320 15764 32360
rect 15916 32320 15956 32360
rect 15724 32152 15764 32192
rect 15916 31648 15956 31688
rect 15724 31144 15764 31184
rect 15436 30640 15476 30680
rect 14668 30388 14708 30428
rect 15148 30388 15188 30428
rect 14572 30220 14612 30260
rect 14668 30136 14708 30176
rect 15244 30304 15284 30344
rect 14860 29884 14900 29924
rect 14956 29296 14996 29336
rect 14860 29128 14900 29168
rect 14668 28120 14708 28160
rect 14572 27448 14612 27488
rect 14476 26776 14516 26816
rect 15052 29128 15092 29168
rect 16204 31816 16244 31856
rect 16588 35848 16628 35888
rect 16588 34840 16628 34880
rect 16876 38200 16916 38240
rect 16780 36856 16820 36896
rect 17164 39712 17204 39752
rect 18028 39964 18068 40004
rect 17836 39880 17876 39920
rect 18220 39628 18260 39668
rect 17548 39040 17588 39080
rect 17068 38200 17108 38240
rect 16972 37612 17012 37652
rect 17260 38620 17300 38660
rect 17260 37948 17300 37988
rect 17644 38200 17684 38240
rect 17164 37444 17204 37484
rect 17068 37276 17108 37316
rect 16972 37192 17012 37232
rect 17356 37612 17396 37652
rect 17260 37360 17300 37400
rect 16972 36940 17012 36980
rect 17164 36688 17204 36728
rect 16972 36604 17012 36644
rect 17356 37276 17396 37316
rect 17548 37108 17588 37148
rect 18124 38620 18164 38660
rect 18220 38032 18260 38072
rect 18604 42064 18644 42104
rect 18508 41980 18548 42020
rect 18508 41140 18548 41180
rect 18892 42652 18932 42692
rect 18892 42484 18932 42524
rect 18700 41392 18740 41432
rect 19948 42736 19988 42776
rect 19468 42568 19508 42608
rect 19276 42400 19316 42440
rect 19564 42148 19604 42188
rect 20048 41560 20088 41600
rect 20130 41560 20170 41600
rect 20212 41560 20252 41600
rect 20294 41560 20334 41600
rect 20376 41560 20416 41600
rect 19084 41308 19124 41348
rect 19180 41056 19220 41096
rect 18700 40972 18740 41012
rect 18604 40888 18644 40928
rect 18808 40804 18848 40844
rect 18890 40804 18930 40844
rect 18972 40804 19012 40844
rect 19054 40804 19094 40844
rect 19136 40804 19176 40844
rect 18796 40636 18836 40676
rect 18988 40636 19028 40676
rect 18604 40468 18644 40508
rect 19180 40300 19220 40340
rect 18604 40216 18644 40256
rect 19756 41140 19796 41180
rect 19372 40300 19412 40340
rect 19276 39880 19316 39920
rect 18412 39460 18452 39500
rect 19180 39628 19220 39668
rect 18988 39460 19028 39500
rect 18700 39292 18740 39332
rect 18808 39292 18848 39332
rect 18890 39292 18930 39332
rect 18972 39292 19012 39332
rect 19054 39292 19094 39332
rect 19136 39292 19176 39332
rect 18412 39208 18452 39248
rect 18604 39208 18644 39248
rect 19756 40384 19796 40424
rect 19660 40216 19700 40256
rect 19564 39124 19604 39164
rect 19468 39040 19508 39080
rect 19084 38956 19124 38996
rect 19276 38956 19316 38996
rect 18604 38872 18644 38912
rect 18412 38704 18452 38744
rect 18604 38452 18644 38492
rect 18316 37024 18356 37064
rect 17836 36940 17876 36980
rect 18028 36940 18068 36980
rect 17644 36856 17684 36896
rect 17932 36772 17972 36812
rect 17260 36520 17300 36560
rect 17068 35512 17108 35552
rect 16780 35428 16820 35468
rect 16396 33160 16436 33200
rect 16910 35008 16950 35048
rect 17164 35008 17204 35048
rect 17068 34756 17108 34796
rect 16780 33496 16820 33536
rect 16684 33244 16724 33284
rect 16588 32992 16628 33032
rect 16684 32404 16724 32444
rect 16684 31312 16724 31352
rect 16396 31144 16436 31184
rect 16876 32824 16916 32864
rect 16012 30640 16052 30680
rect 15916 30052 15956 30092
rect 15820 29968 15860 30008
rect 15436 29884 15476 29924
rect 15916 29884 15956 29924
rect 15820 29800 15860 29840
rect 15340 29212 15380 29252
rect 15244 28456 15284 28496
rect 15532 29128 15572 29168
rect 15820 29128 15860 29168
rect 15436 29044 15476 29084
rect 15628 28960 15668 29000
rect 15532 28372 15572 28412
rect 15340 27784 15380 27824
rect 14860 27532 14900 27572
rect 15148 27532 15188 27572
rect 15052 27448 15092 27488
rect 14860 27112 14900 27152
rect 14284 26608 14324 26648
rect 13804 23836 13844 23876
rect 13804 23080 13844 23120
rect 13516 22492 13556 22532
rect 13516 22156 13556 22196
rect 13420 20728 13460 20768
rect 13612 21988 13652 22028
rect 13228 19468 13268 19508
rect 13516 20056 13556 20096
rect 13036 19132 13076 19172
rect 13132 17956 13172 17996
rect 12364 15772 12404 15812
rect 12268 15520 12308 15560
rect 13420 19300 13460 19340
rect 13324 19132 13364 19172
rect 13420 18208 13460 18248
rect 13996 24760 14036 24800
rect 14572 25264 14612 25304
rect 14380 24592 14420 24632
rect 14284 24508 14324 24548
rect 14380 23836 14420 23876
rect 13996 21652 14036 21692
rect 13900 19804 13940 19844
rect 13900 19468 13940 19508
rect 13804 19132 13844 19172
rect 13900 18964 13940 19004
rect 13708 18712 13748 18752
rect 14380 22996 14420 23036
rect 14284 22324 14324 22364
rect 14188 22240 14228 22280
rect 14188 20644 14228 20684
rect 14188 19804 14228 19844
rect 15052 26524 15092 26564
rect 15244 26356 15284 26396
rect 15436 26272 15476 26312
rect 15340 26188 15380 26228
rect 15820 28540 15860 28580
rect 16204 28456 16244 28496
rect 15724 28288 15764 28328
rect 16204 28120 16244 28160
rect 15820 27616 15860 27656
rect 15628 27112 15668 27152
rect 15436 26104 15476 26144
rect 15244 25684 15284 25724
rect 15820 26356 15860 26396
rect 15724 26272 15764 26312
rect 15820 26020 15860 26060
rect 15532 25516 15572 25556
rect 15436 25432 15476 25472
rect 15436 25264 15476 25304
rect 15244 25012 15284 25052
rect 14860 24592 14900 24632
rect 14956 24340 14996 24380
rect 14764 22996 14804 23036
rect 15052 23752 15092 23792
rect 14860 22156 14900 22196
rect 14668 21064 14708 21104
rect 14476 20476 14516 20516
rect 14476 20224 14516 20264
rect 14380 20056 14420 20096
rect 14380 19552 14420 19592
rect 14380 19384 14420 19424
rect 14092 18712 14132 18752
rect 13996 18544 14036 18584
rect 13900 18460 13940 18500
rect 14092 18460 14132 18500
rect 13708 18292 13748 18332
rect 13612 18124 13652 18164
rect 13228 17704 13268 17744
rect 12940 17116 12980 17156
rect 12748 16360 12788 16400
rect 12748 15268 12788 15308
rect 12460 15100 12500 15140
rect 12172 14848 12212 14888
rect 11980 14512 12020 14552
rect 11980 14344 12020 14384
rect 11596 14176 11636 14216
rect 11788 13840 11828 13880
rect 11500 13420 11540 13460
rect 11500 13252 11540 13292
rect 11116 13168 11156 13208
rect 11404 13168 11444 13208
rect 11116 12496 11156 12536
rect 11308 12496 11348 12536
rect 11116 12328 11156 12368
rect 11116 11824 11156 11864
rect 11020 11068 11060 11108
rect 11020 10396 11060 10436
rect 10828 10228 10868 10268
rect 11308 11404 11348 11444
rect 11500 13000 11540 13040
rect 11692 13252 11732 13292
rect 11788 13168 11828 13208
rect 11980 13924 12020 13964
rect 12172 13840 12212 13880
rect 12364 13924 12404 13964
rect 11692 12496 11732 12536
rect 11596 11908 11636 11948
rect 11404 11068 11444 11108
rect 11692 11152 11732 11192
rect 11692 10816 11732 10856
rect 12268 13168 12308 13208
rect 12364 12496 12404 12536
rect 11980 12244 12020 12284
rect 12364 12244 12404 12284
rect 12268 11656 12308 11696
rect 11980 10732 12020 10772
rect 11596 10312 11636 10352
rect 11596 10060 11636 10100
rect 11404 9976 11444 10016
rect 11404 9808 11444 9848
rect 11500 9640 11540 9680
rect 10828 8716 10868 8756
rect 11116 9472 11156 9512
rect 11020 9388 11060 9428
rect 11116 9304 11156 9344
rect 11020 9136 11060 9176
rect 11308 8968 11348 9008
rect 11116 8800 11156 8840
rect 11020 8464 11060 8504
rect 10924 8128 10964 8168
rect 10924 7876 10964 7916
rect 11020 7624 11060 7664
rect 10924 7372 10964 7412
rect 10924 6280 10964 6320
rect 10732 5356 10772 5396
rect 10636 5188 10676 5228
rect 10540 4264 10580 4304
rect 10540 4096 10580 4136
rect 10636 3928 10676 3968
rect 10924 3928 10964 3968
rect 10444 3844 10484 3884
rect 11308 8464 11348 8504
rect 11596 8632 11636 8672
rect 11404 7960 11444 8000
rect 11500 7540 11540 7580
rect 11500 7372 11540 7412
rect 11884 10564 11924 10604
rect 12076 9976 12116 10016
rect 11788 9724 11828 9764
rect 12076 9808 12116 9848
rect 11884 8716 11924 8756
rect 11884 8044 11924 8084
rect 11788 7540 11828 7580
rect 11212 7288 11252 7328
rect 11500 6868 11540 6908
rect 11212 5608 11252 5648
rect 11116 5188 11156 5228
rect 11116 4971 11156 4976
rect 11116 4936 11156 4971
rect 11404 5440 11444 5480
rect 11404 5188 11444 5228
rect 11308 5104 11348 5144
rect 11212 4096 11252 4136
rect 12268 11068 12308 11108
rect 12556 14764 12596 14804
rect 12748 14680 12788 14720
rect 13612 17788 13652 17828
rect 13516 17704 13556 17744
rect 13900 18208 13940 18248
rect 13804 18124 13844 18164
rect 13708 17704 13748 17744
rect 13516 16360 13556 16400
rect 13420 15688 13460 15728
rect 13228 15604 13268 15644
rect 13324 15352 13364 15392
rect 13612 16108 13652 16148
rect 13612 15520 13652 15560
rect 13228 15268 13268 15308
rect 13132 15100 13172 15140
rect 12940 14848 12980 14888
rect 12844 13924 12884 13964
rect 12652 13840 12692 13880
rect 12748 12160 12788 12200
rect 12652 11824 12692 11864
rect 13132 14260 13172 14300
rect 13228 13924 13268 13964
rect 13228 13504 13268 13544
rect 13036 12496 13076 12536
rect 12940 11572 12980 11612
rect 12556 11068 12596 11108
rect 13228 11656 13268 11696
rect 13708 15268 13748 15308
rect 13516 14260 13556 14300
rect 13420 13420 13460 13460
rect 14188 18124 14228 18164
rect 13996 17032 14036 17072
rect 13900 16024 13940 16064
rect 13900 15268 13940 15308
rect 13804 13840 13844 13880
rect 13612 13420 13652 13460
rect 13996 14596 14036 14636
rect 13900 13168 13940 13208
rect 13612 13084 13652 13124
rect 14188 16192 14228 16232
rect 14188 15688 14228 15728
rect 14188 13084 14228 13124
rect 14092 13000 14132 13040
rect 13900 12496 13940 12536
rect 14092 12496 14132 12536
rect 13708 12244 13748 12284
rect 13516 12160 13556 12200
rect 13420 11992 13460 12032
rect 13324 11320 13364 11360
rect 13132 11068 13172 11108
rect 12460 10648 12500 10688
rect 12364 10144 12404 10184
rect 12268 9556 12308 9596
rect 12172 8884 12212 8924
rect 12268 8548 12308 8588
rect 12172 8044 12212 8084
rect 12268 7876 12308 7916
rect 11980 7456 12020 7496
rect 11692 6448 11732 6488
rect 11596 5188 11636 5228
rect 11500 4432 11540 4472
rect 11596 4180 11636 4220
rect 11116 3844 11156 3884
rect 10636 3676 10676 3716
rect 11020 3676 11060 3716
rect 10540 3508 10580 3548
rect 11404 3844 11444 3884
rect 11020 3424 11060 3464
rect 10540 3256 10580 3296
rect 10060 2500 10100 2540
rect 11116 3172 11156 3212
rect 11404 3172 11444 3212
rect 11308 3004 11348 3044
rect 10540 2668 10580 2708
rect 11116 2668 11156 2708
rect 10636 2500 10676 2540
rect 10252 2416 10292 2456
rect 9868 2248 9908 2288
rect 9484 1156 9524 1196
rect 9388 1072 9428 1112
rect 9388 484 9428 524
rect 9580 1072 9620 1112
rect 10252 1996 10292 2036
rect 10060 1828 10100 1868
rect 10540 2416 10580 2456
rect 10444 1576 10484 1616
rect 9964 988 10004 1028
rect 10252 820 10292 860
rect 10540 1492 10580 1532
rect 10540 1240 10580 1280
rect 10924 2584 10964 2624
rect 10828 2164 10868 2204
rect 11020 2500 11060 2540
rect 10924 1828 10964 1868
rect 11404 2416 11444 2456
rect 11596 2416 11636 2456
rect 11500 2332 11540 2372
rect 11308 2164 11348 2204
rect 11212 1828 11252 1868
rect 11212 1240 11252 1280
rect 11500 1156 11540 1196
rect 11212 1072 11252 1112
rect 10924 820 10964 860
rect 11116 820 11156 860
rect 11212 568 11252 608
rect 11116 484 11156 524
rect 11404 820 11444 860
rect 11308 148 11348 188
rect 11884 6196 11924 6236
rect 11788 5608 11828 5648
rect 11884 5188 11924 5228
rect 12076 6616 12116 6656
rect 11788 5104 11828 5144
rect 11980 4936 12020 4976
rect 12268 5860 12308 5900
rect 13324 10900 13364 10940
rect 13036 10732 13076 10772
rect 12940 10564 12980 10604
rect 12556 8968 12596 9008
rect 12556 8548 12596 8588
rect 12556 8128 12596 8168
rect 12748 10060 12788 10100
rect 13132 10144 13172 10184
rect 13996 12160 14036 12200
rect 13804 11572 13844 11612
rect 13228 9976 13268 10016
rect 13708 10648 13748 10688
rect 13612 9976 13652 10016
rect 13324 9472 13364 9512
rect 13516 9472 13556 9512
rect 13036 9052 13076 9092
rect 13036 8800 13076 8840
rect 12748 8548 12788 8588
rect 12844 7960 12884 8000
rect 13132 8632 13172 8672
rect 13228 8464 13268 8504
rect 13516 8968 13556 9008
rect 13420 8716 13460 8756
rect 13324 8212 13364 8252
rect 13228 8128 13268 8168
rect 12556 7876 12596 7916
rect 12364 5692 12404 5732
rect 12460 5608 12500 5648
rect 12748 7288 12788 7328
rect 13324 7960 13364 8000
rect 13708 9472 13748 9512
rect 13900 11236 13940 11276
rect 14188 12244 14228 12284
rect 14380 18124 14420 18164
rect 14380 17872 14420 17912
rect 14380 16276 14420 16316
rect 14380 14092 14420 14132
rect 14668 20644 14708 20684
rect 15148 21484 15188 21524
rect 14860 20980 14900 21020
rect 14764 19972 14804 20012
rect 14860 19804 14900 19844
rect 15244 19804 15284 19844
rect 15244 19216 15284 19256
rect 14860 19048 14900 19088
rect 15052 19048 15092 19088
rect 14668 18796 14708 18836
rect 14764 18124 14804 18164
rect 14572 17872 14612 17912
rect 14764 17788 14804 17828
rect 14956 18880 14996 18920
rect 15148 18880 15188 18920
rect 15820 25096 15860 25136
rect 15820 23332 15860 23372
rect 15724 23164 15764 23204
rect 15628 22660 15668 22700
rect 15532 22576 15572 22616
rect 15724 22576 15764 22616
rect 15820 21232 15860 21272
rect 16396 30220 16436 30260
rect 16780 30556 16820 30596
rect 16780 29296 16820 29336
rect 16492 29212 16532 29252
rect 16684 29212 16724 29252
rect 16396 29128 16436 29168
rect 16588 28960 16628 29000
rect 16396 28288 16436 28328
rect 16300 27784 16340 27824
rect 16300 27616 16340 27656
rect 16684 28120 16724 28160
rect 17452 36604 17492 36644
rect 17356 35932 17396 35972
rect 17452 35512 17492 35552
rect 17356 35344 17396 35384
rect 17452 35176 17492 35216
rect 18028 35596 18068 35636
rect 17836 35428 17876 35468
rect 17740 35176 17780 35216
rect 18028 35260 18068 35300
rect 17932 35092 17972 35132
rect 17356 34924 17396 34964
rect 17260 33244 17300 33284
rect 17068 32740 17108 32780
rect 16972 32152 17012 32192
rect 17068 31732 17108 31772
rect 17260 32992 17300 33032
rect 17644 34588 17684 34628
rect 17452 34336 17492 34376
rect 17932 34840 17972 34880
rect 17836 34084 17876 34124
rect 18028 34588 18068 34628
rect 18028 34000 18068 34040
rect 17836 33664 17876 33704
rect 17932 33076 17972 33116
rect 18316 35260 18356 35300
rect 18124 33832 18164 33872
rect 18124 33580 18164 33620
rect 18028 32908 18068 32948
rect 17836 32740 17876 32780
rect 18124 32488 18164 32528
rect 18316 34924 18356 34964
rect 18604 38200 18644 38240
rect 18988 38872 19028 38912
rect 19468 38872 19508 38912
rect 19564 38704 19604 38744
rect 19948 40720 19988 40760
rect 20121 40468 20161 40508
rect 20048 40048 20088 40088
rect 20130 40048 20170 40088
rect 20212 40048 20252 40088
rect 20294 40048 20334 40088
rect 20376 40048 20416 40088
rect 19948 39712 19988 39752
rect 19756 38620 19796 38660
rect 20812 39544 20852 39584
rect 20716 39376 20756 39416
rect 20140 39208 20180 39248
rect 20044 38956 20084 38996
rect 20620 38956 20660 38996
rect 19943 38704 19983 38744
rect 20044 38704 20084 38744
rect 19852 38536 19892 38576
rect 20048 38536 20088 38576
rect 20130 38536 20170 38576
rect 20212 38536 20252 38576
rect 20294 38536 20334 38576
rect 20376 38536 20416 38576
rect 18892 38368 18932 38408
rect 19276 38368 19316 38408
rect 19468 38368 19508 38408
rect 20236 38368 20276 38408
rect 19084 38284 19124 38324
rect 18892 38200 18932 38240
rect 20140 38284 20180 38324
rect 20524 38284 20564 38324
rect 19468 38200 19508 38240
rect 19564 37948 19604 37988
rect 18808 37780 18848 37820
rect 18890 37780 18930 37820
rect 18972 37780 19012 37820
rect 19054 37780 19094 37820
rect 19136 37780 19176 37820
rect 19276 37780 19316 37820
rect 18796 37612 18836 37652
rect 19852 37780 19892 37820
rect 18988 37528 19028 37568
rect 20044 38200 20084 38240
rect 19948 37696 19988 37736
rect 18892 37360 18932 37400
rect 19084 37360 19124 37400
rect 19276 37360 19316 37400
rect 18700 37276 18740 37316
rect 18796 37108 18836 37148
rect 18604 36688 18644 36728
rect 18988 37192 19028 37232
rect 19084 36940 19124 36980
rect 19564 37276 19604 37316
rect 19564 36940 19604 36980
rect 19468 36856 19508 36896
rect 19660 36772 19700 36812
rect 18892 36604 18932 36644
rect 19276 36604 19316 36644
rect 18796 36520 18836 36560
rect 19276 36352 19316 36392
rect 18808 36268 18848 36308
rect 18890 36268 18930 36308
rect 18972 36268 19012 36308
rect 19054 36268 19094 36308
rect 19136 36268 19176 36308
rect 19180 35848 19220 35888
rect 18700 35428 18740 35468
rect 18508 34756 18548 34796
rect 18508 34588 18548 34628
rect 18412 34504 18452 34544
rect 18412 34252 18452 34292
rect 18316 34000 18356 34040
rect 18808 34756 18848 34796
rect 18890 34756 18930 34796
rect 18972 34756 19012 34796
rect 19054 34756 19094 34796
rect 19136 34756 19176 34796
rect 18700 34504 18740 34544
rect 19084 34420 19124 34460
rect 19372 36184 19412 36224
rect 20620 37780 20660 37820
rect 20034 37360 20074 37400
rect 20140 37276 20180 37316
rect 19948 37108 19988 37148
rect 20048 37024 20088 37064
rect 20130 37024 20170 37064
rect 20212 37024 20252 37064
rect 20294 37024 20334 37064
rect 20376 37024 20416 37064
rect 19948 36688 19988 36728
rect 20140 36688 20180 36728
rect 20044 36520 20084 36560
rect 19756 36436 19796 36476
rect 20620 36100 20660 36140
rect 19468 35848 19508 35888
rect 19468 34924 19508 34964
rect 19372 34840 19412 34880
rect 19372 34672 19412 34712
rect 18796 33664 18836 33704
rect 19276 34336 19316 34376
rect 19852 35764 19892 35804
rect 19756 35596 19796 35636
rect 19660 35512 19700 35552
rect 19756 35176 19796 35216
rect 20524 35848 20564 35888
rect 20044 35764 20084 35804
rect 20048 35512 20088 35552
rect 20130 35512 20170 35552
rect 20212 35512 20252 35552
rect 20294 35512 20334 35552
rect 20376 35512 20416 35552
rect 19948 34924 19988 34964
rect 19852 34672 19892 34712
rect 19756 34420 19796 34460
rect 19660 34336 19700 34376
rect 19948 34504 19988 34544
rect 20048 34000 20088 34040
rect 20130 34000 20170 34040
rect 20212 34000 20252 34040
rect 20294 34000 20334 34040
rect 20376 34000 20416 34040
rect 19948 33916 19988 33956
rect 21388 39292 21428 39332
rect 21388 39040 21428 39080
rect 20908 37696 20948 37736
rect 20812 35848 20852 35888
rect 20812 35680 20852 35720
rect 20716 35512 20756 35552
rect 20620 34504 20660 34544
rect 20812 34000 20852 34040
rect 20524 33748 20564 33788
rect 19468 33496 19508 33536
rect 19852 33580 19892 33620
rect 20044 33412 20084 33452
rect 18700 33244 18740 33284
rect 18808 33244 18848 33284
rect 18890 33244 18930 33284
rect 18972 33244 19012 33284
rect 19054 33244 19094 33284
rect 19136 33244 19176 33284
rect 18604 33160 18644 33200
rect 20044 33160 20084 33200
rect 19276 33076 19316 33116
rect 18604 32824 18644 32864
rect 18316 32740 18356 32780
rect 17452 32152 17492 32192
rect 17356 31060 17396 31100
rect 17164 30976 17204 31016
rect 17836 31900 17876 31940
rect 17644 31228 17684 31268
rect 17260 30052 17300 30092
rect 17740 30724 17780 30764
rect 17836 30640 17876 30680
rect 18604 32572 18644 32612
rect 18412 32320 18452 32360
rect 18028 31564 18068 31604
rect 18028 31228 18068 31268
rect 18124 31144 18164 31184
rect 18124 30808 18164 30848
rect 18124 30472 18164 30512
rect 17068 29884 17108 29924
rect 17452 29800 17492 29840
rect 17740 30220 17780 30260
rect 17548 29716 17588 29756
rect 16972 29380 17012 29420
rect 16876 27700 16916 27740
rect 16588 27616 16628 27656
rect 16780 27616 16820 27656
rect 17068 29296 17108 29336
rect 17164 29212 17204 29252
rect 17452 29128 17492 29168
rect 17260 28288 17300 28328
rect 16300 27196 16340 27236
rect 17452 27616 17492 27656
rect 17356 27448 17396 27488
rect 16012 27112 16052 27152
rect 17260 27112 17300 27152
rect 17644 27868 17684 27908
rect 17836 30052 17876 30092
rect 18028 29632 18068 29672
rect 17836 29548 17876 29588
rect 17836 27952 17876 27992
rect 17932 27868 17972 27908
rect 17740 27532 17780 27572
rect 16204 27028 16244 27068
rect 17452 27028 17492 27068
rect 17740 27028 17780 27068
rect 16012 26356 16052 26396
rect 16012 26188 16052 26228
rect 16108 26104 16148 26144
rect 17644 26944 17684 26984
rect 16780 26860 16820 26900
rect 17548 26860 17588 26900
rect 16492 26440 16532 26480
rect 16972 26776 17012 26816
rect 17068 26608 17108 26648
rect 16588 26272 16628 26312
rect 16876 26272 16916 26312
rect 16687 26188 16727 26228
rect 16780 26020 16820 26060
rect 17260 26776 17300 26816
rect 17164 26524 17204 26564
rect 17164 26356 17204 26396
rect 16492 25348 16532 25388
rect 16108 25264 16148 25304
rect 16204 25096 16244 25136
rect 16108 24508 16148 24548
rect 17164 25684 17204 25724
rect 16780 25348 16820 25388
rect 16492 25180 16532 25220
rect 16684 25096 16724 25136
rect 16492 24592 16532 24632
rect 16012 24004 16052 24044
rect 16588 24508 16628 24548
rect 16012 23668 16052 23708
rect 16204 23584 16244 23624
rect 16588 23500 16628 23540
rect 16300 23164 16340 23204
rect 16108 22240 16148 22280
rect 16012 21904 16052 21944
rect 15436 19972 15476 20012
rect 15724 19216 15764 19256
rect 15340 18460 15380 18500
rect 15628 18880 15668 18920
rect 15532 18460 15572 18500
rect 15436 18376 15476 18416
rect 15340 18292 15380 18332
rect 15244 18040 15284 18080
rect 14956 17956 14996 17996
rect 15916 19804 15956 19844
rect 15148 17788 15188 17828
rect 15820 17788 15860 17828
rect 14860 17536 14900 17576
rect 14572 17116 14612 17156
rect 14668 17032 14708 17072
rect 14572 16192 14612 16232
rect 14572 16024 14612 16064
rect 14092 11992 14132 12032
rect 14092 11488 14132 11528
rect 14092 10396 14132 10436
rect 14092 9892 14132 9932
rect 13804 9220 13844 9260
rect 13708 9136 13748 9176
rect 13612 7792 13652 7832
rect 13516 7288 13556 7328
rect 12844 6616 12884 6656
rect 12556 4936 12596 4976
rect 12748 4936 12788 4976
rect 12460 4852 12500 4892
rect 12460 4600 12500 4640
rect 12364 4516 12404 4556
rect 12748 4768 12788 4808
rect 12556 4432 12596 4472
rect 12748 4096 12788 4136
rect 12460 4012 12500 4052
rect 12172 3844 12212 3884
rect 12652 3508 12692 3548
rect 11788 3424 11828 3464
rect 11788 3088 11828 3128
rect 11884 2752 11924 2792
rect 11788 2584 11828 2624
rect 12940 5944 12980 5984
rect 14092 7456 14132 7496
rect 13708 6448 13748 6488
rect 13612 5776 13652 5816
rect 13036 5440 13076 5480
rect 13516 4936 13556 4976
rect 12940 4768 12980 4808
rect 13420 4684 13460 4724
rect 13324 4348 13364 4388
rect 13036 3508 13076 3548
rect 13324 3508 13364 3548
rect 12844 3256 12884 3296
rect 13516 4348 13556 4388
rect 13708 4684 13748 4724
rect 13996 7036 14036 7076
rect 14092 6952 14132 6992
rect 14284 11656 14324 11696
rect 14764 16864 14804 16904
rect 14764 14596 14804 14636
rect 14956 16864 14996 16904
rect 14956 16360 14996 16400
rect 15244 16024 15284 16064
rect 14956 15604 14996 15644
rect 14956 15268 14996 15308
rect 15052 15100 15092 15140
rect 15244 14008 15284 14048
rect 15244 13336 15284 13376
rect 14476 12076 14516 12116
rect 14860 12244 14900 12284
rect 14476 11908 14516 11948
rect 14476 11656 14516 11696
rect 14572 11488 14612 11528
rect 14476 11320 14516 11360
rect 14380 11152 14420 11192
rect 14572 11236 14612 11276
rect 15052 11824 15092 11864
rect 14764 11488 14804 11528
rect 14284 10900 14324 10940
rect 14668 10900 14708 10940
rect 14476 10816 14516 10856
rect 14380 10648 14420 10688
rect 14380 9472 14420 9512
rect 14380 7456 14420 7496
rect 14284 7372 14324 7412
rect 14668 10732 14708 10772
rect 14668 9976 14708 10016
rect 14572 8716 14612 8756
rect 15052 11068 15092 11108
rect 15820 17032 15860 17072
rect 15724 16360 15764 16400
rect 15724 15940 15764 15980
rect 15724 15772 15764 15812
rect 15532 15436 15572 15476
rect 15532 15268 15572 15308
rect 15628 14512 15668 14552
rect 15532 13840 15572 13880
rect 15436 13672 15476 13712
rect 15436 12580 15476 12620
rect 15340 12412 15380 12452
rect 15820 14260 15860 14300
rect 15724 13756 15764 13796
rect 15628 11824 15668 11864
rect 15532 11656 15572 11696
rect 15244 10984 15284 11024
rect 15052 10144 15092 10184
rect 15340 10396 15380 10436
rect 15148 10060 15188 10100
rect 15340 9976 15380 10016
rect 15244 9892 15284 9932
rect 14956 9724 14996 9764
rect 14764 9472 14804 9512
rect 14860 8716 14900 8756
rect 15148 9472 15188 9512
rect 15052 9388 15092 9428
rect 15244 9304 15284 9344
rect 15052 8716 15092 8756
rect 14764 8044 14804 8084
rect 14668 7876 14708 7916
rect 14572 7708 14612 7748
rect 14764 7456 14804 7496
rect 14284 7122 14285 7160
rect 14285 7122 14324 7160
rect 14284 7120 14324 7122
rect 14476 7204 14516 7244
rect 14476 6952 14516 6992
rect 14092 6448 14132 6488
rect 14284 6196 14324 6236
rect 14188 5776 14228 5816
rect 14092 5440 14132 5480
rect 13996 5020 14036 5060
rect 13900 4936 13940 4976
rect 13804 4348 13844 4388
rect 14092 4348 14132 4388
rect 13900 4264 13940 4304
rect 14188 4264 14228 4304
rect 13505 3844 13545 3884
rect 13804 3508 13844 3548
rect 14092 3928 14132 3968
rect 13996 3844 14036 3884
rect 13804 3256 13844 3296
rect 13516 3004 13556 3044
rect 13036 2752 13076 2792
rect 11692 2248 11732 2288
rect 11692 2080 11732 2120
rect 12172 1996 12212 2036
rect 12172 1744 12212 1784
rect 11788 1660 11828 1700
rect 11980 1660 12020 1700
rect 12556 1240 12596 1280
rect 12748 1240 12788 1280
rect 12460 1072 12500 1112
rect 12364 484 12404 524
rect 12940 1240 12980 1280
rect 12844 1156 12884 1196
rect 13036 316 13076 356
rect 13420 2248 13460 2288
rect 13996 2752 14036 2792
rect 13996 1744 14036 1784
rect 13900 1492 13940 1532
rect 13516 1240 13556 1280
rect 13708 1240 13748 1280
rect 13324 988 13364 1028
rect 14188 3256 14228 3296
rect 14188 3004 14228 3044
rect 14572 5860 14612 5900
rect 14572 5608 14612 5648
rect 14476 4852 14516 4892
rect 14380 4516 14420 4556
rect 14476 4348 14516 4388
rect 14380 3340 14420 3380
rect 14380 2836 14420 2876
rect 14284 1156 14324 1196
rect 14188 988 14228 1028
rect 14284 904 14324 944
rect 14668 3928 14708 3968
rect 14572 3004 14612 3044
rect 14572 2332 14612 2372
rect 14956 7708 14996 7748
rect 15052 7540 15092 7580
rect 15532 9640 15572 9680
rect 15820 13504 15860 13544
rect 16204 21904 16244 21944
rect 16780 23500 16820 23540
rect 17356 26440 17396 26480
rect 17452 26272 17492 26312
rect 17548 26104 17588 26144
rect 17356 26020 17396 26060
rect 17932 26860 17972 26900
rect 17836 26524 17876 26564
rect 17740 26020 17780 26060
rect 17260 25516 17300 25556
rect 17740 25852 17780 25892
rect 17548 25768 17588 25808
rect 17548 25432 17588 25472
rect 17452 25264 17492 25304
rect 17452 25012 17492 25052
rect 17260 24592 17300 24632
rect 16780 22240 16820 22280
rect 16684 21904 16724 21944
rect 16588 21568 16628 21608
rect 16492 20728 16532 20768
rect 16396 20308 16436 20348
rect 16108 18796 16148 18836
rect 16108 18460 16148 18500
rect 16204 18208 16244 18248
rect 16876 21484 16916 21524
rect 16780 21400 16820 21440
rect 17164 22240 17204 22280
rect 17452 23584 17492 23624
rect 17356 22072 17396 22112
rect 17260 21232 17300 21272
rect 17164 21064 17204 21104
rect 17068 20980 17108 21020
rect 17260 20980 17300 21020
rect 17740 25180 17780 25220
rect 18412 31480 18452 31520
rect 19756 32824 19796 32864
rect 19276 32740 19316 32780
rect 18808 31732 18848 31772
rect 18890 31732 18930 31772
rect 18972 31732 19012 31772
rect 19054 31732 19094 31772
rect 19136 31732 19176 31772
rect 19084 31144 19124 31184
rect 18892 31060 18932 31100
rect 19276 31312 19316 31352
rect 19468 32152 19508 32192
rect 20140 32908 20180 32948
rect 20044 32824 20084 32864
rect 20908 32908 20948 32948
rect 20620 32824 20660 32864
rect 20140 32740 20180 32780
rect 20048 32488 20088 32528
rect 20130 32488 20170 32528
rect 20212 32488 20252 32528
rect 20294 32488 20334 32528
rect 20376 32488 20416 32528
rect 19468 31480 19508 31520
rect 19564 31312 19604 31352
rect 19468 31144 19508 31184
rect 19180 30808 19220 30848
rect 18808 30220 18848 30260
rect 18890 30220 18930 30260
rect 18972 30220 19012 30260
rect 19054 30220 19094 30260
rect 19136 30220 19176 30260
rect 19372 30640 19412 30680
rect 19564 30640 19604 30680
rect 18316 29128 18356 29168
rect 18604 29128 18644 29168
rect 19084 29128 19124 29168
rect 19852 32068 19892 32108
rect 20044 31900 20084 31940
rect 20044 31396 20084 31436
rect 19756 30892 19796 30932
rect 20048 30976 20088 31016
rect 20130 30976 20170 31016
rect 20212 30976 20252 31016
rect 20294 30976 20334 31016
rect 20376 30976 20416 31016
rect 19852 30640 19892 30680
rect 20044 30556 20084 30596
rect 20236 29968 20276 30008
rect 18508 28288 18548 28328
rect 18892 28960 18932 29000
rect 18808 28708 18848 28748
rect 18890 28708 18930 28748
rect 18972 28708 19012 28748
rect 19054 28708 19094 28748
rect 19136 28708 19176 28748
rect 18700 28624 18740 28664
rect 18604 27952 18644 27992
rect 18604 27532 18644 27572
rect 18412 27448 18452 27488
rect 18316 27280 18356 27320
rect 18220 26524 18260 26564
rect 18220 25432 18260 25472
rect 18028 25180 18068 25220
rect 18412 26608 18452 26648
rect 18892 27616 18932 27656
rect 19852 28960 19892 29000
rect 19372 28876 19412 28916
rect 19372 28036 19412 28076
rect 19468 27952 19508 27992
rect 19372 27868 19412 27908
rect 19276 27700 19316 27740
rect 19852 28372 19892 28412
rect 20048 29464 20088 29504
rect 20130 29464 20170 29504
rect 20212 29464 20252 29504
rect 20294 29464 20334 29504
rect 20376 29464 20416 29504
rect 21004 32236 21044 32276
rect 20620 31060 20660 31100
rect 20524 28456 20564 28496
rect 20048 27952 20088 27992
rect 20130 27952 20170 27992
rect 20212 27952 20252 27992
rect 20294 27952 20334 27992
rect 20376 27952 20416 27992
rect 19756 27532 19796 27572
rect 19948 27532 19988 27572
rect 18808 27196 18848 27236
rect 18890 27196 18930 27236
rect 18972 27196 19012 27236
rect 19054 27196 19094 27236
rect 19136 27196 19176 27236
rect 19276 27112 19316 27152
rect 20127 27364 20167 27404
rect 20236 27364 20276 27404
rect 18700 27028 18740 27068
rect 19948 27028 19988 27068
rect 18796 26944 18836 26984
rect 18700 26860 18740 26900
rect 18412 26440 18452 26480
rect 18316 25012 18356 25052
rect 18028 24844 18068 24884
rect 17932 24592 17972 24632
rect 17836 24508 17876 24548
rect 17932 23920 17972 23960
rect 17740 23836 17780 23876
rect 17644 23164 17684 23204
rect 17644 22576 17684 22616
rect 17836 23752 17876 23792
rect 17836 23164 17876 23204
rect 18220 24676 18260 24716
rect 18028 23752 18068 23792
rect 18508 26356 18548 26396
rect 18508 25600 18548 25640
rect 19564 26776 19604 26816
rect 19372 26692 19412 26732
rect 18988 26272 19028 26312
rect 18988 26104 19028 26144
rect 18892 25852 18932 25892
rect 19180 25852 19220 25892
rect 18808 25684 18848 25724
rect 18890 25684 18930 25724
rect 18972 25684 19012 25724
rect 19054 25684 19094 25724
rect 19136 25684 19176 25724
rect 18700 25516 18740 25556
rect 18988 25516 19028 25556
rect 18892 25432 18932 25472
rect 19756 26272 19796 26312
rect 18604 24676 18644 24716
rect 18412 23920 18452 23960
rect 18508 23836 18548 23876
rect 18412 23752 18452 23792
rect 18508 23668 18548 23708
rect 18316 23584 18356 23624
rect 18412 23080 18452 23120
rect 18220 22912 18260 22952
rect 18028 22576 18068 22616
rect 17548 21736 17588 21776
rect 17452 21568 17492 21608
rect 18316 22408 18356 22448
rect 18316 22072 18356 22112
rect 17836 21988 17876 22028
rect 18508 22240 18548 22280
rect 18412 21568 18452 21608
rect 19276 25432 19316 25472
rect 19468 25852 19508 25892
rect 19948 26524 19988 26564
rect 20048 26440 20088 26480
rect 20130 26440 20170 26480
rect 20212 26440 20252 26480
rect 20294 26440 20334 26480
rect 20376 26440 20416 26480
rect 19948 26020 19988 26060
rect 19852 25936 19892 25976
rect 20524 25936 20564 25976
rect 19564 25684 19604 25724
rect 19660 25516 19700 25556
rect 19852 25432 19892 25472
rect 20130 25516 20170 25556
rect 19276 25264 19316 25304
rect 19372 25096 19412 25136
rect 19564 25180 19604 25220
rect 18988 24592 19028 24632
rect 19276 24592 19316 24632
rect 19948 25348 19988 25388
rect 20236 25264 20276 25304
rect 20332 25096 20372 25136
rect 20048 24928 20088 24968
rect 20130 24928 20170 24968
rect 20212 24928 20252 24968
rect 20294 24928 20334 24968
rect 20376 24928 20416 24968
rect 19948 24592 19988 24632
rect 19852 24508 19892 24548
rect 20044 24424 20084 24464
rect 18808 24172 18848 24212
rect 18890 24172 18930 24212
rect 18972 24172 19012 24212
rect 19054 24172 19094 24212
rect 19136 24172 19176 24212
rect 20812 27700 20852 27740
rect 20716 27364 20756 27404
rect 19468 23920 19508 23960
rect 20140 23920 20180 23960
rect 19276 23752 19316 23792
rect 19756 23836 19796 23876
rect 19180 23080 19220 23120
rect 18808 22660 18848 22700
rect 18890 22660 18930 22700
rect 18972 22660 19012 22700
rect 19054 22660 19094 22700
rect 19136 22660 19176 22700
rect 19084 22492 19124 22532
rect 18796 22408 18836 22448
rect 18028 21400 18068 21440
rect 18220 21400 18260 21440
rect 17836 21316 17876 21356
rect 17740 21148 17780 21188
rect 17548 20980 17588 21020
rect 17644 20728 17684 20768
rect 17740 20560 17780 20600
rect 17356 20308 17396 20348
rect 17644 20308 17684 20348
rect 16492 20140 16532 20180
rect 16492 19972 16532 20012
rect 16492 17956 16532 17996
rect 16204 17032 16244 17072
rect 16396 17032 16436 17072
rect 16300 16780 16340 16820
rect 16012 16360 16052 16400
rect 16204 16192 16244 16232
rect 16012 15688 16052 15728
rect 16300 16024 16340 16064
rect 16204 14932 16244 14972
rect 16108 14764 16148 14804
rect 16012 14092 16052 14132
rect 15916 12160 15956 12200
rect 15820 11152 15860 11192
rect 16204 14512 16244 14552
rect 16204 13756 16244 13796
rect 15916 10984 15956 11024
rect 15724 10396 15764 10436
rect 16108 11068 16148 11108
rect 16012 10228 16052 10268
rect 15820 9808 15860 9848
rect 15532 9220 15572 9260
rect 15724 9220 15764 9260
rect 15628 8800 15668 8840
rect 15436 8548 15476 8588
rect 15628 8380 15668 8420
rect 15340 7792 15380 7832
rect 15148 7456 15188 7496
rect 15052 6196 15092 6236
rect 15052 5020 15092 5060
rect 15244 5608 15284 5648
rect 14956 4264 14996 4304
rect 14956 3760 14996 3800
rect 14860 3004 14900 3044
rect 14764 2920 14804 2960
rect 15916 9640 15956 9680
rect 15916 8716 15956 8756
rect 15916 8464 15956 8504
rect 15820 6448 15860 6488
rect 16108 9724 16148 9764
rect 16108 8716 16148 8756
rect 16012 8380 16052 8420
rect 16012 8212 16052 8252
rect 15532 6196 15572 6236
rect 15436 5776 15476 5816
rect 15820 5608 15860 5648
rect 15532 5356 15572 5396
rect 15436 5020 15476 5060
rect 15340 3844 15380 3884
rect 15340 3676 15380 3716
rect 15052 3004 15092 3044
rect 15052 2668 15092 2708
rect 14764 1912 14804 1952
rect 15436 3172 15476 3212
rect 15532 2920 15572 2960
rect 14956 2332 14996 2372
rect 14860 1828 14900 1868
rect 14668 1240 14708 1280
rect 14572 904 14612 944
rect 14764 484 14804 524
rect 15436 2080 15476 2120
rect 15052 1912 15092 1952
rect 15820 4600 15860 4640
rect 16396 15184 16436 15224
rect 16780 19636 16820 19676
rect 16684 19384 16724 19424
rect 16780 18628 16820 18668
rect 16780 18040 16820 18080
rect 16684 17956 16724 17996
rect 16780 16612 16820 16652
rect 16972 19972 17012 20012
rect 17260 19804 17300 19844
rect 17932 21064 17972 21104
rect 18508 20812 18548 20852
rect 18028 20728 18068 20768
rect 18028 20392 18068 20432
rect 18316 20728 18356 20768
rect 18220 20476 18260 20516
rect 17644 19636 17684 19676
rect 17356 19552 17396 19592
rect 17740 19468 17780 19508
rect 17644 19300 17684 19340
rect 17260 19216 17300 19256
rect 17068 18880 17108 18920
rect 17260 18712 17300 18752
rect 17068 18628 17108 18668
rect 17153 18460 17193 18500
rect 17260 18460 17300 18500
rect 18124 20140 18164 20180
rect 18124 19216 18164 19256
rect 18412 20140 18452 20180
rect 18316 19804 18356 19844
rect 17932 18880 17972 18920
rect 17644 18796 17684 18836
rect 17836 18796 17876 18836
rect 17740 18712 17780 18752
rect 17452 18460 17492 18500
rect 16972 17368 17012 17408
rect 17068 17116 17108 17156
rect 16972 17032 17012 17072
rect 16876 16528 16916 16568
rect 16684 16360 16724 16400
rect 16588 15184 16628 15224
rect 17260 17788 17300 17828
rect 17644 18544 17684 18584
rect 17836 18460 17876 18500
rect 18028 18460 18068 18500
rect 17644 18292 17684 18332
rect 17260 17368 17300 17408
rect 17356 17284 17396 17324
rect 17356 17116 17396 17156
rect 18028 18040 18068 18080
rect 17740 17956 17780 17996
rect 17740 17536 17780 17576
rect 17260 16780 17300 16820
rect 17164 16276 17204 16316
rect 16780 15436 16820 15476
rect 16684 15016 16724 15056
rect 16492 14848 16532 14888
rect 16780 14848 16820 14888
rect 16396 14596 16436 14636
rect 16684 14596 16724 14636
rect 16588 14512 16628 14552
rect 16396 14260 16436 14300
rect 16396 13756 16436 13796
rect 16588 13672 16628 13712
rect 17356 16612 17396 16652
rect 17644 16444 17684 16484
rect 17164 15268 17204 15308
rect 17068 15184 17108 15224
rect 16972 14008 17012 14048
rect 17164 14092 17204 14132
rect 17548 15940 17588 15980
rect 17356 15520 17396 15560
rect 17452 15100 17492 15140
rect 17356 15016 17396 15056
rect 17260 13840 17300 13880
rect 17068 13756 17108 13796
rect 16780 13252 16820 13292
rect 16492 13168 16532 13208
rect 16588 12496 16628 12536
rect 16396 11152 16436 11192
rect 16300 8632 16340 8672
rect 16204 7960 16244 8000
rect 16108 7372 16148 7412
rect 16108 7204 16148 7244
rect 16108 6784 16148 6824
rect 16300 6952 16340 6992
rect 16204 6616 16244 6656
rect 16108 6448 16148 6488
rect 17164 12664 17204 12704
rect 17260 12580 17300 12620
rect 17452 13924 17492 13964
rect 17452 12664 17492 12704
rect 17164 12412 17204 12452
rect 17356 12412 17396 12452
rect 16780 11656 16820 11696
rect 16780 11488 16820 11528
rect 16972 11488 17012 11528
rect 16972 11320 17012 11360
rect 17068 11152 17108 11192
rect 16492 11068 16532 11108
rect 16876 10900 16916 10940
rect 16588 10732 16628 10772
rect 16972 10480 17012 10520
rect 16588 10396 16628 10436
rect 17452 10732 17492 10772
rect 17164 10564 17204 10604
rect 17260 10396 17300 10436
rect 16492 10060 16532 10100
rect 17068 10144 17108 10184
rect 16588 9640 16628 9680
rect 17452 9976 17492 10016
rect 16780 9640 16820 9680
rect 16684 9472 16724 9512
rect 16972 9388 17012 9428
rect 16492 8548 16532 8588
rect 16492 8296 16532 8336
rect 17164 9472 17204 9512
rect 17836 17116 17876 17156
rect 17932 15604 17972 15644
rect 17836 15520 17876 15560
rect 17740 15268 17780 15308
rect 17740 15100 17780 15140
rect 17836 14932 17876 14972
rect 17644 14512 17684 14552
rect 17644 14344 17684 14384
rect 18412 18880 18452 18920
rect 18412 17704 18452 17744
rect 18988 22072 19028 22112
rect 18892 21568 18932 21608
rect 19948 23584 19988 23624
rect 20048 23416 20088 23456
rect 20130 23416 20170 23456
rect 20212 23416 20252 23456
rect 20294 23416 20334 23456
rect 20376 23416 20416 23456
rect 19660 23164 19700 23204
rect 19372 22744 19412 22784
rect 19564 22660 19604 22700
rect 19564 22324 19604 22364
rect 19948 23080 19988 23120
rect 19756 22744 19796 22784
rect 19852 22660 19892 22700
rect 20236 23080 20276 23120
rect 20140 22996 20180 23036
rect 20044 22660 20084 22700
rect 19564 21568 19604 21608
rect 19852 21736 19892 21776
rect 19276 21400 19316 21440
rect 19468 21400 19508 21440
rect 20236 22072 20276 22112
rect 20048 21904 20088 21944
rect 20130 21904 20170 21944
rect 20212 21904 20252 21944
rect 20294 21904 20334 21944
rect 20376 21904 20416 21944
rect 20140 21736 20180 21776
rect 20044 21652 20084 21692
rect 18808 21148 18848 21188
rect 18890 21148 18930 21188
rect 18972 21148 19012 21188
rect 19054 21148 19094 21188
rect 19136 21148 19176 21188
rect 18892 20728 18932 20768
rect 18988 20560 19028 20600
rect 18892 19972 18932 20012
rect 19084 20056 19124 20096
rect 18988 19888 19028 19928
rect 19084 19804 19124 19844
rect 19564 20728 19604 20768
rect 20140 20560 20180 20600
rect 19276 20056 19316 20096
rect 18808 19636 18848 19676
rect 18890 19636 18930 19676
rect 18972 19636 19012 19676
rect 19054 19636 19094 19676
rect 19136 19636 19176 19676
rect 19468 19636 19508 19676
rect 19756 20224 19796 20264
rect 20048 20392 20088 20432
rect 20130 20392 20170 20432
rect 20212 20392 20252 20432
rect 20294 20392 20334 20432
rect 20376 20392 20416 20432
rect 19852 19804 19892 19844
rect 19660 19636 19700 19676
rect 19564 19300 19604 19340
rect 19852 19384 19892 19424
rect 20140 19384 20180 19424
rect 20044 19216 20084 19256
rect 19468 18796 19508 18836
rect 19276 18712 19316 18752
rect 18796 18460 18836 18500
rect 18892 18292 18932 18332
rect 19372 18292 19412 18332
rect 19276 18208 19316 18248
rect 18808 18124 18848 18164
rect 18890 18124 18930 18164
rect 18972 18124 19012 18164
rect 19054 18124 19094 18164
rect 19136 18124 19176 18164
rect 19180 17956 19220 17996
rect 18700 17620 18740 17660
rect 18700 17032 18740 17072
rect 19180 17032 19220 17072
rect 18124 16948 18164 16988
rect 18808 16612 18848 16652
rect 18890 16612 18930 16652
rect 18972 16612 19012 16652
rect 19054 16612 19094 16652
rect 19136 16612 19176 16652
rect 19084 16444 19124 16484
rect 19660 18040 19700 18080
rect 19468 17956 19508 17996
rect 20048 18880 20088 18920
rect 20130 18880 20170 18920
rect 20212 18880 20252 18920
rect 20294 18880 20334 18920
rect 20376 18880 20416 18920
rect 20044 18712 20084 18752
rect 20236 18712 20276 18752
rect 21292 28876 21332 28916
rect 21100 25684 21140 25724
rect 21004 23920 21044 23960
rect 20812 21904 20852 21944
rect 19372 17032 19412 17072
rect 18988 16192 19028 16232
rect 19180 16360 19220 16400
rect 18700 15856 18740 15896
rect 18412 15688 18452 15728
rect 18700 15688 18740 15728
rect 18124 15436 18164 15476
rect 18316 15268 18356 15308
rect 18124 15016 18164 15056
rect 17836 14008 17876 14048
rect 17932 13840 17972 13880
rect 17740 13420 17780 13460
rect 17740 13252 17780 13292
rect 17740 13000 17780 13040
rect 17740 11488 17780 11528
rect 17644 10648 17684 10688
rect 17447 9640 17487 9680
rect 17548 9640 17588 9680
rect 17644 9472 17684 9512
rect 17452 9220 17492 9260
rect 17068 8800 17108 8840
rect 17260 8800 17300 8840
rect 16876 8632 16916 8672
rect 17452 8716 17492 8756
rect 16684 8044 16724 8084
rect 16492 7540 16532 7580
rect 17356 8632 17396 8672
rect 18220 14680 18260 14720
rect 18508 15016 18548 15056
rect 18508 14764 18548 14804
rect 19276 16024 19316 16064
rect 19084 15688 19124 15728
rect 18988 15520 19028 15560
rect 18796 15436 18836 15476
rect 18700 15268 18740 15308
rect 19084 15268 19124 15308
rect 18604 14680 18644 14720
rect 18808 15100 18848 15140
rect 18890 15100 18930 15140
rect 18972 15100 19012 15140
rect 19054 15100 19094 15140
rect 19136 15100 19176 15140
rect 19756 17032 19796 17072
rect 19756 16780 19796 16820
rect 20048 17368 20088 17408
rect 20130 17368 20170 17408
rect 20212 17368 20252 17408
rect 20294 17368 20334 17408
rect 20376 17368 20416 17408
rect 19948 16444 19988 16484
rect 19468 16276 19508 16316
rect 19468 15688 19508 15728
rect 19468 15520 19508 15560
rect 19468 15268 19508 15308
rect 19372 15184 19412 15224
rect 19660 16192 19700 16232
rect 19756 16024 19796 16064
rect 20044 16024 20084 16064
rect 20716 17956 20756 17996
rect 20620 15940 20660 15980
rect 20048 15856 20088 15896
rect 20130 15856 20170 15896
rect 20212 15856 20252 15896
rect 20294 15856 20334 15896
rect 20376 15856 20416 15896
rect 20044 15688 20084 15728
rect 19948 15268 19988 15308
rect 19660 15184 19700 15224
rect 19852 15184 19892 15224
rect 19372 15016 19412 15056
rect 18892 14848 18932 14888
rect 18412 14596 18452 14636
rect 19084 14764 19124 14804
rect 19276 14680 19316 14720
rect 19468 14932 19508 14972
rect 19660 15016 19700 15056
rect 20236 15016 20276 15056
rect 19564 14848 19604 14888
rect 19564 14512 19604 14552
rect 18124 13420 18164 13460
rect 18028 12580 18068 12620
rect 18028 10732 18068 10772
rect 18028 10144 18068 10184
rect 17932 9640 17972 9680
rect 18412 14428 18452 14468
rect 19084 14428 19124 14468
rect 18220 13168 18260 13208
rect 19276 13840 19316 13880
rect 18808 13588 18848 13628
rect 18890 13588 18930 13628
rect 18972 13588 19012 13628
rect 19054 13588 19094 13628
rect 19136 13588 19176 13628
rect 18604 13420 18644 13460
rect 18892 13420 18932 13460
rect 18988 13336 19028 13376
rect 19180 13336 19220 13376
rect 18988 12664 19028 12704
rect 19084 12580 19124 12620
rect 19276 12496 19316 12536
rect 20044 14848 20084 14888
rect 19852 14764 19892 14804
rect 19948 14680 19988 14720
rect 19756 14596 19796 14636
rect 20044 14596 20084 14636
rect 19948 14428 19988 14468
rect 19660 14092 19700 14132
rect 19852 14008 19892 14048
rect 20048 14344 20088 14384
rect 20130 14344 20170 14384
rect 20212 14344 20252 14384
rect 20294 14344 20334 14384
rect 20376 14344 20416 14384
rect 20140 14092 20180 14132
rect 19468 13840 19508 13880
rect 19468 13168 19508 13208
rect 19276 12244 19316 12284
rect 18808 12076 18848 12116
rect 18890 12076 18930 12116
rect 18972 12076 19012 12116
rect 19054 12076 19094 12116
rect 19136 12076 19176 12116
rect 18700 11992 18740 12032
rect 21196 24760 21236 24800
rect 21196 22408 21236 22448
rect 21388 26608 21428 26648
rect 21388 26440 21428 26480
rect 21388 25768 21428 25808
rect 21388 25432 21428 25472
rect 21388 25096 21428 25136
rect 21388 24928 21428 24968
rect 21100 17368 21140 17408
rect 21388 19720 21428 19760
rect 21388 18880 21428 18920
rect 21196 15352 21236 15392
rect 21196 14344 21236 14384
rect 19948 13840 19988 13880
rect 19852 13336 19892 13376
rect 19852 13000 19892 13040
rect 19468 11908 19508 11948
rect 19084 11824 19124 11864
rect 19468 11656 19508 11696
rect 18796 11572 18836 11612
rect 19372 11488 19412 11528
rect 18412 11152 18452 11192
rect 18700 11152 18740 11192
rect 18508 10984 18548 11024
rect 18220 10060 18260 10100
rect 18316 9472 18356 9512
rect 17836 8800 17876 8840
rect 18028 8800 18068 8840
rect 16972 8548 17012 8588
rect 17260 8296 17300 8336
rect 17164 8128 17204 8168
rect 16972 8044 17012 8084
rect 16876 7960 16916 8000
rect 17068 7960 17108 8000
rect 17932 8464 17972 8504
rect 17836 8380 17876 8420
rect 17452 8296 17492 8336
rect 17644 8296 17684 8336
rect 17548 8128 17588 8168
rect 17644 7960 17684 8000
rect 18604 10900 18644 10940
rect 19852 12664 19892 12704
rect 18988 11236 19028 11276
rect 19180 11236 19220 11276
rect 19180 11068 19220 11108
rect 19084 10816 19124 10856
rect 18808 10564 18848 10604
rect 18890 10564 18930 10604
rect 18972 10564 19012 10604
rect 19054 10564 19094 10604
rect 19136 10564 19176 10604
rect 18796 10396 18836 10436
rect 18700 9472 18740 9512
rect 19084 10144 19124 10184
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 18316 8632 18356 8672
rect 18220 8212 18260 8252
rect 18028 8128 18068 8168
rect 17932 7960 17972 8000
rect 17068 7540 17108 7580
rect 16684 7456 16724 7496
rect 16588 7372 16628 7412
rect 16972 6952 17012 6992
rect 16396 6364 16436 6404
rect 16204 6196 16244 6236
rect 16108 5776 16148 5816
rect 16108 5356 16148 5396
rect 15724 3844 15764 3884
rect 15820 3508 15860 3548
rect 16396 6112 16436 6152
rect 16300 5776 16340 5816
rect 16396 4096 16436 4136
rect 16588 6532 16628 6572
rect 16684 6448 16724 6488
rect 16588 6280 16628 6320
rect 16588 5440 16628 5480
rect 16108 3424 16148 3464
rect 15916 2920 15956 2960
rect 16300 3424 16340 3464
rect 16204 2752 16244 2792
rect 15820 2668 15860 2708
rect 16012 2584 16052 2624
rect 15724 2164 15764 2204
rect 16012 1996 16052 2036
rect 15628 1576 15668 1616
rect 14956 904 14996 944
rect 15436 1240 15476 1280
rect 15628 1240 15668 1280
rect 15244 1072 15284 1112
rect 15244 568 15284 608
rect 15820 316 15860 356
rect 16108 232 16148 272
rect 16588 2836 16628 2876
rect 16972 5104 17012 5144
rect 17644 7708 17684 7748
rect 17548 7204 17588 7244
rect 17548 6700 17588 6740
rect 17548 6532 17588 6572
rect 17260 6448 17300 6488
rect 17164 6028 17204 6068
rect 17164 4936 17204 4976
rect 17164 3844 17204 3884
rect 17452 6448 17492 6488
rect 17356 5104 17396 5144
rect 17356 3760 17396 3800
rect 18220 7624 18260 7664
rect 17932 7288 17972 7328
rect 17644 6112 17684 6152
rect 18028 6532 18068 6572
rect 17836 6448 17876 6488
rect 18028 6112 18068 6152
rect 17932 5776 17972 5816
rect 17836 5692 17876 5732
rect 17836 5440 17876 5480
rect 17836 5104 17876 5144
rect 17740 4936 17780 4976
rect 17740 4180 17780 4220
rect 17740 3844 17780 3884
rect 17644 3760 17684 3800
rect 17836 3760 17876 3800
rect 17644 3592 17684 3632
rect 16876 2416 16916 2456
rect 17068 3172 17108 3212
rect 16588 2080 16628 2120
rect 17164 2080 17204 2120
rect 16492 1744 16532 1784
rect 16972 1912 17012 1952
rect 16492 904 16532 944
rect 16780 904 16820 944
rect 17836 3508 17876 3548
rect 17452 2668 17492 2708
rect 18604 8632 18644 8672
rect 18508 8548 18548 8588
rect 18604 7960 18644 8000
rect 18604 7540 18644 7580
rect 18604 7120 18644 7160
rect 18412 6700 18452 6740
rect 18508 6616 18548 6656
rect 18412 6112 18452 6152
rect 18220 5776 18260 5816
rect 18124 5608 18164 5648
rect 18124 5356 18164 5396
rect 18028 4936 18068 4976
rect 18508 5188 18548 5228
rect 18220 5104 18260 5144
rect 18412 5104 18452 5144
rect 18028 4516 18068 4556
rect 18220 4936 18260 4976
rect 18604 4936 18644 4976
rect 19180 8800 19220 8840
rect 19756 12412 19796 12452
rect 19852 12244 19892 12284
rect 19756 11236 19796 11276
rect 20140 13084 20180 13124
rect 20044 13000 20084 13040
rect 20048 12832 20088 12872
rect 20130 12832 20170 12872
rect 20212 12832 20252 12872
rect 20294 12832 20334 12872
rect 20376 12832 20416 12872
rect 20044 12244 20084 12284
rect 20524 12160 20564 12200
rect 19948 11908 19988 11948
rect 20716 11908 20756 11948
rect 19948 11572 19988 11612
rect 20044 11488 20084 11528
rect 20048 11320 20088 11360
rect 20130 11320 20170 11360
rect 20212 11320 20252 11360
rect 20294 11320 20334 11360
rect 20376 11320 20416 11360
rect 20044 11152 20084 11192
rect 20236 11152 20276 11192
rect 19660 11068 19700 11108
rect 19564 10984 19604 11024
rect 19660 10900 19700 10940
rect 19372 10396 19412 10436
rect 19468 10228 19508 10268
rect 19756 10480 19796 10520
rect 19564 9472 19604 9512
rect 19468 9136 19508 9176
rect 19756 9388 19796 9428
rect 20140 10732 20180 10772
rect 20044 10480 20084 10520
rect 20236 10228 20276 10268
rect 20044 10060 20084 10100
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 19948 9640 19988 9680
rect 19948 9472 19988 9512
rect 20236 9472 20276 9512
rect 19756 8968 19796 9008
rect 19468 8800 19508 8840
rect 19756 8800 19796 8840
rect 19468 8632 19508 8672
rect 19372 8464 19412 8504
rect 19276 8296 19316 8336
rect 18892 8128 18932 8168
rect 19276 8128 19316 8168
rect 18796 8044 18836 8084
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 18892 7288 18932 7328
rect 18988 7204 19028 7244
rect 19084 7120 19124 7160
rect 19180 6280 19220 6320
rect 19084 6196 19124 6236
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 18316 4768 18356 4808
rect 18700 4768 18740 4808
rect 18700 4600 18740 4640
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 19660 8632 19700 8672
rect 19852 8716 19892 8756
rect 20236 9220 20276 9260
rect 20140 9136 20180 9176
rect 20127 8968 20167 9008
rect 20127 8464 20167 8504
rect 20236 8464 20276 8504
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 19852 8044 19892 8084
rect 19468 7960 19508 8000
rect 20140 8128 20180 8168
rect 19660 7540 19700 7580
rect 19468 7456 19508 7496
rect 19660 7372 19700 7412
rect 20140 7372 20180 7412
rect 19564 7036 19604 7076
rect 19468 6868 19508 6908
rect 19660 6868 19700 6908
rect 19468 6532 19508 6572
rect 19564 6448 19604 6488
rect 19948 7120 19988 7160
rect 20236 7120 20276 7160
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 20236 6616 20276 6656
rect 19372 5188 19412 5228
rect 19372 4432 19412 4472
rect 18700 4348 18740 4388
rect 18412 4264 18452 4304
rect 18316 3844 18356 3884
rect 18028 3760 18068 3800
rect 18124 3676 18164 3716
rect 18028 3256 18068 3296
rect 17932 2920 17972 2960
rect 18220 3424 18260 3464
rect 18124 2668 18164 2708
rect 17164 1408 17204 1448
rect 17068 988 17108 1028
rect 16876 652 16916 692
rect 16588 148 16628 188
rect 16780 64 16820 104
rect 18508 4096 18548 4136
rect 19180 4096 19220 4136
rect 18796 3424 18836 3464
rect 19372 3928 19412 3968
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 19084 2584 19124 2624
rect 17932 1912 17972 1952
rect 17356 1660 17396 1700
rect 17452 1576 17492 1616
rect 17548 1240 17588 1280
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 17740 1240 17780 1280
rect 18316 1240 18356 1280
rect 18988 1240 19028 1280
rect 17836 988 17876 1028
rect 17932 400 17972 440
rect 18124 232 18164 272
rect 18508 1156 18548 1196
rect 18700 820 18740 860
rect 18892 820 18932 860
rect 19084 1072 19124 1112
rect 19852 6280 19892 6320
rect 20044 6196 20084 6236
rect 20140 5860 20180 5900
rect 19756 5608 19796 5648
rect 19756 4096 19796 4136
rect 19660 3592 19700 3632
rect 19948 5524 19988 5564
rect 20236 5524 20276 5564
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 20428 4768 20468 4808
rect 19948 4432 19988 4472
rect 20428 4012 20468 4052
rect 19948 3928 19988 3968
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 20044 3592 20084 3632
rect 19756 3508 19796 3548
rect 19852 3340 19892 3380
rect 19660 3256 19700 3296
rect 19660 2920 19700 2960
rect 20140 3340 20180 3380
rect 20236 2836 20276 2876
rect 20044 2752 20084 2792
rect 20140 2584 20180 2624
rect 19660 2080 19700 2120
rect 20620 11068 20660 11108
rect 20812 9556 20852 9596
rect 20716 9472 20756 9512
rect 20620 9220 20660 9260
rect 20716 8464 20756 8504
rect 20620 5524 20660 5564
rect 20524 2332 20564 2372
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 19756 1912 19796 1952
rect 20044 2080 20084 2120
rect 19948 1912 19988 1952
rect 21004 11740 21044 11780
rect 21100 10816 21140 10856
rect 21004 8296 21044 8336
rect 20908 7708 20948 7748
rect 20812 7120 20852 7160
rect 20908 6868 20948 6908
rect 20812 5776 20852 5816
rect 20812 5188 20852 5228
rect 20716 4600 20756 4640
rect 20812 4264 20852 4304
rect 20812 3844 20852 3884
rect 20716 2836 20756 2876
rect 21004 5776 21044 5816
rect 21004 3424 21044 3464
rect 21196 4852 21236 4892
rect 21388 4096 21428 4136
rect 21388 3760 21428 3800
rect 21100 2668 21140 2708
rect 20044 1744 20084 1784
rect 19276 988 19316 1028
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 19276 652 19316 692
rect 19468 484 19508 524
<< metal3 >>
rect 2179 42904 2188 42944
rect 2228 42904 14996 42944
rect 1219 42860 1277 42861
rect 14956 42860 14996 42904
rect 1219 42820 1228 42860
rect 1268 42820 5452 42860
rect 5492 42820 5501 42860
rect 14947 42820 14956 42860
rect 14996 42820 15005 42860
rect 1219 42819 1277 42820
rect 0 42776 80 42796
rect 0 42736 76 42776
rect 116 42736 125 42776
rect 8323 42736 8332 42776
rect 8372 42736 19948 42776
rect 19988 42736 19997 42776
rect 0 42716 80 42736
rect 4771 42692 4829 42693
rect 18499 42692 18557 42693
rect 4771 42652 4780 42692
rect 4820 42652 9676 42692
rect 9716 42652 9725 42692
rect 18499 42652 18508 42692
rect 18548 42652 18892 42692
rect 18932 42652 18941 42692
rect 4771 42651 4829 42652
rect 18499 42651 18557 42652
rect 1603 42568 1612 42608
rect 1652 42568 5068 42608
rect 5108 42568 5117 42608
rect 14563 42568 14572 42608
rect 14612 42568 19468 42608
rect 19508 42568 19517 42608
rect 2467 42484 2476 42524
rect 2516 42484 2764 42524
rect 2804 42484 2813 42524
rect 6691 42484 6700 42524
rect 6740 42484 12364 42524
rect 12404 42484 12413 42524
rect 15235 42484 15244 42524
rect 15284 42484 18892 42524
rect 18932 42484 18941 42524
rect 0 42440 80 42460
rect 0 42400 748 42440
rect 788 42400 797 42440
rect 1891 42400 1900 42440
rect 1940 42400 4108 42440
rect 4148 42400 4157 42440
rect 14371 42400 14380 42440
rect 14420 42400 19276 42440
rect 19316 42400 19325 42440
rect 0 42380 80 42400
rect 10243 42356 10301 42357
rect 3715 42316 3724 42356
rect 3764 42316 10252 42356
rect 10292 42316 10301 42356
rect 14275 42316 14284 42356
rect 14324 42316 17836 42356
rect 17876 42316 17885 42356
rect 10243 42315 10301 42316
rect 2851 42272 2909 42273
rect 15043 42272 15101 42273
rect 1795 42232 1804 42272
rect 1844 42232 2860 42272
rect 2900 42232 2909 42272
rect 9091 42232 9100 42272
rect 9140 42232 11360 42272
rect 2851 42231 2909 42232
rect 4675 42188 4733 42189
rect 10147 42188 10205 42189
rect 4675 42148 4684 42188
rect 4724 42148 9484 42188
rect 9524 42148 9533 42188
rect 10051 42148 10060 42188
rect 10100 42148 10156 42188
rect 10196 42148 10205 42188
rect 11320 42188 11360 42232
rect 15043 42232 15052 42272
rect 15092 42232 17548 42272
rect 17588 42232 17597 42272
rect 17731 42232 17740 42272
rect 17780 42232 18412 42272
rect 18452 42232 18461 42272
rect 15043 42231 15101 42232
rect 11320 42148 11692 42188
rect 11732 42148 11741 42188
rect 16003 42148 16012 42188
rect 16052 42148 19564 42188
rect 19604 42148 19613 42188
rect 4675 42147 4733 42148
rect 10147 42147 10205 42148
rect 0 42104 80 42124
rect 0 42064 268 42104
rect 308 42064 317 42104
rect 9187 42064 9196 42104
rect 9236 42064 11980 42104
rect 12020 42064 12029 42104
rect 15043 42064 15052 42104
rect 15092 42064 18604 42104
rect 18644 42064 18653 42104
rect 0 42044 80 42064
rect 17539 42020 17597 42021
rect 2179 41980 2188 42020
rect 2228 41980 7756 42020
rect 7796 41980 7805 42020
rect 14659 41980 14668 42020
rect 14708 41980 17548 42020
rect 17588 41980 17597 42020
rect 17539 41979 17597 41980
rect 17731 42020 17789 42021
rect 17731 41980 17740 42020
rect 17780 41980 18508 42020
rect 18548 41980 18557 42020
rect 17731 41979 17789 41980
rect 4195 41936 4253 41937
rect 4195 41896 4204 41936
rect 4244 41896 8524 41936
rect 8564 41896 8573 41936
rect 13699 41896 13708 41936
rect 13748 41896 17740 41936
rect 17780 41896 17789 41936
rect 4195 41895 4253 41896
rect 2947 41852 3005 41853
rect 7843 41852 7901 41853
rect 15619 41852 15677 41853
rect 2947 41812 2956 41852
rect 2996 41812 6028 41852
rect 6068 41812 6077 41852
rect 7843 41812 7852 41852
rect 7892 41812 8716 41852
rect 8756 41812 8765 41852
rect 11320 41812 14764 41852
rect 14804 41812 14813 41852
rect 15619 41812 15628 41852
rect 15668 41812 17356 41852
rect 17396 41812 17405 41852
rect 2947 41811 3005 41812
rect 7843 41811 7901 41812
rect 0 41768 80 41788
rect 0 41728 1420 41768
rect 1460 41728 1469 41768
rect 4387 41728 4396 41768
rect 4436 41728 4876 41768
rect 4916 41728 4925 41768
rect 5635 41728 5644 41768
rect 5684 41728 5932 41768
rect 5972 41728 5981 41768
rect 6307 41728 6316 41768
rect 6356 41728 11020 41768
rect 11060 41728 11069 41768
rect 0 41708 80 41728
rect 5443 41644 5452 41684
rect 5492 41644 6796 41684
rect 6836 41644 6845 41684
rect 11320 41600 11360 41812
rect 15619 41811 15677 41812
rect 17827 41768 17885 41769
rect 14083 41728 14092 41768
rect 14132 41728 17260 41768
rect 17300 41728 17309 41768
rect 17827 41728 17836 41768
rect 17876 41728 18316 41768
rect 18356 41728 18365 41768
rect 17827 41727 17885 41728
rect 12163 41684 12221 41685
rect 12163 41644 12172 41684
rect 12212 41644 13132 41684
rect 13172 41644 13181 41684
rect 14467 41644 14476 41684
rect 14516 41644 16876 41684
rect 16916 41644 16925 41684
rect 12163 41643 12221 41644
rect 12547 41600 12605 41601
rect 16771 41600 16829 41601
rect 1507 41560 1516 41600
rect 1556 41560 4492 41600
rect 4532 41560 4541 41600
rect 4919 41560 4928 41600
rect 4968 41560 5010 41600
rect 5050 41560 5092 41600
rect 5132 41560 5174 41600
rect 5214 41560 5256 41600
rect 5296 41560 5305 41600
rect 5827 41560 5836 41600
rect 5876 41560 8140 41600
rect 8180 41560 8189 41600
rect 10348 41560 11308 41600
rect 11348 41560 11360 41600
rect 12462 41560 12556 41600
rect 12596 41560 12605 41600
rect 13315 41560 13324 41600
rect 13364 41560 16588 41600
rect 16628 41560 16637 41600
rect 16686 41560 16780 41600
rect 16820 41560 16829 41600
rect 4579 41476 4588 41516
rect 4628 41476 5356 41516
rect 5396 41476 7276 41516
rect 7316 41476 7325 41516
rect 0 41432 80 41452
rect 1603 41432 1661 41433
rect 0 41392 1612 41432
rect 1652 41392 1661 41432
rect 0 41372 80 41392
rect 1603 41391 1661 41392
rect 2563 41432 2621 41433
rect 6220 41432 6260 41476
rect 9379 41432 9437 41433
rect 2563 41392 2572 41432
rect 2612 41392 5740 41432
rect 5780 41392 5789 41432
rect 6211 41392 6220 41432
rect 6260 41392 6269 41432
rect 6595 41392 6604 41432
rect 6644 41392 7660 41432
rect 7700 41392 7709 41432
rect 9379 41392 9388 41432
rect 9428 41392 10252 41432
rect 10292 41392 10301 41432
rect 2563 41391 2621 41392
rect 9379 41391 9437 41392
rect 2371 41348 2429 41349
rect 10348 41348 10388 41560
rect 12547 41559 12605 41560
rect 16771 41559 16829 41560
rect 16963 41600 17021 41601
rect 18115 41600 18173 41601
rect 16963 41560 16972 41600
rect 17012 41560 17106 41600
rect 18030 41560 18124 41600
rect 18164 41560 18173 41600
rect 20039 41560 20048 41600
rect 20088 41560 20130 41600
rect 20170 41560 20212 41600
rect 20252 41560 20294 41600
rect 20334 41560 20376 41600
rect 20416 41560 20425 41600
rect 16963 41559 17021 41560
rect 18115 41559 18173 41560
rect 10435 41476 10444 41516
rect 10484 41476 10828 41516
rect 10868 41476 10877 41516
rect 13507 41476 13516 41516
rect 13556 41476 17356 41516
rect 17396 41476 17405 41516
rect 17923 41476 17932 41516
rect 17972 41476 18220 41516
rect 18260 41476 18269 41516
rect 13891 41432 13949 41433
rect 2371 41308 2380 41348
rect 2420 41308 6028 41348
rect 6068 41308 6077 41348
rect 7180 41308 10388 41348
rect 10636 41392 12652 41432
rect 12692 41392 12701 41432
rect 13806 41392 13900 41432
rect 13940 41392 13949 41432
rect 2371 41307 2429 41308
rect 3331 41264 3389 41265
rect 3246 41224 3340 41264
rect 3380 41224 3389 41264
rect 3331 41223 3389 41224
rect 4099 41264 4157 41265
rect 4099 41224 4108 41264
rect 4148 41224 6604 41264
rect 6644 41224 6653 41264
rect 4099 41223 4157 41224
rect 1315 41180 1373 41181
rect 1230 41140 1324 41180
rect 1364 41140 1373 41180
rect 1507 41140 1516 41180
rect 1556 41140 3916 41180
rect 3956 41140 3965 41180
rect 1315 41139 1373 41140
rect 0 41096 80 41116
rect 7180 41096 7220 41308
rect 10636 41264 10676 41392
rect 13891 41391 13949 41392
rect 15235 41432 15293 41433
rect 15235 41392 15244 41432
rect 15284 41392 18700 41432
rect 18740 41392 18749 41432
rect 15235 41391 15293 41392
rect 17539 41348 17597 41349
rect 18019 41348 18077 41349
rect 11875 41308 11884 41348
rect 11924 41308 12556 41348
rect 12596 41308 15476 41348
rect 16771 41308 16780 41348
rect 16820 41308 17164 41348
rect 17204 41308 17213 41348
rect 17539 41308 17548 41348
rect 17588 41308 17644 41348
rect 17684 41308 17693 41348
rect 18019 41308 18028 41348
rect 18068 41308 19084 41348
rect 19124 41308 19133 41348
rect 11884 41264 11924 41308
rect 7267 41224 7276 41264
rect 7316 41224 7852 41264
rect 7892 41224 7901 41264
rect 8227 41224 8236 41264
rect 8276 41224 10636 41264
rect 10676 41224 10685 41264
rect 10732 41224 11924 41264
rect 12355 41264 12413 41265
rect 15331 41264 15389 41265
rect 12355 41224 12364 41264
rect 12404 41224 12460 41264
rect 12500 41224 12509 41264
rect 13699 41224 13708 41264
rect 13748 41224 15340 41264
rect 15380 41224 15389 41264
rect 15436 41264 15476 41308
rect 17539 41307 17597 41308
rect 18019 41307 18077 41308
rect 15436 41224 19796 41264
rect 7852 41180 7892 41224
rect 7852 41140 9484 41180
rect 9524 41140 9533 41180
rect 10147 41140 10156 41180
rect 10196 41140 10540 41180
rect 10580 41140 10589 41180
rect 10732 41096 10772 41224
rect 12355 41223 12413 41224
rect 15331 41223 15389 41224
rect 19756 41180 19796 41224
rect 11011 41140 11020 41180
rect 11060 41140 12172 41180
rect 12212 41140 12221 41180
rect 14851 41140 14860 41180
rect 14900 41140 18508 41180
rect 18548 41140 18557 41180
rect 19747 41140 19756 41180
rect 19796 41140 19805 41180
rect 14755 41096 14813 41097
rect 0 41056 7220 41096
rect 9091 41056 9100 41096
rect 9140 41056 10772 41096
rect 14179 41056 14188 41096
rect 14228 41056 14764 41096
rect 14804 41056 14813 41096
rect 14947 41056 14956 41096
rect 14996 41056 19180 41096
rect 19220 41056 19229 41096
rect 0 41036 80 41056
rect 14755 41055 14813 41056
rect 3523 41012 3581 41013
rect 3139 40972 3148 41012
rect 3188 40972 3532 41012
rect 3572 40972 3581 41012
rect 3523 40971 3581 40972
rect 4867 41012 4925 41013
rect 17155 41012 17213 41013
rect 17539 41012 17597 41013
rect 17923 41012 17981 41013
rect 18307 41012 18365 41013
rect 18691 41012 18749 41013
rect 4867 40972 4876 41012
rect 4916 40972 7372 41012
rect 7412 40972 7421 41012
rect 9667 40972 9676 41012
rect 9716 40972 11500 41012
rect 11540 40972 11549 41012
rect 12259 40972 12268 41012
rect 12308 40972 12317 41012
rect 12652 40972 13900 41012
rect 13940 40972 13949 41012
rect 17070 40972 17164 41012
rect 17204 40972 17213 41012
rect 17454 40972 17548 41012
rect 17588 40972 17597 41012
rect 17838 40972 17932 41012
rect 17972 40972 17981 41012
rect 18222 40972 18316 41012
rect 18356 40972 18365 41012
rect 18606 40972 18700 41012
rect 18740 40972 18749 41012
rect 4867 40971 4925 40972
rect 12268 40928 12308 40972
rect 3148 40888 12308 40928
rect 0 40760 80 40780
rect 3148 40760 3188 40888
rect 12652 40844 12692 40972
rect 17155 40971 17213 40972
rect 17539 40971 17597 40972
rect 17923 40971 17981 40972
rect 18307 40971 18365 40972
rect 18691 40971 18749 40972
rect 17635 40928 17693 40929
rect 3679 40804 3688 40844
rect 3728 40804 3770 40844
rect 3810 40804 3852 40844
rect 3892 40804 3934 40844
rect 3974 40804 4016 40844
rect 4056 40804 4065 40844
rect 5539 40804 5548 40844
rect 5588 40804 12692 40844
rect 13228 40888 17644 40928
rect 17684 40888 17693 40928
rect 18115 40888 18124 40928
rect 18164 40888 18604 40928
rect 18644 40888 18653 40928
rect 13228 40760 13268 40888
rect 17635 40887 17693 40888
rect 17251 40844 17309 40845
rect 16963 40804 16972 40844
rect 17012 40804 17260 40844
rect 17300 40804 17309 40844
rect 18799 40804 18808 40844
rect 18848 40804 18890 40844
rect 18930 40804 18972 40844
rect 19012 40804 19054 40844
rect 19094 40804 19136 40844
rect 19176 40804 19185 40844
rect 17251 40803 17309 40804
rect 14563 40760 14621 40761
rect 0 40720 2540 40760
rect 3139 40720 3148 40760
rect 3188 40720 3197 40760
rect 3244 40720 4148 40760
rect 4483 40720 4492 40760
rect 4532 40720 4972 40760
rect 5012 40720 8180 40760
rect 10147 40720 10156 40760
rect 10196 40720 13268 40760
rect 14478 40720 14572 40760
rect 14612 40720 14621 40760
rect 16675 40720 16684 40760
rect 16724 40720 19948 40760
rect 19988 40720 19997 40760
rect 0 40700 80 40720
rect 2500 40676 2540 40720
rect 3244 40676 3284 40720
rect 4108 40676 4148 40720
rect 8140 40676 8180 40720
rect 14563 40719 14621 40720
rect 14371 40676 14429 40677
rect 2500 40636 3284 40676
rect 3331 40636 3340 40676
rect 3380 40636 3532 40676
rect 3572 40636 3581 40676
rect 4099 40636 4108 40676
rect 4148 40636 4157 40676
rect 4588 40636 7564 40676
rect 7604 40636 7613 40676
rect 8131 40636 8140 40676
rect 8180 40636 13036 40676
rect 13076 40636 13085 40676
rect 14275 40636 14284 40676
rect 14324 40636 14380 40676
rect 14420 40636 14429 40676
rect 15811 40636 15820 40676
rect 15860 40636 18796 40676
rect 18836 40636 18845 40676
rect 18979 40636 18988 40676
rect 19028 40636 19037 40676
rect 4588 40592 4628 40636
rect 14371 40635 14429 40636
rect 14755 40592 14813 40593
rect 17059 40592 17117 40593
rect 17539 40592 17597 40593
rect 17923 40592 17981 40593
rect 18988 40592 19028 40636
rect 2083 40552 2092 40592
rect 2132 40552 4628 40592
rect 4684 40552 5068 40592
rect 5108 40552 5117 40592
rect 8035 40552 8044 40592
rect 8084 40552 9580 40592
rect 9620 40552 9629 40592
rect 9676 40552 14572 40592
rect 14612 40552 14621 40592
rect 14755 40552 14764 40592
rect 14804 40552 16628 40592
rect 1411 40508 1469 40509
rect 4684 40508 4724 40552
rect 5635 40508 5693 40509
rect 9676 40508 9716 40552
rect 14755 40551 14813 40552
rect 1326 40468 1420 40508
rect 1460 40468 1469 40508
rect 3523 40468 3532 40508
rect 3572 40468 4724 40508
rect 5550 40468 5644 40508
rect 5684 40468 5693 40508
rect 6979 40468 6988 40508
rect 7028 40468 7756 40508
rect 7796 40468 7805 40508
rect 8323 40468 8332 40508
rect 8372 40468 9716 40508
rect 10723 40508 10781 40509
rect 16588 40508 16628 40552
rect 17059 40552 17068 40592
rect 17108 40552 17164 40592
rect 17204 40552 17213 40592
rect 17454 40552 17548 40592
rect 17588 40552 17597 40592
rect 17838 40552 17932 40592
rect 17972 40552 17981 40592
rect 17059 40551 17117 40552
rect 17539 40551 17597 40552
rect 17923 40551 17981 40552
rect 18028 40552 19028 40592
rect 18028 40508 18068 40552
rect 18595 40508 18653 40509
rect 10723 40468 10732 40508
rect 10772 40468 10866 40508
rect 16588 40468 18068 40508
rect 18510 40468 18604 40508
rect 18644 40468 18653 40508
rect 1411 40467 1469 40468
rect 5635 40467 5693 40468
rect 10723 40467 10781 40468
rect 18595 40467 18653 40468
rect 18700 40468 20121 40508
rect 20161 40468 20170 40508
rect 0 40424 80 40444
rect 1795 40424 1853 40425
rect 0 40384 364 40424
rect 404 40384 413 40424
rect 1795 40384 1804 40424
rect 1844 40384 2284 40424
rect 2324 40384 2333 40424
rect 3427 40384 3436 40424
rect 3476 40384 3485 40424
rect 6403 40384 6412 40424
rect 6452 40384 9964 40424
rect 10004 40384 10013 40424
rect 10434 40398 10443 40438
rect 10483 40425 10492 40438
rect 10483 40424 10493 40425
rect 16387 40424 16445 40425
rect 18700 40424 18740 40468
rect 10435 40384 10444 40398
rect 10484 40384 10564 40424
rect 11683 40384 11692 40424
rect 11732 40384 11741 40424
rect 13603 40384 13612 40424
rect 13652 40384 13900 40424
rect 13940 40384 13949 40424
rect 14947 40384 14956 40424
rect 14996 40384 15628 40424
rect 15668 40384 15677 40424
rect 16387 40384 16396 40424
rect 16436 40384 18740 40424
rect 18883 40424 18941 40425
rect 19747 40424 19805 40425
rect 18883 40384 18892 40424
rect 18932 40384 19756 40424
rect 19796 40384 19805 40424
rect 0 40364 80 40384
rect 1795 40383 1853 40384
rect 1027 40340 1085 40341
rect 3436 40340 3476 40384
rect 10435 40383 10493 40384
rect 7267 40340 7325 40341
rect 11587 40340 11645 40341
rect 1027 40300 1036 40340
rect 1076 40300 1900 40340
rect 1940 40300 1949 40340
rect 2083 40300 2092 40340
rect 2132 40300 3476 40340
rect 3724 40300 3916 40340
rect 3956 40300 3965 40340
rect 5347 40300 5356 40340
rect 5396 40300 6988 40340
rect 7028 40300 7037 40340
rect 7267 40300 7276 40340
rect 7316 40300 7410 40340
rect 9091 40300 9100 40340
rect 9140 40300 9292 40340
rect 9332 40300 9341 40340
rect 9475 40300 9484 40340
rect 9524 40300 10732 40340
rect 10772 40300 10781 40340
rect 11320 40300 11596 40340
rect 11636 40300 11645 40340
rect 1027 40299 1085 40300
rect 1891 40256 1949 40257
rect 3427 40256 3485 40257
rect 3724 40256 3764 40300
rect 7267 40299 7325 40300
rect 4867 40256 4925 40257
rect 11320 40256 11360 40300
rect 11587 40299 11645 40300
rect 11692 40256 11732 40384
rect 16387 40383 16445 40384
rect 18883 40383 18941 40384
rect 19747 40383 19805 40384
rect 20611 40340 20669 40341
rect 12643 40300 12652 40340
rect 12692 40300 13460 40340
rect 13507 40300 13516 40340
rect 13556 40300 14092 40340
rect 14132 40300 14804 40340
rect 1891 40216 1900 40256
rect 1940 40216 2540 40256
rect 1891 40215 1949 40216
rect 1411 40172 1469 40173
rect 2500 40172 2540 40216
rect 3427 40216 3436 40256
rect 3476 40216 3764 40256
rect 3820 40216 4492 40256
rect 4532 40216 4541 40256
rect 4675 40216 4684 40256
rect 4724 40216 4876 40256
rect 4916 40216 4925 40256
rect 7363 40216 7372 40256
rect 7412 40216 11360 40256
rect 11491 40216 11500 40256
rect 11540 40216 11732 40256
rect 13420 40256 13460 40300
rect 14764 40256 14804 40300
rect 15148 40300 16684 40340
rect 16724 40300 16733 40340
rect 17155 40300 17164 40340
rect 17204 40300 19180 40340
rect 19220 40300 19229 40340
rect 19363 40300 19372 40340
rect 19412 40300 20620 40340
rect 20660 40300 20669 40340
rect 13420 40216 13804 40256
rect 13844 40216 13853 40256
rect 14275 40216 14284 40256
rect 14324 40216 14572 40256
rect 14612 40216 14621 40256
rect 14755 40216 14764 40256
rect 14804 40216 14813 40256
rect 3427 40215 3485 40216
rect 3820 40172 3860 40216
rect 4867 40215 4925 40216
rect 7363 40172 7421 40173
rect 10051 40172 10109 40173
rect 15148 40172 15188 40300
rect 20611 40299 20669 40300
rect 19459 40256 19517 40257
rect 15235 40216 15244 40256
rect 15284 40216 18604 40256
rect 18644 40216 18653 40256
rect 19459 40216 19468 40256
rect 19508 40216 19660 40256
rect 19700 40216 19709 40256
rect 19459 40215 19517 40216
rect 1411 40132 1420 40172
rect 1460 40132 1996 40172
rect 2036 40132 2045 40172
rect 2500 40132 3860 40172
rect 3907 40132 3916 40172
rect 3956 40132 5396 40172
rect 1411 40131 1469 40132
rect 0 40088 80 40108
rect 3427 40088 3485 40089
rect 4291 40088 4349 40089
rect 5356 40088 5396 40132
rect 7363 40132 7372 40172
rect 7412 40132 9676 40172
rect 9716 40132 9725 40172
rect 9966 40132 10060 40172
rect 10100 40132 10109 40172
rect 11011 40132 11020 40172
rect 11060 40132 15188 40172
rect 17251 40132 17260 40172
rect 17300 40132 20852 40172
rect 7363 40131 7421 40132
rect 10051 40131 10109 40132
rect 8323 40088 8381 40089
rect 10915 40088 10973 40089
rect 14275 40088 14333 40089
rect 16675 40088 16733 40089
rect 18499 40088 18557 40089
rect 20812 40088 20852 40132
rect 21424 40088 21504 40108
rect 0 40048 3436 40088
rect 3476 40048 3485 40088
rect 4206 40048 4300 40088
rect 4340 40048 4349 40088
rect 4919 40048 4928 40088
rect 4968 40048 5010 40088
rect 5050 40048 5092 40088
rect 5132 40048 5174 40088
rect 5214 40048 5256 40088
rect 5296 40048 5305 40088
rect 5356 40048 7276 40088
rect 7316 40048 7325 40088
rect 7843 40048 7852 40088
rect 7892 40048 8332 40088
rect 8372 40048 10348 40088
rect 10388 40048 10397 40088
rect 10915 40048 10924 40088
rect 10964 40048 11212 40088
rect 11252 40048 11261 40088
rect 11320 40048 14284 40088
rect 14324 40048 15148 40088
rect 15188 40048 15197 40088
rect 15244 40048 16396 40088
rect 16436 40048 16445 40088
rect 16675 40048 16684 40088
rect 16724 40048 18508 40088
rect 18548 40048 18557 40088
rect 20039 40048 20048 40088
rect 20088 40048 20130 40088
rect 20170 40048 20212 40088
rect 20252 40048 20294 40088
rect 20334 40048 20376 40088
rect 20416 40048 20425 40088
rect 20812 40048 21504 40088
rect 0 40028 80 40048
rect 3427 40047 3485 40048
rect 4291 40047 4349 40048
rect 8323 40047 8381 40048
rect 10915 40047 10973 40048
rect 11320 40004 11360 40048
rect 14275 40047 14333 40048
rect 2659 39964 2668 40004
rect 2708 39964 11360 40004
rect 12451 40004 12509 40005
rect 15244 40004 15284 40048
rect 16675 40047 16733 40048
rect 18499 40047 18557 40048
rect 21424 40028 21504 40048
rect 12451 39964 12460 40004
rect 12500 39964 15284 40004
rect 16291 39964 16300 40004
rect 16340 39964 18028 40004
rect 18068 39964 18077 40004
rect 12451 39963 12509 39964
rect 16579 39920 16637 39921
rect 4972 39880 7604 39920
rect 7843 39880 7852 39920
rect 7892 39880 8524 39920
rect 8564 39880 8573 39920
rect 9283 39880 9292 39920
rect 9332 39880 9484 39920
rect 9524 39880 9533 39920
rect 9667 39880 9676 39920
rect 9716 39880 10156 39920
rect 10196 39880 10205 39920
rect 10339 39880 10348 39920
rect 10388 39880 10540 39920
rect 10580 39880 10589 39920
rect 11320 39880 11404 39920
rect 11444 39880 11453 39920
rect 13987 39880 13996 39920
rect 14036 39880 15340 39920
rect 15380 39880 15389 39920
rect 16579 39880 16588 39920
rect 16628 39880 16780 39920
rect 16820 39880 16829 39920
rect 17827 39880 17836 39920
rect 17876 39880 19276 39920
rect 19316 39880 19325 39920
rect 3619 39836 3677 39837
rect 3523 39796 3532 39836
rect 3572 39796 3628 39836
rect 3668 39796 3677 39836
rect 3619 39795 3677 39796
rect 0 39752 80 39772
rect 1699 39752 1757 39753
rect 4972 39752 5012 39880
rect 5068 39796 6220 39836
rect 6260 39796 6269 39836
rect 5068 39752 5108 39796
rect 6211 39752 6269 39753
rect 7564 39752 7604 39880
rect 11320 39836 11360 39880
rect 16579 39879 16637 39880
rect 7651 39796 7660 39836
rect 7700 39796 9964 39836
rect 10004 39796 11360 39836
rect 11587 39836 11645 39837
rect 17827 39836 17885 39837
rect 11587 39796 11596 39836
rect 11636 39796 17836 39836
rect 17876 39796 17885 39836
rect 11587 39795 11645 39796
rect 17827 39795 17885 39796
rect 12931 39752 12989 39753
rect 15907 39752 15965 39753
rect 16867 39752 16925 39753
rect 18499 39752 18557 39753
rect 0 39712 1708 39752
rect 1748 39712 1757 39752
rect 2083 39712 2092 39752
rect 2132 39712 5012 39752
rect 5059 39712 5068 39752
rect 5108 39712 5117 39752
rect 5731 39712 5740 39752
rect 5780 39712 6220 39752
rect 6260 39712 6269 39752
rect 6979 39712 6988 39752
rect 7028 39712 7180 39752
rect 7220 39712 7229 39752
rect 7564 39712 9100 39752
rect 9140 39712 9149 39752
rect 10051 39712 10060 39752
rect 10100 39712 10109 39752
rect 11395 39712 11404 39752
rect 11444 39712 12940 39752
rect 12980 39712 12989 39752
rect 13699 39712 13708 39752
rect 13748 39712 14380 39752
rect 14420 39712 14860 39752
rect 14900 39712 15052 39752
rect 15092 39712 15101 39752
rect 15907 39712 15916 39752
rect 15956 39712 16204 39752
rect 16244 39712 16253 39752
rect 16867 39712 16876 39752
rect 16916 39712 17164 39752
rect 17204 39712 17213 39752
rect 18499 39712 18508 39752
rect 18548 39712 19948 39752
rect 19988 39712 19997 39752
rect 0 39692 80 39712
rect 1699 39711 1757 39712
rect 6211 39711 6269 39712
rect 3139 39668 3197 39669
rect 4483 39668 4541 39669
rect 163 39628 172 39668
rect 212 39628 2668 39668
rect 2708 39628 2717 39668
rect 3139 39628 3148 39668
rect 3188 39628 3724 39668
rect 3764 39628 3773 39668
rect 4398 39628 4492 39668
rect 4532 39628 4541 39668
rect 3139 39627 3197 39628
rect 4483 39627 4541 39628
rect 4675 39668 4733 39669
rect 5731 39668 5789 39669
rect 6115 39668 6173 39669
rect 10060 39668 10100 39712
rect 12931 39711 12989 39712
rect 15907 39711 15965 39712
rect 16867 39711 16925 39712
rect 18499 39711 18557 39712
rect 13891 39668 13949 39669
rect 16579 39668 16637 39669
rect 18211 39668 18269 39669
rect 4675 39628 4684 39668
rect 4724 39628 4818 39668
rect 4867 39628 4876 39668
rect 4916 39628 5740 39668
rect 5780 39628 5789 39668
rect 6030 39628 6124 39668
rect 6164 39628 6173 39668
rect 4675 39627 4733 39628
rect 5731 39627 5789 39628
rect 6115 39627 6173 39628
rect 6220 39628 9292 39668
rect 9332 39628 9341 39668
rect 10060 39628 13324 39668
rect 13364 39628 13373 39668
rect 13891 39628 13900 39668
rect 13940 39628 15724 39668
rect 15764 39628 15773 39668
rect 16494 39628 16588 39668
rect 16628 39628 16637 39668
rect 18126 39628 18220 39668
rect 18260 39628 18269 39668
rect 19171 39628 19180 39668
rect 19220 39628 19229 39668
rect 6220 39584 6260 39628
rect 13891 39627 13949 39628
rect 16579 39627 16637 39628
rect 18211 39627 18269 39628
rect 14755 39584 14813 39585
rect 19180 39584 19220 39628
rect 21424 39584 21504 39604
rect 2500 39544 6260 39584
rect 8227 39544 8236 39584
rect 8276 39544 11980 39584
rect 12020 39544 12556 39584
rect 12596 39544 12605 39584
rect 12940 39544 13420 39584
rect 13460 39544 14188 39584
rect 14228 39544 14764 39584
rect 14804 39544 14813 39584
rect 1219 39460 1228 39500
rect 1268 39460 2092 39500
rect 2132 39460 2141 39500
rect 0 39416 80 39436
rect 2500 39416 2540 39544
rect 9859 39500 9917 39501
rect 12940 39500 12980 39544
rect 14755 39543 14813 39544
rect 15148 39544 19220 39584
rect 20803 39544 20812 39584
rect 20852 39544 21504 39584
rect 14563 39500 14621 39501
rect 15148 39500 15188 39544
rect 21424 39524 21504 39544
rect 16099 39500 16157 39501
rect 18403 39500 18461 39501
rect 19363 39500 19421 39501
rect 2668 39460 4244 39500
rect 5251 39460 5260 39500
rect 5300 39460 7988 39500
rect 9667 39460 9676 39500
rect 9716 39460 9725 39500
rect 9859 39460 9868 39500
rect 9908 39460 10002 39500
rect 10339 39460 10348 39500
rect 10388 39460 11360 39500
rect 12931 39460 12940 39500
rect 12980 39460 12989 39500
rect 14083 39460 14092 39500
rect 14132 39460 14572 39500
rect 14612 39460 14621 39500
rect 14755 39460 14764 39500
rect 14804 39460 15188 39500
rect 15523 39460 15532 39500
rect 15572 39460 16108 39500
rect 16148 39460 16157 39500
rect 18318 39460 18412 39500
rect 18452 39460 18461 39500
rect 18979 39460 18988 39500
rect 19028 39460 19372 39500
rect 19412 39460 19421 39500
rect 2668 39416 2708 39460
rect 4204 39416 4244 39460
rect 7171 39416 7229 39417
rect 0 39376 1556 39416
rect 1603 39376 1612 39416
rect 1652 39376 2540 39416
rect 2659 39376 2668 39416
rect 2708 39376 2717 39416
rect 3532 39376 4148 39416
rect 4204 39376 7180 39416
rect 7220 39376 7229 39416
rect 7948 39416 7988 39460
rect 9676 39416 9716 39460
rect 9859 39459 9917 39460
rect 11320 39416 11360 39460
rect 14563 39459 14621 39460
rect 16099 39459 16157 39460
rect 18403 39459 18461 39460
rect 19363 39459 19421 39460
rect 7948 39376 8428 39416
rect 8468 39376 8477 39416
rect 9676 39376 11116 39416
rect 11156 39376 11165 39416
rect 11320 39376 20716 39416
rect 20756 39376 20765 39416
rect 0 39356 80 39376
rect 1516 39332 1556 39376
rect 1987 39332 2045 39333
rect 3532 39332 3572 39376
rect 4108 39332 4148 39376
rect 7171 39375 7229 39376
rect 11491 39332 11549 39333
rect 19267 39332 19325 39333
rect 1516 39292 1996 39332
rect 2036 39292 3572 39332
rect 3679 39292 3688 39332
rect 3728 39292 3770 39332
rect 3810 39292 3852 39332
rect 3892 39292 3934 39332
rect 3974 39292 4016 39332
rect 4056 39292 4065 39332
rect 4108 39292 8140 39332
rect 8180 39292 8189 39332
rect 9091 39292 9100 39332
rect 9140 39292 9868 39332
rect 9908 39292 9917 39332
rect 10732 39292 11360 39332
rect 1987 39291 2045 39292
rect 1699 39248 1757 39249
rect 6019 39248 6077 39249
rect 10627 39248 10685 39249
rect 1614 39208 1708 39248
rect 1748 39208 1757 39248
rect 1699 39207 1757 39208
rect 2500 39208 5836 39248
rect 5876 39208 5885 39248
rect 6019 39208 6028 39248
rect 6068 39208 6220 39248
rect 6260 39208 6269 39248
rect 6700 39208 10636 39248
rect 10676 39208 10685 39248
rect 1891 39164 1949 39165
rect 1516 39124 1900 39164
rect 1940 39124 1949 39164
rect 0 39080 80 39100
rect 1516 39080 1556 39124
rect 1891 39123 1949 39124
rect 0 39040 1556 39080
rect 2083 39080 2141 39081
rect 2500 39080 2540 39208
rect 6019 39207 6077 39208
rect 2755 39164 2813 39165
rect 3043 39164 3101 39165
rect 4003 39164 4061 39165
rect 6700 39164 6740 39208
rect 10627 39207 10685 39208
rect 10732 39164 10772 39292
rect 11107 39248 11165 39249
rect 2670 39124 2764 39164
rect 2804 39124 2813 39164
rect 2947 39124 2956 39164
rect 2996 39124 3052 39164
rect 3092 39124 3101 39164
rect 3918 39124 4012 39164
rect 4052 39124 4061 39164
rect 4195 39124 4204 39164
rect 4244 39124 4588 39164
rect 4628 39124 4637 39164
rect 5347 39124 5356 39164
rect 5396 39124 6740 39164
rect 6787 39124 6796 39164
rect 6836 39124 10772 39164
rect 10828 39208 10924 39248
rect 10964 39208 10973 39248
rect 11107 39208 11116 39248
rect 11156 39208 11212 39248
rect 11252 39208 11261 39248
rect 2755 39123 2813 39124
rect 3043 39123 3101 39124
rect 4003 39123 4061 39124
rect 3331 39080 3389 39081
rect 4291 39080 4349 39081
rect 7267 39080 7325 39081
rect 10828 39080 10868 39208
rect 11107 39207 11165 39208
rect 11320 39164 11360 39292
rect 11491 39292 11500 39332
rect 11540 39292 12980 39332
rect 13027 39292 13036 39332
rect 13076 39292 14380 39332
rect 14420 39292 14429 39332
rect 16291 39292 16300 39332
rect 16340 39292 18700 39332
rect 18740 39292 18749 39332
rect 18799 39292 18808 39332
rect 18848 39292 18890 39332
rect 18930 39292 18972 39332
rect 19012 39292 19054 39332
rect 19094 39292 19136 39332
rect 19176 39292 19185 39332
rect 19267 39292 19276 39332
rect 19316 39292 21388 39332
rect 21428 39292 21437 39332
rect 11491 39291 11549 39292
rect 12835 39248 12893 39249
rect 12750 39208 12844 39248
rect 12884 39208 12893 39248
rect 12940 39248 12980 39292
rect 19267 39291 19325 39292
rect 18115 39248 18173 39249
rect 18403 39248 18461 39249
rect 12940 39208 18124 39248
rect 18164 39208 18173 39248
rect 18318 39208 18412 39248
rect 18452 39208 18461 39248
rect 18595 39208 18604 39248
rect 18644 39208 20140 39248
rect 20180 39208 20189 39248
rect 12835 39207 12893 39208
rect 18115 39207 18173 39208
rect 18403 39207 18461 39208
rect 11320 39124 19564 39164
rect 19604 39124 19613 39164
rect 15811 39080 15869 39081
rect 17923 39080 17981 39081
rect 19267 39080 19325 39081
rect 19555 39080 19613 39081
rect 20995 39080 21053 39081
rect 21424 39080 21504 39100
rect 2083 39040 2092 39080
rect 2132 39040 2540 39080
rect 3139 39040 3148 39080
rect 3188 39040 3340 39080
rect 3380 39040 3628 39080
rect 3668 39040 3677 39080
rect 4099 39040 4108 39080
rect 4148 39040 4300 39080
rect 4340 39040 4349 39080
rect 7171 39040 7180 39080
rect 7220 39040 7276 39080
rect 7316 39040 7325 39080
rect 8035 39040 8044 39080
rect 8084 39040 8716 39080
rect 8756 39040 10868 39080
rect 10915 39040 10924 39080
rect 10964 39040 11212 39080
rect 11252 39040 14572 39080
rect 14612 39040 14621 39080
rect 15811 39040 15820 39080
rect 15860 39040 16012 39080
rect 16052 39040 17548 39080
rect 17588 39040 17597 39080
rect 17923 39040 17932 39080
rect 17972 39040 19276 39080
rect 19316 39040 19325 39080
rect 19459 39040 19468 39080
rect 19508 39040 19564 39080
rect 19604 39040 19613 39080
rect 0 39020 80 39040
rect 2083 39039 2141 39040
rect 3331 39039 3389 39040
rect 4291 39039 4349 39040
rect 7267 39039 7325 39040
rect 547 38996 605 38997
rect 2371 38996 2429 38997
rect 4099 38996 4157 38997
rect 547 38956 556 38996
rect 596 38956 1996 38996
rect 2036 38956 2045 38996
rect 2286 38956 2380 38996
rect 2420 38956 2429 38996
rect 547 38955 605 38956
rect 2371 38955 2429 38956
rect 2500 38956 3532 38996
rect 3572 38956 4108 38996
rect 4148 38956 4157 38996
rect 1507 38872 1516 38912
rect 1556 38872 1708 38912
rect 1748 38872 1757 38912
rect 0 38744 80 38764
rect 1123 38744 1181 38745
rect 2500 38744 2540 38956
rect 4099 38955 4157 38956
rect 6691 38996 6749 38997
rect 8035 38996 8093 38997
rect 6691 38956 6700 38996
rect 6740 38956 8044 38996
rect 8084 38956 8093 38996
rect 6691 38955 6749 38956
rect 8035 38955 8093 38956
rect 8227 38996 8285 38997
rect 10243 38996 10301 38997
rect 10828 38996 10868 39040
rect 15811 39039 15869 39040
rect 17923 39039 17981 39040
rect 19267 39039 19325 39040
rect 19555 39039 19613 39040
rect 19756 39040 21004 39080
rect 21044 39040 21053 39080
rect 21379 39040 21388 39080
rect 21428 39040 21504 39080
rect 11011 38996 11069 38997
rect 8227 38956 8236 38996
rect 8276 38956 8370 38996
rect 9475 38956 9484 38996
rect 9524 38956 9533 38996
rect 10243 38956 10252 38996
rect 10292 38956 10444 38996
rect 10484 38956 10493 38996
rect 10828 38956 11020 38996
rect 11060 38956 11069 38996
rect 8227 38955 8285 38956
rect 6403 38912 6461 38913
rect 8611 38912 8669 38913
rect 9484 38912 9524 38956
rect 10243 38955 10301 38956
rect 11011 38955 11069 38956
rect 11203 38996 11261 38997
rect 14851 38996 14909 38997
rect 17251 38996 17309 38997
rect 19756 38996 19796 39040
rect 20995 39039 21053 39040
rect 21424 39020 21504 39040
rect 11203 38956 11212 38996
rect 11252 38956 13036 38996
rect 13076 38956 13085 38996
rect 14851 38956 14860 38996
rect 14900 38956 17260 38996
rect 17300 38956 19084 38996
rect 19124 38956 19133 38996
rect 19267 38956 19276 38996
rect 19316 38956 19796 38996
rect 20035 38956 20044 38996
rect 20084 38956 20620 38996
rect 20660 38956 20669 38996
rect 11203 38955 11261 38956
rect 14851 38955 14909 38956
rect 17251 38955 17309 38956
rect 3148 38872 3340 38912
rect 3380 38872 3389 38912
rect 3820 38872 4108 38912
rect 4148 38872 4157 38912
rect 4483 38872 4492 38912
rect 4532 38872 6412 38912
rect 6452 38872 6461 38912
rect 7459 38872 7468 38912
rect 7508 38872 8140 38912
rect 8180 38872 8189 38912
rect 8526 38872 8620 38912
rect 8660 38872 8669 38912
rect 8995 38872 9004 38912
rect 9044 38872 10252 38912
rect 10292 38872 10301 38912
rect 11875 38872 11884 38912
rect 11924 38872 12172 38912
rect 12212 38872 13132 38912
rect 13172 38872 13181 38912
rect 15043 38872 15052 38912
rect 15092 38872 15628 38912
rect 15668 38872 15677 38912
rect 18412 38872 18604 38912
rect 18644 38872 18653 38912
rect 18979 38872 18988 38912
rect 19028 38872 19468 38912
rect 19508 38872 19517 38912
rect 3148 38828 3188 38872
rect 3820 38828 3860 38872
rect 6403 38871 6461 38872
rect 8611 38871 8669 38872
rect 4003 38828 4061 38829
rect 13987 38828 14045 38829
rect 3139 38788 3148 38828
rect 3188 38788 3197 38828
rect 3811 38788 3820 38828
rect 3860 38788 3869 38828
rect 4003 38788 4012 38828
rect 4052 38788 11360 38828
rect 11971 38788 11980 38828
rect 12020 38788 12940 38828
rect 12980 38788 12989 38828
rect 13987 38788 13996 38828
rect 14036 38788 16300 38828
rect 16340 38788 16349 38828
rect 4003 38787 4061 38788
rect 7075 38744 7133 38745
rect 8227 38744 8285 38745
rect 10243 38744 10301 38745
rect 0 38704 1132 38744
rect 1172 38704 2540 38744
rect 2947 38704 2956 38744
rect 2996 38704 3284 38744
rect 3331 38704 3340 38744
rect 3380 38704 7084 38744
rect 7124 38704 7133 38744
rect 7555 38704 7564 38744
rect 7604 38704 7852 38744
rect 7892 38704 7901 38744
rect 8227 38704 8236 38744
rect 8276 38704 10060 38744
rect 10100 38704 10252 38744
rect 10292 38704 10301 38744
rect 11320 38744 11360 38788
rect 13987 38787 14045 38788
rect 18019 38744 18077 38745
rect 18412 38744 18452 38872
rect 21283 38828 21341 38829
rect 19564 38788 21292 38828
rect 21332 38788 21341 38828
rect 19564 38744 19604 38788
rect 21283 38787 21341 38788
rect 21379 38744 21437 38745
rect 11320 38704 12748 38744
rect 12788 38704 12797 38744
rect 13603 38704 13612 38744
rect 13652 38704 18028 38744
rect 18068 38704 18077 38744
rect 18403 38704 18412 38744
rect 18452 38704 18461 38744
rect 19555 38704 19564 38744
rect 19604 38704 19613 38744
rect 19660 38704 19943 38744
rect 19983 38704 19992 38744
rect 20035 38704 20044 38744
rect 20084 38704 21388 38744
rect 21428 38704 21437 38744
rect 0 38684 80 38704
rect 1123 38703 1181 38704
rect 1699 38620 1708 38660
rect 1748 38620 2284 38660
rect 2324 38620 2333 38660
rect 2083 38576 2141 38577
rect 2947 38576 3005 38577
rect 1795 38536 1804 38576
rect 1844 38536 2092 38576
rect 2132 38536 2141 38576
rect 2862 38536 2956 38576
rect 2996 38536 3005 38576
rect 3244 38576 3284 38704
rect 7075 38703 7133 38704
rect 8227 38703 8285 38704
rect 10243 38703 10301 38704
rect 18019 38703 18077 38704
rect 11203 38660 11261 38661
rect 19660 38660 19700 38704
rect 21379 38703 21437 38704
rect 20899 38660 20957 38661
rect 4003 38620 4012 38660
rect 4052 38620 4396 38660
rect 4436 38620 4445 38660
rect 4492 38620 11212 38660
rect 11252 38620 11261 38660
rect 11587 38620 11596 38660
rect 11636 38620 11884 38660
rect 11924 38620 11933 38660
rect 12547 38620 12556 38660
rect 12596 38620 13708 38660
rect 13748 38620 13757 38660
rect 15532 38620 17260 38660
rect 17300 38620 17309 38660
rect 18115 38620 18124 38660
rect 18164 38620 19700 38660
rect 19747 38620 19756 38660
rect 19796 38620 20908 38660
rect 20948 38620 20957 38660
rect 4195 38576 4253 38577
rect 4492 38576 4532 38620
rect 11203 38619 11261 38620
rect 8707 38576 8765 38577
rect 10051 38576 10109 38577
rect 12643 38576 12701 38577
rect 15532 38576 15572 38620
rect 20899 38619 20957 38620
rect 21424 38576 21504 38596
rect 3244 38536 4204 38576
rect 4244 38536 4253 38576
rect 2083 38535 2141 38536
rect 2947 38535 3005 38536
rect 4195 38535 4253 38536
rect 4300 38536 4532 38576
rect 4919 38536 4928 38576
rect 4968 38536 5010 38576
rect 5050 38536 5092 38576
rect 5132 38536 5174 38576
rect 5214 38536 5256 38576
rect 5296 38536 5305 38576
rect 7171 38536 7180 38576
rect 7220 38536 8468 38576
rect 4300 38492 4340 38536
rect 7180 38492 7220 38536
rect 8428 38492 8468 38536
rect 8707 38536 8716 38576
rect 8756 38536 10060 38576
rect 10100 38536 10109 38576
rect 10243 38536 10252 38576
rect 10292 38536 11020 38576
rect 11060 38536 11069 38576
rect 12643 38536 12652 38576
rect 12692 38536 15572 38576
rect 15628 38536 19852 38576
rect 19892 38536 19901 38576
rect 20039 38536 20048 38576
rect 20088 38536 20130 38576
rect 20170 38536 20212 38576
rect 20252 38536 20294 38576
rect 20334 38536 20376 38576
rect 20416 38536 20425 38576
rect 20812 38536 21504 38576
rect 8707 38535 8765 38536
rect 10051 38535 10109 38536
rect 12643 38535 12701 38536
rect 15235 38492 15293 38493
rect 1603 38452 1612 38492
rect 1652 38452 3572 38492
rect 3619 38452 3628 38492
rect 3668 38452 4340 38492
rect 4387 38452 4396 38492
rect 4436 38452 7220 38492
rect 7843 38452 7852 38492
rect 7892 38452 8044 38492
rect 8084 38452 8093 38492
rect 8419 38452 8428 38492
rect 8468 38452 9580 38492
rect 9620 38452 11980 38492
rect 12020 38452 12029 38492
rect 12163 38452 12172 38492
rect 12212 38452 12556 38492
rect 12596 38452 12605 38492
rect 13219 38452 13228 38492
rect 13268 38452 15244 38492
rect 15284 38452 15293 38492
rect 0 38408 80 38428
rect 3532 38408 3572 38452
rect 15235 38451 15293 38452
rect 0 38368 1748 38408
rect 1795 38368 1804 38408
rect 1844 38368 3148 38408
rect 3188 38368 3197 38408
rect 3532 38368 7700 38408
rect 8131 38368 8140 38408
rect 8180 38368 14476 38408
rect 14516 38368 14525 38408
rect 0 38348 80 38368
rect 1708 38324 1748 38368
rect 2179 38324 2237 38325
rect 7363 38324 7421 38325
rect 1708 38284 2188 38324
rect 2228 38284 2237 38324
rect 2563 38284 2572 38324
rect 2612 38284 7372 38324
rect 7412 38284 7421 38324
rect 2179 38283 2237 38284
rect 7363 38283 7421 38284
rect 7660 38241 7700 38368
rect 8035 38324 8093 38325
rect 9763 38324 9821 38325
rect 15628 38324 15668 38536
rect 16867 38492 16925 38493
rect 19651 38492 19709 38493
rect 16675 38452 16684 38492
rect 16724 38452 16876 38492
rect 16916 38452 16925 38492
rect 18595 38452 18604 38492
rect 18644 38452 19660 38492
rect 19700 38452 19709 38492
rect 16867 38451 16925 38452
rect 19651 38451 19709 38452
rect 19843 38492 19901 38493
rect 20812 38492 20852 38536
rect 21424 38516 21504 38536
rect 19843 38452 19852 38492
rect 19892 38452 20852 38492
rect 19843 38451 19901 38452
rect 16003 38408 16061 38409
rect 15918 38368 16012 38408
rect 16052 38368 16061 38408
rect 16579 38368 16588 38408
rect 16628 38368 16637 38408
rect 18883 38368 18892 38408
rect 18932 38368 19276 38408
rect 19316 38368 19325 38408
rect 19459 38368 19468 38408
rect 19508 38368 20236 38408
rect 20276 38368 20285 38408
rect 16003 38367 16061 38368
rect 7950 38284 8044 38324
rect 8084 38284 8093 38324
rect 8323 38284 8332 38324
rect 8372 38284 9772 38324
rect 9812 38284 15668 38324
rect 8035 38283 8093 38284
rect 9763 38283 9821 38284
rect 4579 38240 4637 38241
rect 5539 38240 5597 38241
rect 1516 38200 4588 38240
rect 4628 38200 4637 38240
rect 5059 38200 5068 38240
rect 5108 38200 5548 38240
rect 5588 38200 5597 38240
rect 1516 38156 1556 38200
rect 4579 38199 4637 38200
rect 5539 38199 5597 38200
rect 7651 38240 7709 38241
rect 8707 38240 8765 38241
rect 16588 38240 16628 38368
rect 19075 38284 19084 38324
rect 19124 38284 20140 38324
rect 20180 38284 20524 38324
rect 20564 38284 20573 38324
rect 17635 38240 17693 38241
rect 19267 38240 19325 38241
rect 19939 38240 19997 38241
rect 7651 38200 7660 38240
rect 7700 38200 8716 38240
rect 8756 38200 8765 38240
rect 9283 38200 9292 38240
rect 9332 38200 9868 38240
rect 9908 38200 9917 38240
rect 10051 38200 10060 38240
rect 10100 38200 13652 38240
rect 14659 38200 14668 38240
rect 14708 38200 15052 38240
rect 15092 38200 15101 38240
rect 15907 38200 15916 38240
rect 15956 38200 16876 38240
rect 16916 38200 17068 38240
rect 17108 38200 17117 38240
rect 17550 38200 17644 38240
rect 17684 38200 17693 38240
rect 18595 38200 18604 38240
rect 18644 38200 18892 38240
rect 18932 38200 18941 38240
rect 19267 38200 19276 38240
rect 19316 38200 19468 38240
rect 19508 38200 19517 38240
rect 19939 38200 19948 38240
rect 19988 38200 20044 38240
rect 20084 38200 20093 38240
rect 7651 38199 7709 38200
rect 8707 38199 8765 38200
rect 2371 38156 2429 38157
rect 1507 38116 1516 38156
rect 1556 38116 1565 38156
rect 2179 38116 2188 38156
rect 2228 38116 2380 38156
rect 2420 38116 2429 38156
rect 2371 38115 2429 38116
rect 2563 38156 2621 38157
rect 3331 38156 3389 38157
rect 9955 38156 10013 38157
rect 13411 38156 13469 38157
rect 2563 38116 2572 38156
rect 2612 38116 2706 38156
rect 2755 38116 2764 38156
rect 2804 38116 3340 38156
rect 3380 38116 3389 38156
rect 3715 38116 3724 38156
rect 3764 38116 9964 38156
rect 10004 38116 10013 38156
rect 11299 38116 11308 38156
rect 11348 38116 11596 38156
rect 11636 38116 11980 38156
rect 12020 38116 12029 38156
rect 13326 38116 13420 38156
rect 13460 38116 13469 38156
rect 2563 38115 2621 38116
rect 3331 38115 3389 38116
rect 9955 38115 10013 38116
rect 13411 38115 13469 38116
rect 0 38072 80 38092
rect 4867 38072 4925 38073
rect 8803 38072 8861 38073
rect 11491 38072 11549 38073
rect 0 38032 3628 38072
rect 3668 38032 3677 38072
rect 4782 38032 4876 38072
rect 4916 38032 4925 38072
rect 7555 38032 7564 38072
rect 7604 38032 7756 38072
rect 7796 38032 8812 38072
rect 8852 38032 8861 38072
rect 9571 38032 9580 38072
rect 9620 38032 11500 38072
rect 11540 38032 11549 38072
rect 13612 38072 13652 38200
rect 17635 38199 17693 38200
rect 19267 38199 19325 38200
rect 19939 38199 19997 38200
rect 16291 38156 16349 38157
rect 19843 38156 19901 38157
rect 13699 38116 13708 38156
rect 13748 38116 16052 38156
rect 13612 38032 14860 38072
rect 14900 38032 15532 38072
rect 15572 38032 15581 38072
rect 0 38012 80 38032
rect 4867 38031 4925 38032
rect 8803 38031 8861 38032
rect 11491 38031 11549 38032
rect 1507 37988 1565 37989
rect 16012 37988 16052 38116
rect 16291 38116 16300 38156
rect 16340 38116 19852 38156
rect 19892 38116 19901 38156
rect 16291 38115 16349 38116
rect 19843 38115 19901 38116
rect 19363 38072 19421 38073
rect 21424 38072 21504 38092
rect 16387 38032 16396 38072
rect 16436 38032 18220 38072
rect 18260 38032 18269 38072
rect 19363 38032 19372 38072
rect 19412 38032 21504 38072
rect 19363 38031 19421 38032
rect 21424 38012 21504 38032
rect 1507 37948 1516 37988
rect 1556 37948 3148 37988
rect 3188 37948 3197 37988
rect 3811 37948 3820 37988
rect 3860 37948 3869 37988
rect 4579 37948 4588 37988
rect 4628 37948 5740 37988
rect 5780 37948 5789 37988
rect 6307 37948 6316 37988
rect 6356 37948 9004 37988
rect 9044 37948 9053 37988
rect 9763 37948 9772 37988
rect 9812 37948 9821 37988
rect 9955 37948 9964 37988
rect 10004 37948 15916 37988
rect 15956 37948 15965 37988
rect 16012 37948 16628 37988
rect 17251 37948 17260 37988
rect 17300 37948 19564 37988
rect 19604 37948 19613 37988
rect 1507 37947 1565 37948
rect 2947 37904 3005 37905
rect 3820 37904 3860 37948
rect 7660 37904 7700 37948
rect 9772 37904 9812 37948
rect 12835 37904 12893 37905
rect 15715 37904 15773 37905
rect 2862 37864 2956 37904
rect 2996 37864 3005 37904
rect 2947 37863 3005 37864
rect 3052 37864 3860 37904
rect 7564 37864 7700 37904
rect 7843 37864 7852 37904
rect 7892 37864 8428 37904
rect 8468 37864 8477 37904
rect 9772 37864 10060 37904
rect 10100 37864 10109 37904
rect 11203 37864 11212 37904
rect 11252 37864 11596 37904
rect 11636 37864 11645 37904
rect 11692 37864 12212 37904
rect 2755 37820 2813 37821
rect 3052 37820 3092 37864
rect 7564 37820 7604 37864
rect 9475 37820 9533 37821
rect 11107 37820 11165 37821
rect 11692 37820 11732 37864
rect 1188 37780 1228 37820
rect 1268 37780 1277 37820
rect 2670 37780 2764 37820
rect 2804 37780 2813 37820
rect 0 37736 80 37756
rect 931 37736 989 37737
rect 0 37696 940 37736
rect 980 37696 989 37736
rect 1228 37736 1268 37780
rect 2755 37779 2813 37780
rect 2956 37780 3092 37820
rect 3679 37780 3688 37820
rect 3728 37780 3770 37820
rect 3810 37780 3852 37820
rect 3892 37780 3934 37820
rect 3974 37780 4016 37820
rect 4056 37780 4065 37820
rect 7555 37780 7564 37820
rect 7604 37780 7613 37820
rect 9390 37780 9484 37820
rect 9524 37780 9533 37820
rect 10500 37780 10540 37820
rect 10580 37780 10589 37820
rect 11022 37780 11116 37820
rect 11156 37780 11165 37820
rect 1228 37696 1900 37736
rect 1940 37696 1949 37736
rect 0 37676 80 37696
rect 931 37695 989 37696
rect 2563 37652 2621 37653
rect 2956 37652 2996 37780
rect 9475 37779 9533 37780
rect 3043 37736 3101 37737
rect 10540 37736 10580 37780
rect 11107 37779 11165 37780
rect 11212 37780 11732 37820
rect 11212 37736 11252 37780
rect 3043 37696 3052 37736
rect 3092 37696 4588 37736
rect 4628 37696 4637 37736
rect 5251 37696 5260 37736
rect 5300 37696 5932 37736
rect 5972 37696 6164 37736
rect 6211 37696 6220 37736
rect 6260 37696 9908 37736
rect 10540 37696 11252 37736
rect 11299 37736 11357 37737
rect 12172 37736 12212 37864
rect 12835 37864 12844 37904
rect 12884 37864 12940 37904
rect 12980 37864 12989 37904
rect 15619 37864 15628 37904
rect 15668 37864 15724 37904
rect 15764 37864 15773 37904
rect 16588 37904 16628 37948
rect 17443 37904 17501 37905
rect 16588 37864 17452 37904
rect 17492 37864 17501 37904
rect 12835 37863 12893 37864
rect 15715 37863 15773 37864
rect 17443 37863 17501 37864
rect 13027 37820 13085 37821
rect 14179 37820 14237 37821
rect 16483 37820 16541 37821
rect 12942 37780 13036 37820
rect 13076 37780 13085 37820
rect 14094 37780 14188 37820
rect 14228 37780 14237 37820
rect 15235 37780 15244 37820
rect 15284 37780 16108 37820
rect 16148 37780 16157 37820
rect 16398 37780 16492 37820
rect 16532 37780 16541 37820
rect 18799 37780 18808 37820
rect 18848 37780 18890 37820
rect 18930 37780 18972 37820
rect 19012 37780 19054 37820
rect 19094 37780 19136 37820
rect 19176 37780 19185 37820
rect 19267 37780 19276 37820
rect 19316 37780 19852 37820
rect 19892 37780 19901 37820
rect 20580 37780 20620 37820
rect 20660 37780 20669 37820
rect 13027 37779 13085 37780
rect 14179 37779 14237 37780
rect 16483 37779 16541 37780
rect 16483 37736 16541 37737
rect 16867 37736 16925 37737
rect 20620 37736 20660 37780
rect 11299 37696 11308 37736
rect 11348 37696 12076 37736
rect 12116 37696 12125 37736
rect 12172 37696 13748 37736
rect 13987 37696 13996 37736
rect 14036 37696 16436 37736
rect 3043 37695 3101 37696
rect 6124 37652 6164 37696
rect 9763 37652 9821 37653
rect 1219 37612 1228 37652
rect 1268 37612 2572 37652
rect 2612 37612 2996 37652
rect 4291 37612 4300 37652
rect 4340 37612 6028 37652
rect 6068 37612 6077 37652
rect 6124 37612 7372 37652
rect 7412 37612 7421 37652
rect 7651 37612 7660 37652
rect 7700 37612 8140 37652
rect 8180 37612 9004 37652
rect 9044 37612 9053 37652
rect 9187 37612 9196 37652
rect 9236 37612 9484 37652
rect 9524 37612 9533 37652
rect 9678 37612 9772 37652
rect 9812 37612 9821 37652
rect 9868 37652 9908 37696
rect 11299 37695 11357 37696
rect 12643 37652 12701 37653
rect 9868 37612 12652 37652
rect 12692 37612 12701 37652
rect 13708 37652 13748 37696
rect 15427 37652 15485 37653
rect 13708 37612 15052 37652
rect 15092 37612 15101 37652
rect 15342 37612 15436 37652
rect 15476 37612 15485 37652
rect 2563 37611 2621 37612
rect 9763 37611 9821 37612
rect 12643 37611 12701 37612
rect 15427 37611 15485 37612
rect 3715 37568 3773 37569
rect 11299 37568 11357 37569
rect 13315 37568 13373 37569
rect 16396 37568 16436 37696
rect 16483 37696 16492 37736
rect 16532 37696 16684 37736
rect 16724 37696 16733 37736
rect 16867 37696 16876 37736
rect 16916 37696 16925 37736
rect 19939 37696 19948 37736
rect 19988 37696 19997 37736
rect 20620 37696 20908 37736
rect 20948 37696 20957 37736
rect 16483 37695 16541 37696
rect 16867 37695 16925 37696
rect 16876 37652 16916 37695
rect 19948 37652 19988 37696
rect 16579 37612 16588 37652
rect 16628 37612 16916 37652
rect 16963 37612 16972 37652
rect 17012 37612 17356 37652
rect 17396 37612 17405 37652
rect 18787 37612 18796 37652
rect 18836 37612 19988 37652
rect 19267 37568 19325 37569
rect 2083 37528 2092 37568
rect 2132 37528 3724 37568
rect 3764 37528 3773 37568
rect 3715 37527 3773 37528
rect 3916 37528 5260 37568
rect 5300 37528 5309 37568
rect 5443 37528 5452 37568
rect 5492 37528 11308 37568
rect 11348 37528 11357 37568
rect 11683 37528 11692 37568
rect 11732 37528 12076 37568
rect 12116 37528 12125 37568
rect 12739 37528 12748 37568
rect 12788 37528 13324 37568
rect 13364 37528 15532 37568
rect 15572 37528 15581 37568
rect 16396 37528 18988 37568
rect 19028 37528 19276 37568
rect 19316 37528 19325 37568
rect 1315 37484 1373 37485
rect 3916 37484 3956 37528
rect 11299 37527 11357 37528
rect 13315 37527 13373 37528
rect 19267 37527 19325 37528
rect 21187 37568 21245 37569
rect 21424 37568 21504 37588
rect 21187 37528 21196 37568
rect 21236 37528 21504 37568
rect 21187 37527 21245 37528
rect 21424 37508 21504 37528
rect 4099 37484 4157 37485
rect 4483 37484 4541 37485
rect 1230 37444 1324 37484
rect 1364 37444 1373 37484
rect 1315 37443 1373 37444
rect 2764 37444 3956 37484
rect 4014 37444 4108 37484
rect 4148 37444 4157 37484
rect 4398 37444 4492 37484
rect 4532 37444 4541 37484
rect 0 37400 80 37420
rect 2764 37401 2804 37444
rect 4099 37443 4157 37444
rect 4483 37443 4541 37444
rect 5635 37484 5693 37485
rect 8707 37484 8765 37485
rect 12355 37484 12413 37485
rect 15235 37484 15293 37485
rect 19363 37484 19421 37485
rect 5635 37444 5644 37484
rect 5684 37444 7084 37484
rect 7124 37444 7133 37484
rect 8707 37444 8716 37484
rect 8756 37444 9388 37484
rect 9428 37444 9437 37484
rect 10915 37444 10924 37484
rect 10964 37444 12364 37484
rect 12404 37444 14668 37484
rect 14708 37444 14717 37484
rect 15235 37444 15244 37484
rect 15284 37444 15293 37484
rect 16195 37444 16204 37484
rect 16244 37444 17164 37484
rect 17204 37444 17213 37484
rect 19363 37444 19372 37484
rect 19412 37444 19796 37484
rect 5635 37443 5693 37444
rect 8707 37443 8765 37444
rect 12355 37443 12413 37444
rect 15235 37443 15293 37444
rect 19363 37443 19421 37444
rect 2755 37400 2813 37401
rect 3235 37400 3293 37401
rect 9475 37400 9533 37401
rect 11683 37400 11741 37401
rect 15244 37400 15284 37443
rect 17443 37400 17501 37401
rect 19756 37400 19796 37444
rect 0 37360 2764 37400
rect 2804 37360 2813 37400
rect 3139 37360 3148 37400
rect 3188 37360 3244 37400
rect 3284 37360 3293 37400
rect 3811 37360 3820 37400
rect 3860 37360 6412 37400
rect 6452 37360 6461 37400
rect 8995 37360 9004 37400
rect 9044 37360 9484 37400
rect 9524 37360 9533 37400
rect 11587 37360 11596 37400
rect 11636 37360 11692 37400
rect 11732 37360 11741 37400
rect 12643 37360 12652 37400
rect 12692 37360 13420 37400
rect 13460 37360 13469 37400
rect 14851 37360 14860 37400
rect 14900 37360 15148 37400
rect 15188 37360 15197 37400
rect 15244 37360 15436 37400
rect 15476 37360 15485 37400
rect 15907 37360 15916 37400
rect 15956 37360 16108 37400
rect 16148 37360 17260 37400
rect 17300 37360 17309 37400
rect 17443 37360 17452 37400
rect 17492 37360 18892 37400
rect 18932 37360 19084 37400
rect 19124 37360 19133 37400
rect 19267 37360 19276 37400
rect 19316 37360 19700 37400
rect 19756 37360 20034 37400
rect 20074 37360 20083 37400
rect 0 37340 80 37360
rect 2755 37359 2813 37360
rect 3235 37359 3293 37360
rect 9475 37359 9533 37360
rect 11683 37359 11741 37360
rect 17443 37359 17501 37360
rect 5635 37316 5693 37317
rect 5923 37316 5981 37317
rect 8899 37316 8957 37317
rect 15523 37316 15581 37317
rect 16483 37316 16541 37317
rect 17347 37316 17405 37317
rect 19660 37316 19700 37360
rect 2563 37276 2572 37316
rect 2612 37276 5644 37316
rect 5684 37276 5693 37316
rect 5838 37276 5932 37316
rect 5972 37276 5981 37316
rect 7363 37276 7372 37316
rect 7412 37276 8908 37316
rect 8948 37276 8957 37316
rect 12451 37276 12460 37316
rect 12500 37276 12748 37316
rect 12788 37276 12797 37316
rect 13219 37276 13228 37316
rect 13268 37276 15532 37316
rect 15572 37276 16492 37316
rect 16532 37276 16541 37316
rect 17059 37276 17068 37316
rect 17108 37276 17117 37316
rect 17262 37276 17356 37316
rect 17396 37276 17405 37316
rect 18691 37276 18700 37316
rect 18740 37276 19564 37316
rect 19604 37276 19613 37316
rect 19660 37276 20140 37316
rect 20180 37276 20189 37316
rect 5635 37275 5693 37276
rect 5923 37275 5981 37276
rect 8899 37275 8957 37276
rect 15523 37275 15581 37276
rect 16483 37275 16541 37276
rect 1123 37232 1181 37233
rect 16867 37232 16925 37233
rect 17068 37232 17108 37276
rect 17347 37275 17405 37276
rect 1123 37192 1132 37232
rect 1172 37192 1324 37232
rect 1364 37192 1373 37232
rect 1699 37192 1708 37232
rect 1748 37192 3820 37232
rect 3860 37192 3869 37232
rect 3916 37192 6892 37232
rect 6932 37192 6941 37232
rect 15523 37192 15532 37232
rect 15572 37192 16436 37232
rect 1123 37191 1181 37192
rect 3916 37148 3956 37192
rect 5827 37148 5885 37149
rect 6019 37148 6077 37149
rect 3523 37108 3532 37148
rect 3572 37108 3956 37148
rect 4483 37108 4492 37148
rect 4532 37108 5836 37148
rect 5876 37108 5885 37148
rect 5934 37108 6028 37148
rect 6068 37108 6077 37148
rect 10819 37108 10828 37148
rect 10868 37108 15628 37148
rect 15668 37108 16340 37148
rect 5827 37107 5885 37108
rect 6019 37107 6077 37108
rect 0 37064 80 37084
rect 16195 37064 16253 37065
rect 0 37024 212 37064
rect 1411 37024 1420 37064
rect 1460 37024 1900 37064
rect 1940 37024 1949 37064
rect 4919 37024 4928 37064
rect 4968 37024 5010 37064
rect 5050 37024 5092 37064
rect 5132 37024 5174 37064
rect 5214 37024 5256 37064
rect 5296 37024 5305 37064
rect 5452 37024 6508 37064
rect 6548 37024 6796 37064
rect 6836 37024 6845 37064
rect 7555 37024 7564 37064
rect 7604 37024 8140 37064
rect 8180 37024 8189 37064
rect 11011 37024 11020 37064
rect 11060 37024 13036 37064
rect 13076 37024 13085 37064
rect 13411 37024 13420 37064
rect 13460 37024 16204 37064
rect 16244 37024 16253 37064
rect 0 37004 80 37024
rect 172 36896 212 37024
rect 5452 36980 5492 37024
rect 16195 37023 16253 37024
rect 16300 36980 16340 37108
rect 16396 37064 16436 37192
rect 16867 37192 16876 37232
rect 16916 37192 16972 37232
rect 17012 37192 17021 37232
rect 17068 37192 18988 37232
rect 19028 37192 19037 37232
rect 16867 37191 16925 37192
rect 17539 37108 17548 37148
rect 17588 37108 18796 37148
rect 18836 37108 19948 37148
rect 19988 37108 19997 37148
rect 20803 37064 20861 37065
rect 21424 37064 21504 37084
rect 16396 37024 18316 37064
rect 18356 37024 18365 37064
rect 20039 37024 20048 37064
rect 20088 37024 20130 37064
rect 20170 37024 20212 37064
rect 20252 37024 20294 37064
rect 20334 37024 20376 37064
rect 20416 37024 20425 37064
rect 20803 37024 20812 37064
rect 20852 37024 21504 37064
rect 20803 37023 20861 37024
rect 21424 37004 21504 37024
rect 19939 36980 19997 36981
rect 2500 36940 5492 36980
rect 5548 36940 7180 36980
rect 7220 36940 7229 36980
rect 8803 36940 8812 36980
rect 8852 36940 9772 36980
rect 9812 36940 9821 36980
rect 10243 36940 10252 36980
rect 10292 36940 14860 36980
rect 14900 36940 16108 36980
rect 16148 36940 16157 36980
rect 16300 36940 16396 36980
rect 16436 36940 16445 36980
rect 16963 36940 16972 36980
rect 17012 36940 17836 36980
rect 17876 36940 17885 36980
rect 18019 36940 18028 36980
rect 18068 36940 19084 36980
rect 19124 36940 19133 36980
rect 19555 36940 19564 36980
rect 19604 36940 19948 36980
rect 19988 36940 19997 36980
rect 2275 36896 2333 36897
rect 2500 36896 2540 36940
rect 2947 36896 3005 36897
rect 172 36856 2284 36896
rect 2324 36856 2540 36896
rect 2851 36856 2860 36896
rect 2900 36856 2956 36896
rect 2996 36856 3532 36896
rect 3572 36856 3581 36896
rect 2275 36855 2333 36856
rect 2947 36855 3005 36856
rect 5548 36812 5588 36940
rect 5635 36856 5644 36896
rect 5684 36856 6700 36896
rect 6740 36856 6749 36896
rect 7180 36812 7220 36940
rect 19939 36939 19997 36940
rect 8131 36896 8189 36897
rect 15619 36896 15677 36897
rect 8046 36856 8140 36896
rect 8180 36856 9004 36896
rect 9044 36856 9053 36896
rect 11203 36856 11212 36896
rect 11252 36856 15628 36896
rect 15668 36856 15677 36896
rect 15811 36856 15820 36896
rect 15860 36856 16780 36896
rect 16820 36856 16829 36896
rect 17635 36856 17644 36896
rect 17684 36856 19468 36896
rect 19508 36856 19517 36896
rect 8131 36855 8189 36856
rect 15619 36855 15677 36856
rect 16291 36812 16349 36813
rect 2500 36772 5588 36812
rect 5923 36772 5932 36812
rect 5972 36772 6220 36812
rect 6260 36772 6269 36812
rect 7180 36772 10196 36812
rect 10243 36772 10252 36812
rect 10292 36772 10828 36812
rect 10868 36772 10877 36812
rect 13315 36772 13324 36812
rect 13364 36772 16300 36812
rect 16340 36772 16349 36812
rect 0 36728 80 36748
rect 2500 36728 2540 36772
rect 5827 36728 5885 36729
rect 7459 36728 7517 36729
rect 0 36688 2540 36728
rect 5742 36688 5836 36728
rect 5876 36688 5885 36728
rect 0 36668 80 36688
rect 5827 36687 5885 36688
rect 6316 36688 7468 36728
rect 7508 36688 7517 36728
rect 5443 36644 5501 36645
rect 6316 36644 6356 36688
rect 7459 36687 7517 36688
rect 8035 36728 8093 36729
rect 8611 36728 8669 36729
rect 8035 36688 8044 36728
rect 8084 36688 8620 36728
rect 8660 36688 8669 36728
rect 8035 36687 8093 36688
rect 8611 36687 8669 36688
rect 9091 36728 9149 36729
rect 9091 36688 9100 36728
rect 9140 36688 9234 36728
rect 9091 36687 9149 36688
rect 10156 36644 10196 36772
rect 16291 36771 16349 36772
rect 16483 36812 16541 36813
rect 17443 36812 17501 36813
rect 16483 36772 16492 36812
rect 16532 36772 17300 36812
rect 16483 36771 16541 36772
rect 15427 36728 15485 36729
rect 16867 36728 16925 36729
rect 10435 36688 10444 36728
rect 10484 36688 15052 36728
rect 15092 36688 15101 36728
rect 15147 36688 15156 36728
rect 15196 36688 15436 36728
rect 15476 36688 15485 36728
rect 15715 36688 15724 36728
rect 15764 36688 16300 36728
rect 16340 36688 16349 36728
rect 16867 36688 16876 36728
rect 16916 36688 17164 36728
rect 17204 36688 17213 36728
rect 14851 36644 14909 36645
rect 2083 36604 2092 36644
rect 2132 36604 2476 36644
rect 2516 36604 2525 36644
rect 5358 36604 5452 36644
rect 5492 36604 5501 36644
rect 6307 36604 6316 36644
rect 6356 36604 6365 36644
rect 6508 36604 8908 36644
rect 8948 36604 8957 36644
rect 10156 36604 11788 36644
rect 11828 36604 14860 36644
rect 14900 36604 14909 36644
rect 15052 36644 15092 36688
rect 15427 36687 15485 36688
rect 16867 36687 16925 36688
rect 17260 36644 17300 36772
rect 17443 36772 17452 36812
rect 17492 36772 17932 36812
rect 17972 36772 19660 36812
rect 19700 36772 20180 36812
rect 17443 36771 17501 36772
rect 20140 36728 20180 36772
rect 18595 36688 18604 36728
rect 18644 36688 19948 36728
rect 19988 36688 19997 36728
rect 20131 36688 20140 36728
rect 20180 36688 20189 36728
rect 19267 36644 19325 36645
rect 15052 36604 16972 36644
rect 17012 36604 17021 36644
rect 17260 36604 17452 36644
rect 17492 36604 17501 36644
rect 18883 36604 18892 36644
rect 18932 36604 18941 36644
rect 19182 36604 19276 36644
rect 19316 36604 19325 36644
rect 5443 36603 5501 36604
rect 1315 36560 1373 36561
rect 5251 36560 5309 36561
rect 6508 36560 6548 36604
rect 14851 36603 14909 36604
rect 9283 36560 9341 36561
rect 10819 36560 10877 36561
rect 1315 36520 1324 36560
rect 1364 36520 1612 36560
rect 1652 36520 1661 36560
rect 1891 36520 1900 36560
rect 1940 36520 3052 36560
rect 3092 36520 3101 36560
rect 3331 36520 3340 36560
rect 3380 36520 4300 36560
rect 4340 36520 4349 36560
rect 5166 36520 5260 36560
rect 5300 36520 5309 36560
rect 6499 36520 6508 36560
rect 6548 36520 6557 36560
rect 6883 36520 6892 36560
rect 6932 36520 7180 36560
rect 7220 36520 7229 36560
rect 7939 36520 7948 36560
rect 7988 36520 8812 36560
rect 8852 36520 8861 36560
rect 9187 36520 9196 36560
rect 9236 36520 9292 36560
rect 9332 36520 9341 36560
rect 10734 36520 10828 36560
rect 10868 36520 10877 36560
rect 1315 36519 1373 36520
rect 5251 36519 5309 36520
rect 9283 36519 9341 36520
rect 10819 36519 10877 36520
rect 11875 36560 11933 36561
rect 15235 36560 15293 36561
rect 18892 36560 18932 36604
rect 19267 36603 19325 36604
rect 20611 36560 20669 36561
rect 21424 36560 21504 36580
rect 11875 36520 11884 36560
rect 11924 36520 13516 36560
rect 13556 36520 13565 36560
rect 14851 36520 14860 36560
rect 14900 36520 15052 36560
rect 15092 36520 15101 36560
rect 15235 36520 15244 36560
rect 15284 36520 15436 36560
rect 15476 36520 15485 36560
rect 15811 36520 15820 36560
rect 15860 36520 16532 36560
rect 16579 36520 16588 36560
rect 16628 36520 17260 36560
rect 17300 36520 18796 36560
rect 18836 36520 18845 36560
rect 18892 36520 20044 36560
rect 20084 36520 20093 36560
rect 20611 36520 20620 36560
rect 20660 36520 21504 36560
rect 11875 36519 11933 36520
rect 15235 36519 15293 36520
rect 1891 36476 1949 36477
rect 10915 36476 10973 36477
rect 16492 36476 16532 36520
rect 20611 36519 20669 36520
rect 21424 36500 21504 36520
rect 16867 36476 16925 36477
rect 1891 36436 1900 36476
rect 1940 36436 5068 36476
rect 5108 36436 5117 36476
rect 5347 36436 5356 36476
rect 5396 36436 10924 36476
rect 10964 36436 10973 36476
rect 15331 36436 15340 36476
rect 15380 36436 15532 36476
rect 15572 36436 15581 36476
rect 15907 36436 15916 36476
rect 15956 36436 15965 36476
rect 16483 36436 16492 36476
rect 16532 36436 16541 36476
rect 16867 36436 16876 36476
rect 16916 36436 19756 36476
rect 19796 36436 19805 36476
rect 1891 36435 1949 36436
rect 10915 36435 10973 36436
rect 0 36392 80 36412
rect 5731 36392 5789 36393
rect 15916 36392 15956 36436
rect 16867 36435 16925 36436
rect 17347 36392 17405 36393
rect 19459 36392 19517 36393
rect 0 36352 5740 36392
rect 5780 36352 8332 36392
rect 8372 36352 8381 36392
rect 14755 36352 14764 36392
rect 14804 36352 15956 36392
rect 16003 36352 16012 36392
rect 16052 36352 17356 36392
rect 17396 36352 17405 36392
rect 19267 36352 19276 36392
rect 19316 36352 19468 36392
rect 19508 36352 19517 36392
rect 0 36332 80 36352
rect 5731 36351 5789 36352
rect 17347 36351 17405 36352
rect 19459 36351 19517 36352
rect 17635 36308 17693 36309
rect 3679 36268 3688 36308
rect 3728 36268 3770 36308
rect 3810 36268 3852 36308
rect 3892 36268 3934 36308
rect 3974 36268 4016 36308
rect 4056 36268 4065 36308
rect 7747 36268 7756 36308
rect 7796 36268 8140 36308
rect 8180 36268 8189 36308
rect 12163 36268 12172 36308
rect 12212 36268 17644 36308
rect 17684 36268 17693 36308
rect 18799 36268 18808 36308
rect 18848 36268 18890 36308
rect 18930 36268 18972 36308
rect 19012 36268 19054 36308
rect 19094 36268 19136 36308
rect 19176 36268 19185 36308
rect 17635 36267 17693 36268
rect 8227 36224 8285 36225
rect 3139 36184 3148 36224
rect 3188 36184 8236 36224
rect 8276 36184 8285 36224
rect 15523 36184 15532 36224
rect 15572 36184 16396 36224
rect 16436 36184 19372 36224
rect 19412 36184 19421 36224
rect 8227 36183 8285 36184
rect 2851 36140 2909 36141
rect 4771 36140 4829 36141
rect 8323 36140 8381 36141
rect 1699 36100 1708 36140
rect 1748 36100 1996 36140
rect 2036 36100 2045 36140
rect 2371 36100 2380 36140
rect 2420 36100 2708 36140
rect 0 36056 80 36076
rect 1507 36056 1565 36057
rect 0 36016 1516 36056
rect 1556 36016 1565 36056
rect 0 35996 80 36016
rect 1507 36015 1565 36016
rect 2668 35972 2708 36100
rect 2851 36100 2860 36140
rect 2900 36100 4780 36140
rect 4820 36100 4876 36140
rect 4916 36100 4925 36140
rect 8323 36100 8332 36140
rect 8372 36100 20620 36140
rect 20660 36100 20669 36140
rect 2851 36099 2909 36100
rect 4771 36099 4829 36100
rect 8323 36099 8381 36100
rect 7555 36056 7613 36057
rect 21424 36056 21504 36076
rect 3811 36016 3820 36056
rect 3860 36016 7372 36056
rect 7412 36016 7421 36056
rect 7555 36016 7564 36056
rect 7604 36016 7852 36056
rect 7892 36016 7901 36056
rect 9379 36016 9388 36056
rect 9428 36016 10348 36056
rect 10388 36016 10397 36056
rect 11587 36016 11596 36056
rect 11636 36016 21504 36056
rect 7555 36015 7613 36016
rect 21424 35996 21504 36016
rect 4771 35972 4829 35973
rect 10147 35972 10205 35973
rect 17443 35972 17501 35973
rect 931 35932 940 35972
rect 980 35932 2540 35972
rect 2668 35932 2860 35972
rect 2900 35932 4780 35972
rect 4820 35932 4829 35972
rect 7747 35932 7756 35972
rect 7796 35932 10156 35972
rect 10196 35932 10205 35972
rect 11203 35932 11212 35972
rect 11252 35932 12844 35972
rect 12884 35932 12893 35972
rect 14563 35932 14572 35972
rect 14612 35932 16204 35972
rect 16244 35932 16253 35972
rect 17347 35932 17356 35972
rect 17396 35932 17452 35972
rect 17492 35932 17501 35972
rect 2500 35888 2540 35932
rect 4771 35931 4829 35932
rect 10147 35931 10205 35932
rect 17443 35931 17501 35932
rect 7363 35888 7421 35889
rect 13123 35888 13181 35889
rect 19267 35888 19325 35889
rect 19555 35888 19613 35889
rect 2500 35848 4204 35888
rect 4244 35848 4396 35888
rect 4436 35848 4445 35888
rect 4579 35848 4588 35888
rect 4628 35848 6892 35888
rect 6932 35848 6941 35888
rect 7363 35848 7372 35888
rect 7412 35848 7852 35888
rect 7892 35848 7901 35888
rect 8323 35848 8332 35888
rect 8372 35848 9580 35888
rect 9620 35848 11884 35888
rect 11924 35848 11933 35888
rect 13123 35848 13132 35888
rect 13172 35848 13324 35888
rect 13364 35848 13373 35888
rect 13891 35848 13900 35888
rect 13940 35848 16588 35888
rect 16628 35848 16637 35888
rect 19171 35848 19180 35888
rect 19220 35848 19276 35888
rect 19316 35848 19325 35888
rect 19459 35848 19468 35888
rect 19508 35848 19564 35888
rect 19604 35848 19613 35888
rect 20515 35848 20524 35888
rect 20564 35848 20812 35888
rect 20852 35848 20861 35888
rect 7363 35847 7421 35848
rect 13123 35847 13181 35848
rect 19267 35847 19325 35848
rect 19555 35847 19613 35848
rect 835 35804 893 35805
rect 13219 35804 13277 35805
rect 835 35764 844 35804
rect 884 35764 3820 35804
rect 3860 35764 3869 35804
rect 6316 35764 9004 35804
rect 9044 35764 9053 35804
rect 13134 35764 13228 35804
rect 13268 35764 13277 35804
rect 835 35763 893 35764
rect 0 35720 80 35740
rect 451 35720 509 35721
rect 6316 35720 6356 35764
rect 13219 35763 13277 35764
rect 14755 35804 14813 35805
rect 18691 35804 18749 35805
rect 14755 35764 14764 35804
rect 14804 35764 18700 35804
rect 18740 35764 18749 35804
rect 19843 35764 19852 35804
rect 19892 35764 20044 35804
rect 20084 35764 20093 35804
rect 14755 35763 14813 35764
rect 18691 35763 18749 35764
rect 9955 35720 10013 35721
rect 0 35680 212 35720
rect 0 35660 80 35680
rect 172 35468 212 35680
rect 451 35680 460 35720
rect 500 35680 4780 35720
rect 4820 35680 4829 35720
rect 4876 35680 6356 35720
rect 6403 35680 6412 35720
rect 6452 35680 8812 35720
rect 8852 35680 8861 35720
rect 9955 35680 9964 35720
rect 10004 35680 20812 35720
rect 20852 35680 20861 35720
rect 451 35679 509 35680
rect 1315 35636 1373 35637
rect 4387 35636 4445 35637
rect 4876 35636 4916 35680
rect 6316 35636 6356 35680
rect 9955 35679 10013 35680
rect 8227 35636 8285 35637
rect 13315 35636 13373 35637
rect 16003 35636 16061 35637
rect 17827 35636 17885 35637
rect 18115 35636 18173 35637
rect 19843 35636 19901 35637
rect 1230 35596 1324 35636
rect 1364 35596 1373 35636
rect 2563 35596 2572 35636
rect 2612 35596 3764 35636
rect 4291 35596 4300 35636
rect 4340 35596 4396 35636
rect 4436 35596 4445 35636
rect 1315 35595 1373 35596
rect 3427 35552 3485 35553
rect 3724 35552 3764 35596
rect 4387 35595 4445 35596
rect 4492 35596 4916 35636
rect 6211 35596 6220 35636
rect 6260 35596 6269 35636
rect 6316 35596 6892 35636
rect 6932 35596 6941 35636
rect 8227 35596 8236 35636
rect 8276 35596 9388 35636
rect 9428 35596 9437 35636
rect 13230 35596 13324 35636
rect 13364 35596 13373 35636
rect 14275 35596 14284 35636
rect 14324 35596 14764 35636
rect 14804 35596 14813 35636
rect 15331 35596 15340 35636
rect 15380 35596 16012 35636
rect 16052 35596 16061 35636
rect 16195 35596 16204 35636
rect 16244 35596 17836 35636
rect 17876 35596 17885 35636
rect 18019 35596 18028 35636
rect 18068 35596 18124 35636
rect 18164 35596 18173 35636
rect 19747 35596 19756 35636
rect 19796 35596 19852 35636
rect 19892 35596 19901 35636
rect 4492 35552 4532 35596
rect 6220 35552 6260 35596
rect 8227 35595 8285 35596
rect 13315 35595 13373 35596
rect 16003 35595 16061 35596
rect 17827 35595 17885 35596
rect 18115 35595 18173 35596
rect 19843 35595 19901 35596
rect 21424 35552 21504 35572
rect 1891 35512 1900 35552
rect 1940 35512 3148 35552
rect 3188 35512 3197 35552
rect 3427 35512 3436 35552
rect 3476 35512 3628 35552
rect 3668 35512 3677 35552
rect 3724 35512 4532 35552
rect 4919 35512 4928 35552
rect 4968 35512 5010 35552
rect 5050 35512 5092 35552
rect 5132 35512 5174 35552
rect 5214 35512 5256 35552
rect 5296 35512 5305 35552
rect 6220 35512 6412 35552
rect 6452 35512 6461 35552
rect 10627 35512 10636 35552
rect 10676 35512 11116 35552
rect 11156 35512 13900 35552
rect 13940 35512 13949 35552
rect 17059 35512 17068 35552
rect 17108 35512 17452 35552
rect 17492 35512 17501 35552
rect 17620 35512 19660 35552
rect 19700 35512 19709 35552
rect 20039 35512 20048 35552
rect 20088 35512 20130 35552
rect 20170 35512 20212 35552
rect 20252 35512 20294 35552
rect 20334 35512 20376 35552
rect 20416 35512 20425 35552
rect 20707 35512 20716 35552
rect 20756 35512 21504 35552
rect 3427 35511 3485 35512
rect 1795 35468 1853 35469
rect 2083 35468 2141 35469
rect 3043 35468 3101 35469
rect 15043 35468 15101 35469
rect 17620 35468 17660 35512
rect 21424 35492 21504 35512
rect 18019 35468 18077 35469
rect 172 35428 1804 35468
rect 1844 35428 2092 35468
rect 2132 35428 2141 35468
rect 2947 35428 2956 35468
rect 2996 35428 3052 35468
rect 3092 35428 3101 35468
rect 3523 35428 3532 35468
rect 3572 35428 3581 35468
rect 4387 35428 4396 35468
rect 4436 35428 8236 35468
rect 8276 35428 8285 35468
rect 10147 35428 10156 35468
rect 10196 35428 13172 35468
rect 13699 35428 13708 35468
rect 13748 35428 15052 35468
rect 15092 35428 15101 35468
rect 1795 35427 1853 35428
rect 2083 35427 2141 35428
rect 3043 35427 3101 35428
rect 0 35384 80 35404
rect 3331 35384 3389 35385
rect 0 35344 3340 35384
rect 3380 35344 3389 35384
rect 0 35324 80 35344
rect 3331 35343 3389 35344
rect 1795 35300 1853 35301
rect 2467 35300 2525 35301
rect 1710 35260 1804 35300
rect 1844 35260 1853 35300
rect 2371 35260 2380 35300
rect 2420 35260 2476 35300
rect 2516 35260 2525 35300
rect 1795 35259 1853 35260
rect 2467 35259 2525 35260
rect 2371 35216 2429 35217
rect 3532 35216 3572 35428
rect 3619 35384 3677 35385
rect 13132 35384 13172 35428
rect 15043 35427 15101 35428
rect 16108 35428 16780 35468
rect 16820 35428 17660 35468
rect 17827 35428 17836 35468
rect 17876 35428 18028 35468
rect 18068 35428 18700 35468
rect 18740 35428 18749 35468
rect 16108 35384 16148 35428
rect 18019 35427 18077 35428
rect 16291 35384 16349 35385
rect 17347 35384 17405 35385
rect 3619 35344 3628 35384
rect 3668 35344 3820 35384
rect 3860 35344 3869 35384
rect 4483 35344 4492 35384
rect 4532 35344 4541 35384
rect 6307 35344 6316 35384
rect 6356 35344 10060 35384
rect 10100 35344 10109 35384
rect 11011 35344 11020 35384
rect 11060 35344 11596 35384
rect 11636 35344 11645 35384
rect 13132 35344 16148 35384
rect 16206 35344 16300 35384
rect 16340 35344 16349 35384
rect 17262 35344 17356 35384
rect 17396 35344 17405 35384
rect 3619 35343 3677 35344
rect 4492 35300 4532 35344
rect 16291 35343 16349 35344
rect 17347 35343 17405 35344
rect 5347 35300 5405 35301
rect 15139 35300 15197 35301
rect 15619 35300 15677 35301
rect 18403 35300 18461 35301
rect 4492 35260 5356 35300
rect 5396 35260 5405 35300
rect 6019 35260 6028 35300
rect 6068 35260 6796 35300
rect 6836 35260 6845 35300
rect 6979 35260 6988 35300
rect 7028 35260 10156 35300
rect 10196 35260 10205 35300
rect 10723 35260 10732 35300
rect 10772 35260 12364 35300
rect 12404 35260 12413 35300
rect 13324 35260 13804 35300
rect 13844 35260 13853 35300
rect 14659 35260 14668 35300
rect 14708 35260 14956 35300
rect 14996 35260 15005 35300
rect 15108 35260 15148 35300
rect 15188 35260 15197 35300
rect 15534 35260 15628 35300
rect 15668 35260 15677 35300
rect 16099 35260 16108 35300
rect 16148 35260 18028 35300
rect 18068 35260 18077 35300
rect 18307 35260 18316 35300
rect 18356 35260 18412 35300
rect 18452 35260 18461 35300
rect 5347 35259 5405 35260
rect 6307 35216 6365 35217
rect 6499 35216 6557 35217
rect 9667 35216 9725 35217
rect 11203 35216 11261 35217
rect 11683 35216 11741 35217
rect 2179 35176 2188 35216
rect 2228 35176 2380 35216
rect 2420 35176 2429 35216
rect 3139 35176 3148 35216
rect 3188 35176 3572 35216
rect 4195 35176 4204 35216
rect 4244 35176 4972 35216
rect 5012 35176 5021 35216
rect 6115 35176 6124 35216
rect 6164 35176 6316 35216
rect 6356 35176 6365 35216
rect 6414 35176 6508 35216
rect 6548 35176 6557 35216
rect 7747 35176 7756 35216
rect 7796 35176 8332 35216
rect 8372 35176 8381 35216
rect 9571 35176 9580 35216
rect 9620 35176 9676 35216
rect 9716 35176 9725 35216
rect 11118 35176 11212 35216
rect 11252 35176 11261 35216
rect 11587 35176 11596 35216
rect 11636 35176 11692 35216
rect 11732 35176 11741 35216
rect 2371 35175 2429 35176
rect 6307 35175 6365 35176
rect 6499 35175 6557 35176
rect 9667 35175 9725 35176
rect 11203 35175 11261 35176
rect 11683 35175 11741 35176
rect 4099 35132 4157 35133
rect 13324 35132 13364 35260
rect 15139 35259 15197 35260
rect 15619 35259 15677 35260
rect 18403 35259 18461 35260
rect 13507 35216 13565 35217
rect 14083 35216 14141 35217
rect 15148 35216 15188 35259
rect 18211 35216 18269 35217
rect 13411 35176 13420 35216
rect 13460 35176 13516 35216
rect 13556 35176 13565 35216
rect 13987 35176 13996 35216
rect 14036 35176 14092 35216
rect 14132 35176 14141 35216
rect 14467 35176 14476 35216
rect 14516 35176 15188 35216
rect 16387 35176 16396 35216
rect 16436 35176 17452 35216
rect 17492 35176 17740 35216
rect 17780 35176 17789 35216
rect 18211 35176 18220 35216
rect 18260 35176 19756 35216
rect 19796 35176 19805 35216
rect 13507 35175 13565 35176
rect 14083 35175 14141 35176
rect 18211 35175 18269 35176
rect 14563 35132 14621 35133
rect 3043 35092 3052 35132
rect 3092 35092 3724 35132
rect 3764 35092 3773 35132
rect 3818 35092 3827 35132
rect 3867 35092 4108 35132
rect 4148 35092 4157 35132
rect 4483 35092 4492 35132
rect 4532 35092 6700 35132
rect 6740 35092 7948 35132
rect 7988 35092 8908 35132
rect 8948 35092 9196 35132
rect 9236 35092 9245 35132
rect 9955 35092 9964 35132
rect 10004 35092 10444 35132
rect 10484 35092 10924 35132
rect 10964 35092 10973 35132
rect 13315 35092 13324 35132
rect 13364 35092 13373 35132
rect 14478 35092 14572 35132
rect 14612 35092 14621 35132
rect 15235 35092 15244 35132
rect 15284 35092 17932 35132
rect 17972 35092 17981 35132
rect 4099 35091 4157 35092
rect 14563 35091 14621 35092
rect 0 35048 80 35068
rect 13219 35048 13277 35049
rect 18115 35048 18173 35049
rect 21424 35048 21504 35068
rect 0 35008 2540 35048
rect 2659 35008 2668 35048
rect 2708 35008 4060 35048
rect 4100 35008 4109 35048
rect 4675 35008 4684 35048
rect 4724 35008 7852 35048
rect 7892 35008 8140 35048
rect 8180 35008 8189 35048
rect 13219 35008 13228 35048
rect 13268 35008 15532 35048
rect 15572 35008 15581 35048
rect 15715 35008 15724 35048
rect 15764 35008 16910 35048
rect 16950 35008 16959 35048
rect 17155 35008 17164 35048
rect 17204 35008 18124 35048
rect 18164 35008 18173 35048
rect 0 34988 80 35008
rect 67 34880 125 34881
rect 2500 34880 2540 35008
rect 13219 35007 13277 35008
rect 18115 35007 18173 35008
rect 20140 35008 21504 35048
rect 6115 34964 6173 34965
rect 16675 34964 16733 34965
rect 18499 34964 18557 34965
rect 3331 34924 3340 34964
rect 3380 34924 3532 34964
rect 3572 34924 3581 34964
rect 3907 34924 3916 34964
rect 3956 34924 4396 34964
rect 4436 34924 4445 34964
rect 5740 34924 6124 34964
rect 6164 34924 6173 34964
rect 14755 34924 14764 34964
rect 14804 34924 16684 34964
rect 16724 34924 16733 34964
rect 17347 34924 17356 34964
rect 17396 34924 18316 34964
rect 18356 34924 18365 34964
rect 18499 34924 18508 34964
rect 18548 34924 18557 34964
rect 19459 34924 19468 34964
rect 19508 34924 19948 34964
rect 19988 34924 19997 34964
rect 5740 34880 5780 34924
rect 6115 34923 6173 34924
rect 16675 34923 16733 34924
rect 18499 34923 18557 34924
rect 67 34840 76 34880
rect 116 34840 1804 34880
rect 1844 34840 1853 34880
rect 2500 34840 5780 34880
rect 6307 34880 6365 34881
rect 18508 34880 18548 34923
rect 19459 34880 19517 34881
rect 6307 34840 6316 34880
rect 6356 34840 7756 34880
rect 7796 34840 7805 34880
rect 7939 34840 7948 34880
rect 7988 34840 8236 34880
rect 8276 34840 8285 34880
rect 15139 34840 15148 34880
rect 15188 34840 16588 34880
rect 16628 34840 16637 34880
rect 17923 34840 17932 34880
rect 17972 34840 18548 34880
rect 19363 34840 19372 34880
rect 19412 34840 19468 34880
rect 19508 34840 19517 34880
rect 67 34839 125 34840
rect 6307 34839 6365 34840
rect 19459 34839 19517 34840
rect 18499 34796 18557 34797
rect 1315 34756 1324 34796
rect 1364 34756 2540 34796
rect 3679 34756 3688 34796
rect 3728 34756 3770 34796
rect 3810 34756 3852 34796
rect 3892 34756 3934 34796
rect 3974 34756 4016 34796
rect 4056 34756 4065 34796
rect 4675 34756 4684 34796
rect 4724 34756 4876 34796
rect 4916 34756 7372 34796
rect 7412 34756 7421 34796
rect 9379 34756 9388 34796
rect 9428 34756 14668 34796
rect 14708 34756 14717 34796
rect 16492 34756 17068 34796
rect 17108 34756 17117 34796
rect 18414 34756 18508 34796
rect 18548 34756 18557 34796
rect 18799 34756 18808 34796
rect 18848 34756 18890 34796
rect 18930 34756 18972 34796
rect 19012 34756 19054 34796
rect 19094 34756 19136 34796
rect 19176 34756 19185 34796
rect 0 34712 80 34732
rect 2500 34712 2540 34756
rect 6595 34712 6653 34713
rect 15427 34712 15485 34713
rect 16492 34712 16532 34756
rect 18499 34755 18557 34756
rect 0 34672 2188 34712
rect 2228 34672 2237 34712
rect 2500 34672 5356 34712
rect 5396 34672 5405 34712
rect 6595 34672 6604 34712
rect 6644 34672 6892 34712
rect 6932 34672 6941 34712
rect 8419 34672 8428 34712
rect 8468 34672 14572 34712
rect 14612 34672 14621 34712
rect 15427 34672 15436 34712
rect 15476 34672 15724 34712
rect 15764 34672 16532 34712
rect 16588 34672 19372 34712
rect 19412 34672 19852 34712
rect 19892 34672 19901 34712
rect 0 34652 80 34672
rect 6595 34671 6653 34672
rect 15427 34671 15485 34672
rect 16588 34629 16628 34672
rect 4003 34628 4061 34629
rect 4483 34628 4541 34629
rect 16579 34628 16637 34629
rect 19555 34628 19613 34629
rect 1603 34588 1612 34628
rect 1652 34588 2764 34628
rect 2804 34588 2813 34628
rect 3235 34588 3244 34628
rect 3284 34588 4012 34628
rect 4052 34588 4492 34628
rect 4532 34588 4541 34628
rect 4003 34587 4061 34588
rect 4483 34587 4541 34588
rect 6892 34588 7180 34628
rect 7220 34588 7229 34628
rect 9571 34588 9580 34628
rect 9620 34588 16588 34628
rect 16628 34588 16637 34628
rect 17635 34588 17644 34628
rect 17684 34588 18028 34628
rect 18068 34588 18508 34628
rect 18548 34588 19564 34628
rect 19604 34588 19613 34628
rect 1699 34544 1757 34545
rect 6499 34544 6557 34545
rect 940 34504 1708 34544
rect 1748 34504 6508 34544
rect 6548 34504 6557 34544
rect 0 34376 80 34396
rect 940 34376 980 34504
rect 1699 34503 1757 34504
rect 6499 34503 6557 34504
rect 6892 34460 6932 34588
rect 16579 34587 16637 34588
rect 19555 34587 19613 34588
rect 6979 34504 6988 34544
rect 7028 34504 8140 34544
rect 8180 34504 8189 34544
rect 8323 34504 8332 34544
rect 8372 34504 10924 34544
rect 10964 34504 10973 34544
rect 11779 34504 11788 34544
rect 11828 34504 12076 34544
rect 12116 34504 12125 34544
rect 13699 34504 13708 34544
rect 13748 34504 18412 34544
rect 18452 34504 18461 34544
rect 18691 34504 18700 34544
rect 18740 34504 19948 34544
rect 19988 34504 19997 34544
rect 8899 34460 8957 34461
rect 19747 34460 19805 34461
rect 1027 34420 1036 34460
rect 1076 34420 1420 34460
rect 1460 34420 1469 34460
rect 2380 34420 3148 34460
rect 3188 34420 3197 34460
rect 6691 34420 6700 34460
rect 6740 34420 8908 34460
rect 8948 34420 8957 34460
rect 11011 34420 11020 34460
rect 11060 34420 16244 34460
rect 19075 34420 19084 34460
rect 19124 34420 19756 34460
rect 19796 34420 19805 34460
rect 1603 34376 1661 34377
rect 2380 34376 2420 34420
rect 8899 34419 8957 34420
rect 4099 34376 4157 34377
rect 6883 34376 6941 34377
rect 7363 34376 7421 34377
rect 7651 34376 7709 34377
rect 9187 34376 9245 34377
rect 0 34336 980 34376
rect 1518 34336 1612 34376
rect 1652 34336 1661 34376
rect 2371 34336 2380 34376
rect 2420 34336 2429 34376
rect 2659 34336 2668 34376
rect 2708 34336 3436 34376
rect 3476 34336 3485 34376
rect 3907 34336 3916 34376
rect 3956 34336 4108 34376
rect 4148 34336 4157 34376
rect 4579 34336 4588 34376
rect 4628 34336 6220 34376
rect 6260 34336 6508 34376
rect 6548 34336 6557 34376
rect 6883 34336 6892 34376
rect 6932 34336 7180 34376
rect 7220 34336 7372 34376
rect 7412 34336 7421 34376
rect 7566 34336 7660 34376
rect 7700 34336 7709 34376
rect 8227 34336 8236 34376
rect 8276 34336 8285 34376
rect 9102 34336 9196 34376
rect 9236 34336 9245 34376
rect 0 34316 80 34336
rect 1603 34335 1661 34336
rect 4099 34335 4157 34336
rect 6883 34335 6941 34336
rect 7363 34335 7421 34336
rect 7651 34335 7709 34336
rect 5347 34292 5405 34293
rect 8236 34292 8276 34336
rect 9187 34335 9245 34336
rect 12355 34376 12413 34377
rect 13507 34376 13565 34377
rect 14467 34376 14525 34377
rect 12355 34336 12364 34376
rect 12404 34336 12460 34376
rect 12500 34336 12509 34376
rect 13123 34336 13132 34376
rect 13172 34336 13516 34376
rect 13556 34336 13565 34376
rect 14382 34336 14476 34376
rect 14516 34336 14525 34376
rect 12355 34335 12413 34336
rect 13507 34335 13565 34336
rect 14467 34335 14525 34336
rect 15619 34376 15677 34377
rect 16204 34376 16244 34420
rect 19747 34419 19805 34420
rect 18211 34376 18269 34377
rect 15619 34336 15628 34376
rect 15668 34336 15916 34376
rect 15956 34336 15965 34376
rect 16195 34336 16204 34376
rect 16244 34336 16253 34376
rect 17443 34336 17452 34376
rect 17492 34336 18220 34376
rect 18260 34336 18269 34376
rect 19267 34336 19276 34376
rect 19316 34336 19660 34376
rect 19700 34336 19709 34376
rect 15619 34335 15677 34336
rect 18211 34335 18269 34336
rect 18403 34292 18461 34293
rect 1507 34252 1516 34292
rect 1556 34252 2188 34292
rect 2228 34252 2237 34292
rect 2851 34252 2860 34292
rect 2900 34252 5356 34292
rect 5396 34252 5405 34292
rect 6883 34252 6892 34292
rect 6932 34252 8276 34292
rect 8803 34252 8812 34292
rect 8852 34252 10444 34292
rect 10484 34252 10493 34292
rect 12067 34252 12076 34292
rect 12116 34252 15820 34292
rect 15860 34252 15869 34292
rect 18318 34252 18412 34292
rect 18452 34252 18461 34292
rect 5347 34251 5405 34252
rect 18403 34251 18461 34252
rect 10051 34208 10109 34209
rect 13315 34208 13373 34209
rect 20140 34208 20180 35008
rect 21424 34988 21504 35008
rect 21424 34544 21504 34564
rect 20611 34504 20620 34544
rect 20660 34504 21504 34544
rect 21424 34484 21504 34504
rect 4195 34168 4204 34208
rect 4244 34168 4492 34208
rect 4532 34168 4541 34208
rect 4963 34168 4972 34208
rect 5012 34168 8716 34208
rect 8756 34168 8765 34208
rect 10051 34168 10060 34208
rect 10100 34168 10828 34208
rect 10868 34168 13324 34208
rect 13364 34168 13373 34208
rect 13603 34168 13612 34208
rect 13652 34168 20180 34208
rect 10051 34167 10109 34168
rect 13315 34167 13373 34168
rect 14179 34124 14237 34125
rect 16003 34124 16061 34125
rect 17827 34124 17885 34125
rect 1795 34084 1804 34124
rect 1844 34084 2284 34124
rect 2324 34084 2333 34124
rect 2500 34084 4684 34124
rect 4724 34084 4733 34124
rect 6211 34084 6220 34124
rect 6260 34084 6412 34124
rect 6452 34084 7756 34124
rect 7796 34084 10100 34124
rect 10435 34084 10444 34124
rect 10484 34084 12076 34124
rect 12116 34084 12125 34124
rect 12643 34084 12652 34124
rect 12692 34084 13708 34124
rect 13748 34084 13757 34124
rect 14094 34084 14188 34124
rect 14228 34084 14237 34124
rect 0 34040 80 34060
rect 2500 34040 2540 34084
rect 7267 34040 7325 34041
rect 0 34000 2540 34040
rect 3139 34000 3148 34040
rect 3188 34000 4780 34040
rect 4820 34000 4829 34040
rect 4919 34000 4928 34040
rect 4968 34000 5010 34040
rect 5050 34000 5092 34040
rect 5132 34000 5174 34040
rect 5214 34000 5256 34040
rect 5296 34000 5305 34040
rect 5443 34000 5452 34040
rect 5492 34000 7124 34040
rect 7182 34000 7276 34040
rect 7316 34000 7325 34040
rect 7939 34000 7948 34040
rect 7988 34000 8028 34040
rect 8995 34000 9004 34040
rect 9044 34000 9292 34040
rect 9332 34000 9341 34040
rect 0 33980 80 34000
rect 2947 33956 3005 33957
rect 7084 33956 7124 34000
rect 7267 33999 7325 34000
rect 7948 33956 7988 34000
rect 2179 33916 2188 33956
rect 2228 33916 2572 33956
rect 2612 33916 2621 33956
rect 2947 33916 2956 33956
rect 2996 33916 3628 33956
rect 3668 33916 3677 33956
rect 3811 33916 3820 33956
rect 3860 33916 4684 33956
rect 4724 33916 6316 33956
rect 6356 33916 6365 33956
rect 7084 33916 8332 33956
rect 8372 33916 8381 33956
rect 8611 33916 8620 33956
rect 8660 33916 8812 33956
rect 8852 33916 8861 33956
rect 2947 33915 3005 33916
rect 1411 33872 1469 33873
rect 10060 33872 10100 34084
rect 14179 34083 14237 34084
rect 14284 34084 14900 34124
rect 14947 34084 14956 34124
rect 14996 34084 15340 34124
rect 15380 34084 15572 34124
rect 14284 34040 14324 34084
rect 14860 34040 14900 34084
rect 15043 34040 15101 34041
rect 15427 34040 15485 34041
rect 13891 34000 13900 34040
rect 13940 34000 14324 34040
rect 14572 34000 14668 34040
rect 14708 34000 14717 34040
rect 14860 34000 15052 34040
rect 15092 34000 15101 34040
rect 15342 34000 15436 34040
rect 15476 34000 15485 34040
rect 15532 34040 15572 34084
rect 16003 34084 16012 34124
rect 16052 34084 16396 34124
rect 16436 34084 16445 34124
rect 17742 34084 17836 34124
rect 17876 34084 17885 34124
rect 16003 34083 16061 34084
rect 17827 34083 17885 34084
rect 17932 34084 18452 34124
rect 16483 34040 16541 34041
rect 15532 34000 16492 34040
rect 16532 34000 16541 34040
rect 11107 33956 11165 33957
rect 14572 33956 14612 34000
rect 15043 33999 15101 34000
rect 15427 33999 15485 34000
rect 16483 33999 16541 34000
rect 17635 34040 17693 34041
rect 17932 34040 17972 34084
rect 18412 34040 18452 34084
rect 21424 34040 21504 34060
rect 17635 34000 17644 34040
rect 17684 34000 17972 34040
rect 18019 34000 18028 34040
rect 18068 34000 18316 34040
rect 18356 34000 18365 34040
rect 18412 34000 18644 34040
rect 20039 34000 20048 34040
rect 20088 34000 20130 34040
rect 20170 34000 20212 34040
rect 20252 34000 20294 34040
rect 20334 34000 20376 34040
rect 20416 34000 20425 34040
rect 20803 34000 20812 34040
rect 20852 34000 21504 34040
rect 17635 33999 17693 34000
rect 18499 33956 18557 33957
rect 11107 33916 11116 33956
rect 11156 33916 12844 33956
rect 12884 33916 12893 33956
rect 13795 33916 13804 33956
rect 13844 33916 14612 33956
rect 14764 33916 18508 33956
rect 18548 33916 18557 33956
rect 18604 33956 18644 34000
rect 21424 33980 21504 34000
rect 18604 33916 19948 33956
rect 19988 33916 19997 33956
rect 11107 33915 11165 33916
rect 14764 33872 14804 33916
rect 18499 33915 18557 33916
rect 1326 33832 1420 33872
rect 1460 33832 1469 33872
rect 2275 33832 2284 33872
rect 2324 33832 4108 33872
rect 4148 33832 4157 33872
rect 6499 33832 6508 33872
rect 6548 33832 7564 33872
rect 7604 33832 7756 33872
rect 7796 33832 7805 33872
rect 10051 33832 10060 33872
rect 10100 33832 10109 33872
rect 10243 33832 10252 33872
rect 10292 33832 10301 33872
rect 11587 33832 11596 33872
rect 11636 33832 14804 33872
rect 14851 33832 14860 33872
rect 14900 33832 18124 33872
rect 18164 33832 18173 33872
rect 1411 33831 1469 33832
rect 2755 33788 2813 33789
rect 8707 33788 8765 33789
rect 1324 33748 2764 33788
rect 2804 33748 2813 33788
rect 2947 33748 2956 33788
rect 2996 33748 8428 33788
rect 8468 33748 8477 33788
rect 8707 33748 8716 33788
rect 8756 33748 8812 33788
rect 8852 33748 9868 33788
rect 9908 33748 9917 33788
rect 0 33704 80 33724
rect 1219 33704 1277 33705
rect 0 33664 1228 33704
rect 1268 33664 1277 33704
rect 0 33644 80 33664
rect 1219 33663 1277 33664
rect 1324 33620 1364 33748
rect 2755 33747 2813 33748
rect 8707 33747 8765 33748
rect 9955 33704 10013 33705
rect 10252 33704 10292 33832
rect 10540 33748 11020 33788
rect 11060 33748 11069 33788
rect 12835 33748 12844 33788
rect 12884 33748 16436 33788
rect 10540 33704 10580 33748
rect 11779 33704 11837 33705
rect 14275 33704 14333 33705
rect 5251 33664 5260 33704
rect 5300 33664 5644 33704
rect 5684 33664 9580 33704
rect 9620 33664 9629 33704
rect 9955 33664 9964 33704
rect 10004 33664 10292 33704
rect 10531 33664 10540 33704
rect 10580 33664 10589 33704
rect 11683 33664 11692 33704
rect 11732 33664 11788 33704
rect 11828 33664 11837 33704
rect 14190 33664 14284 33704
rect 14324 33664 14333 33704
rect 9955 33663 10013 33664
rect 11779 33663 11837 33664
rect 14275 33663 14333 33664
rect 15235 33704 15293 33705
rect 16003 33704 16061 33705
rect 15235 33664 15244 33704
rect 15284 33664 15532 33704
rect 15572 33664 16012 33704
rect 16052 33664 16061 33704
rect 16396 33704 16436 33748
rect 18892 33748 20524 33788
rect 20564 33748 20573 33788
rect 18115 33704 18173 33705
rect 16396 33664 17836 33704
rect 17876 33664 17885 33704
rect 18115 33664 18124 33704
rect 18164 33664 18796 33704
rect 18836 33664 18845 33704
rect 15235 33663 15293 33664
rect 16003 33663 16061 33664
rect 18115 33663 18173 33664
rect 259 33580 268 33620
rect 308 33580 1132 33620
rect 1172 33580 1364 33620
rect 2755 33620 2813 33621
rect 5539 33620 5597 33621
rect 13891 33620 13949 33621
rect 16291 33620 16349 33621
rect 2755 33580 2764 33620
rect 2804 33580 3764 33620
rect 3811 33580 3820 33620
rect 3860 33580 4876 33620
rect 4916 33580 4925 33620
rect 5347 33580 5356 33620
rect 5396 33580 5548 33620
rect 5588 33580 5597 33620
rect 2755 33579 2813 33580
rect 3619 33536 3677 33537
rect 3523 33496 3532 33536
rect 3572 33496 3628 33536
rect 3668 33496 3677 33536
rect 3724 33536 3764 33580
rect 5539 33579 5597 33580
rect 5644 33580 6412 33620
rect 6452 33580 6461 33620
rect 6787 33580 6796 33620
rect 6836 33580 11212 33620
rect 11252 33580 13900 33620
rect 13940 33580 13949 33620
rect 14179 33580 14188 33620
rect 14228 33580 14380 33620
rect 14420 33580 15148 33620
rect 15188 33580 15197 33620
rect 16291 33580 16300 33620
rect 16340 33580 18124 33620
rect 18164 33580 18173 33620
rect 5644 33536 5684 33580
rect 13891 33579 13949 33580
rect 16291 33579 16349 33580
rect 7171 33536 7229 33537
rect 18892 33536 18932 33748
rect 19843 33620 19901 33621
rect 19758 33580 19852 33620
rect 19892 33580 19901 33620
rect 19843 33579 19901 33580
rect 19459 33536 19517 33537
rect 3724 33496 5684 33536
rect 5731 33496 5740 33536
rect 5780 33496 6700 33536
rect 6740 33496 6749 33536
rect 7171 33496 7180 33536
rect 7220 33496 7276 33536
rect 7316 33496 7325 33536
rect 9859 33496 9868 33536
rect 9908 33496 11596 33536
rect 11636 33496 11645 33536
rect 14563 33496 14572 33536
rect 14612 33496 14621 33536
rect 16771 33496 16780 33536
rect 16820 33496 18932 33536
rect 19374 33496 19468 33536
rect 19508 33496 19517 33536
rect 3619 33495 3677 33496
rect 7171 33495 7229 33496
rect 2947 33452 3005 33453
rect 11299 33452 11357 33453
rect 2947 33412 2956 33452
rect 2996 33412 6988 33452
rect 7028 33412 7037 33452
rect 8227 33412 8236 33452
rect 8276 33412 10060 33452
rect 10100 33412 10109 33452
rect 11107 33412 11116 33452
rect 11156 33412 11308 33452
rect 11348 33412 11357 33452
rect 12835 33412 12844 33452
rect 12884 33412 13804 33452
rect 13844 33412 14380 33452
rect 14420 33412 14429 33452
rect 2947 33411 3005 33412
rect 11299 33411 11357 33412
rect 0 33368 80 33388
rect 3427 33368 3485 33369
rect 0 33328 3436 33368
rect 3476 33328 3485 33368
rect 0 33308 80 33328
rect 3427 33327 3485 33328
rect 3532 33328 4396 33368
rect 4436 33328 4445 33368
rect 4771 33328 4780 33368
rect 4820 33328 6220 33368
rect 6260 33328 11596 33368
rect 11636 33328 11645 33368
rect 3532 33284 3572 33328
rect 13123 33284 13181 33285
rect 14467 33284 14525 33285
rect 2851 33244 2860 33284
rect 2900 33244 3052 33284
rect 3092 33244 3101 33284
rect 3427 33244 3436 33284
rect 3476 33244 3572 33284
rect 3679 33244 3688 33284
rect 3728 33244 3770 33284
rect 3810 33244 3852 33284
rect 3892 33244 3934 33284
rect 3974 33244 4016 33284
rect 4056 33244 4065 33284
rect 4204 33244 9004 33284
rect 9044 33244 9053 33284
rect 9667 33244 9676 33284
rect 9716 33244 13132 33284
rect 13172 33244 13181 33284
rect 14179 33244 14188 33284
rect 14228 33244 14476 33284
rect 14516 33244 14525 33284
rect 14572 33284 14612 33496
rect 19459 33495 19517 33496
rect 20803 33536 20861 33537
rect 21424 33536 21504 33556
rect 20803 33496 20812 33536
rect 20852 33496 21504 33536
rect 20803 33495 20861 33496
rect 21424 33476 21504 33496
rect 20611 33452 20669 33453
rect 20035 33412 20044 33452
rect 20084 33412 20620 33452
rect 20660 33412 20669 33452
rect 20611 33411 20669 33412
rect 18211 33284 18269 33285
rect 14572 33244 15340 33284
rect 15380 33244 15389 33284
rect 16675 33244 16684 33284
rect 16724 33244 17260 33284
rect 17300 33244 17309 33284
rect 18211 33244 18220 33284
rect 18260 33244 18700 33284
rect 18740 33244 18749 33284
rect 18799 33244 18808 33284
rect 18848 33244 18890 33284
rect 18930 33244 18972 33284
rect 19012 33244 19054 33284
rect 19094 33244 19136 33284
rect 19176 33244 19185 33284
rect 1219 33200 1277 33201
rect 1134 33160 1228 33200
rect 1268 33160 1277 33200
rect 1219 33159 1277 33160
rect 4204 33116 4244 33244
rect 13123 33243 13181 33244
rect 14467 33243 14525 33244
rect 18211 33243 18269 33244
rect 10627 33200 10685 33201
rect 6307 33160 6316 33200
rect 6356 33160 8620 33200
rect 8660 33160 8669 33200
rect 10627 33160 10636 33200
rect 10676 33160 12652 33200
rect 12692 33160 16396 33200
rect 16436 33160 16445 33200
rect 18595 33160 18604 33200
rect 18644 33160 20044 33200
rect 20084 33160 20093 33200
rect 10627 33159 10685 33160
rect 15907 33116 15965 33117
rect 19267 33116 19325 33117
rect 1228 33076 3764 33116
rect 3811 33076 3820 33116
rect 3860 33076 4244 33116
rect 4291 33076 4300 33116
rect 4340 33076 5972 33116
rect 6595 33076 6604 33116
rect 6644 33076 7756 33116
rect 7796 33076 7805 33116
rect 7939 33076 7948 33116
rect 7988 33076 8332 33116
rect 8372 33076 9004 33116
rect 9044 33076 9053 33116
rect 10243 33076 10252 33116
rect 10292 33076 10301 33116
rect 14467 33076 14476 33116
rect 14516 33076 15436 33116
rect 15476 33076 15485 33116
rect 15907 33076 15916 33116
rect 15956 33076 17932 33116
rect 17972 33076 17981 33116
rect 19182 33076 19276 33116
rect 19316 33076 19325 33116
rect 0 33032 80 33052
rect 1228 33032 1268 33076
rect 3331 33032 3389 33033
rect 0 32992 1268 33032
rect 2947 32992 2956 33032
rect 2996 32992 3036 33032
rect 3235 32992 3244 33032
rect 3284 32992 3340 33032
rect 3380 32992 3389 33032
rect 3724 33032 3764 33076
rect 4195 33032 4253 33033
rect 5932 33032 5972 33076
rect 10252 33032 10292 33076
rect 15907 33075 15965 33076
rect 19267 33075 19325 33076
rect 17635 33032 17693 33033
rect 3724 32992 4204 33032
rect 4244 32992 4253 33032
rect 5923 32992 5932 33032
rect 5972 32992 5981 33032
rect 6028 32992 10292 33032
rect 14659 32992 14668 33032
rect 14708 32992 16588 33032
rect 16628 32992 16637 33032
rect 17251 32992 17260 33032
rect 17300 32992 17644 33032
rect 17684 32992 17693 33032
rect 0 32972 80 32992
rect 2956 32948 2996 32992
rect 3331 32991 3389 32992
rect 4195 32991 4253 32992
rect 3907 32948 3965 32949
rect 2500 32908 3916 32948
rect 3956 32908 3965 32948
rect 931 32864 989 32865
rect 2500 32864 2540 32908
rect 3907 32907 3965 32908
rect 4099 32948 4157 32949
rect 6028 32948 6068 32992
rect 17635 32991 17693 32992
rect 20707 33032 20765 33033
rect 21424 33032 21504 33052
rect 20707 32992 20716 33032
rect 20756 32992 21504 33032
rect 20707 32991 20765 32992
rect 21424 32972 21504 32992
rect 15139 32948 15197 32949
rect 16675 32948 16733 32949
rect 4099 32908 4108 32948
rect 4148 32908 4242 32948
rect 4291 32908 4300 32948
rect 4340 32908 6068 32948
rect 7363 32908 7372 32948
rect 7412 32908 9812 32948
rect 10339 32908 10348 32948
rect 10388 32908 13804 32948
rect 13844 32908 13853 32948
rect 15139 32908 15148 32948
rect 15188 32908 15820 32948
rect 15860 32908 15869 32948
rect 16675 32908 16684 32948
rect 16724 32908 18028 32948
rect 18068 32908 18077 32948
rect 20131 32908 20140 32948
rect 20180 32908 20908 32948
rect 20948 32908 20957 32948
rect 4099 32907 4157 32908
rect 4771 32864 4829 32865
rect 7555 32864 7613 32865
rect 9187 32864 9245 32865
rect 9772 32864 9812 32908
rect 15139 32907 15197 32908
rect 16675 32907 16733 32908
rect 19555 32864 19613 32865
rect 931 32824 940 32864
rect 980 32824 2540 32864
rect 3427 32824 3436 32864
rect 3476 32824 4588 32864
rect 4628 32824 4637 32864
rect 4771 32824 4780 32864
rect 4820 32824 5740 32864
rect 5780 32824 6316 32864
rect 6356 32824 6365 32864
rect 7470 32824 7564 32864
rect 7604 32824 7613 32864
rect 9102 32824 9196 32864
rect 9236 32824 9388 32864
rect 9428 32824 9437 32864
rect 9667 32824 9676 32864
rect 9716 32824 9725 32864
rect 9772 32824 10540 32864
rect 10580 32824 10589 32864
rect 10828 32824 11884 32864
rect 11924 32824 11933 32864
rect 13987 32824 13996 32864
rect 14036 32824 15052 32864
rect 15092 32824 15244 32864
rect 15284 32824 15916 32864
rect 15956 32824 15965 32864
rect 16867 32824 16876 32864
rect 16916 32824 18604 32864
rect 18644 32824 18653 32864
rect 19555 32824 19564 32864
rect 19604 32824 19756 32864
rect 19796 32824 19805 32864
rect 20035 32824 20044 32864
rect 20084 32824 20620 32864
rect 20660 32824 20669 32864
rect 931 32823 989 32824
rect 4771 32823 4829 32824
rect 7555 32823 7613 32824
rect 9187 32823 9245 32824
rect 4291 32780 4349 32781
rect 9676 32780 9716 32824
rect 4291 32740 4300 32780
rect 4340 32740 4492 32780
rect 4532 32740 4541 32780
rect 4771 32740 4780 32780
rect 4820 32740 9716 32780
rect 4291 32739 4349 32740
rect 0 32696 80 32716
rect 2947 32696 3005 32697
rect 10828 32696 10868 32824
rect 19555 32823 19613 32824
rect 10915 32780 10973 32781
rect 12355 32780 12413 32781
rect 13027 32780 13085 32781
rect 10915 32740 10924 32780
rect 10964 32740 11020 32780
rect 11060 32740 11069 32780
rect 12355 32740 12364 32780
rect 12404 32740 12460 32780
rect 12500 32740 12509 32780
rect 13027 32740 13036 32780
rect 13076 32740 17068 32780
rect 17108 32740 17117 32780
rect 17827 32740 17836 32780
rect 17876 32740 18316 32780
rect 18356 32740 18365 32780
rect 19267 32740 19276 32780
rect 19316 32740 20140 32780
rect 20180 32740 20189 32780
rect 10915 32739 10973 32740
rect 12355 32739 12413 32740
rect 13027 32739 13085 32740
rect 0 32656 1268 32696
rect 2275 32656 2284 32696
rect 2324 32656 2764 32696
rect 2804 32656 2813 32696
rect 2862 32656 2956 32696
rect 2996 32656 3005 32696
rect 3619 32656 3628 32696
rect 3668 32656 4204 32696
rect 4244 32656 4396 32696
rect 4436 32656 4445 32696
rect 4867 32656 4876 32696
rect 4916 32656 8428 32696
rect 8468 32656 8477 32696
rect 10051 32656 10060 32696
rect 10100 32656 10444 32696
rect 10484 32656 10868 32696
rect 11779 32696 11837 32697
rect 15427 32696 15485 32697
rect 16291 32696 16349 32697
rect 11779 32656 11788 32696
rect 11828 32656 11884 32696
rect 11924 32656 11933 32696
rect 14659 32656 14668 32696
rect 14708 32656 15436 32696
rect 15476 32656 15485 32696
rect 15619 32656 15628 32696
rect 15668 32656 16300 32696
rect 16340 32656 16349 32696
rect 0 32636 80 32656
rect 1228 32528 1268 32656
rect 2947 32655 3005 32656
rect 11779 32655 11837 32656
rect 15427 32655 15485 32656
rect 16291 32655 16349 32656
rect 10051 32612 10109 32613
rect 15619 32612 15677 32613
rect 1315 32572 1324 32612
rect 1364 32572 8524 32612
rect 8564 32572 8573 32612
rect 10051 32572 10060 32612
rect 10100 32572 15628 32612
rect 15668 32572 15677 32612
rect 10051 32571 10109 32572
rect 15619 32571 15677 32572
rect 18019 32612 18077 32613
rect 18019 32572 18028 32612
rect 18068 32572 18604 32612
rect 18644 32572 18653 32612
rect 18019 32571 18077 32572
rect 4291 32528 4349 32529
rect 15811 32528 15869 32529
rect 19555 32528 19613 32529
rect 20995 32528 21053 32529
rect 21424 32528 21504 32548
rect 1228 32488 4300 32528
rect 4340 32488 4349 32528
rect 4919 32488 4928 32528
rect 4968 32488 5010 32528
rect 5050 32488 5092 32528
rect 5132 32488 5174 32528
rect 5214 32488 5256 32528
rect 5296 32488 5305 32528
rect 8611 32488 8620 32528
rect 8660 32488 9580 32528
rect 9620 32488 9868 32528
rect 9908 32488 9917 32528
rect 10723 32488 10732 32528
rect 10772 32488 15820 32528
rect 15860 32488 15869 32528
rect 18115 32488 18124 32528
rect 18164 32488 19564 32528
rect 19604 32488 19613 32528
rect 20039 32488 20048 32528
rect 20088 32488 20130 32528
rect 20170 32488 20212 32528
rect 20252 32488 20294 32528
rect 20334 32488 20376 32528
rect 20416 32488 20425 32528
rect 20995 32488 21004 32528
rect 21044 32488 21504 32528
rect 4291 32487 4349 32488
rect 15811 32487 15869 32488
rect 19555 32487 19613 32488
rect 20995 32487 21053 32488
rect 21424 32468 21504 32488
rect 1123 32444 1181 32445
rect 8419 32444 8477 32445
rect 8707 32444 8765 32445
rect 1123 32404 1132 32444
rect 1172 32404 1708 32444
rect 1748 32404 1757 32444
rect 3043 32404 3052 32444
rect 3092 32404 3101 32444
rect 3235 32404 3244 32444
rect 3284 32404 6220 32444
rect 6260 32404 7564 32444
rect 7604 32404 7613 32444
rect 8419 32404 8428 32444
rect 8468 32404 8716 32444
rect 8756 32404 10772 32444
rect 11299 32404 11308 32444
rect 11348 32404 12692 32444
rect 12739 32404 12748 32444
rect 12788 32404 16684 32444
rect 16724 32404 16733 32444
rect 1123 32403 1181 32404
rect 0 32360 80 32380
rect 2083 32360 2141 32361
rect 0 32320 2092 32360
rect 2132 32320 2141 32360
rect 2563 32320 2572 32360
rect 2612 32320 2956 32360
rect 2996 32320 3005 32360
rect 0 32300 80 32320
rect 2083 32319 2141 32320
rect 3052 32276 3092 32404
rect 8419 32403 8477 32404
rect 8707 32403 8765 32404
rect 3907 32360 3965 32361
rect 10732 32360 10772 32404
rect 12652 32361 12692 32404
rect 12643 32360 12701 32361
rect 12931 32360 12989 32361
rect 14947 32360 15005 32361
rect 3139 32320 3148 32360
rect 3188 32320 3724 32360
rect 3764 32320 3773 32360
rect 3888 32320 3916 32360
rect 3956 32320 4012 32360
rect 4052 32320 4780 32360
rect 4820 32320 4829 32360
rect 6691 32320 6700 32360
rect 6740 32320 10636 32360
rect 10676 32320 10685 32360
rect 10732 32320 12460 32360
rect 12500 32320 12509 32360
rect 12643 32320 12652 32360
rect 12692 32320 12940 32360
rect 12980 32320 12989 32360
rect 14755 32320 14764 32360
rect 14804 32320 14956 32360
rect 14996 32320 15005 32360
rect 3907 32319 3965 32320
rect 12643 32319 12701 32320
rect 12931 32319 12989 32320
rect 14947 32319 15005 32320
rect 15427 32360 15485 32361
rect 15907 32360 15965 32361
rect 18499 32360 18557 32361
rect 15427 32320 15436 32360
rect 15476 32320 15724 32360
rect 15764 32320 15773 32360
rect 15822 32320 15916 32360
rect 15956 32320 15965 32360
rect 18403 32320 18412 32360
rect 18452 32320 18508 32360
rect 18548 32320 18557 32360
rect 15427 32319 15485 32320
rect 15907 32319 15965 32320
rect 18499 32319 18557 32320
rect 12259 32276 12317 32277
rect 3052 32236 5356 32276
rect 5396 32236 5405 32276
rect 6403 32236 6412 32276
rect 6452 32236 11308 32276
rect 11348 32236 11357 32276
rect 12174 32236 12268 32276
rect 12308 32236 12317 32276
rect 13795 32236 13804 32276
rect 13844 32236 21004 32276
rect 21044 32236 21053 32276
rect 12259 32235 12317 32236
rect 2083 32192 2141 32193
rect 8323 32192 8381 32193
rect 9571 32192 9629 32193
rect 14467 32192 14525 32193
rect 1998 32152 2092 32192
rect 2132 32152 2141 32192
rect 2755 32152 2764 32192
rect 2804 32152 3916 32192
rect 3956 32152 3965 32192
rect 8238 32152 8332 32192
rect 8372 32152 8381 32192
rect 8515 32152 8524 32192
rect 8564 32152 9388 32192
rect 9428 32152 9437 32192
rect 9571 32152 9580 32192
rect 9620 32152 11500 32192
rect 11540 32152 12364 32192
rect 12404 32152 12413 32192
rect 14382 32152 14476 32192
rect 14516 32152 14525 32192
rect 2083 32151 2141 32152
rect 8323 32151 8381 32152
rect 9571 32151 9629 32152
rect 14467 32151 14525 32152
rect 15523 32192 15581 32193
rect 18691 32192 18749 32193
rect 15523 32152 15532 32192
rect 15572 32152 15724 32192
rect 15764 32152 15773 32192
rect 16963 32152 16972 32192
rect 17012 32152 17452 32192
rect 17492 32152 18700 32192
rect 18740 32152 19468 32192
rect 19508 32152 19517 32192
rect 15523 32151 15581 32152
rect 18691 32151 18749 32152
rect 1507 32108 1565 32109
rect 10915 32108 10973 32109
rect 18211 32108 18269 32109
rect 1422 32068 1516 32108
rect 1556 32068 1565 32108
rect 7843 32068 7852 32108
rect 7892 32068 8140 32108
rect 8180 32068 8189 32108
rect 10627 32068 10636 32108
rect 10676 32068 10924 32108
rect 10964 32068 18220 32108
rect 18260 32068 18269 32108
rect 1507 32067 1565 32068
rect 10915 32067 10973 32068
rect 18211 32067 18269 32068
rect 18892 32068 19852 32108
rect 19892 32068 19901 32108
rect 0 32024 80 32044
rect 739 32024 797 32025
rect 4099 32024 4157 32025
rect 14947 32024 15005 32025
rect 15139 32024 15197 32025
rect 0 31984 748 32024
rect 788 31984 797 32024
rect 1411 31984 1420 32024
rect 1460 31984 1708 32024
rect 1748 31984 1757 32024
rect 4099 31984 4108 32024
rect 4148 31984 8044 32024
rect 8084 31984 8093 32024
rect 8611 31984 8620 32024
rect 8660 31984 9580 32024
rect 9620 31984 9629 32024
rect 14862 31984 14956 32024
rect 14996 31984 15005 32024
rect 15054 31984 15148 32024
rect 15188 31984 15197 32024
rect 0 31964 80 31984
rect 739 31983 797 31984
rect 4099 31983 4157 31984
rect 14947 31983 15005 31984
rect 15139 31983 15197 31984
rect 15331 32024 15389 32025
rect 18892 32024 18932 32068
rect 15331 31984 15340 32024
rect 15380 31984 18932 32024
rect 19651 32024 19709 32025
rect 21424 32024 21504 32044
rect 19651 31984 19660 32024
rect 19700 31984 21504 32024
rect 15331 31983 15389 31984
rect 19651 31983 19709 31984
rect 21424 31964 21504 31984
rect 6979 31940 7037 31941
rect 19939 31940 19997 31941
rect 355 31900 364 31940
rect 404 31900 4780 31940
rect 4820 31900 4916 31940
rect 2659 31856 2717 31857
rect 4876 31856 4916 31900
rect 6979 31900 6988 31940
rect 7028 31900 17836 31940
rect 17876 31900 17885 31940
rect 19939 31900 19948 31940
rect 19988 31900 20044 31940
rect 20084 31900 20093 31940
rect 6979 31899 7037 31900
rect 19939 31899 19997 31900
rect 9091 31856 9149 31857
rect 10051 31856 10109 31857
rect 2563 31816 2572 31856
rect 2612 31816 2668 31856
rect 2708 31816 2717 31856
rect 3043 31816 3052 31856
rect 3092 31816 4820 31856
rect 4876 31816 9100 31856
rect 9140 31816 10060 31856
rect 10100 31816 10109 31856
rect 2659 31815 2717 31816
rect 4780 31772 4820 31816
rect 9091 31815 9149 31816
rect 10051 31815 10109 31816
rect 12643 31856 12701 31857
rect 12643 31816 12652 31856
rect 12692 31816 16204 31856
rect 16244 31816 16253 31856
rect 12643 31815 12701 31816
rect 9955 31772 10013 31773
rect 14947 31772 15005 31773
rect 1219 31732 1228 31772
rect 1268 31732 2956 31772
rect 2996 31732 3005 31772
rect 3679 31732 3688 31772
rect 3728 31732 3770 31772
rect 3810 31732 3852 31772
rect 3892 31732 3934 31772
rect 3974 31732 4016 31772
rect 4056 31732 4065 31772
rect 4780 31732 9964 31772
rect 10004 31732 10636 31772
rect 10676 31732 10685 31772
rect 11587 31732 11596 31772
rect 11636 31732 14956 31772
rect 14996 31732 17068 31772
rect 17108 31732 17117 31772
rect 18799 31732 18808 31772
rect 18848 31732 18890 31772
rect 18930 31732 18972 31772
rect 19012 31732 19054 31772
rect 19094 31732 19136 31772
rect 19176 31732 19185 31772
rect 9955 31731 10013 31732
rect 14947 31731 15005 31732
rect 0 31688 80 31708
rect 3523 31688 3581 31689
rect 12931 31688 12989 31689
rect 0 31648 3532 31688
rect 3572 31648 3581 31688
rect 5731 31648 5740 31688
rect 5780 31648 6124 31688
rect 6164 31648 6173 31688
rect 7651 31648 7660 31688
rect 7700 31648 11308 31688
rect 11348 31648 11357 31688
rect 11683 31648 11692 31688
rect 11732 31648 12460 31688
rect 12500 31648 12509 31688
rect 12846 31648 12940 31688
rect 12980 31648 12989 31688
rect 14275 31648 14284 31688
rect 14324 31648 14572 31688
rect 14612 31648 14621 31688
rect 15139 31648 15148 31688
rect 15188 31648 15916 31688
rect 15956 31648 15965 31688
rect 0 31628 80 31648
rect 3523 31647 3581 31648
rect 12931 31647 12989 31648
rect 2371 31604 2429 31605
rect 3043 31604 3101 31605
rect 3619 31604 3677 31605
rect 12067 31604 12125 31605
rect 15139 31604 15197 31605
rect 2371 31564 2380 31604
rect 2420 31564 2572 31604
rect 2612 31564 2621 31604
rect 3043 31564 3052 31604
rect 3092 31564 3628 31604
rect 3668 31564 12076 31604
rect 12116 31564 12125 31604
rect 12355 31564 12364 31604
rect 12404 31564 15148 31604
rect 15188 31564 15197 31604
rect 18019 31564 18028 31604
rect 18068 31564 18077 31604
rect 2371 31563 2429 31564
rect 3043 31563 3101 31564
rect 3619 31563 3677 31564
rect 12067 31563 12125 31564
rect 15139 31563 15197 31564
rect 9283 31520 9341 31521
rect 16867 31520 16925 31521
rect 1411 31480 1420 31520
rect 1460 31480 2188 31520
rect 2228 31480 2237 31520
rect 3619 31480 3628 31520
rect 3668 31480 4684 31520
rect 4724 31480 4733 31520
rect 5443 31480 5452 31520
rect 5492 31480 5836 31520
rect 5876 31480 5885 31520
rect 6403 31480 6412 31520
rect 6452 31480 6836 31520
rect 7459 31480 7468 31520
rect 7508 31480 7660 31520
rect 7700 31480 7709 31520
rect 9091 31480 9100 31520
rect 9140 31480 9292 31520
rect 9332 31480 9341 31520
rect 11587 31480 11596 31520
rect 11636 31480 13612 31520
rect 13652 31480 13661 31520
rect 13795 31480 13804 31520
rect 13844 31480 14188 31520
rect 14228 31480 14237 31520
rect 14371 31480 14380 31520
rect 14420 31480 14668 31520
rect 14708 31480 14717 31520
rect 14851 31480 14860 31520
rect 14900 31480 16876 31520
rect 16916 31480 16925 31520
rect 6796 31436 6836 31480
rect 9283 31479 9341 31480
rect 16867 31479 16925 31480
rect 18028 31436 18068 31564
rect 20899 31520 20957 31521
rect 21424 31520 21504 31540
rect 18403 31480 18412 31520
rect 18452 31480 19468 31520
rect 19508 31480 19517 31520
rect 20899 31480 20908 31520
rect 20948 31480 21504 31520
rect 20899 31479 20957 31480
rect 21424 31460 21504 31480
rect 1123 31396 1132 31436
rect 1172 31396 5644 31436
rect 5684 31396 5693 31436
rect 6787 31396 6796 31436
rect 6836 31396 6845 31436
rect 8131 31396 8140 31436
rect 8180 31396 10156 31436
rect 10196 31396 10205 31436
rect 11299 31396 11308 31436
rect 11348 31396 12980 31436
rect 13507 31396 13516 31436
rect 13556 31396 13565 31436
rect 13987 31396 13996 31436
rect 14036 31396 18068 31436
rect 18124 31396 20044 31436
rect 20084 31396 20093 31436
rect 0 31352 80 31372
rect 12940 31352 12980 31396
rect 0 31312 8372 31352
rect 11683 31312 11692 31352
rect 11732 31312 12172 31352
rect 12212 31312 12221 31352
rect 12931 31312 12940 31352
rect 12980 31312 13132 31352
rect 13172 31312 13181 31352
rect 13411 31312 13420 31352
rect 13460 31312 13469 31352
rect 0 31292 80 31312
rect 2851 31268 2909 31269
rect 4003 31268 4061 31269
rect 4579 31268 4637 31269
rect 1603 31228 1612 31268
rect 1652 31228 2860 31268
rect 2900 31228 2909 31268
rect 3139 31228 3148 31268
rect 3188 31228 3820 31268
rect 3860 31228 3869 31268
rect 4003 31228 4012 31268
rect 4052 31228 4204 31268
rect 4244 31228 4253 31268
rect 4579 31228 4588 31268
rect 4628 31228 7852 31268
rect 7892 31228 7901 31268
rect 2851 31227 2909 31228
rect 4003 31227 4061 31228
rect 4579 31227 4637 31228
rect 1315 31184 1373 31185
rect 2755 31184 2813 31185
rect 3331 31184 3389 31185
rect 8332 31184 8372 31312
rect 9955 31268 10013 31269
rect 13219 31268 13277 31269
rect 9187 31228 9196 31268
rect 9236 31228 9676 31268
rect 9716 31228 9725 31268
rect 9870 31228 9964 31268
rect 10004 31228 10013 31268
rect 10435 31228 10444 31268
rect 10484 31228 13228 31268
rect 13268 31228 13277 31268
rect 9955 31227 10013 31228
rect 13219 31227 13277 31228
rect 13420 31184 13460 31312
rect 13516 31268 13556 31396
rect 17251 31352 17309 31353
rect 18124 31352 18164 31396
rect 14179 31312 14188 31352
rect 14228 31312 16684 31352
rect 16724 31312 16733 31352
rect 17251 31312 17260 31352
rect 17300 31312 18164 31352
rect 19267 31312 19276 31352
rect 19316 31312 19564 31352
rect 19604 31312 19613 31352
rect 17251 31311 17309 31312
rect 18211 31268 18269 31269
rect 13516 31228 17644 31268
rect 17684 31228 17693 31268
rect 18019 31228 18028 31268
rect 18068 31228 18220 31268
rect 18260 31228 18269 31268
rect 18211 31227 18269 31228
rect 16387 31184 16445 31185
rect 18115 31184 18173 31185
rect 1230 31144 1324 31184
rect 1364 31144 1373 31184
rect 2563 31144 2572 31184
rect 2612 31144 2764 31184
rect 2804 31144 3340 31184
rect 3380 31144 3389 31184
rect 4003 31144 4012 31184
rect 4052 31144 6316 31184
rect 6356 31144 6365 31184
rect 8332 31144 11116 31184
rect 11156 31144 12364 31184
rect 12404 31144 12413 31184
rect 12931 31144 12940 31184
rect 12980 31144 13460 31184
rect 14083 31144 14092 31184
rect 14132 31144 14956 31184
rect 14996 31144 15724 31184
rect 15764 31144 15773 31184
rect 16302 31144 16396 31184
rect 16436 31144 16445 31184
rect 18030 31144 18124 31184
rect 18164 31144 18173 31184
rect 19075 31144 19084 31184
rect 19124 31144 19468 31184
rect 19508 31144 19517 31184
rect 1315 31143 1373 31144
rect 2755 31143 2813 31144
rect 3331 31143 3389 31144
rect 16387 31143 16445 31144
rect 18115 31143 18173 31144
rect 1987 31100 2045 31101
rect 6979 31100 7037 31101
rect 11779 31100 11837 31101
rect 1987 31060 1996 31100
rect 2036 31060 2188 31100
rect 2228 31060 2237 31100
rect 2500 31060 6604 31100
rect 6644 31060 6653 31100
rect 6979 31060 6988 31100
rect 7028 31060 8428 31100
rect 8468 31060 8477 31100
rect 11320 31060 11692 31100
rect 11732 31060 11788 31100
rect 11828 31060 11856 31100
rect 13699 31060 13708 31100
rect 13748 31060 17356 31100
rect 17396 31060 17405 31100
rect 18883 31060 18892 31100
rect 18932 31060 20620 31100
rect 20660 31060 20669 31100
rect 1987 31059 2045 31060
rect 0 31016 80 31036
rect 2500 31016 2540 31060
rect 6979 31059 7037 31060
rect 11320 31016 11360 31060
rect 11779 31059 11837 31060
rect 0 30976 844 31016
rect 884 30976 893 31016
rect 1228 30976 2540 31016
rect 4919 30976 4928 31016
rect 4968 30976 5010 31016
rect 5050 30976 5092 31016
rect 5132 30976 5174 31016
rect 5214 30976 5256 31016
rect 5296 30976 5305 31016
rect 5443 30976 5452 31016
rect 5492 30976 7468 31016
rect 7508 30976 7517 31016
rect 8332 30976 11360 31016
rect 12067 31016 12125 31017
rect 21283 31016 21341 31017
rect 21424 31016 21504 31036
rect 12067 30976 12076 31016
rect 12116 30976 12980 31016
rect 13027 30976 13036 31016
rect 13076 30976 13228 31016
rect 13268 30976 13277 31016
rect 14179 30976 14188 31016
rect 14228 30976 17164 31016
rect 17204 30976 17213 31016
rect 20039 30976 20048 31016
rect 20088 30976 20130 31016
rect 20170 30976 20212 31016
rect 20252 30976 20294 31016
rect 20334 30976 20376 31016
rect 20416 30976 20425 31016
rect 21283 30976 21292 31016
rect 21332 30976 21504 31016
rect 0 30956 80 30976
rect 0 30680 80 30700
rect 1228 30680 1268 30976
rect 2659 30932 2717 30933
rect 4003 30932 4061 30933
rect 4387 30932 4445 30933
rect 8332 30932 8372 30976
rect 12067 30975 12125 30976
rect 12940 30932 12980 30976
rect 21283 30975 21341 30976
rect 21424 30956 21504 30976
rect 19747 30932 19805 30933
rect 1315 30892 1324 30932
rect 1364 30892 2668 30932
rect 2708 30892 4012 30932
rect 4052 30892 4061 30932
rect 4195 30892 4204 30932
rect 4244 30892 4396 30932
rect 4436 30892 8372 30932
rect 8419 30892 8428 30932
rect 8468 30892 12748 30932
rect 12788 30892 12797 30932
rect 12940 30892 14380 30932
rect 14420 30892 14429 30932
rect 14668 30892 19756 30932
rect 19796 30892 19805 30932
rect 2659 30891 2717 30892
rect 4003 30891 4061 30892
rect 4387 30891 4445 30892
rect 3043 30848 3101 30849
rect 7363 30848 7421 30849
rect 14668 30848 14708 30892
rect 19747 30891 19805 30892
rect 17443 30848 17501 30849
rect 18787 30848 18845 30849
rect 2083 30808 2092 30848
rect 2132 30808 2476 30848
rect 2516 30808 2525 30848
rect 2572 30808 3052 30848
rect 3092 30808 4300 30848
rect 4340 30808 4349 30848
rect 5059 30808 5068 30848
rect 5108 30808 5452 30848
rect 5492 30808 5501 30848
rect 7267 30808 7276 30848
rect 7316 30808 7372 30848
rect 7412 30808 9868 30848
rect 9908 30808 9917 30848
rect 11971 30808 11980 30848
rect 12020 30808 14668 30848
rect 14708 30808 14717 30848
rect 17443 30808 17452 30848
rect 17492 30808 18124 30848
rect 18164 30808 18173 30848
rect 18787 30808 18796 30848
rect 18836 30808 19180 30848
rect 19220 30808 19229 30848
rect 2572 30764 2612 30808
rect 3043 30807 3101 30808
rect 7363 30807 7421 30808
rect 17443 30807 17501 30808
rect 18787 30807 18845 30808
rect 11107 30764 11165 30765
rect 14275 30764 14333 30765
rect 1795 30724 1804 30764
rect 1844 30724 2612 30764
rect 2659 30724 2668 30764
rect 2708 30724 2860 30764
rect 2900 30724 3340 30764
rect 3380 30724 5932 30764
rect 5972 30724 5981 30764
rect 6028 30724 11116 30764
rect 11156 30724 11165 30764
rect 11875 30724 11884 30764
rect 11924 30724 12172 30764
rect 12212 30724 12221 30764
rect 13219 30724 13228 30764
rect 13268 30724 13612 30764
rect 13652 30724 13661 30764
rect 13891 30724 13900 30764
rect 13940 30724 14284 30764
rect 14324 30724 14333 30764
rect 17731 30724 17740 30764
rect 17780 30724 19508 30764
rect 2755 30680 2813 30681
rect 4003 30680 4061 30681
rect 6028 30680 6068 30724
rect 11107 30723 11165 30724
rect 14275 30723 14333 30724
rect 17251 30680 17309 30681
rect 18403 30680 18461 30681
rect 18691 30680 18749 30681
rect 0 30640 1652 30680
rect 0 30620 80 30640
rect 1612 30428 1652 30640
rect 2755 30640 2764 30680
rect 2804 30640 3724 30680
rect 3764 30640 3773 30680
rect 4003 30640 4012 30680
rect 4052 30640 6068 30680
rect 6307 30640 6316 30680
rect 6356 30640 7756 30680
rect 7796 30640 7805 30680
rect 9379 30640 9388 30680
rect 9428 30640 9676 30680
rect 9716 30640 9725 30680
rect 11320 30640 14860 30680
rect 14900 30640 14909 30680
rect 15427 30640 15436 30680
rect 15476 30640 16012 30680
rect 16052 30640 16061 30680
rect 17251 30640 17260 30680
rect 17300 30640 17836 30680
rect 17876 30640 17885 30680
rect 18403 30640 18412 30680
rect 18452 30640 18700 30680
rect 18740 30640 19372 30680
rect 19412 30640 19421 30680
rect 2755 30639 2813 30640
rect 4003 30639 4061 30640
rect 4099 30596 4157 30597
rect 11320 30596 11360 30640
rect 17251 30639 17309 30640
rect 18403 30639 18461 30640
rect 18691 30639 18749 30640
rect 2467 30556 2476 30596
rect 2516 30556 2572 30596
rect 2612 30556 4108 30596
rect 4148 30556 4157 30596
rect 8899 30556 8908 30596
rect 8948 30556 11360 30596
rect 11491 30596 11549 30597
rect 17443 30596 17501 30597
rect 11491 30556 11500 30596
rect 11540 30556 12268 30596
rect 12308 30556 12317 30596
rect 12739 30556 12748 30596
rect 12788 30556 16780 30596
rect 16820 30556 17452 30596
rect 17492 30556 17501 30596
rect 19468 30596 19508 30724
rect 20515 30680 20573 30681
rect 19555 30640 19564 30680
rect 19604 30640 19852 30680
rect 19892 30640 20524 30680
rect 20564 30640 20573 30680
rect 20515 30639 20573 30640
rect 19468 30556 20044 30596
rect 20084 30556 20093 30596
rect 4099 30555 4157 30556
rect 11491 30555 11549 30556
rect 17443 30555 17501 30556
rect 21424 30513 21504 30532
rect 17923 30512 17981 30513
rect 21379 30512 21504 30513
rect 2275 30472 2284 30512
rect 2324 30472 2668 30512
rect 2708 30472 2717 30512
rect 3331 30472 3340 30512
rect 3380 30472 3628 30512
rect 3668 30472 3677 30512
rect 3811 30472 3820 30512
rect 3860 30472 5452 30512
rect 5492 30472 6028 30512
rect 6068 30472 6077 30512
rect 7939 30472 7948 30512
rect 7988 30472 10444 30512
rect 10484 30472 10493 30512
rect 11395 30472 11404 30512
rect 11444 30472 11596 30512
rect 11636 30472 11645 30512
rect 13699 30472 13708 30512
rect 13748 30472 13996 30512
rect 14036 30472 14045 30512
rect 17923 30472 17932 30512
rect 17972 30472 18124 30512
rect 18164 30472 18173 30512
rect 21379 30472 21388 30512
rect 21428 30472 21504 30512
rect 17923 30471 17981 30472
rect 21379 30471 21504 30472
rect 21424 30452 21504 30471
rect 15139 30428 15197 30429
rect 1315 30388 1324 30428
rect 1364 30388 1516 30428
rect 1556 30388 1565 30428
rect 1612 30388 2572 30428
rect 2612 30388 2621 30428
rect 4003 30388 4012 30428
rect 4052 30388 4396 30428
rect 4436 30388 4445 30428
rect 10147 30388 10156 30428
rect 10196 30388 14668 30428
rect 14708 30388 14717 30428
rect 15054 30388 15148 30428
rect 15188 30388 15197 30428
rect 15139 30387 15197 30388
rect 0 30344 80 30364
rect 5347 30344 5405 30345
rect 7747 30344 7805 30345
rect 14083 30344 14141 30345
rect 0 30304 1132 30344
rect 1172 30304 1181 30344
rect 2572 30304 2804 30344
rect 3043 30304 3052 30344
rect 3092 30304 4204 30344
rect 4244 30304 4253 30344
rect 5347 30304 5356 30344
rect 5396 30304 7756 30344
rect 7796 30304 7805 30344
rect 9091 30304 9100 30344
rect 9140 30304 11308 30344
rect 11348 30304 11357 30344
rect 13987 30304 13996 30344
rect 14036 30304 14092 30344
rect 14132 30304 14141 30344
rect 15235 30304 15244 30344
rect 15284 30304 19316 30344
rect 0 30284 80 30304
rect 2572 30260 2612 30304
rect 1699 30220 1708 30260
rect 1748 30220 2380 30260
rect 2420 30220 2429 30260
rect 2500 30220 2612 30260
rect 2500 30176 2540 30220
rect 2764 30176 2804 30304
rect 5347 30303 5405 30304
rect 7747 30303 7805 30304
rect 14083 30303 14141 30304
rect 2851 30220 2860 30260
rect 2900 30220 3532 30260
rect 3572 30220 3581 30260
rect 3679 30220 3688 30260
rect 3728 30220 3770 30260
rect 3810 30220 3852 30260
rect 3892 30220 3934 30260
rect 3974 30220 4016 30260
rect 4056 30220 4065 30260
rect 4771 30220 4780 30260
rect 4820 30220 5356 30260
rect 5396 30220 5644 30260
rect 5684 30220 9716 30260
rect 10243 30220 10252 30260
rect 10292 30220 14572 30260
rect 14612 30220 14621 30260
rect 16387 30220 16396 30260
rect 16436 30220 17740 30260
rect 17780 30220 17789 30260
rect 18799 30220 18808 30260
rect 18848 30220 18890 30260
rect 18930 30220 18972 30260
rect 19012 30220 19054 30260
rect 19094 30220 19136 30260
rect 19176 30220 19185 30260
rect 7075 30176 7133 30177
rect 9571 30176 9629 30177
rect 1795 30136 1804 30176
rect 1844 30136 2540 30176
rect 2659 30136 2668 30176
rect 2708 30136 2717 30176
rect 2764 30136 4492 30176
rect 4532 30136 4541 30176
rect 7075 30136 7084 30176
rect 7124 30136 7948 30176
rect 7988 30136 7997 30176
rect 9475 30136 9484 30176
rect 9524 30136 9580 30176
rect 9620 30136 9629 30176
rect 9676 30176 9716 30220
rect 14851 30176 14909 30177
rect 9676 30136 11020 30176
rect 11060 30136 11069 30176
rect 14659 30136 14668 30176
rect 14708 30136 14860 30176
rect 14900 30136 14909 30176
rect 19276 30176 19316 30304
rect 21379 30176 21437 30177
rect 19276 30136 21388 30176
rect 21428 30136 21437 30176
rect 2668 30092 2708 30136
rect 7075 30135 7133 30136
rect 9571 30135 9629 30136
rect 14851 30135 14909 30136
rect 21379 30135 21437 30136
rect 3139 30092 3197 30093
rect 14083 30092 14141 30093
rect 1699 30052 1708 30092
rect 1748 30052 2708 30092
rect 2755 30052 2764 30092
rect 2804 30052 3148 30092
rect 3188 30052 3197 30092
rect 6691 30052 6700 30092
rect 6740 30052 6988 30092
rect 7028 30052 7037 30092
rect 9091 30052 9100 30092
rect 9140 30052 9964 30092
rect 10004 30052 10013 30092
rect 11320 30052 12076 30092
rect 12116 30052 12125 30092
rect 13315 30052 13324 30092
rect 13364 30052 13612 30092
rect 13652 30052 13661 30092
rect 14083 30052 14092 30092
rect 14132 30052 15916 30092
rect 15956 30052 15965 30092
rect 17251 30052 17260 30092
rect 17300 30052 17836 30092
rect 17876 30052 17885 30092
rect 3139 30051 3197 30052
rect 0 30008 80 30028
rect 11320 30008 11360 30052
rect 14083 30051 14141 30052
rect 20707 30008 20765 30009
rect 21424 30008 21504 30028
rect 0 29968 2092 30008
rect 2132 29968 11360 30008
rect 11683 29968 11692 30008
rect 11732 29968 15820 30008
rect 15860 29968 15869 30008
rect 20227 29968 20236 30008
rect 20276 29968 20716 30008
rect 20756 29968 20765 30008
rect 0 29948 80 29968
rect 20707 29967 20765 29968
rect 20812 29968 21504 30008
rect 4195 29924 4253 29925
rect 8995 29924 9053 29925
rect 14467 29924 14525 29925
rect 20812 29924 20852 29968
rect 21424 29948 21504 29968
rect 739 29884 748 29924
rect 788 29884 1228 29924
rect 1268 29884 1277 29924
rect 4195 29884 4204 29924
rect 4244 29884 4300 29924
rect 4340 29884 4349 29924
rect 5731 29884 5740 29924
rect 5780 29884 9004 29924
rect 9044 29884 9524 29924
rect 12163 29884 12172 29924
rect 12212 29884 12460 29924
rect 12500 29884 13228 29924
rect 13268 29884 13277 29924
rect 13603 29884 13612 29924
rect 13652 29884 14188 29924
rect 14228 29884 14237 29924
rect 14467 29884 14476 29924
rect 14516 29884 14860 29924
rect 14900 29884 15436 29924
rect 15476 29884 15485 29924
rect 15907 29884 15916 29924
rect 15956 29884 17068 29924
rect 17108 29884 17117 29924
rect 20140 29884 20852 29924
rect 4195 29883 4253 29884
rect 8995 29883 9053 29884
rect 2755 29840 2813 29841
rect 6595 29840 6653 29841
rect 7267 29840 7325 29841
rect 9484 29840 9524 29884
rect 14467 29883 14525 29884
rect 10627 29840 10685 29841
rect 2755 29800 2764 29840
rect 2804 29800 5836 29840
rect 5876 29800 5885 29840
rect 6595 29800 6604 29840
rect 6644 29800 6988 29840
rect 7028 29800 7276 29840
rect 7316 29800 7325 29840
rect 7651 29800 7660 29840
rect 7700 29800 8332 29840
rect 8372 29800 8381 29840
rect 8515 29800 8524 29840
rect 8564 29800 8812 29840
rect 8852 29800 8861 29840
rect 9475 29800 9484 29840
rect 9524 29800 9533 29840
rect 10435 29800 10444 29840
rect 10484 29800 10493 29840
rect 10627 29800 10636 29840
rect 10676 29800 10770 29840
rect 13411 29800 13420 29840
rect 13460 29800 13900 29840
rect 13940 29800 13949 29840
rect 14371 29800 14380 29840
rect 14420 29800 15820 29840
rect 15860 29800 15869 29840
rect 17443 29800 17452 29840
rect 17492 29800 17501 29840
rect 2755 29799 2813 29800
rect 6595 29799 6653 29800
rect 7267 29799 7325 29800
rect 10444 29756 10484 29800
rect 10627 29799 10685 29800
rect 13315 29756 13373 29757
rect 16291 29756 16349 29757
rect 17452 29756 17492 29800
rect 20140 29756 20180 29884
rect 1132 29716 2284 29756
rect 2324 29716 2333 29756
rect 3235 29716 3244 29756
rect 3284 29716 5068 29756
rect 5108 29716 5117 29756
rect 5443 29716 5452 29756
rect 5492 29716 7084 29756
rect 7124 29716 10484 29756
rect 13230 29716 13324 29756
rect 13364 29716 13373 29756
rect 13795 29716 13804 29756
rect 13844 29716 16300 29756
rect 16340 29716 17492 29756
rect 17539 29716 17548 29756
rect 17588 29716 20180 29756
rect 0 29673 80 29692
rect 0 29672 125 29673
rect 1132 29672 1172 29716
rect 13315 29715 13373 29716
rect 16291 29715 16349 29716
rect 7075 29672 7133 29673
rect 10051 29672 10109 29673
rect 11107 29672 11165 29673
rect 0 29632 76 29672
rect 116 29632 1172 29672
rect 1219 29632 1228 29672
rect 1268 29632 7084 29672
rect 7124 29632 7133 29672
rect 7843 29632 7852 29672
rect 7892 29632 8716 29672
rect 8756 29632 8765 29672
rect 8995 29632 9004 29672
rect 9044 29632 9196 29672
rect 9236 29632 9245 29672
rect 9966 29632 10060 29672
rect 10100 29632 10109 29672
rect 10435 29632 10444 29672
rect 10484 29632 11020 29672
rect 11060 29632 11116 29672
rect 11156 29632 11165 29672
rect 12067 29632 12076 29672
rect 12116 29632 18028 29672
rect 18068 29632 18077 29672
rect 0 29631 125 29632
rect 7075 29631 7133 29632
rect 10051 29631 10109 29632
rect 11107 29631 11165 29632
rect 0 29612 80 29631
rect 451 29548 460 29588
rect 500 29548 14284 29588
rect 14324 29548 14333 29588
rect 14380 29548 17836 29588
rect 17876 29548 17885 29588
rect 3043 29504 3101 29505
rect 6499 29504 6557 29505
rect 8419 29504 8477 29505
rect 13315 29504 13373 29505
rect 14380 29504 14420 29548
rect 3043 29464 3052 29504
rect 3092 29464 3148 29504
rect 3188 29464 3197 29504
rect 4919 29464 4928 29504
rect 4968 29464 5010 29504
rect 5050 29464 5092 29504
rect 5132 29464 5174 29504
rect 5214 29464 5256 29504
rect 5296 29464 5305 29504
rect 6499 29464 6508 29504
rect 6548 29464 6892 29504
rect 6932 29464 8428 29504
rect 8468 29464 8477 29504
rect 12835 29464 12844 29504
rect 12884 29464 13324 29504
rect 13364 29464 13612 29504
rect 13652 29464 14420 29504
rect 15427 29504 15485 29505
rect 20611 29504 20669 29505
rect 21424 29504 21504 29524
rect 15427 29464 15436 29504
rect 15476 29464 17108 29504
rect 20039 29464 20048 29504
rect 20088 29464 20130 29504
rect 20170 29464 20212 29504
rect 20252 29464 20294 29504
rect 20334 29464 20376 29504
rect 20416 29464 20425 29504
rect 20611 29464 20620 29504
rect 20660 29464 21504 29504
rect 3043 29463 3101 29464
rect 6499 29463 6557 29464
rect 8419 29463 8477 29464
rect 13315 29463 13373 29464
rect 15427 29463 15485 29464
rect 16867 29420 16925 29421
rect 2947 29380 2956 29420
rect 2996 29380 5356 29420
rect 5396 29380 5836 29420
rect 5876 29380 5885 29420
rect 13315 29380 13324 29420
rect 13364 29380 13804 29420
rect 13844 29380 13853 29420
rect 16867 29380 16876 29420
rect 16916 29380 16972 29420
rect 17012 29380 17021 29420
rect 16867 29379 16925 29380
rect 0 29336 80 29356
rect 931 29336 989 29337
rect 5731 29336 5789 29337
rect 6019 29336 6077 29337
rect 17068 29336 17108 29464
rect 20611 29463 20669 29464
rect 21424 29444 21504 29464
rect 0 29296 940 29336
rect 980 29296 989 29336
rect 0 29276 80 29296
rect 931 29295 989 29296
rect 2500 29296 3244 29336
rect 3284 29296 3293 29336
rect 5059 29296 5068 29336
rect 5108 29296 5740 29336
rect 5780 29296 6028 29336
rect 6068 29296 6077 29336
rect 6691 29296 6700 29336
rect 6740 29296 8428 29336
rect 8468 29296 8716 29336
rect 8756 29296 10348 29336
rect 10388 29296 10397 29336
rect 14947 29296 14956 29336
rect 14996 29296 16780 29336
rect 16820 29296 16829 29336
rect 17059 29296 17068 29336
rect 17108 29296 17117 29336
rect 1987 29168 2045 29169
rect 2500 29168 2540 29296
rect 5731 29295 5789 29296
rect 6019 29295 6077 29296
rect 14275 29252 14333 29253
rect 2851 29212 2860 29252
rect 2900 29212 5684 29252
rect 9187 29212 9196 29252
rect 9236 29212 9964 29252
rect 10004 29212 10540 29252
rect 10580 29212 10589 29252
rect 11299 29212 11308 29252
rect 11348 29212 12460 29252
rect 12500 29212 12509 29252
rect 14190 29212 14284 29252
rect 14324 29212 14333 29252
rect 15331 29212 15340 29252
rect 15380 29212 16492 29252
rect 16532 29212 16541 29252
rect 16675 29212 16684 29252
rect 16724 29212 17164 29252
rect 17204 29212 17213 29252
rect 5644 29168 5684 29212
rect 14275 29211 14333 29212
rect 11203 29168 11261 29169
rect 12835 29168 12893 29169
rect 1603 29128 1612 29168
rect 1652 29128 1996 29168
rect 2036 29128 2045 29168
rect 2467 29128 2476 29168
rect 2516 29128 2540 29168
rect 5635 29128 5644 29168
rect 5684 29128 5693 29168
rect 8227 29128 8236 29168
rect 8276 29128 8524 29168
rect 8564 29128 8573 29168
rect 8899 29128 8908 29168
rect 8948 29128 10636 29168
rect 10676 29128 10685 29168
rect 11118 29128 11212 29168
rect 11252 29128 11261 29168
rect 12750 29128 12844 29168
rect 12884 29128 12893 29168
rect 1987 29127 2045 29128
rect 451 29084 509 29085
rect 451 29044 460 29084
rect 500 29044 884 29084
rect 931 29044 940 29084
rect 980 29044 1172 29084
rect 1507 29044 1516 29084
rect 1556 29044 4108 29084
rect 4148 29044 4157 29084
rect 451 29043 509 29044
rect 0 29000 80 29020
rect 844 29001 884 29044
rect 835 29000 893 29001
rect 1132 29000 1172 29044
rect 8332 29000 8372 29128
rect 11203 29127 11261 29128
rect 12835 29127 12893 29128
rect 13123 29168 13181 29169
rect 15811 29168 15869 29169
rect 16579 29168 16637 29169
rect 13123 29128 13132 29168
rect 13172 29128 13324 29168
rect 13364 29128 13373 29168
rect 13987 29128 13996 29168
rect 14036 29128 14860 29168
rect 14900 29128 14909 29168
rect 15043 29128 15052 29168
rect 15092 29128 15532 29168
rect 15572 29128 15581 29168
rect 15726 29128 15820 29168
rect 15860 29128 15869 29168
rect 16387 29128 16396 29168
rect 16436 29128 16445 29168
rect 16579 29128 16588 29168
rect 16628 29128 17452 29168
rect 17492 29128 18316 29168
rect 18356 29128 18604 29168
rect 18644 29128 19084 29168
rect 19124 29128 19133 29168
rect 13123 29127 13181 29128
rect 15811 29127 15869 29128
rect 16396 29084 16436 29128
rect 16579 29127 16637 29128
rect 19939 29084 19997 29085
rect 9379 29044 9388 29084
rect 9428 29044 9580 29084
rect 9620 29044 10196 29084
rect 9955 29000 10013 29001
rect 10156 29000 10196 29044
rect 10252 29044 11348 29084
rect 14179 29044 14188 29084
rect 14228 29044 15380 29084
rect 15427 29044 15436 29084
rect 15476 29044 16436 29084
rect 16588 29044 19604 29084
rect 0 28960 172 29000
rect 212 28960 221 29000
rect 804 28960 844 29000
rect 884 28960 893 29000
rect 1092 28960 1132 29000
rect 1172 28960 1181 29000
rect 1987 28960 1996 29000
rect 2036 28960 2668 29000
rect 2708 28960 2717 29000
rect 3043 28960 3052 29000
rect 3092 28960 3820 29000
rect 3860 28960 4684 29000
rect 4724 28960 4733 29000
rect 8332 28960 9772 29000
rect 9812 28960 9964 29000
rect 10004 28960 10013 29000
rect 10116 28960 10156 29000
rect 10196 28960 10205 29000
rect 0 28940 80 28960
rect 835 28959 893 28960
rect 9955 28959 10013 28960
rect 1795 28916 1853 28917
rect 10252 28916 10292 29044
rect 10819 29000 10877 29001
rect 10734 28960 10828 29000
rect 10868 28960 10877 29000
rect 11308 29000 11348 29044
rect 15340 29000 15380 29044
rect 15427 29000 15485 29001
rect 16588 29000 16628 29044
rect 11308 28960 11404 29000
rect 11444 28960 11453 29000
rect 15340 28960 15436 29000
rect 15476 28960 15628 29000
rect 15668 28960 15677 29000
rect 16548 28960 16588 29000
rect 16628 28960 16637 29000
rect 18883 28960 18892 29000
rect 18932 28960 18941 29000
rect 10819 28959 10877 28960
rect 15427 28959 15485 28960
rect 18892 28916 18932 28960
rect 19564 28916 19604 29044
rect 19939 29044 19948 29084
rect 19988 29044 21236 29084
rect 19939 29043 19997 29044
rect 19843 29000 19901 29001
rect 19758 28960 19852 29000
rect 19892 28960 19901 29000
rect 21196 29000 21236 29044
rect 21424 29000 21504 29020
rect 21196 28960 21504 29000
rect 19843 28959 19901 28960
rect 21424 28940 21504 28960
rect 1699 28876 1708 28916
rect 1748 28876 1804 28916
rect 1844 28876 1853 28916
rect 7555 28876 7564 28916
rect 7604 28876 10292 28916
rect 12643 28876 12652 28916
rect 12692 28876 13228 28916
rect 13268 28876 13277 28916
rect 18892 28876 19372 28916
rect 19412 28876 19421 28916
rect 19564 28876 21292 28916
rect 21332 28876 21341 28916
rect 1795 28875 1853 28876
rect 6979 28832 7037 28833
rect 67 28792 76 28832
rect 116 28792 2092 28832
rect 2132 28792 4492 28832
rect 4532 28792 6988 28832
rect 7028 28792 7037 28832
rect 6979 28791 7037 28792
rect 10627 28832 10685 28833
rect 10627 28792 10636 28832
rect 10676 28792 10828 28832
rect 10868 28792 10877 28832
rect 10627 28791 10685 28792
rect 3427 28748 3485 28749
rect 3342 28708 3436 28748
rect 3476 28708 3485 28748
rect 3679 28708 3688 28748
rect 3728 28708 3770 28748
rect 3810 28708 3852 28748
rect 3892 28708 3934 28748
rect 3974 28708 4016 28748
rect 4056 28708 4065 28748
rect 8803 28708 8812 28748
rect 8852 28708 9484 28748
rect 9524 28708 9533 28748
rect 9667 28708 9676 28748
rect 9716 28708 10732 28748
rect 10772 28708 10781 28748
rect 18799 28708 18808 28748
rect 18848 28708 18890 28748
rect 18930 28708 18972 28748
rect 19012 28708 19054 28748
rect 19094 28708 19136 28748
rect 19176 28708 19185 28748
rect 3427 28707 3485 28708
rect 0 28664 80 28684
rect 7939 28664 7997 28665
rect 0 28624 7948 28664
rect 7988 28624 7997 28664
rect 0 28604 80 28624
rect 7939 28623 7997 28624
rect 8419 28664 8477 28665
rect 9484 28664 9524 28708
rect 8419 28624 8428 28664
rect 8468 28624 8716 28664
rect 8756 28624 8765 28664
rect 9484 28624 9868 28664
rect 9908 28624 9917 28664
rect 11320 28624 18700 28664
rect 18740 28624 18749 28664
rect 8419 28623 8477 28624
rect 3907 28540 3916 28580
rect 3956 28540 4204 28580
rect 4244 28540 4253 28580
rect 6307 28540 6316 28580
rect 6356 28540 10540 28580
rect 10580 28540 10589 28580
rect 1891 28456 1900 28496
rect 1940 28456 2380 28496
rect 2420 28456 2429 28496
rect 6595 28456 6604 28496
rect 6644 28456 10924 28496
rect 10964 28456 10973 28496
rect 9667 28412 9725 28413
rect 11320 28412 11360 28624
rect 15427 28580 15485 28581
rect 12835 28540 12844 28580
rect 12884 28540 13132 28580
rect 13172 28540 13521 28580
rect 13561 28540 13570 28580
rect 15427 28540 15436 28580
rect 15476 28540 15820 28580
rect 15860 28540 15869 28580
rect 15427 28539 15485 28540
rect 21424 28496 21504 28516
rect 12643 28456 12652 28496
rect 12692 28456 12884 28496
rect 15235 28456 15244 28496
rect 15284 28456 16204 28496
rect 16244 28456 16253 28496
rect 20515 28456 20524 28496
rect 20564 28456 21504 28496
rect 3139 28372 3148 28412
rect 3188 28372 4012 28412
rect 4052 28372 4061 28412
rect 4195 28372 4204 28412
rect 4244 28372 5260 28412
rect 5300 28372 5309 28412
rect 5923 28372 5932 28412
rect 5972 28372 6508 28412
rect 6548 28372 7276 28412
rect 7316 28372 7325 28412
rect 8419 28372 8428 28412
rect 8468 28372 9388 28412
rect 9428 28372 9437 28412
rect 9667 28372 9676 28412
rect 9716 28372 11360 28412
rect 9667 28371 9725 28372
rect 0 28328 80 28348
rect 9475 28328 9533 28329
rect 12844 28328 12884 28456
rect 21424 28436 21504 28456
rect 13603 28412 13661 28413
rect 19555 28412 19613 28413
rect 13603 28372 13612 28412
rect 13652 28372 15532 28412
rect 15572 28372 15581 28412
rect 19555 28372 19564 28412
rect 19604 28372 19852 28412
rect 19892 28372 19901 28412
rect 13603 28371 13661 28372
rect 19555 28371 19613 28372
rect 0 28288 1708 28328
rect 1748 28288 1757 28328
rect 4291 28288 4300 28328
rect 4340 28288 5452 28328
rect 5492 28288 5501 28328
rect 6019 28288 6028 28328
rect 6068 28288 6220 28328
rect 6260 28288 6269 28328
rect 6787 28288 6796 28328
rect 6836 28288 8620 28328
rect 8660 28288 8669 28328
rect 8899 28288 8908 28328
rect 8948 28288 9100 28328
rect 9140 28288 9149 28328
rect 9475 28288 9484 28328
rect 9524 28288 9618 28328
rect 9859 28288 9868 28328
rect 9908 28288 10444 28328
rect 10484 28288 10493 28328
rect 12835 28288 12844 28328
rect 12884 28288 12893 28328
rect 13315 28288 13324 28328
rect 13364 28288 13708 28328
rect 13748 28288 13757 28328
rect 15715 28288 15724 28328
rect 15764 28288 16396 28328
rect 16436 28288 16445 28328
rect 17251 28288 17260 28328
rect 17300 28288 18508 28328
rect 18548 28288 18557 28328
rect 0 28268 80 28288
rect 9475 28287 9533 28288
rect 6691 28244 6749 28245
rect 13987 28244 14045 28245
rect 1027 28204 1036 28244
rect 1076 28204 3724 28244
rect 3764 28204 3773 28244
rect 6691 28204 6700 28244
rect 6740 28204 6892 28244
rect 6932 28204 6941 28244
rect 8515 28204 8524 28244
rect 8564 28204 8660 28244
rect 11395 28204 11404 28244
rect 11444 28204 13996 28244
rect 14036 28204 14045 28244
rect 6691 28203 6749 28204
rect 1219 28160 1277 28161
rect 8620 28160 8660 28204
rect 13987 28203 14045 28204
rect 1200 28120 1228 28160
rect 1268 28120 1324 28160
rect 1364 28120 1612 28160
rect 1652 28120 1661 28160
rect 3043 28120 3052 28160
rect 3092 28120 4492 28160
rect 4532 28120 5644 28160
rect 5684 28120 5693 28160
rect 8620 28120 10060 28160
rect 10100 28120 10109 28160
rect 13027 28120 13036 28160
rect 13076 28120 13612 28160
rect 13652 28120 13661 28160
rect 13795 28120 13804 28160
rect 13844 28120 14668 28160
rect 14708 28120 14717 28160
rect 16195 28120 16204 28160
rect 16244 28120 16684 28160
rect 16724 28120 16733 28160
rect 1219 28119 1277 28120
rect 14947 28076 15005 28077
rect 2500 28036 6356 28076
rect 6403 28036 6412 28076
rect 6452 28036 14956 28076
rect 14996 28036 15005 28076
rect 19363 28036 19372 28076
rect 19412 28036 20852 28076
rect 0 27992 80 28012
rect 2500 27992 2540 28036
rect 3235 27992 3293 27993
rect 5635 27992 5693 27993
rect 0 27952 2540 27992
rect 3150 27952 3244 27992
rect 3284 27952 3293 27992
rect 4919 27952 4928 27992
rect 4968 27952 5010 27992
rect 5050 27952 5092 27992
rect 5132 27952 5174 27992
rect 5214 27952 5256 27992
rect 5296 27952 5305 27992
rect 5347 27952 5356 27992
rect 5396 27952 5644 27992
rect 5684 27952 5693 27992
rect 6316 27992 6356 28036
rect 14947 28035 15005 28036
rect 9475 27992 9533 27993
rect 20812 27992 20852 28036
rect 21424 27992 21504 28012
rect 6316 27952 8140 27992
rect 8180 27952 8428 27992
rect 8468 27952 8477 27992
rect 8800 27952 9484 27992
rect 9524 27952 9533 27992
rect 17827 27952 17836 27992
rect 17876 27952 18604 27992
rect 18644 27952 19468 27992
rect 19508 27952 19517 27992
rect 20039 27952 20048 27992
rect 20088 27952 20130 27992
rect 20170 27952 20212 27992
rect 20252 27952 20294 27992
rect 20334 27952 20376 27992
rect 20416 27952 20425 27992
rect 20812 27952 21504 27992
rect 0 27932 80 27952
rect 3235 27951 3293 27952
rect 5635 27951 5693 27952
rect 2659 27908 2717 27909
rect 8800 27908 8840 27952
rect 9475 27951 9533 27952
rect 21424 27932 21504 27952
rect 17251 27908 17309 27909
rect 2659 27868 2668 27908
rect 2708 27868 2764 27908
rect 2804 27868 2813 27908
rect 5356 27868 5548 27908
rect 5588 27868 5597 27908
rect 5827 27868 5836 27908
rect 5876 27868 8840 27908
rect 12163 27868 12172 27908
rect 12212 27868 17260 27908
rect 17300 27868 17309 27908
rect 17635 27868 17644 27908
rect 17684 27868 17932 27908
rect 17972 27868 19372 27908
rect 19412 27868 19421 27908
rect 2659 27867 2717 27868
rect 4483 27824 4541 27825
rect 4771 27824 4829 27825
rect 1795 27784 1804 27824
rect 1844 27784 2476 27824
rect 2516 27784 2525 27824
rect 2851 27784 2860 27824
rect 2900 27784 3244 27824
rect 3284 27784 3293 27824
rect 4291 27784 4300 27824
rect 4340 27784 4492 27824
rect 4532 27784 4780 27824
rect 4820 27784 4829 27824
rect 4483 27783 4541 27784
rect 4771 27783 4829 27784
rect 1891 27740 1949 27741
rect 5356 27740 5396 27868
rect 17251 27867 17309 27868
rect 5539 27824 5597 27825
rect 13891 27824 13949 27825
rect 5443 27784 5452 27824
rect 5492 27784 5548 27824
rect 5588 27784 5597 27824
rect 6115 27784 6124 27824
rect 6164 27784 6604 27824
rect 6644 27784 6653 27824
rect 7372 27784 8044 27824
rect 8084 27784 8093 27824
rect 8323 27784 8332 27824
rect 8372 27784 8812 27824
rect 8852 27784 11116 27824
rect 11156 27784 11165 27824
rect 12643 27784 12652 27824
rect 12692 27784 13708 27824
rect 13748 27784 13757 27824
rect 13891 27784 13900 27824
rect 13940 27784 15340 27824
rect 15380 27784 15389 27824
rect 16291 27784 16300 27824
rect 16340 27784 17396 27824
rect 5539 27783 5597 27784
rect 7372 27740 7412 27784
rect 13891 27783 13949 27784
rect 9763 27740 9821 27741
rect 13603 27740 13661 27741
rect 15331 27740 15389 27741
rect 1315 27700 1324 27740
rect 1364 27700 1900 27740
rect 1940 27700 1949 27740
rect 2563 27700 2572 27740
rect 2612 27700 3148 27740
rect 3188 27700 5396 27740
rect 5731 27700 5740 27740
rect 5780 27700 7372 27740
rect 7412 27700 7421 27740
rect 7555 27700 7564 27740
rect 7604 27700 8908 27740
rect 8948 27700 9388 27740
rect 9428 27700 9437 27740
rect 9763 27700 9772 27740
rect 9812 27700 10060 27740
rect 10100 27700 10109 27740
rect 11395 27700 11404 27740
rect 11444 27700 13172 27740
rect 13518 27700 13612 27740
rect 13652 27700 13661 27740
rect 1891 27699 1949 27700
rect 0 27656 80 27676
rect 2467 27656 2525 27657
rect 0 27616 2476 27656
rect 2516 27616 2525 27656
rect 2755 27616 2764 27656
rect 2804 27616 3916 27656
rect 3956 27616 3965 27656
rect 4099 27616 4108 27656
rect 4148 27616 4780 27656
rect 4820 27616 4829 27656
rect 0 27596 80 27616
rect 2467 27615 2525 27616
rect 4108 27572 4148 27616
rect 3148 27532 3532 27572
rect 3572 27532 4148 27572
rect 7372 27572 7412 27700
rect 9763 27699 9821 27700
rect 12643 27656 12701 27657
rect 13132 27656 13172 27700
rect 13603 27699 13661 27700
rect 14188 27700 15340 27740
rect 15380 27700 15389 27740
rect 14083 27656 14141 27657
rect 7459 27616 7468 27656
rect 7508 27616 8044 27656
rect 8084 27616 8093 27656
rect 8515 27616 8524 27656
rect 8564 27616 11020 27656
rect 11060 27616 11069 27656
rect 11875 27616 11884 27656
rect 11924 27616 12652 27656
rect 12692 27616 12701 27656
rect 13123 27616 13132 27656
rect 13172 27616 14092 27656
rect 14132 27616 14141 27656
rect 12643 27615 12701 27616
rect 8995 27572 9053 27573
rect 7372 27532 8428 27572
rect 8468 27532 8477 27572
rect 8910 27532 9004 27572
rect 9044 27532 9053 27572
rect 3148 27488 3188 27532
rect 8995 27531 9053 27532
rect 9571 27572 9629 27573
rect 9571 27532 9580 27572
rect 9620 27532 9908 27572
rect 9571 27531 9629 27532
rect 7267 27488 7325 27489
rect 7747 27488 7805 27489
rect 9868 27488 9908 27532
rect 13516 27488 13556 27616
rect 14083 27615 14141 27616
rect 14188 27572 14228 27700
rect 15331 27699 15389 27700
rect 15619 27740 15677 27741
rect 15619 27700 15628 27740
rect 15668 27700 16876 27740
rect 16916 27700 16925 27740
rect 15619 27699 15677 27700
rect 15811 27616 15820 27656
rect 15860 27616 16300 27656
rect 16340 27616 16588 27656
rect 16628 27616 16637 27656
rect 16771 27616 16780 27656
rect 16820 27616 16829 27656
rect 16780 27572 16820 27616
rect 13795 27532 13804 27572
rect 13844 27532 14228 27572
rect 14851 27532 14860 27572
rect 14900 27532 15148 27572
rect 15188 27532 16820 27572
rect 17356 27572 17396 27784
rect 19267 27700 19276 27740
rect 19316 27700 20812 27740
rect 20852 27700 20861 27740
rect 17443 27656 17501 27657
rect 17443 27616 17452 27656
rect 17492 27616 18892 27656
rect 18932 27616 18941 27656
rect 17443 27615 17501 27616
rect 17356 27532 17684 27572
rect 17731 27532 17740 27572
rect 17780 27532 18604 27572
rect 18644 27532 19756 27572
rect 19796 27532 19805 27572
rect 19939 27532 19948 27572
rect 19988 27532 20180 27572
rect 14851 27488 14909 27489
rect 15715 27488 15773 27489
rect 16291 27488 16349 27489
rect 17644 27488 17684 27532
rect 20140 27488 20180 27532
rect 21424 27488 21504 27508
rect 2659 27448 2668 27488
rect 2708 27448 3148 27488
rect 3188 27448 3197 27488
rect 3811 27448 3820 27488
rect 3860 27448 7276 27488
rect 7316 27448 7325 27488
rect 7662 27448 7756 27488
rect 7796 27448 7805 27488
rect 8515 27448 8524 27488
rect 8564 27448 9484 27488
rect 9524 27448 9533 27488
rect 9859 27448 9868 27488
rect 9908 27448 9917 27488
rect 13507 27448 13516 27488
rect 13556 27448 13565 27488
rect 14563 27448 14572 27488
rect 14612 27448 14860 27488
rect 14900 27448 15052 27488
rect 15092 27448 15101 27488
rect 15715 27448 15724 27488
rect 15764 27448 16300 27488
rect 16340 27448 17356 27488
rect 17396 27448 17405 27488
rect 17644 27448 18412 27488
rect 18452 27448 18461 27488
rect 20140 27448 21504 27488
rect 7267 27447 7325 27448
rect 7747 27447 7805 27448
rect 14851 27447 14909 27448
rect 15715 27447 15773 27448
rect 16291 27447 16349 27448
rect 21424 27428 21504 27448
rect 9379 27404 9437 27405
rect 9667 27404 9725 27405
rect 1315 27364 1324 27404
rect 1364 27364 2764 27404
rect 2804 27364 2813 27404
rect 2856 27364 2865 27404
rect 2905 27364 3052 27404
rect 3092 27364 3101 27404
rect 6115 27364 6124 27404
rect 6164 27364 9388 27404
rect 9428 27364 9676 27404
rect 9716 27364 9725 27404
rect 12835 27364 12844 27404
rect 12884 27364 13420 27404
rect 13460 27364 20127 27404
rect 20167 27364 20176 27404
rect 20227 27364 20236 27404
rect 20276 27364 20716 27404
rect 20756 27364 20765 27404
rect 9379 27363 9437 27364
rect 9667 27363 9725 27364
rect 0 27320 80 27340
rect 19363 27320 19421 27321
rect 0 27280 18316 27320
rect 18356 27280 19372 27320
rect 19412 27280 19421 27320
rect 0 27260 80 27280
rect 19363 27279 19421 27280
rect 13411 27236 13469 27237
rect 16675 27236 16733 27237
rect 2851 27196 2860 27236
rect 2900 27196 3244 27236
rect 3284 27196 3293 27236
rect 3679 27196 3688 27236
rect 3728 27196 3770 27236
rect 3810 27196 3852 27236
rect 3892 27196 3934 27236
rect 3974 27196 4016 27236
rect 4056 27196 4065 27236
rect 5452 27196 8620 27236
rect 8660 27196 8669 27236
rect 12835 27196 12844 27236
rect 12884 27196 13420 27236
rect 13460 27196 13469 27236
rect 5452 27152 5492 27196
rect 13411 27195 13469 27196
rect 13996 27196 16300 27236
rect 16340 27196 16349 27236
rect 16675 27196 16684 27236
rect 16724 27196 18740 27236
rect 18799 27196 18808 27236
rect 18848 27196 18890 27236
rect 18930 27196 18972 27236
rect 19012 27196 19054 27236
rect 19094 27196 19136 27236
rect 19176 27196 19185 27236
rect 7939 27152 7997 27153
rect 172 27112 5492 27152
rect 5731 27112 5740 27152
rect 5780 27112 6220 27152
rect 6260 27112 6269 27152
rect 6403 27112 6412 27152
rect 6452 27112 7028 27152
rect 7075 27112 7084 27152
rect 7124 27112 7948 27152
rect 7988 27112 7997 27152
rect 0 26984 80 27004
rect 172 26984 212 27112
rect 3619 27068 3677 27069
rect 6307 27068 6365 27069
rect 6988 27068 7028 27112
rect 7939 27111 7997 27112
rect 3427 27028 3436 27068
rect 3476 27028 3628 27068
rect 3668 27028 3677 27068
rect 5635 27028 5644 27068
rect 5684 27028 6316 27068
rect 6356 27028 6644 27068
rect 6988 27028 7180 27068
rect 7220 27028 7229 27068
rect 8803 27028 8812 27068
rect 8852 27028 9100 27068
rect 9140 27028 9149 27068
rect 3619 27027 3677 27028
rect 6307 27027 6365 27028
rect 0 26944 212 26984
rect 3043 26984 3101 26985
rect 6604 26984 6644 27028
rect 13996 26984 14036 27196
rect 16675 27195 16733 27196
rect 18700 27152 18740 27196
rect 14371 27112 14380 27152
rect 14420 27112 14860 27152
rect 14900 27112 14909 27152
rect 15619 27112 15628 27152
rect 15668 27112 16012 27152
rect 16052 27112 17260 27152
rect 17300 27112 17309 27152
rect 18700 27112 19276 27152
rect 19316 27112 19325 27152
rect 14083 27068 14141 27069
rect 17731 27068 17789 27069
rect 18691 27068 18749 27069
rect 14083 27028 14092 27068
rect 14132 27028 14226 27068
rect 16195 27028 16204 27068
rect 16244 27028 17452 27068
rect 17492 27028 17501 27068
rect 17646 27028 17740 27068
rect 17780 27028 17789 27068
rect 18606 27028 18700 27068
rect 18740 27028 18749 27068
rect 14083 27027 14141 27028
rect 17731 27027 17789 27028
rect 18691 27027 18749 27028
rect 3043 26944 3052 26984
rect 3092 26944 3244 26984
rect 3284 26944 3293 26984
rect 4195 26944 4204 26984
rect 4244 26944 6508 26984
rect 6548 26944 6557 26984
rect 6604 26944 8840 26984
rect 11395 26944 11404 26984
rect 11444 26944 12076 26984
rect 12116 26944 12125 26984
rect 13987 26944 13996 26984
rect 14036 26944 14045 26984
rect 14371 26944 14380 26984
rect 14420 26944 17644 26984
rect 17684 26944 18796 26984
rect 18836 26944 18845 26984
rect 0 26924 80 26944
rect 3043 26943 3101 26944
rect 4291 26900 4349 26901
rect 6403 26900 6461 26901
rect 8800 26900 8840 26944
rect 16771 26900 16829 26901
rect 17347 26900 17405 26901
rect 18019 26900 18077 26901
rect 18892 26900 18932 27112
rect 19939 27028 19948 27068
rect 19988 27028 20180 27068
rect 20140 26984 20180 27028
rect 21424 26984 21504 27004
rect 20140 26944 21504 26984
rect 21424 26924 21504 26944
rect 19555 26900 19613 26901
rect 1795 26860 1804 26900
rect 1844 26860 4244 26900
rect 4204 26816 4244 26860
rect 4291 26860 4300 26900
rect 4340 26860 4396 26900
rect 4436 26860 4445 26900
rect 5932 26860 6412 26900
rect 6452 26860 7276 26900
rect 7316 26860 7325 26900
rect 8800 26860 13748 26900
rect 14275 26860 14284 26900
rect 14324 26860 16400 26900
rect 4291 26859 4349 26860
rect 5932 26816 5972 26860
rect 6403 26859 6461 26860
rect 6499 26816 6557 26817
rect 9283 26816 9341 26817
rect 9667 26816 9725 26817
rect 9955 26816 10013 26817
rect 1219 26776 1228 26816
rect 1268 26776 2188 26816
rect 2228 26776 2237 26816
rect 4204 26776 5972 26816
rect 6115 26776 6124 26816
rect 6164 26776 6508 26816
rect 6548 26776 6557 26816
rect 6787 26776 6796 26816
rect 6836 26776 7564 26816
rect 7604 26776 7613 26816
rect 8707 26776 8716 26816
rect 8756 26776 9292 26816
rect 9332 26776 9676 26816
rect 9716 26776 9725 26816
rect 9870 26776 9964 26816
rect 10004 26776 10013 26816
rect 11011 26776 11020 26816
rect 11060 26776 11212 26816
rect 11252 26776 11261 26816
rect 12739 26776 12748 26816
rect 12788 26776 13420 26816
rect 13460 26776 13469 26816
rect 6499 26775 6557 26776
rect 9283 26775 9341 26776
rect 9667 26775 9725 26776
rect 9955 26775 10013 26776
rect 2755 26732 2813 26733
rect 6307 26732 6365 26733
rect 11971 26732 12029 26733
rect 643 26692 652 26732
rect 692 26692 2764 26732
rect 2804 26692 3532 26732
rect 3572 26692 3581 26732
rect 4003 26692 4012 26732
rect 4052 26692 5932 26732
rect 5972 26692 5981 26732
rect 6307 26692 6316 26732
rect 6356 26692 6412 26732
rect 6452 26692 6461 26732
rect 6504 26692 6513 26732
rect 6553 26692 7180 26732
rect 7220 26692 7229 26732
rect 11683 26692 11692 26732
rect 11732 26692 11980 26732
rect 12020 26692 12029 26732
rect 2755 26691 2813 26692
rect 6307 26691 6365 26692
rect 11971 26691 12029 26692
rect 0 26648 80 26668
rect 4291 26648 4349 26649
rect 7171 26648 7229 26649
rect 9571 26648 9629 26649
rect 0 26608 2572 26648
rect 2612 26608 2621 26648
rect 4291 26608 4300 26648
rect 4340 26608 7180 26648
rect 7220 26608 7229 26648
rect 9486 26608 9580 26648
rect 9620 26608 9629 26648
rect 0 26588 80 26608
rect 4291 26607 4349 26608
rect 7171 26607 7229 26608
rect 9571 26607 9629 26608
rect 12931 26648 12989 26649
rect 13411 26648 13469 26649
rect 12931 26608 12940 26648
rect 12980 26608 13228 26648
rect 13268 26608 13277 26648
rect 13326 26608 13420 26648
rect 13460 26608 13469 26648
rect 13708 26648 13748 26860
rect 13795 26776 13804 26816
rect 13844 26776 14476 26816
rect 14516 26776 14525 26816
rect 16360 26732 16400 26860
rect 16771 26860 16780 26900
rect 16820 26860 16914 26900
rect 17347 26860 17356 26900
rect 17396 26860 17548 26900
rect 17588 26860 17597 26900
rect 17923 26860 17932 26900
rect 17972 26860 18028 26900
rect 18068 26860 18077 26900
rect 18691 26860 18700 26900
rect 18740 26860 19564 26900
rect 19604 26860 19613 26900
rect 16771 26859 16829 26860
rect 17347 26859 17405 26860
rect 18019 26859 18077 26860
rect 19555 26859 19613 26860
rect 17443 26816 17501 26817
rect 16963 26776 16972 26816
rect 17012 26776 17260 26816
rect 17300 26776 17309 26816
rect 17443 26776 17452 26816
rect 17492 26776 19564 26816
rect 19604 26776 19613 26816
rect 17443 26775 17501 26776
rect 19939 26732 19997 26733
rect 16360 26692 19372 26732
rect 19412 26692 19948 26732
rect 19988 26692 19997 26732
rect 19939 26691 19997 26692
rect 16675 26648 16733 26649
rect 17251 26648 17309 26649
rect 13708 26608 14284 26648
rect 14324 26608 14333 26648
rect 14956 26608 16684 26648
rect 16724 26608 16733 26648
rect 17059 26608 17068 26648
rect 17108 26608 17260 26648
rect 17300 26608 17309 26648
rect 18403 26608 18412 26648
rect 18452 26608 21388 26648
rect 21428 26608 21437 26648
rect 12931 26607 12989 26608
rect 13411 26607 13469 26608
rect 14956 26564 14996 26608
rect 16675 26607 16733 26608
rect 17251 26607 17309 26608
rect 4195 26524 4204 26564
rect 4244 26524 5396 26564
rect 5443 26524 5452 26564
rect 5492 26524 7372 26564
rect 7412 26524 7421 26564
rect 9859 26524 9868 26564
rect 9908 26524 14996 26564
rect 15043 26524 15052 26564
rect 15092 26524 17164 26564
rect 17204 26524 17836 26564
rect 17876 26524 17885 26564
rect 18211 26524 18220 26564
rect 18260 26524 19948 26564
rect 19988 26524 19997 26564
rect 1315 26480 1373 26481
rect 5356 26480 5396 26524
rect 5635 26480 5693 26481
rect 6499 26480 6557 26481
rect 7267 26480 7325 26481
rect 19651 26480 19709 26481
rect 21424 26480 21504 26500
rect 1315 26440 1324 26480
rect 1364 26440 1420 26480
rect 1460 26440 1469 26480
rect 3427 26440 3436 26480
rect 3476 26440 3485 26480
rect 4919 26440 4928 26480
rect 4968 26440 5010 26480
rect 5050 26440 5092 26480
rect 5132 26440 5174 26480
rect 5214 26440 5256 26480
rect 5296 26440 5305 26480
rect 5356 26440 5644 26480
rect 5684 26440 5693 26480
rect 6414 26440 6508 26480
rect 6548 26440 6557 26480
rect 7182 26440 7276 26480
rect 7316 26440 7325 26480
rect 16483 26440 16492 26480
rect 16532 26440 17356 26480
rect 17396 26440 17405 26480
rect 18403 26440 18412 26480
rect 18452 26440 19660 26480
rect 19700 26440 19709 26480
rect 20039 26440 20048 26480
rect 20088 26440 20130 26480
rect 20170 26440 20212 26480
rect 20252 26440 20294 26480
rect 20334 26440 20376 26480
rect 20416 26440 20425 26480
rect 21379 26440 21388 26480
rect 21428 26440 21504 26480
rect 1315 26439 1373 26440
rect 2467 26396 2525 26397
rect 2083 26356 2092 26396
rect 2132 26356 2476 26396
rect 2516 26356 2525 26396
rect 2467 26355 2525 26356
rect 2947 26396 3005 26397
rect 3331 26396 3389 26397
rect 2947 26356 2956 26396
rect 2996 26356 3340 26396
rect 3380 26356 3389 26396
rect 3436 26396 3476 26440
rect 5635 26439 5693 26440
rect 6499 26439 6557 26440
rect 7267 26439 7325 26440
rect 19651 26439 19709 26440
rect 21424 26420 21504 26440
rect 3715 26396 3773 26397
rect 7747 26396 7805 26397
rect 8611 26396 8669 26397
rect 18691 26396 18749 26397
rect 3436 26356 3724 26396
rect 3764 26356 3773 26396
rect 6307 26356 6316 26396
rect 6356 26356 6604 26396
rect 6644 26356 6653 26396
rect 7747 26356 7756 26396
rect 7796 26356 8620 26396
rect 8660 26356 11360 26396
rect 15235 26356 15244 26396
rect 15284 26356 15820 26396
rect 15860 26356 15869 26396
rect 16003 26356 16012 26396
rect 16052 26356 17164 26396
rect 17204 26356 17213 26396
rect 18499 26356 18508 26396
rect 18548 26356 18700 26396
rect 18740 26356 18749 26396
rect 2947 26355 3005 26356
rect 3331 26355 3389 26356
rect 3715 26355 3773 26356
rect 7747 26355 7805 26356
rect 8611 26355 8669 26356
rect 0 26312 80 26332
rect 3427 26312 3485 26313
rect 6403 26312 6461 26313
rect 10051 26312 10109 26313
rect 11107 26312 11165 26313
rect 0 26272 3436 26312
rect 3476 26272 3485 26312
rect 3619 26272 3628 26312
rect 3668 26272 4012 26312
rect 4052 26272 4061 26312
rect 6318 26272 6412 26312
rect 6452 26272 6461 26312
rect 0 26252 80 26272
rect 3427 26271 3485 26272
rect 6403 26271 6461 26272
rect 6508 26272 6892 26312
rect 6932 26272 6941 26312
rect 7363 26272 7372 26312
rect 7412 26272 7852 26312
rect 7892 26272 7901 26312
rect 8419 26272 8428 26312
rect 8468 26272 10060 26312
rect 10100 26272 10109 26312
rect 11022 26272 11116 26312
rect 11156 26272 11165 26312
rect 11320 26312 11360 26356
rect 18691 26355 18749 26356
rect 11875 26312 11933 26313
rect 11320 26272 11500 26312
rect 11540 26272 11549 26312
rect 11790 26272 11884 26312
rect 11924 26272 11933 26312
rect 15427 26272 15436 26312
rect 15476 26272 15724 26312
rect 15764 26272 15773 26312
rect 16579 26272 16588 26312
rect 16628 26272 16876 26312
rect 16916 26272 17452 26312
rect 17492 26272 17501 26312
rect 18979 26272 18988 26312
rect 19028 26272 19756 26312
rect 19796 26272 19805 26312
rect 3204 26188 3241 26228
rect 3281 26188 3290 26228
rect 4675 26188 4684 26228
rect 4724 26188 4876 26228
rect 4916 26188 4925 26228
rect 2467 26144 2525 26145
rect 3244 26144 3284 26188
rect 4483 26144 4541 26145
rect 6508 26144 6548 26272
rect 10051 26271 10109 26272
rect 11107 26271 11165 26272
rect 11875 26271 11933 26272
rect 10243 26228 10301 26229
rect 15139 26228 15197 26229
rect 16771 26228 16829 26229
rect 10243 26188 10252 26228
rect 10292 26188 10540 26228
rect 10580 26188 12076 26228
rect 12116 26188 12125 26228
rect 13804 26188 15148 26228
rect 15188 26188 15197 26228
rect 15331 26188 15340 26228
rect 15380 26188 16012 26228
rect 16052 26188 16061 26228
rect 16678 26188 16687 26228
rect 16727 26188 16780 26228
rect 16820 26188 16829 26228
rect 10243 26187 10301 26188
rect 8419 26144 8477 26145
rect 2381 26104 2476 26144
rect 2516 26104 2764 26144
rect 2804 26104 2813 26144
rect 2947 26104 2956 26144
rect 2996 26104 4108 26144
rect 4148 26104 4157 26144
rect 4483 26104 4492 26144
rect 4532 26104 5356 26144
rect 5396 26104 6548 26144
rect 6595 26104 6604 26144
rect 6644 26104 7852 26144
rect 7892 26104 7901 26144
rect 8334 26104 8428 26144
rect 8468 26104 8477 26144
rect 2467 26103 2525 26104
rect 4483 26103 4541 26104
rect 6508 26061 6548 26104
rect 8419 26103 8477 26104
rect 8611 26144 8669 26145
rect 13804 26144 13844 26188
rect 15139 26187 15197 26188
rect 16771 26187 16829 26188
rect 16675 26144 16733 26145
rect 17731 26144 17789 26145
rect 18403 26144 18461 26145
rect 8611 26104 8620 26144
rect 8660 26104 9868 26144
rect 9908 26104 9917 26144
rect 10051 26104 10060 26144
rect 10100 26104 13844 26144
rect 13987 26104 13996 26144
rect 14036 26104 14045 26144
rect 15427 26104 15436 26144
rect 15476 26104 16108 26144
rect 16148 26104 16157 26144
rect 16204 26104 16684 26144
rect 16724 26104 17548 26144
rect 17588 26104 17597 26144
rect 17731 26104 17740 26144
rect 17780 26104 18412 26144
rect 18452 26104 18988 26144
rect 19028 26104 19037 26144
rect 8611 26103 8669 26104
rect 6499 26060 6557 26061
rect 13996 26060 14036 26104
rect 16204 26060 16244 26104
rect 16675 26103 16733 26104
rect 17731 26103 17789 26104
rect 18403 26103 18461 26104
rect 1219 26020 1228 26060
rect 1268 26020 3628 26060
rect 3668 26020 4588 26060
rect 4628 26020 4637 26060
rect 5059 26020 5068 26060
rect 5108 26020 5932 26060
rect 5972 26020 5981 26060
rect 6499 26020 6508 26060
rect 6548 26020 6557 26060
rect 0 25976 80 25996
rect 0 25936 212 25976
rect 0 25916 80 25936
rect 172 25808 212 25936
rect 3340 25892 3380 26020
rect 6499 26019 6557 26020
rect 7468 26020 14036 26060
rect 15811 26020 15820 26060
rect 15860 26020 16244 26060
rect 16771 26020 16780 26060
rect 16820 26020 17356 26060
rect 17396 26020 17405 26060
rect 17731 26020 17740 26060
rect 17780 26020 19948 26060
rect 19988 26020 19997 26060
rect 4195 25976 4253 25977
rect 4110 25936 4204 25976
rect 4244 25936 4253 25976
rect 4195 25935 4253 25936
rect 6211 25892 6269 25893
rect 7468 25892 7508 26020
rect 13027 25976 13085 25977
rect 21424 25976 21504 25996
rect 8803 25936 8812 25976
rect 8852 25936 9676 25976
rect 9716 25936 9725 25976
rect 9859 25936 9868 25976
rect 9908 25936 13036 25976
rect 13076 25936 13085 25976
rect 19843 25936 19852 25976
rect 19892 25936 20180 25976
rect 20515 25936 20524 25976
rect 20564 25936 21504 25976
rect 13027 25935 13085 25936
rect 3331 25852 3340 25892
rect 3380 25852 3389 25892
rect 3619 25852 3628 25892
rect 3668 25852 4588 25892
rect 4628 25852 4637 25892
rect 6211 25852 6220 25892
rect 6260 25852 7564 25892
rect 7604 25852 7632 25892
rect 9100 25852 17740 25892
rect 17780 25852 17789 25892
rect 18700 25852 18892 25892
rect 18932 25852 18941 25892
rect 19171 25852 19180 25892
rect 19220 25852 19468 25892
rect 19508 25852 19517 25892
rect 6211 25851 6269 25852
rect 6307 25808 6365 25809
rect 172 25768 2540 25808
rect 3427 25768 3436 25808
rect 3476 25768 6316 25808
rect 6356 25768 6365 25808
rect 6499 25768 6508 25808
rect 6548 25768 6988 25808
rect 7028 25768 7037 25808
rect 7171 25768 7180 25808
rect 7220 25768 8236 25808
rect 8276 25768 9004 25808
rect 9044 25768 9053 25808
rect 0 25640 80 25660
rect 2500 25640 2540 25768
rect 6307 25767 6365 25768
rect 7171 25724 7229 25725
rect 9100 25724 9140 25852
rect 12355 25768 12364 25808
rect 12404 25768 17548 25808
rect 17588 25768 17597 25808
rect 3679 25684 3688 25724
rect 3728 25684 3770 25724
rect 3810 25684 3852 25724
rect 3892 25684 3934 25724
rect 3974 25684 4016 25724
rect 4056 25684 4065 25724
rect 7171 25684 7180 25724
rect 7220 25684 9140 25724
rect 10051 25724 10109 25725
rect 16771 25724 16829 25725
rect 10051 25684 10060 25724
rect 10100 25684 15244 25724
rect 15284 25684 15293 25724
rect 16771 25684 16780 25724
rect 16820 25684 17164 25724
rect 17204 25684 17213 25724
rect 7171 25683 7229 25684
rect 10051 25683 10109 25684
rect 16771 25683 16829 25684
rect 18700 25640 18740 25852
rect 20140 25808 20180 25936
rect 21424 25916 21504 25936
rect 20140 25768 21388 25808
rect 21428 25768 21437 25808
rect 18799 25684 18808 25724
rect 18848 25684 18890 25724
rect 18930 25684 18972 25724
rect 19012 25684 19054 25724
rect 19094 25684 19136 25724
rect 19176 25684 19185 25724
rect 19555 25684 19564 25724
rect 19604 25684 21100 25724
rect 21140 25684 21149 25724
rect 0 25600 940 25640
rect 980 25600 989 25640
rect 2500 25600 11360 25640
rect 12259 25600 12268 25640
rect 12308 25600 13900 25640
rect 13940 25600 18508 25640
rect 18548 25600 18557 25640
rect 18700 25600 19028 25640
rect 0 25580 80 25600
rect 3331 25556 3389 25557
rect 4675 25556 4733 25557
rect 3331 25516 3340 25556
rect 3380 25516 3628 25556
rect 3668 25516 3677 25556
rect 4675 25516 4684 25556
rect 4724 25516 8812 25556
rect 8852 25516 8861 25556
rect 3331 25515 3389 25516
rect 4675 25515 4733 25516
rect 11320 25472 11360 25600
rect 14083 25556 14141 25557
rect 18019 25556 18077 25557
rect 18988 25556 19028 25600
rect 13987 25516 13996 25556
rect 14036 25516 14092 25556
rect 14132 25516 14141 25556
rect 15523 25516 15532 25556
rect 15572 25516 17260 25556
rect 17300 25516 17309 25556
rect 18019 25516 18028 25556
rect 18068 25516 18700 25556
rect 18740 25516 18749 25556
rect 18979 25516 18988 25556
rect 19028 25516 19037 25556
rect 19651 25516 19660 25556
rect 19700 25516 20130 25556
rect 20170 25516 20179 25556
rect 14083 25515 14141 25516
rect 18019 25515 18077 25516
rect 16195 25472 16253 25473
rect 16771 25472 16829 25473
rect 21424 25472 21504 25492
rect 3235 25432 3244 25472
rect 3284 25432 4300 25472
rect 4340 25432 4349 25472
rect 6796 25432 8276 25472
rect 11320 25432 15436 25472
rect 15476 25432 15485 25472
rect 16195 25432 16204 25472
rect 16244 25432 16780 25472
rect 16820 25432 16829 25472
rect 17539 25432 17548 25472
rect 17588 25432 18220 25472
rect 18260 25432 18892 25472
rect 18932 25432 18941 25472
rect 19267 25432 19276 25472
rect 19316 25432 19852 25472
rect 19892 25432 19901 25472
rect 21379 25432 21388 25472
rect 21428 25432 21504 25472
rect 2275 25388 2333 25389
rect 5443 25388 5501 25389
rect 1315 25348 1324 25388
rect 1364 25348 2284 25388
rect 2324 25348 2333 25388
rect 4867 25348 4876 25388
rect 4916 25348 5452 25388
rect 5492 25348 5501 25388
rect 2275 25347 2333 25348
rect 5443 25347 5501 25348
rect 5731 25388 5789 25389
rect 6796 25388 6836 25432
rect 5731 25348 5740 25388
rect 5780 25348 6836 25388
rect 5731 25347 5789 25348
rect 0 25304 80 25324
rect 6979 25304 7037 25305
rect 8236 25304 8276 25432
rect 16195 25431 16253 25432
rect 16771 25431 16829 25432
rect 21424 25412 21504 25432
rect 11587 25388 11645 25389
rect 13123 25388 13181 25389
rect 11502 25348 11596 25388
rect 11636 25348 11645 25388
rect 11587 25347 11645 25348
rect 12172 25348 12364 25388
rect 12404 25348 12413 25388
rect 12739 25348 12748 25388
rect 12788 25348 13132 25388
rect 13172 25348 13181 25388
rect 12172 25304 12212 25348
rect 13123 25347 13181 25348
rect 13603 25388 13661 25389
rect 15523 25388 15581 25389
rect 18499 25388 18557 25389
rect 19939 25388 19997 25389
rect 13603 25348 13612 25388
rect 13652 25348 15532 25388
rect 15572 25348 15581 25388
rect 16483 25348 16492 25388
rect 16532 25348 16780 25388
rect 16820 25348 16829 25388
rect 18499 25348 18508 25388
rect 18548 25348 19316 25388
rect 19854 25348 19948 25388
rect 19988 25348 19997 25388
rect 13603 25347 13661 25348
rect 15523 25347 15581 25348
rect 18499 25347 18557 25348
rect 12835 25304 12893 25305
rect 15811 25304 15869 25305
rect 17731 25304 17789 25305
rect 19276 25304 19316 25348
rect 19939 25347 19997 25348
rect 0 25264 5164 25304
rect 5204 25264 5213 25304
rect 5539 25264 5548 25304
rect 5588 25264 5932 25304
rect 5972 25264 5981 25304
rect 6595 25264 6604 25304
rect 6644 25264 6988 25304
rect 7028 25264 7468 25304
rect 7508 25264 7517 25304
rect 8236 25264 12212 25304
rect 12259 25264 12268 25304
rect 12308 25264 12844 25304
rect 12884 25264 14572 25304
rect 14612 25264 14621 25304
rect 15427 25264 15436 25304
rect 15476 25264 15820 25304
rect 15860 25264 16108 25304
rect 16148 25264 16157 25304
rect 17443 25264 17452 25304
rect 17492 25264 17740 25304
rect 17780 25264 17789 25304
rect 19267 25264 19276 25304
rect 19316 25264 19325 25304
rect 20140 25264 20236 25304
rect 20276 25264 20285 25304
rect 0 25244 80 25264
rect 6979 25263 7037 25264
rect 12835 25263 12893 25264
rect 15811 25263 15869 25264
rect 17731 25263 17789 25264
rect 5923 25220 5981 25221
rect 8227 25220 8285 25221
rect 14083 25220 14141 25221
rect 2500 25180 3572 25220
rect 4003 25180 4012 25220
rect 4052 25180 5068 25220
rect 5108 25180 5260 25220
rect 5300 25180 5309 25220
rect 5836 25180 5932 25220
rect 5972 25180 5981 25220
rect 2500 25136 2540 25180
rect 3235 25136 3293 25137
rect 3532 25136 3572 25180
rect 5836 25136 5876 25180
rect 5923 25179 5981 25180
rect 6220 25180 7660 25220
rect 7700 25180 7709 25220
rect 8227 25180 8236 25220
rect 8276 25180 8620 25220
rect 8660 25180 8669 25220
rect 13998 25180 14092 25220
rect 14132 25180 14141 25220
rect 6220 25136 6260 25180
rect 8227 25179 8285 25180
rect 14083 25179 14141 25180
rect 15139 25220 15197 25221
rect 16195 25220 16253 25221
rect 16579 25220 16637 25221
rect 17059 25220 17117 25221
rect 17740 25220 17780 25263
rect 15139 25180 15148 25220
rect 15188 25180 16204 25220
rect 16244 25180 16253 25220
rect 16483 25180 16492 25220
rect 16532 25180 16588 25220
rect 16628 25180 16637 25220
rect 15139 25179 15197 25180
rect 16195 25179 16253 25180
rect 16579 25179 16637 25180
rect 16684 25180 17068 25220
rect 17108 25180 17117 25220
rect 17731 25180 17740 25220
rect 17780 25180 17789 25220
rect 18019 25180 18028 25220
rect 18068 25180 19564 25220
rect 19604 25180 19613 25220
rect 1699 25096 1708 25136
rect 1748 25096 2540 25136
rect 2659 25096 2668 25136
rect 2708 25096 2717 25136
rect 3150 25096 3244 25136
rect 3284 25096 3293 25136
rect 3523 25096 3532 25136
rect 3572 25096 3581 25136
rect 5347 25096 5356 25136
rect 5396 25096 5644 25136
rect 5684 25096 5693 25136
rect 5827 25096 5836 25136
rect 5876 25096 5885 25136
rect 6211 25096 6220 25136
rect 6260 25096 6269 25136
rect 2668 25052 2708 25096
rect 3235 25095 3293 25096
rect 2467 25012 2476 25052
rect 2516 25012 2708 25052
rect 0 24968 80 24988
rect 163 24968 221 24969
rect 8236 24968 8276 25179
rect 10435 25136 10493 25137
rect 12163 25136 12221 25137
rect 15427 25136 15485 25137
rect 16684 25136 16724 25180
rect 17059 25179 17117 25180
rect 19363 25136 19421 25137
rect 10435 25096 10444 25136
rect 10484 25096 12172 25136
rect 12212 25096 12221 25136
rect 13987 25096 13996 25136
rect 14036 25096 14045 25136
rect 15427 25096 15436 25136
rect 15476 25096 15820 25136
rect 15860 25096 16204 25136
rect 16244 25096 16253 25136
rect 16675 25096 16684 25136
rect 16724 25096 16733 25136
rect 19278 25096 19372 25136
rect 19412 25096 19421 25136
rect 10435 25095 10493 25096
rect 12163 25095 12221 25096
rect 8611 25052 8669 25053
rect 11971 25052 12029 25053
rect 13996 25052 14036 25096
rect 15427 25095 15485 25096
rect 19363 25095 19421 25096
rect 20140 25052 20180 25264
rect 20323 25096 20332 25136
rect 20372 25096 21388 25136
rect 21428 25096 21437 25136
rect 8611 25012 8620 25052
rect 8660 25012 9196 25052
rect 9236 25012 10060 25052
rect 10100 25012 10109 25052
rect 11971 25012 11980 25052
rect 12020 25012 14036 25052
rect 15235 25012 15244 25052
rect 15284 25012 17452 25052
rect 17492 25012 17501 25052
rect 18307 25012 18316 25052
rect 18356 25012 20180 25052
rect 8611 25011 8669 25012
rect 11971 25011 12029 25012
rect 14083 24968 14141 24969
rect 21424 24968 21504 24988
rect 0 24928 172 24968
rect 212 24928 221 24968
rect 4919 24928 4928 24968
rect 4968 24928 5010 24968
rect 5050 24928 5092 24968
rect 5132 24928 5174 24968
rect 5214 24928 5256 24968
rect 5296 24928 5305 24968
rect 8227 24928 8236 24968
rect 8276 24928 8285 24968
rect 8611 24928 8620 24968
rect 8660 24928 9388 24968
rect 9428 24928 9437 24968
rect 9676 24928 14092 24968
rect 14132 24928 14141 24968
rect 20039 24928 20048 24968
rect 20088 24928 20130 24968
rect 20170 24928 20212 24968
rect 20252 24928 20294 24968
rect 20334 24928 20376 24968
rect 20416 24928 20425 24968
rect 21379 24928 21388 24968
rect 21428 24928 21504 24968
rect 0 24908 80 24928
rect 163 24927 221 24928
rect 9676 24884 9716 24928
rect 14083 24927 14141 24928
rect 21424 24908 21504 24928
rect 3619 24844 3628 24884
rect 3668 24844 9716 24884
rect 9763 24884 9821 24885
rect 9763 24844 9772 24884
rect 9812 24844 9868 24884
rect 9908 24844 9917 24884
rect 11779 24844 11788 24884
rect 11828 24844 11837 24884
rect 14860 24844 18028 24884
rect 18068 24844 18077 24884
rect 9763 24843 9821 24844
rect 5443 24800 5501 24801
rect 10819 24800 10877 24801
rect 2659 24760 2668 24800
rect 2708 24760 5452 24800
rect 5492 24760 5501 24800
rect 6499 24760 6508 24800
rect 6548 24760 8524 24800
rect 8564 24760 8573 24800
rect 8707 24760 8716 24800
rect 8756 24760 10828 24800
rect 10868 24760 10877 24800
rect 11788 24800 11828 24844
rect 11788 24760 13996 24800
rect 14036 24760 14045 24800
rect 5443 24759 5501 24760
rect 10819 24759 10877 24760
rect 4579 24716 4637 24717
rect 11875 24716 11933 24717
rect 14860 24716 14900 24844
rect 14947 24800 15005 24801
rect 14947 24760 14956 24800
rect 14996 24760 21196 24800
rect 21236 24760 21245 24800
rect 14947 24759 15005 24760
rect 18595 24716 18653 24717
rect 3139 24676 3148 24716
rect 3188 24676 4396 24716
rect 4436 24676 4445 24716
rect 4579 24676 4588 24716
rect 4628 24676 4780 24716
rect 4820 24676 10964 24716
rect 4579 24675 4637 24676
rect 0 24632 80 24652
rect 1219 24632 1277 24633
rect 0 24592 1228 24632
rect 1268 24592 1277 24632
rect 0 24572 80 24592
rect 1219 24591 1277 24592
rect 1411 24632 1469 24633
rect 10924 24632 10964 24676
rect 11875 24676 11884 24716
rect 11924 24676 14900 24716
rect 18211 24676 18220 24716
rect 18260 24676 18300 24716
rect 18510 24676 18604 24716
rect 18644 24676 18653 24716
rect 11875 24675 11933 24676
rect 13027 24632 13085 24633
rect 18220 24632 18260 24676
rect 18595 24675 18653 24676
rect 1411 24592 1420 24632
rect 1460 24592 1996 24632
rect 2036 24592 2045 24632
rect 2467 24592 2476 24632
rect 2516 24592 3820 24632
rect 3860 24592 3869 24632
rect 4099 24592 4108 24632
rect 4148 24592 5548 24632
rect 5588 24592 5597 24632
rect 6307 24592 6316 24632
rect 6356 24592 7180 24632
rect 7220 24592 7229 24632
rect 8323 24592 8332 24632
rect 8372 24592 8524 24632
rect 8564 24592 8573 24632
rect 8995 24592 9004 24632
rect 9044 24592 9292 24632
rect 9332 24592 9341 24632
rect 9859 24592 9868 24632
rect 9908 24592 10444 24632
rect 10484 24592 10493 24632
rect 10915 24592 10924 24632
rect 10964 24592 10973 24632
rect 12942 24592 13036 24632
rect 13076 24592 13085 24632
rect 14371 24592 14380 24632
rect 14420 24592 14860 24632
rect 14900 24592 14909 24632
rect 16483 24592 16492 24632
rect 16532 24592 17260 24632
rect 17300 24592 17309 24632
rect 17923 24592 17932 24632
rect 17972 24592 18988 24632
rect 19028 24592 19037 24632
rect 19267 24592 19276 24632
rect 19316 24592 19948 24632
rect 19988 24592 19997 24632
rect 1411 24591 1469 24592
rect 2467 24548 2525 24549
rect 3820 24548 3860 24592
rect 13027 24591 13085 24592
rect 8419 24548 8477 24549
rect 17731 24548 17789 24549
rect 2467 24508 2476 24548
rect 2516 24508 3764 24548
rect 3820 24508 5356 24548
rect 5396 24508 5405 24548
rect 6412 24508 6892 24548
rect 6932 24508 8428 24548
rect 8468 24508 8477 24548
rect 10339 24508 10348 24548
rect 10388 24508 11308 24548
rect 11348 24508 11980 24548
rect 12020 24508 12029 24548
rect 14275 24508 14284 24548
rect 14324 24508 16108 24548
rect 16148 24508 16588 24548
rect 16628 24508 16637 24548
rect 17731 24508 17740 24548
rect 17780 24508 17836 24548
rect 17876 24508 17885 24548
rect 19843 24508 19852 24548
rect 19892 24508 19901 24548
rect 2467 24507 2525 24508
rect 2371 24464 2429 24465
rect 3724 24464 3764 24508
rect 6412 24464 6452 24508
rect 8419 24507 8477 24508
rect 17731 24507 17789 24508
rect 19852 24464 19892 24508
rect 21424 24464 21504 24484
rect 2371 24424 2380 24464
rect 2420 24424 2668 24464
rect 2708 24424 2717 24464
rect 2851 24424 2860 24464
rect 2900 24424 3052 24464
rect 3092 24424 3436 24464
rect 3476 24424 3485 24464
rect 3724 24424 6452 24464
rect 6499 24424 6508 24464
rect 6548 24424 9772 24464
rect 9812 24424 9821 24464
rect 11320 24424 19892 24464
rect 20035 24424 20044 24464
rect 20084 24424 21504 24464
rect 2371 24423 2429 24424
rect 11320 24380 11360 24424
rect 21424 24404 21504 24424
rect 3619 24340 3628 24380
rect 3668 24340 4396 24380
rect 4436 24340 4445 24380
rect 8131 24340 8140 24380
rect 8180 24340 11360 24380
rect 12643 24340 12652 24380
rect 12692 24340 14956 24380
rect 14996 24340 15005 24380
rect 0 24296 80 24316
rect 0 24256 8908 24296
rect 8948 24256 9196 24296
rect 9236 24256 9245 24296
rect 10723 24256 10732 24296
rect 10772 24256 13420 24296
rect 13460 24256 13469 24296
rect 0 24236 80 24256
rect 4771 24212 4829 24213
rect 10627 24212 10685 24213
rect 2275 24172 2284 24212
rect 2324 24172 3572 24212
rect 3679 24172 3688 24212
rect 3728 24172 3770 24212
rect 3810 24172 3852 24212
rect 3892 24172 3934 24212
rect 3974 24172 4016 24212
rect 4056 24172 4065 24212
rect 4771 24172 4780 24212
rect 4820 24172 8140 24212
rect 8180 24172 8189 24212
rect 8707 24172 8716 24212
rect 8756 24172 9292 24212
rect 9332 24172 9341 24212
rect 10627 24172 10636 24212
rect 10676 24172 11020 24212
rect 11060 24172 11069 24212
rect 12835 24172 12844 24212
rect 12884 24172 13324 24212
rect 13364 24172 13373 24212
rect 18799 24172 18808 24212
rect 18848 24172 18890 24212
rect 18930 24172 18972 24212
rect 19012 24172 19054 24212
rect 19094 24172 19136 24212
rect 19176 24172 19185 24212
rect 3532 24128 3572 24172
rect 4771 24171 4829 24172
rect 10627 24171 10685 24172
rect 3532 24088 4876 24128
rect 4916 24088 9868 24128
rect 9908 24088 9917 24128
rect 10435 24088 10444 24128
rect 10484 24088 11212 24128
rect 11252 24088 11884 24128
rect 11924 24088 11933 24128
rect 13507 24044 13565 24045
rect 835 24004 844 24044
rect 884 24004 2540 24044
rect 3427 24004 3436 24044
rect 3476 24004 4012 24044
rect 4052 24004 4061 24044
rect 4108 24004 5644 24044
rect 5684 24004 5693 24044
rect 7747 24004 7756 24044
rect 7796 24004 9388 24044
rect 9428 24004 11404 24044
rect 11444 24004 11453 24044
rect 12835 24004 12844 24044
rect 12884 24004 13516 24044
rect 13556 24004 13565 24044
rect 16003 24004 16012 24044
rect 16052 24004 16061 24044
rect 0 23960 80 23980
rect 2500 23960 2540 24004
rect 4108 23960 4148 24004
rect 9772 23960 9812 24004
rect 13507 24003 13565 24004
rect 10531 23960 10589 23961
rect 0 23920 652 23960
rect 692 23920 701 23960
rect 2500 23920 3340 23960
rect 3380 23920 4148 23960
rect 4195 23920 4204 23960
rect 4244 23920 4972 23960
rect 5012 23920 5021 23960
rect 8707 23920 8716 23960
rect 8756 23920 9676 23960
rect 9716 23920 9725 23960
rect 9772 23920 9841 23960
rect 9881 23920 9890 23960
rect 9955 23920 9964 23960
rect 10004 23920 10013 23960
rect 10446 23920 10540 23960
rect 10580 23920 10589 23960
rect 0 23900 80 23920
rect 1603 23876 1661 23877
rect 1518 23836 1612 23876
rect 1652 23836 1661 23876
rect 1603 23835 1661 23836
rect 4291 23876 4349 23877
rect 9964 23876 10004 23920
rect 10531 23919 10589 23920
rect 10819 23960 10877 23961
rect 10819 23920 10828 23960
rect 10868 23920 10924 23960
rect 10964 23920 10973 23960
rect 10819 23919 10877 23920
rect 4291 23836 4300 23876
rect 4340 23836 4780 23876
rect 4820 23836 4829 23876
rect 6403 23836 6412 23876
rect 6452 23836 7988 23876
rect 8323 23836 8332 23876
rect 8372 23836 10004 23876
rect 10051 23836 10060 23876
rect 10100 23836 11060 23876
rect 11107 23836 11116 23876
rect 11156 23836 11165 23876
rect 13795 23836 13804 23876
rect 13844 23836 14380 23876
rect 14420 23836 14429 23876
rect 4291 23835 4349 23836
rect 1891 23792 1949 23793
rect 3043 23792 3101 23793
rect 7075 23792 7133 23793
rect 1806 23752 1900 23792
rect 1940 23752 1949 23792
rect 2563 23752 2572 23792
rect 2612 23752 2621 23792
rect 2958 23752 3052 23792
rect 3092 23752 3101 23792
rect 3331 23752 3340 23792
rect 3380 23752 4492 23792
rect 4532 23752 4541 23792
rect 6883 23752 6892 23792
rect 6932 23752 7084 23792
rect 7124 23752 7133 23792
rect 7948 23792 7988 23836
rect 10531 23792 10589 23793
rect 11020 23792 11060 23836
rect 11116 23792 11156 23836
rect 12259 23792 12317 23793
rect 7948 23752 8716 23792
rect 8756 23752 8765 23792
rect 9763 23752 9772 23792
rect 9812 23752 10540 23792
rect 10580 23752 10589 23792
rect 11011 23752 11020 23792
rect 11060 23752 11069 23792
rect 11116 23752 12268 23792
rect 12308 23752 12556 23792
rect 12596 23752 12605 23792
rect 12739 23752 12748 23792
rect 12788 23752 15052 23792
rect 15092 23752 15101 23792
rect 1891 23751 1949 23752
rect 2572 23708 2612 23752
rect 3043 23751 3101 23752
rect 7075 23751 7133 23752
rect 10531 23751 10589 23752
rect 12259 23751 12317 23752
rect 11779 23708 11837 23709
rect 15331 23708 15389 23709
rect 16012 23708 16052 24004
rect 17923 23960 17981 23961
rect 18403 23960 18461 23961
rect 17838 23920 17932 23960
rect 17972 23920 17981 23960
rect 18318 23920 18412 23960
rect 18452 23920 18461 23960
rect 17923 23919 17981 23920
rect 18403 23919 18461 23920
rect 19363 23960 19421 23961
rect 20515 23960 20573 23961
rect 21424 23960 21504 23980
rect 19363 23920 19372 23960
rect 19412 23920 19468 23960
rect 19508 23920 19517 23960
rect 20131 23920 20140 23960
rect 20180 23920 20524 23960
rect 20564 23920 20573 23960
rect 20995 23920 21004 23960
rect 21044 23920 21504 23960
rect 19363 23919 19421 23920
rect 20515 23919 20573 23920
rect 21424 23900 21504 23920
rect 19843 23876 19901 23877
rect 17731 23836 17740 23876
rect 17780 23836 18508 23876
rect 18548 23836 18557 23876
rect 19747 23836 19756 23876
rect 19796 23836 19852 23876
rect 19892 23836 19901 23876
rect 19843 23835 19901 23836
rect 16291 23792 16349 23793
rect 19363 23792 19421 23793
rect 16291 23752 16300 23792
rect 16340 23752 17836 23792
rect 17876 23752 17885 23792
rect 18019 23752 18028 23792
rect 18068 23752 18412 23792
rect 18452 23752 18461 23792
rect 19267 23752 19276 23792
rect 19316 23752 19372 23792
rect 19412 23752 19421 23792
rect 16291 23751 16349 23752
rect 19363 23751 19421 23752
rect 16579 23708 16637 23709
rect 18499 23708 18557 23709
rect 2572 23668 4588 23708
rect 4628 23668 10540 23708
rect 10580 23668 10589 23708
rect 11779 23668 11788 23708
rect 11828 23668 15340 23708
rect 15380 23668 15389 23708
rect 16003 23668 16012 23708
rect 16052 23668 16061 23708
rect 16579 23668 16588 23708
rect 16628 23668 18508 23708
rect 18548 23668 18557 23708
rect 0 23624 80 23644
rect 3715 23624 3773 23625
rect 9763 23624 9821 23625
rect 0 23584 460 23624
rect 500 23584 509 23624
rect 2179 23584 2188 23624
rect 2228 23584 3724 23624
rect 3764 23584 3773 23624
rect 8707 23584 8716 23624
rect 8756 23584 9484 23624
rect 9524 23584 9533 23624
rect 9763 23584 9772 23624
rect 9812 23584 9868 23624
rect 9908 23584 9917 23624
rect 0 23564 80 23584
rect 3715 23583 3773 23584
rect 9763 23583 9821 23584
rect 4099 23540 4157 23541
rect 4099 23500 4108 23540
rect 4148 23500 7852 23540
rect 7892 23500 8140 23540
rect 8180 23500 8189 23540
rect 4099 23499 4157 23500
rect 2755 23456 2813 23457
rect 8611 23456 8669 23457
rect 10156 23456 10196 23668
rect 11779 23667 11837 23668
rect 15331 23667 15389 23668
rect 16579 23667 16637 23668
rect 18499 23667 18557 23668
rect 16195 23584 16204 23624
rect 16244 23584 17452 23624
rect 17492 23584 18316 23624
rect 18356 23584 18365 23624
rect 19939 23584 19948 23624
rect 19988 23584 21428 23624
rect 16579 23500 16588 23540
rect 16628 23500 16780 23540
rect 16820 23500 16829 23540
rect 21388 23476 21428 23584
rect 10531 23456 10589 23457
rect 2755 23416 2764 23456
rect 2804 23416 4780 23456
rect 4820 23416 4829 23456
rect 4919 23416 4928 23456
rect 4968 23416 5010 23456
rect 5050 23416 5092 23456
rect 5132 23416 5174 23456
rect 5214 23416 5256 23456
rect 5296 23416 5305 23456
rect 6508 23416 8620 23456
rect 8660 23416 8669 23456
rect 10147 23416 10156 23456
rect 10196 23416 10205 23456
rect 10531 23416 10540 23456
rect 10580 23416 10732 23456
rect 10772 23416 10781 23456
rect 20039 23416 20048 23456
rect 20088 23416 20130 23456
rect 20170 23416 20212 23456
rect 20252 23416 20294 23456
rect 20334 23416 20376 23456
rect 20416 23416 20425 23456
rect 21388 23416 21504 23476
rect 2755 23415 2813 23416
rect 3043 23372 3101 23373
rect 6508 23372 6548 23416
rect 8611 23415 8669 23416
rect 10531 23415 10589 23416
rect 21424 23396 21504 23416
rect 1699 23332 1708 23372
rect 1748 23332 2188 23372
rect 2228 23332 2237 23372
rect 3043 23332 3052 23372
rect 3092 23332 6548 23372
rect 6595 23332 6604 23372
rect 6644 23332 9292 23372
rect 9332 23332 9341 23372
rect 9955 23332 9964 23372
rect 10004 23332 10540 23372
rect 10580 23332 11500 23372
rect 11540 23332 11549 23372
rect 11596 23332 15820 23372
rect 15860 23332 15869 23372
rect 3043 23331 3101 23332
rect 0 23288 80 23308
rect 11596 23288 11636 23332
rect 11779 23288 11837 23289
rect 12643 23288 12701 23289
rect 0 23248 11636 23288
rect 11683 23248 11692 23288
rect 11732 23248 11788 23288
rect 11828 23248 11837 23288
rect 12451 23248 12460 23288
rect 12500 23248 12652 23288
rect 12692 23248 12701 23288
rect 0 23228 80 23248
rect 11779 23247 11837 23248
rect 12643 23247 12701 23248
rect 10051 23204 10109 23205
rect 1507 23164 1516 23204
rect 1556 23164 9236 23204
rect 2755 23120 2813 23121
rect 6691 23120 6749 23121
rect 9091 23120 9149 23121
rect 2755 23080 2764 23120
rect 2804 23080 2860 23120
rect 2900 23080 2909 23120
rect 3235 23080 3244 23120
rect 3284 23080 6124 23120
rect 6164 23080 6173 23120
rect 6606 23080 6700 23120
rect 6740 23080 6749 23120
rect 8035 23080 8044 23120
rect 8084 23080 8524 23120
rect 8564 23080 8573 23120
rect 9006 23080 9100 23120
rect 9140 23080 9149 23120
rect 9196 23120 9236 23164
rect 10051 23164 10060 23204
rect 10100 23164 10348 23204
rect 10388 23164 10397 23204
rect 11107 23164 11116 23204
rect 11156 23164 11596 23204
rect 11636 23164 11645 23204
rect 15715 23164 15724 23204
rect 15764 23164 16300 23204
rect 16340 23164 16349 23204
rect 17635 23164 17644 23204
rect 17684 23164 17836 23204
rect 17876 23164 19660 23204
rect 19700 23164 19709 23204
rect 10051 23163 10109 23164
rect 9571 23120 9629 23121
rect 15331 23120 15389 23121
rect 9196 23080 9580 23120
rect 9620 23080 13804 23120
rect 13844 23080 13853 23120
rect 15331 23080 15340 23120
rect 15380 23080 18412 23120
rect 18452 23080 18461 23120
rect 19171 23080 19180 23120
rect 19220 23080 19948 23120
rect 19988 23080 20236 23120
rect 20276 23080 20285 23120
rect 2755 23079 2813 23080
rect 6691 23079 6749 23080
rect 9091 23079 9149 23080
rect 9571 23079 9629 23080
rect 15331 23079 15389 23080
rect 4291 23036 4349 23037
rect 10819 23036 10877 23037
rect 19363 23036 19421 23037
rect 1027 22996 1036 23036
rect 1076 22996 1708 23036
rect 1748 22996 1757 23036
rect 2947 22996 2956 23036
rect 2996 22996 3036 23036
rect 4099 22996 4108 23036
rect 4148 22996 4300 23036
rect 4340 22996 4349 23036
rect 4483 22996 4492 23036
rect 4532 22996 5356 23036
rect 5396 22996 5405 23036
rect 8323 22996 8332 23036
rect 8372 22996 8812 23036
rect 8852 22996 8861 23036
rect 10734 22996 10828 23036
rect 10868 22996 10877 23036
rect 11299 22996 11308 23036
rect 11348 22996 11692 23036
rect 11732 22996 11741 23036
rect 14371 22996 14380 23036
rect 14420 22996 14764 23036
rect 14804 22996 14813 23036
rect 19363 22996 19372 23036
rect 19412 22996 20140 23036
rect 20180 22996 20189 23036
rect 0 22952 80 22972
rect 2956 22952 2996 22996
rect 4291 22995 4349 22996
rect 10819 22995 10877 22996
rect 19363 22995 19421 22996
rect 3427 22952 3485 22953
rect 8707 22952 8765 22953
rect 21424 22952 21504 22972
rect 0 22912 3436 22952
rect 3476 22912 3485 22952
rect 8622 22912 8716 22952
rect 8756 22912 8765 22952
rect 18211 22912 18220 22952
rect 18260 22912 21504 22952
rect 0 22892 80 22912
rect 3427 22911 3485 22912
rect 8707 22911 8765 22912
rect 21424 22892 21504 22912
rect 4099 22868 4157 22869
rect 12835 22868 12893 22869
rect 547 22828 556 22868
rect 596 22828 1516 22868
rect 1556 22828 1565 22868
rect 2947 22828 2956 22868
rect 2996 22828 3820 22868
rect 3860 22828 3869 22868
rect 4099 22828 4108 22868
rect 4148 22828 4157 22868
rect 4867 22828 4876 22868
rect 4916 22828 8332 22868
rect 8372 22828 8381 22868
rect 8611 22828 8620 22868
rect 8660 22828 10156 22868
rect 10196 22828 11308 22868
rect 11348 22828 11357 22868
rect 12643 22828 12652 22868
rect 12692 22828 12844 22868
rect 12884 22828 12893 22868
rect 4099 22827 4157 22828
rect 12835 22827 12893 22828
rect 4108 22784 4148 22827
rect 10531 22784 10589 22785
rect 2572 22744 4148 22784
rect 5347 22744 5356 22784
rect 5396 22744 6220 22784
rect 6260 22744 10540 22784
rect 10580 22744 10589 22784
rect 19363 22744 19372 22784
rect 19412 22744 19756 22784
rect 19796 22744 19805 22784
rect 2275 22700 2333 22701
rect 1411 22660 1420 22700
rect 1460 22660 2284 22700
rect 2324 22660 2333 22700
rect 2275 22659 2333 22660
rect 0 22616 80 22636
rect 2572 22616 2612 22744
rect 8716 22700 8756 22744
rect 10531 22743 10589 22744
rect 16483 22700 16541 22701
rect 2851 22660 2860 22700
rect 2900 22660 3436 22700
rect 3476 22660 3485 22700
rect 3679 22660 3688 22700
rect 3728 22660 3770 22700
rect 3810 22660 3852 22700
rect 3892 22660 3934 22700
rect 3974 22660 4016 22700
rect 4056 22660 4065 22700
rect 6787 22660 6796 22700
rect 6836 22660 6988 22700
rect 7028 22660 7037 22700
rect 8707 22660 8716 22700
rect 8756 22660 8765 22700
rect 8995 22660 9004 22700
rect 9044 22660 11116 22700
rect 11156 22660 11884 22700
rect 11924 22660 11933 22700
rect 15619 22660 15628 22700
rect 15668 22660 16492 22700
rect 16532 22660 16541 22700
rect 16483 22659 16541 22660
rect 17827 22700 17885 22701
rect 18691 22700 18749 22701
rect 19555 22700 19613 22701
rect 17827 22660 17836 22700
rect 17876 22660 18700 22700
rect 18740 22660 18749 22700
rect 18799 22660 18808 22700
rect 18848 22660 18890 22700
rect 18930 22660 18972 22700
rect 19012 22660 19054 22700
rect 19094 22660 19136 22700
rect 19176 22660 19185 22700
rect 19470 22660 19564 22700
rect 19604 22660 19613 22700
rect 19843 22660 19852 22700
rect 19892 22660 20044 22700
rect 20084 22660 20093 22700
rect 17827 22659 17885 22660
rect 18691 22659 18749 22660
rect 19555 22659 19613 22660
rect 19852 22616 19892 22660
rect 0 22576 1804 22616
rect 1844 22576 1853 22616
rect 2467 22576 2476 22616
rect 2516 22576 2612 22616
rect 3331 22576 3340 22616
rect 3380 22576 4300 22616
rect 4340 22576 4349 22616
rect 4867 22576 4876 22616
rect 4916 22576 4925 22616
rect 9091 22576 9100 22616
rect 9140 22576 11020 22616
rect 11060 22576 11980 22616
rect 12020 22576 12029 22616
rect 12739 22576 12748 22616
rect 12788 22576 13228 22616
rect 13268 22576 15532 22616
rect 15572 22576 15724 22616
rect 15764 22576 15773 22616
rect 17635 22576 17644 22616
rect 17684 22576 18028 22616
rect 18068 22576 19892 22616
rect 0 22556 80 22576
rect 3235 22532 3293 22533
rect 4876 22532 4916 22576
rect 1315 22492 1324 22532
rect 1364 22492 3244 22532
rect 3284 22492 4916 22532
rect 6307 22532 6365 22533
rect 19363 22532 19421 22533
rect 6307 22492 6316 22532
rect 6356 22492 6988 22532
rect 7028 22492 7037 22532
rect 13507 22492 13516 22532
rect 13556 22492 13565 22532
rect 19075 22492 19084 22532
rect 19124 22492 19372 22532
rect 19412 22492 19421 22532
rect 3235 22491 3293 22492
rect 6307 22491 6365 22492
rect 3523 22448 3581 22449
rect 13315 22448 13373 22449
rect 3139 22408 3148 22448
rect 3188 22408 3532 22448
rect 3572 22408 3581 22448
rect 4483 22408 4492 22448
rect 4532 22408 7660 22448
rect 7700 22408 7709 22448
rect 9283 22408 9292 22448
rect 9332 22408 13324 22448
rect 13364 22408 13373 22448
rect 3523 22407 3581 22408
rect 13315 22407 13373 22408
rect 7075 22364 7133 22365
rect 11299 22364 11357 22365
rect 2371 22324 2380 22364
rect 2420 22324 4396 22364
rect 4436 22324 4445 22364
rect 4492 22324 5452 22364
rect 5492 22324 5501 22364
rect 6990 22324 7084 22364
rect 7124 22324 8236 22364
rect 8276 22324 10156 22364
rect 10196 22324 10205 22364
rect 10339 22324 10348 22364
rect 10388 22324 10540 22364
rect 10580 22324 11308 22364
rect 11348 22324 11357 22364
rect 0 22280 80 22300
rect 1219 22280 1277 22281
rect 4492 22280 4532 22324
rect 7075 22323 7133 22324
rect 11299 22323 11357 22324
rect 5347 22280 5405 22281
rect 0 22240 1228 22280
rect 1268 22240 1277 22280
rect 1699 22240 1708 22280
rect 1748 22240 2188 22280
rect 2228 22240 4532 22280
rect 4675 22240 4684 22280
rect 4724 22240 5356 22280
rect 5396 22240 5405 22280
rect 7171 22240 7180 22280
rect 7220 22240 7564 22280
rect 7604 22240 7613 22280
rect 9667 22240 9676 22280
rect 9716 22240 10252 22280
rect 10292 22240 11020 22280
rect 11060 22240 12076 22280
rect 12116 22240 12125 22280
rect 0 22220 80 22240
rect 1219 22239 1277 22240
rect 5347 22239 5405 22240
rect 13516 22196 13556 22492
rect 19363 22491 19421 22492
rect 21424 22448 21504 22468
rect 18307 22408 18316 22448
rect 18356 22408 18796 22448
rect 18836 22408 18845 22448
rect 21187 22408 21196 22448
rect 21236 22408 21504 22448
rect 21424 22388 21504 22408
rect 14275 22324 14284 22364
rect 14324 22324 19564 22364
rect 19604 22324 19613 22364
rect 16483 22280 16541 22281
rect 17155 22280 17213 22281
rect 14179 22240 14188 22280
rect 14228 22240 16108 22280
rect 16148 22240 16492 22280
rect 16532 22240 16780 22280
rect 16820 22240 16829 22280
rect 17070 22240 17164 22280
rect 17204 22240 17213 22280
rect 18499 22240 18508 22280
rect 18548 22240 18557 22280
rect 16483 22239 16541 22240
rect 17155 22239 17213 22240
rect 13891 22196 13949 22197
rect 18508 22196 18548 22240
rect 5731 22156 5740 22196
rect 5780 22156 5789 22196
rect 7564 22156 7948 22196
rect 7988 22156 10100 22196
rect 10147 22156 10156 22196
rect 10196 22156 11404 22196
rect 11444 22156 11453 22196
rect 11683 22156 11692 22196
rect 11732 22156 12556 22196
rect 12596 22156 12605 22196
rect 13507 22156 13516 22196
rect 13556 22156 13565 22196
rect 13891 22156 13900 22196
rect 13940 22156 14860 22196
rect 14900 22156 18548 22196
rect 3331 22112 3389 22113
rect 5740 22112 5780 22156
rect 7564 22112 7604 22156
rect 8227 22112 8285 22113
rect 2659 22072 2668 22112
rect 2708 22072 2860 22112
rect 2900 22072 2909 22112
rect 3331 22072 3340 22112
rect 3380 22072 5780 22112
rect 5827 22072 5836 22112
rect 5876 22072 7564 22112
rect 7604 22072 7613 22112
rect 8142 22072 8236 22112
rect 8276 22072 8285 22112
rect 3331 22071 3389 22072
rect 8227 22071 8285 22072
rect 8419 22112 8477 22113
rect 8611 22112 8669 22113
rect 10060 22112 10100 22156
rect 13891 22155 13949 22156
rect 12259 22112 12317 22113
rect 8419 22072 8428 22112
rect 8468 22072 8562 22112
rect 8611 22072 8620 22112
rect 8660 22072 8716 22112
rect 8756 22072 8765 22112
rect 10060 22072 12268 22112
rect 12308 22072 12317 22112
rect 17347 22072 17356 22112
rect 17396 22072 18316 22112
rect 18356 22072 18365 22112
rect 18979 22072 18988 22112
rect 19028 22072 20236 22112
rect 20276 22072 20285 22112
rect 8419 22071 8477 22072
rect 8611 22071 8669 22072
rect 12259 22071 12317 22072
rect 8428 22028 8468 22071
rect 11779 22028 11837 22029
rect 16483 22028 16541 22029
rect 2083 21988 2092 22028
rect 2132 21988 6604 22028
rect 6644 21988 6653 22028
rect 8428 21988 9772 22028
rect 9812 21988 9821 22028
rect 10243 21988 10252 22028
rect 10292 21988 10732 22028
rect 10772 21988 10781 22028
rect 11694 21988 11788 22028
rect 11828 21988 13612 22028
rect 13652 21988 13661 22028
rect 16483 21988 16492 22028
rect 16532 21988 17836 22028
rect 17876 21988 17885 22028
rect 11779 21987 11837 21988
rect 16483 21987 16541 21988
rect 0 21944 80 21964
rect 3427 21944 3485 21945
rect 6115 21944 6173 21945
rect 21424 21944 21504 21964
rect 0 21904 2572 21944
rect 2612 21904 2621 21944
rect 3342 21904 3436 21944
rect 3476 21904 3485 21944
rect 4919 21904 4928 21944
rect 4968 21904 5010 21944
rect 5050 21904 5092 21944
rect 5132 21904 5174 21944
rect 5214 21904 5256 21944
rect 5296 21904 5305 21944
rect 6030 21904 6124 21944
rect 6164 21904 6173 21944
rect 9187 21904 9196 21944
rect 9236 21904 9580 21944
rect 9620 21904 9629 21944
rect 10339 21904 10348 21944
rect 10388 21904 10636 21944
rect 10676 21904 10685 21944
rect 11320 21904 11500 21944
rect 11540 21904 11549 21944
rect 16003 21904 16012 21944
rect 16052 21904 16204 21944
rect 16244 21904 16253 21944
rect 16675 21904 16684 21944
rect 16724 21904 16733 21944
rect 20039 21904 20048 21944
rect 20088 21904 20130 21944
rect 20170 21904 20212 21944
rect 20252 21904 20294 21944
rect 20334 21904 20376 21944
rect 20416 21904 20425 21944
rect 20803 21904 20812 21944
rect 20852 21904 21504 21944
rect 0 21884 80 21904
rect 3427 21903 3485 21904
rect 6115 21903 6173 21904
rect 11320 21860 11360 21904
rect 3331 21820 3340 21860
rect 3380 21820 3724 21860
rect 3764 21820 3773 21860
rect 4291 21820 4300 21860
rect 4340 21820 11020 21860
rect 11060 21820 11360 21860
rect 4099 21776 4157 21777
rect 3907 21736 3916 21776
rect 3956 21736 4108 21776
rect 4148 21736 4396 21776
rect 4436 21736 4445 21776
rect 6019 21736 6028 21776
rect 6068 21736 6508 21776
rect 6548 21736 6557 21776
rect 6883 21736 6892 21776
rect 6932 21736 11116 21776
rect 11156 21736 11165 21776
rect 4099 21735 4157 21736
rect 16684 21692 16724 21904
rect 21424 21884 21504 21904
rect 16867 21776 16925 21777
rect 18115 21776 18173 21777
rect 16867 21736 16876 21776
rect 16916 21736 17548 21776
rect 17588 21736 18124 21776
rect 18164 21736 18173 21776
rect 19843 21736 19852 21776
rect 19892 21736 20140 21776
rect 20180 21736 20189 21776
rect 16867 21735 16925 21736
rect 18115 21735 18173 21736
rect 1411 21652 1420 21692
rect 1460 21652 13996 21692
rect 14036 21652 14045 21692
rect 16684 21652 20044 21692
rect 20084 21652 20093 21692
rect 0 21608 80 21628
rect 259 21608 317 21609
rect 1795 21608 1853 21609
rect 2179 21608 2237 21609
rect 4483 21608 4541 21609
rect 4675 21608 4733 21609
rect 7363 21608 7421 21609
rect 16867 21608 16925 21609
rect 0 21568 268 21608
rect 308 21568 317 21608
rect 1603 21568 1612 21608
rect 1652 21568 1804 21608
rect 1844 21568 2188 21608
rect 2228 21568 2237 21608
rect 2659 21568 2668 21608
rect 2708 21568 3052 21608
rect 3092 21568 4204 21608
rect 4244 21568 4253 21608
rect 4483 21568 4492 21608
rect 4532 21568 4588 21608
rect 4628 21568 4684 21608
rect 4724 21568 4752 21608
rect 6115 21568 6124 21608
rect 6164 21568 6316 21608
rect 6356 21568 6365 21608
rect 6787 21568 6796 21608
rect 6836 21568 7084 21608
rect 7124 21568 7133 21608
rect 7278 21568 7372 21608
rect 7412 21568 8812 21608
rect 8852 21568 8861 21608
rect 9475 21568 9484 21608
rect 9524 21568 10484 21608
rect 10531 21568 10540 21608
rect 10580 21568 11308 21608
rect 11348 21568 11357 21608
rect 12835 21568 12844 21608
rect 12884 21568 13132 21608
rect 13172 21568 13181 21608
rect 16579 21568 16588 21608
rect 16628 21568 16876 21608
rect 16916 21568 16925 21608
rect 17443 21568 17452 21608
rect 17492 21568 18412 21608
rect 18452 21568 18461 21608
rect 18883 21568 18892 21608
rect 18932 21568 19564 21608
rect 19604 21568 19613 21608
rect 0 21548 80 21568
rect 259 21567 317 21568
rect 1795 21567 1853 21568
rect 2179 21567 2237 21568
rect 4483 21567 4541 21568
rect 4675 21567 4733 21568
rect 7363 21567 7421 21568
rect 3427 21524 3485 21525
rect 3907 21524 3965 21525
rect 6403 21524 6461 21525
rect 8707 21524 8765 21525
rect 10444 21524 10484 21568
rect 16867 21567 16925 21568
rect 11299 21524 11357 21525
rect 2275 21484 2284 21524
rect 2324 21484 2476 21524
rect 2516 21484 2860 21524
rect 2900 21484 2909 21524
rect 3331 21484 3340 21524
rect 3380 21484 3436 21524
rect 3476 21484 3485 21524
rect 3822 21484 3916 21524
rect 3956 21484 6412 21524
rect 6452 21484 6461 21524
rect 8035 21484 8044 21524
rect 8084 21484 8716 21524
rect 8756 21484 8765 21524
rect 8899 21484 8908 21524
rect 8948 21484 10060 21524
rect 10100 21484 10109 21524
rect 10444 21484 11308 21524
rect 11348 21484 11357 21524
rect 12067 21484 12076 21524
rect 12116 21484 12364 21524
rect 12404 21484 15148 21524
rect 15188 21484 15197 21524
rect 16867 21484 16876 21524
rect 16916 21484 19316 21524
rect 3427 21483 3485 21484
rect 3907 21483 3965 21484
rect 6403 21483 6461 21484
rect 8707 21483 8765 21484
rect 11299 21483 11357 21484
rect 3331 21440 3389 21441
rect 6307 21440 6365 21441
rect 3139 21400 3148 21440
rect 3188 21400 3340 21440
rect 3380 21400 3389 21440
rect 3811 21400 3820 21440
rect 3860 21400 4396 21440
rect 4436 21400 4445 21440
rect 5347 21400 5356 21440
rect 5396 21400 6316 21440
rect 6356 21400 6365 21440
rect 3331 21399 3389 21400
rect 6307 21399 6365 21400
rect 7363 21440 7421 21441
rect 8515 21440 8573 21441
rect 7363 21400 7372 21440
rect 7412 21400 8524 21440
rect 8564 21400 8573 21440
rect 7363 21399 7421 21400
rect 8515 21399 8573 21400
rect 9283 21440 9341 21441
rect 11875 21440 11933 21441
rect 12259 21440 12317 21441
rect 19276 21440 19316 21484
rect 21424 21440 21504 21460
rect 9283 21400 9292 21440
rect 9332 21400 9868 21440
rect 9908 21400 9917 21440
rect 11779 21400 11788 21440
rect 11828 21400 11884 21440
rect 11924 21400 11933 21440
rect 12174 21400 12268 21440
rect 12308 21400 12317 21440
rect 16771 21400 16780 21440
rect 16820 21400 17972 21440
rect 18019 21400 18028 21440
rect 18068 21400 18220 21440
rect 18260 21400 18269 21440
rect 19267 21400 19276 21440
rect 19316 21400 19325 21440
rect 19459 21400 19468 21440
rect 19508 21400 21504 21440
rect 9283 21399 9341 21400
rect 11875 21399 11933 21400
rect 12259 21399 12317 21400
rect 2083 21356 2141 21357
rect 7747 21356 7805 21357
rect 8803 21356 8861 21357
rect 163 21316 172 21356
rect 212 21316 1228 21356
rect 1268 21316 1277 21356
rect 2083 21316 2092 21356
rect 2132 21316 6892 21356
rect 6932 21316 6941 21356
rect 7747 21316 7756 21356
rect 7796 21316 8812 21356
rect 8852 21316 8861 21356
rect 2083 21315 2141 21316
rect 7747 21315 7805 21316
rect 8803 21315 8861 21316
rect 17731 21356 17789 21357
rect 17731 21316 17740 21356
rect 17780 21316 17836 21356
rect 17876 21316 17885 21356
rect 17731 21315 17789 21316
rect 0 21272 80 21292
rect 1987 21272 2045 21273
rect 9283 21272 9341 21273
rect 0 21232 1268 21272
rect 0 21212 80 21232
rect 1228 21188 1268 21232
rect 1987 21232 1996 21272
rect 2036 21232 9292 21272
rect 9332 21232 9341 21272
rect 1987 21231 2045 21232
rect 9283 21231 9341 21232
rect 10339 21272 10397 21273
rect 10339 21232 10348 21272
rect 10388 21232 10444 21272
rect 10484 21232 10493 21272
rect 11971 21232 11980 21272
rect 12020 21232 12460 21272
rect 12500 21232 12509 21272
rect 15811 21232 15820 21272
rect 15860 21232 17260 21272
rect 17300 21232 17309 21272
rect 10339 21231 10397 21232
rect 2755 21188 2813 21189
rect 6883 21188 6941 21189
rect 1228 21148 2572 21188
rect 2612 21148 2764 21188
rect 2804 21148 2813 21188
rect 3679 21148 3688 21188
rect 3728 21148 3770 21188
rect 3810 21148 3852 21188
rect 3892 21148 3934 21188
rect 3974 21148 4016 21188
rect 4056 21148 4065 21188
rect 4108 21148 6892 21188
rect 6932 21148 10252 21188
rect 10292 21148 10301 21188
rect 12643 21148 12652 21188
rect 12692 21148 17740 21188
rect 17780 21148 17789 21188
rect 2755 21147 2813 21148
rect 4108 21104 4148 21148
rect 6883 21147 6941 21148
rect 13891 21104 13949 21105
rect 16483 21104 16541 21105
rect 17932 21104 17972 21400
rect 21424 21380 21504 21400
rect 18799 21148 18808 21188
rect 18848 21148 18890 21188
rect 18930 21148 18972 21188
rect 19012 21148 19054 21188
rect 19094 21148 19136 21188
rect 19176 21148 19185 21188
rect 172 21064 4148 21104
rect 4867 21064 4876 21104
rect 4916 21064 13900 21104
rect 13940 21064 13949 21104
rect 14659 21064 14668 21104
rect 14708 21064 14717 21104
rect 16483 21064 16492 21104
rect 16532 21064 17164 21104
rect 17204 21064 17213 21104
rect 17923 21064 17932 21104
rect 17972 21064 17981 21104
rect 0 20936 80 20956
rect 172 20936 212 21064
rect 13891 21063 13949 21064
rect 14668 21020 14708 21064
rect 16483 21063 16541 21064
rect 2947 20980 2956 21020
rect 2996 20980 3005 21020
rect 4108 20980 6836 21020
rect 6883 20980 6892 21020
rect 6932 20980 12652 21020
rect 12692 20980 12701 21020
rect 14668 20980 14860 21020
rect 14900 20980 14909 21020
rect 17059 20980 17068 21020
rect 17108 20980 17260 21020
rect 17300 20980 17548 21020
rect 17588 20980 17597 21020
rect 2851 20936 2909 20937
rect 0 20896 212 20936
rect 2766 20896 2860 20936
rect 2900 20896 2909 20936
rect 2956 20936 2996 20980
rect 2956 20896 4012 20936
rect 4052 20896 4061 20936
rect 0 20876 80 20896
rect 2851 20895 2909 20896
rect 3235 20812 3244 20852
rect 3284 20812 3532 20852
rect 3572 20812 3581 20852
rect 1987 20768 2045 20769
rect 4108 20768 4148 20980
rect 6499 20936 6557 20937
rect 4387 20896 4396 20936
rect 4436 20896 4445 20936
rect 6403 20896 6412 20936
rect 6452 20896 6508 20936
rect 6548 20896 6557 20936
rect 6796 20936 6836 20980
rect 7075 20936 7133 20937
rect 21424 20936 21504 20956
rect 6796 20896 7084 20936
rect 7124 20896 9100 20936
rect 9140 20896 9149 20936
rect 9196 20896 9524 20936
rect 10147 20896 10156 20936
rect 10196 20896 21504 20936
rect 4396 20768 4436 20896
rect 6499 20895 6557 20896
rect 7075 20895 7133 20896
rect 6211 20852 6269 20853
rect 9196 20852 9236 20896
rect 9379 20852 9437 20853
rect 6211 20812 6220 20852
rect 6260 20812 9236 20852
rect 9294 20812 9388 20852
rect 9428 20812 9437 20852
rect 9484 20852 9524 20896
rect 21424 20876 21504 20896
rect 9484 20812 18508 20852
rect 18548 20812 18557 20852
rect 6211 20811 6269 20812
rect 9379 20811 9437 20812
rect 4675 20768 4733 20769
rect 6307 20768 6365 20769
rect 7267 20768 7325 20769
rect 10531 20768 10589 20769
rect 10819 20768 10877 20769
rect 11203 20768 11261 20769
rect 18403 20768 18461 20769
rect 19363 20768 19421 20769
rect 1315 20728 1324 20768
rect 1364 20728 1996 20768
rect 2036 20728 2045 20768
rect 1987 20727 2045 20728
rect 2500 20728 4148 20768
rect 4195 20728 4204 20768
rect 4244 20728 4436 20768
rect 4590 20728 4684 20768
rect 4724 20728 4733 20768
rect 5347 20728 5356 20768
rect 5396 20728 5836 20768
rect 5876 20728 5885 20768
rect 6222 20728 6316 20768
rect 6356 20728 7276 20768
rect 7316 20728 7325 20768
rect 8995 20728 9004 20768
rect 9044 20728 10540 20768
rect 10580 20728 10636 20768
rect 10676 20728 10685 20768
rect 10819 20728 10828 20768
rect 10868 20728 11212 20768
rect 11252 20728 13420 20768
rect 13460 20728 16492 20768
rect 16532 20728 16541 20768
rect 17635 20728 17644 20768
rect 17684 20728 18028 20768
rect 18068 20728 18077 20768
rect 18307 20728 18316 20768
rect 18356 20728 18412 20768
rect 18452 20728 18461 20768
rect 18883 20728 18892 20768
rect 18932 20728 19372 20768
rect 19412 20728 19564 20768
rect 19604 20728 19613 20768
rect 2500 20684 2540 20728
rect 4675 20727 4733 20728
rect 6307 20727 6365 20728
rect 7267 20727 7325 20728
rect 10531 20727 10589 20728
rect 10819 20727 10877 20728
rect 11203 20727 11261 20728
rect 18403 20727 18461 20728
rect 19363 20727 19421 20728
rect 15715 20684 15773 20685
rect 1891 20644 1900 20684
rect 1940 20644 2540 20684
rect 2659 20644 2668 20684
rect 2708 20644 4396 20684
rect 4436 20644 4780 20684
rect 4820 20644 4829 20684
rect 9379 20644 9388 20684
rect 9428 20644 10348 20684
rect 10388 20644 11020 20684
rect 11060 20644 11069 20684
rect 14179 20644 14188 20684
rect 14228 20644 14668 20684
rect 14708 20644 14717 20684
rect 15715 20644 15724 20684
rect 15764 20644 18452 20684
rect 15715 20643 15773 20644
rect 0 20600 80 20620
rect 3427 20600 3485 20601
rect 4483 20600 4541 20601
rect 10915 20600 10973 20601
rect 0 20560 2540 20600
rect 0 20540 80 20560
rect 2500 20516 2540 20560
rect 3427 20560 3436 20600
rect 3476 20560 3820 20600
rect 3860 20560 4492 20600
rect 4532 20560 4541 20600
rect 4675 20560 4684 20600
rect 4724 20560 4876 20600
rect 4916 20560 4925 20600
rect 10915 20560 10924 20600
rect 10964 20560 17740 20600
rect 17780 20560 17789 20600
rect 3427 20559 3485 20560
rect 4483 20559 4541 20560
rect 10915 20559 10973 20560
rect 18412 20516 18452 20644
rect 18691 20600 18749 20601
rect 19651 20600 19709 20601
rect 18691 20560 18700 20600
rect 18740 20560 18988 20600
rect 19028 20560 19037 20600
rect 19651 20560 19660 20600
rect 19700 20560 20140 20600
rect 20180 20560 20189 20600
rect 18691 20559 18749 20560
rect 19651 20559 19709 20560
rect 2500 20476 11404 20516
rect 11444 20476 11453 20516
rect 14467 20476 14476 20516
rect 14516 20476 18220 20516
rect 18260 20476 18269 20516
rect 18412 20476 20852 20516
rect 2659 20432 2717 20433
rect 4099 20432 4157 20433
rect 5443 20432 5501 20433
rect 20812 20432 20852 20476
rect 21424 20432 21504 20452
rect 2563 20392 2572 20432
rect 2612 20392 2668 20432
rect 2708 20392 2717 20432
rect 3043 20392 3052 20432
rect 3092 20392 3340 20432
rect 3380 20392 3389 20432
rect 4014 20392 4108 20432
rect 4148 20392 4406 20432
rect 4446 20392 4455 20432
rect 4919 20392 4928 20432
rect 4968 20392 5010 20432
rect 5050 20392 5092 20432
rect 5132 20392 5174 20432
rect 5214 20392 5256 20432
rect 5296 20392 5305 20432
rect 5443 20392 5452 20432
rect 5492 20392 5836 20432
rect 5876 20392 5885 20432
rect 11320 20392 18028 20432
rect 18068 20392 18077 20432
rect 20039 20392 20048 20432
rect 20088 20392 20130 20432
rect 20170 20392 20212 20432
rect 20252 20392 20294 20432
rect 20334 20392 20376 20432
rect 20416 20392 20425 20432
rect 20812 20392 21504 20432
rect 2659 20391 2717 20392
rect 4099 20391 4157 20392
rect 5443 20391 5501 20392
rect 11320 20348 11360 20392
rect 21424 20372 21504 20392
rect 18019 20348 18077 20349
rect 1507 20308 1516 20348
rect 1556 20308 11360 20348
rect 16387 20308 16396 20348
rect 16436 20308 17356 20348
rect 17396 20308 17405 20348
rect 17635 20308 17644 20348
rect 17684 20308 18028 20348
rect 18068 20308 18077 20348
rect 18019 20307 18077 20308
rect 0 20264 80 20284
rect 0 20224 2900 20264
rect 2947 20224 2956 20264
rect 2996 20224 3436 20264
rect 3476 20224 3628 20264
rect 3668 20224 3677 20264
rect 5539 20224 5548 20264
rect 5588 20224 5972 20264
rect 10339 20224 10348 20264
rect 10388 20224 14476 20264
rect 14516 20224 14525 20264
rect 19747 20224 19756 20264
rect 19796 20224 19805 20264
rect 0 20204 80 20224
rect 2860 20180 2900 20224
rect 2947 20180 3005 20181
rect 2860 20140 2956 20180
rect 2996 20140 3005 20180
rect 2947 20139 3005 20140
rect 2467 20096 2525 20097
rect 4291 20096 4349 20097
rect 5932 20096 5972 20224
rect 11299 20180 11357 20181
rect 11203 20140 11212 20180
rect 11252 20140 11308 20180
rect 11348 20140 11357 20180
rect 16483 20140 16492 20180
rect 16532 20140 17660 20180
rect 18115 20140 18124 20180
rect 18164 20140 18412 20180
rect 18452 20140 18461 20180
rect 11299 20139 11357 20140
rect 6499 20096 6557 20097
rect 8995 20096 9053 20097
rect 10435 20096 10493 20097
rect 17620 20096 17660 20140
rect 2382 20056 2476 20096
rect 2516 20056 2525 20096
rect 2947 20056 2956 20096
rect 2996 20056 3532 20096
rect 3572 20056 3581 20096
rect 4291 20056 4300 20096
rect 4340 20056 5876 20096
rect 5932 20056 6508 20096
rect 6548 20056 6557 20096
rect 8035 20056 8044 20096
rect 8084 20056 9004 20096
rect 9044 20056 9053 20096
rect 10147 20056 10156 20096
rect 10196 20056 10348 20096
rect 10388 20056 10444 20096
rect 10484 20056 10512 20096
rect 12355 20056 12364 20096
rect 12404 20056 12652 20096
rect 12692 20056 12701 20096
rect 13507 20056 13516 20096
rect 13556 20056 14380 20096
rect 14420 20056 14429 20096
rect 17620 20056 19028 20096
rect 19075 20056 19084 20096
rect 19124 20056 19276 20096
rect 19316 20056 19325 20096
rect 2467 20055 2525 20056
rect 4291 20055 4349 20056
rect 2179 20012 2237 20013
rect 5836 20012 5876 20056
rect 6499 20055 6557 20056
rect 8995 20055 9053 20056
rect 10435 20055 10493 20056
rect 9667 20012 9725 20013
rect 13795 20012 13853 20013
rect 14851 20012 14909 20013
rect 15811 20012 15869 20013
rect 18988 20012 19028 20056
rect 19756 20012 19796 20224
rect 2179 19972 2188 20012
rect 2228 19972 4396 20012
rect 4436 19972 4445 20012
rect 5836 19972 7372 20012
rect 7412 19972 7421 20012
rect 9667 19972 9676 20012
rect 9716 19972 9868 20012
rect 9908 19972 9917 20012
rect 12739 19972 12748 20012
rect 12788 19972 13804 20012
rect 13844 19972 13853 20012
rect 14755 19972 14764 20012
rect 14804 19972 14860 20012
rect 14900 19972 14909 20012
rect 15427 19972 15436 20012
rect 15476 19972 15820 20012
rect 15860 19972 16492 20012
rect 16532 19972 16972 20012
rect 17012 19972 18892 20012
rect 18932 19972 18941 20012
rect 18988 19972 19796 20012
rect 2179 19971 2237 19972
rect 9667 19971 9725 19972
rect 13795 19971 13853 19972
rect 14851 19971 14909 19972
rect 15811 19971 15869 19972
rect 0 19928 80 19948
rect 16579 19928 16637 19929
rect 21424 19928 21504 19948
rect 0 19888 3860 19928
rect 3907 19888 3916 19928
rect 3956 19888 4108 19928
rect 4148 19888 4157 19928
rect 5731 19888 5740 19928
rect 5780 19888 6892 19928
rect 6932 19888 6941 19928
rect 12835 19888 12844 19928
rect 12884 19888 16588 19928
rect 16628 19888 16637 19928
rect 18979 19888 18988 19928
rect 19028 19888 21504 19928
rect 0 19868 80 19888
rect 2755 19844 2813 19845
rect 2275 19804 2284 19844
rect 2324 19804 2764 19844
rect 2804 19804 2813 19844
rect 2755 19803 2813 19804
rect 3523 19844 3581 19845
rect 3523 19804 3532 19844
rect 3572 19804 3628 19844
rect 3668 19804 3677 19844
rect 3523 19803 3581 19804
rect 3820 19760 3860 19888
rect 16579 19887 16637 19888
rect 21424 19868 21504 19888
rect 4195 19844 4253 19845
rect 13987 19844 14045 19845
rect 17155 19844 17213 19845
rect 4110 19804 4204 19844
rect 4244 19804 4253 19844
rect 6019 19804 6028 19844
rect 6068 19804 7084 19844
rect 7124 19804 7133 19844
rect 13891 19804 13900 19844
rect 13940 19804 13996 19844
rect 14036 19804 14045 19844
rect 14179 19804 14188 19844
rect 14228 19804 14860 19844
rect 14900 19804 14909 19844
rect 15235 19804 15244 19844
rect 15284 19804 15916 19844
rect 15956 19804 15965 19844
rect 17155 19804 17164 19844
rect 17204 19804 17260 19844
rect 17300 19804 17309 19844
rect 18307 19804 18316 19844
rect 18356 19804 19084 19844
rect 19124 19804 19852 19844
rect 19892 19804 19901 19844
rect 4195 19803 4253 19804
rect 13987 19803 14045 19804
rect 17155 19803 17213 19804
rect 1315 19720 1324 19760
rect 1364 19720 3436 19760
rect 3476 19720 3485 19760
rect 3820 19720 6412 19760
rect 6452 19720 6461 19760
rect 7651 19720 7660 19760
rect 7700 19720 21388 19760
rect 21428 19720 21437 19760
rect 17635 19676 17693 19677
rect 19363 19676 19421 19677
rect 19651 19676 19709 19677
rect 2275 19636 2284 19676
rect 2324 19636 3148 19676
rect 3188 19636 3197 19676
rect 3679 19636 3688 19676
rect 3728 19636 3770 19676
rect 3810 19636 3852 19676
rect 3892 19636 3934 19676
rect 3974 19636 4016 19676
rect 4056 19636 4065 19676
rect 12067 19636 12076 19676
rect 12116 19636 16780 19676
rect 16820 19636 16829 19676
rect 17635 19636 17644 19676
rect 17684 19636 17778 19676
rect 18799 19636 18808 19676
rect 18848 19636 18890 19676
rect 18930 19636 18972 19676
rect 19012 19636 19054 19676
rect 19094 19636 19136 19676
rect 19176 19636 19185 19676
rect 19363 19636 19372 19676
rect 19412 19636 19468 19676
rect 19508 19636 19517 19676
rect 19651 19636 19660 19676
rect 19700 19636 19794 19676
rect 17635 19635 17693 19636
rect 19363 19635 19421 19636
rect 19651 19635 19709 19636
rect 0 19592 80 19612
rect 10915 19592 10973 19593
rect 16771 19592 16829 19593
rect 0 19552 10924 19592
rect 10964 19552 10973 19592
rect 12835 19552 12844 19592
rect 12884 19552 14380 19592
rect 14420 19552 16780 19592
rect 16820 19552 16829 19592
rect 17347 19552 17356 19592
rect 17396 19552 21332 19592
rect 0 19532 80 19552
rect 10915 19551 10973 19552
rect 16771 19551 16829 19552
rect 2659 19508 2717 19509
rect 2574 19468 2668 19508
rect 2708 19468 2717 19508
rect 2947 19468 2956 19508
rect 2996 19468 4012 19508
rect 4052 19468 4492 19508
rect 4532 19468 4541 19508
rect 5251 19468 5260 19508
rect 5300 19468 6316 19508
rect 6356 19468 6365 19508
rect 13219 19468 13228 19508
rect 13268 19468 13900 19508
rect 13940 19468 17740 19508
rect 17780 19468 17789 19508
rect 2659 19467 2717 19468
rect 2755 19424 2813 19425
rect 14371 19424 14429 19425
rect 17251 19424 17309 19425
rect 21292 19424 21332 19552
rect 21424 19424 21504 19444
rect 2670 19384 2764 19424
rect 2804 19384 2813 19424
rect 3427 19384 3436 19424
rect 3476 19384 3485 19424
rect 3619 19384 3628 19424
rect 3668 19384 7852 19424
rect 7892 19384 7901 19424
rect 11587 19384 11596 19424
rect 11636 19384 11884 19424
rect 11924 19384 11933 19424
rect 14286 19384 14380 19424
rect 14420 19384 14429 19424
rect 16675 19384 16684 19424
rect 16724 19384 16733 19424
rect 17251 19384 17260 19424
rect 17300 19384 19852 19424
rect 19892 19384 19901 19424
rect 20131 19384 20140 19424
rect 20180 19384 20189 19424
rect 21292 19384 21504 19424
rect 2755 19383 2813 19384
rect 3436 19340 3476 19384
rect 14371 19383 14429 19384
rect 6019 19340 6077 19341
rect 6211 19340 6269 19341
rect 3436 19300 6028 19340
rect 6068 19300 6220 19340
rect 6260 19300 6269 19340
rect 6019 19299 6077 19300
rect 6211 19299 6269 19300
rect 9475 19340 9533 19341
rect 10627 19340 10685 19341
rect 16003 19340 16061 19341
rect 9475 19300 9484 19340
rect 9524 19300 10636 19340
rect 10676 19300 10828 19340
rect 10868 19300 10877 19340
rect 13411 19300 13420 19340
rect 13460 19300 16012 19340
rect 16052 19300 16061 19340
rect 16684 19340 16724 19384
rect 17251 19383 17309 19384
rect 20140 19340 20180 19384
rect 21424 19364 21504 19384
rect 16684 19300 17644 19340
rect 17684 19300 17693 19340
rect 19555 19300 19564 19340
rect 19604 19300 20180 19340
rect 9475 19299 9533 19300
rect 10627 19299 10685 19300
rect 16003 19299 16061 19300
rect 0 19256 80 19276
rect 2083 19256 2141 19257
rect 4099 19256 4157 19257
rect 4771 19256 4829 19257
rect 6499 19256 6557 19257
rect 9667 19256 9725 19257
rect 17155 19256 17213 19257
rect 0 19216 2092 19256
rect 2132 19216 2141 19256
rect 2467 19216 2476 19256
rect 2516 19216 2956 19256
rect 2996 19216 3005 19256
rect 3052 19216 3436 19256
rect 3476 19216 3485 19256
rect 3811 19216 3820 19256
rect 3860 19216 4108 19256
rect 4148 19216 4780 19256
rect 4820 19216 4829 19256
rect 5731 19216 5740 19256
rect 5780 19216 6028 19256
rect 6068 19216 6077 19256
rect 6499 19216 6508 19256
rect 6548 19216 6604 19256
rect 6644 19216 6653 19256
rect 8323 19216 8332 19256
rect 8372 19216 9100 19256
rect 9140 19216 9149 19256
rect 9582 19216 9676 19256
rect 9716 19216 9725 19256
rect 0 19196 80 19216
rect 2083 19215 2141 19216
rect 1699 19172 1757 19173
rect 3052 19172 3092 19216
rect 4099 19215 4157 19216
rect 4771 19215 4829 19216
rect 6499 19215 6557 19216
rect 9667 19215 9725 19216
rect 11320 19216 15244 19256
rect 15284 19216 15293 19256
rect 15715 19216 15724 19256
rect 15764 19216 17164 19256
rect 17204 19216 17260 19256
rect 17300 19216 17309 19256
rect 18115 19216 18124 19256
rect 18164 19216 20044 19256
rect 20084 19216 20093 19256
rect 8323 19172 8381 19173
rect 1614 19132 1708 19172
rect 1748 19132 1757 19172
rect 2851 19132 2860 19172
rect 2900 19132 3092 19172
rect 3139 19132 3148 19172
rect 3188 19132 6220 19172
rect 6260 19132 7564 19172
rect 7604 19132 7613 19172
rect 8304 19132 8332 19172
rect 8372 19132 8428 19172
rect 8468 19132 9196 19172
rect 9236 19132 9388 19172
rect 9428 19132 9437 19172
rect 1699 19131 1757 19132
rect 8323 19131 8381 19132
rect 4291 19088 4349 19089
rect 10819 19088 10877 19089
rect 3331 19048 3340 19088
rect 3380 19048 4300 19088
rect 4340 19048 4396 19088
rect 4436 19048 4445 19088
rect 7267 19048 7276 19088
rect 7316 19048 10828 19088
rect 10868 19048 10877 19088
rect 4291 19047 4349 19048
rect 10819 19047 10877 19048
rect 9283 19004 9341 19005
rect 11320 19004 11360 19216
rect 17155 19215 17213 19216
rect 13795 19172 13853 19173
rect 13027 19132 13036 19172
rect 13076 19132 13324 19172
rect 13364 19132 13373 19172
rect 13710 19132 13804 19172
rect 13844 19132 13853 19172
rect 13795 19131 13853 19132
rect 14371 19172 14429 19173
rect 20803 19172 20861 19173
rect 14371 19132 14380 19172
rect 14420 19132 20812 19172
rect 20852 19132 20861 19172
rect 14371 19131 14429 19132
rect 20803 19131 20861 19132
rect 14083 19088 14141 19089
rect 17155 19088 17213 19089
rect 14083 19048 14092 19088
rect 14132 19048 14860 19088
rect 14900 19048 14909 19088
rect 15043 19048 15052 19088
rect 15092 19048 17164 19088
rect 17204 19048 17213 19088
rect 14083 19047 14141 19048
rect 17155 19047 17213 19048
rect 5635 18964 5644 19004
rect 5684 18964 8620 19004
rect 8660 18964 8669 19004
rect 9091 18964 9100 19004
rect 9140 18964 9292 19004
rect 9332 18964 11360 19004
rect 13795 19004 13853 19005
rect 16867 19004 16925 19005
rect 13795 18964 13804 19004
rect 13844 18964 13900 19004
rect 13940 18964 13949 19004
rect 15052 18964 16876 19004
rect 16916 18964 16925 19004
rect 9283 18963 9341 18964
rect 13795 18963 13853 18964
rect 0 18920 80 18940
rect 6019 18920 6077 18921
rect 10915 18920 10973 18921
rect 15052 18920 15092 18964
rect 16867 18963 16925 18964
rect 17635 18920 17693 18921
rect 21424 18920 21504 18940
rect 0 18880 2092 18920
rect 2132 18880 2141 18920
rect 4919 18880 4928 18920
rect 4968 18880 5010 18920
rect 5050 18880 5092 18920
rect 5132 18880 5174 18920
rect 5214 18880 5256 18920
rect 5296 18880 5305 18920
rect 6019 18880 6028 18920
rect 6068 18880 6700 18920
rect 6740 18880 6749 18920
rect 6796 18880 10924 18920
rect 10964 18880 10973 18920
rect 11395 18880 11404 18920
rect 11444 18880 14900 18920
rect 14947 18880 14956 18920
rect 14996 18880 15092 18920
rect 15139 18880 15148 18920
rect 15188 18880 15628 18920
rect 15668 18880 17068 18920
rect 17108 18880 17117 18920
rect 17164 18880 17644 18920
rect 17684 18880 17693 18920
rect 17923 18880 17932 18920
rect 17972 18880 17981 18920
rect 18403 18880 18412 18920
rect 18452 18880 19988 18920
rect 20039 18880 20048 18920
rect 20088 18880 20130 18920
rect 20170 18880 20212 18920
rect 20252 18880 20294 18920
rect 20334 18880 20376 18920
rect 20416 18880 20425 18920
rect 21379 18880 21388 18920
rect 21428 18880 21504 18920
rect 0 18860 80 18880
rect 6019 18879 6077 18880
rect 5443 18836 5501 18837
rect 6796 18836 6836 18880
rect 10915 18879 10973 18880
rect 14860 18836 14900 18880
rect 4195 18796 4204 18836
rect 4244 18796 5452 18836
rect 5492 18796 6836 18836
rect 6979 18796 6988 18836
rect 7028 18796 11596 18836
rect 11636 18796 11645 18836
rect 13612 18796 14668 18836
rect 14708 18796 14717 18836
rect 14860 18796 16108 18836
rect 16148 18796 16157 18836
rect 5443 18795 5501 18796
rect 5347 18752 5405 18753
rect 13612 18752 13652 18796
rect 17164 18752 17204 18880
rect 17635 18879 17693 18880
rect 17932 18836 17972 18880
rect 19948 18836 19988 18880
rect 21424 18860 21504 18880
rect 17635 18796 17644 18836
rect 17684 18796 17836 18836
rect 17876 18796 17885 18836
rect 17932 18796 19468 18836
rect 19508 18796 19517 18836
rect 19948 18796 20276 18836
rect 17932 18752 17972 18796
rect 20236 18752 20276 18796
rect 3907 18712 3916 18752
rect 3956 18712 5356 18752
rect 5396 18712 5405 18752
rect 6115 18712 6124 18752
rect 6164 18712 6173 18752
rect 7363 18712 7372 18752
rect 7412 18712 9388 18752
rect 9428 18712 9437 18752
rect 10627 18712 10636 18752
rect 10676 18712 13652 18752
rect 13699 18712 13708 18752
rect 13748 18712 14092 18752
rect 14132 18712 14141 18752
rect 16012 18712 17204 18752
rect 17251 18712 17260 18752
rect 17300 18712 17660 18752
rect 17731 18712 17740 18752
rect 17780 18712 17972 18752
rect 19267 18712 19276 18752
rect 19316 18712 20044 18752
rect 20084 18712 20093 18752
rect 20227 18712 20236 18752
rect 20276 18712 20285 18752
rect 5347 18711 5405 18712
rect 6124 18668 6164 18712
rect 10435 18668 10493 18669
rect 16012 18668 16052 18712
rect 931 18628 940 18668
rect 980 18628 2092 18668
rect 2132 18628 3340 18668
rect 3380 18628 3389 18668
rect 5251 18628 5260 18668
rect 5300 18628 6164 18668
rect 6595 18628 6604 18668
rect 6644 18628 6988 18668
rect 7028 18628 7037 18668
rect 10435 18628 10444 18668
rect 10484 18628 16052 18668
rect 16771 18628 16780 18668
rect 16820 18628 17068 18668
rect 17108 18628 17117 18668
rect 10435 18627 10493 18628
rect 0 18584 80 18604
rect 6115 18584 6173 18585
rect 17620 18584 17660 18712
rect 0 18544 2612 18584
rect 2659 18544 2668 18584
rect 2708 18544 3628 18584
rect 3668 18544 3820 18584
rect 3860 18544 3869 18584
rect 5443 18544 5452 18584
rect 5492 18544 5836 18584
rect 5876 18544 5885 18584
rect 6030 18544 6124 18584
rect 6164 18544 6173 18584
rect 7747 18544 7756 18584
rect 7796 18544 11360 18584
rect 12259 18544 12268 18584
rect 12308 18544 12556 18584
rect 12596 18544 13940 18584
rect 13987 18544 13996 18584
rect 14036 18544 14045 18584
rect 17620 18544 17644 18584
rect 17684 18544 17693 18584
rect 0 18524 80 18544
rect 1507 18500 1565 18501
rect 1219 18460 1228 18500
rect 1268 18460 1516 18500
rect 1556 18460 1565 18500
rect 2572 18500 2612 18544
rect 6115 18543 6173 18544
rect 3139 18500 3197 18501
rect 11320 18500 11360 18544
rect 13900 18500 13940 18544
rect 13996 18500 14036 18544
rect 2572 18460 3148 18500
rect 3188 18460 8140 18500
rect 8180 18460 8189 18500
rect 9763 18460 9772 18500
rect 9812 18460 10636 18500
rect 10676 18460 10685 18500
rect 11320 18460 12652 18500
rect 12692 18460 12701 18500
rect 13891 18460 13900 18500
rect 13940 18460 13949 18500
rect 13996 18460 14092 18500
rect 14132 18460 14141 18500
rect 15331 18460 15340 18500
rect 15380 18460 15532 18500
rect 15572 18460 15581 18500
rect 16099 18460 16108 18500
rect 16148 18460 17153 18500
rect 17193 18460 17202 18500
rect 17251 18460 17260 18500
rect 17300 18460 17452 18500
rect 17492 18460 17836 18500
rect 17876 18460 17885 18500
rect 18019 18460 18028 18500
rect 18068 18460 18796 18500
rect 18836 18460 18845 18500
rect 1507 18459 1565 18460
rect 3139 18459 3197 18460
rect 13219 18416 13277 18417
rect 16675 18416 16733 18417
rect 21424 18416 21504 18436
rect 3619 18376 3628 18416
rect 3668 18376 4108 18416
rect 4148 18376 4157 18416
rect 9379 18376 9388 18416
rect 9428 18376 13228 18416
rect 13268 18376 15436 18416
rect 15476 18376 15485 18416
rect 16675 18376 16684 18416
rect 16724 18376 21504 18416
rect 13219 18375 13277 18376
rect 16675 18375 16733 18376
rect 21424 18356 21504 18376
rect 2947 18332 3005 18333
rect 3139 18332 3197 18333
rect 10627 18332 10685 18333
rect 2947 18292 2956 18332
rect 2996 18292 3148 18332
rect 3188 18292 3244 18332
rect 3284 18292 3293 18332
rect 4003 18292 4012 18332
rect 4052 18292 5452 18332
rect 5492 18292 5501 18332
rect 5923 18292 5932 18332
rect 5972 18292 6892 18332
rect 6932 18292 6941 18332
rect 10627 18292 10636 18332
rect 10676 18292 11020 18332
rect 11060 18292 11069 18332
rect 11299 18292 11308 18332
rect 11348 18292 13708 18332
rect 13748 18292 13757 18332
rect 15331 18292 15340 18332
rect 15380 18292 17644 18332
rect 17684 18292 17693 18332
rect 18883 18292 18892 18332
rect 18932 18292 19372 18332
rect 19412 18292 19421 18332
rect 2947 18291 3005 18292
rect 3139 18291 3197 18292
rect 0 18248 80 18268
rect 3244 18248 3284 18292
rect 10627 18291 10685 18292
rect 5731 18248 5789 18249
rect 13795 18248 13853 18249
rect 0 18208 1228 18248
rect 1268 18208 1277 18248
rect 3244 18208 5684 18248
rect 0 18188 80 18208
rect 5644 18164 5684 18208
rect 5731 18208 5740 18248
rect 5780 18208 10924 18248
rect 10964 18208 13420 18248
rect 13460 18208 13469 18248
rect 13795 18208 13804 18248
rect 13844 18208 13900 18248
rect 13940 18208 13949 18248
rect 16195 18208 16204 18248
rect 16244 18208 19276 18248
rect 19316 18208 19325 18248
rect 5731 18207 5789 18208
rect 13795 18207 13853 18208
rect 3679 18124 3688 18164
rect 3728 18124 3770 18164
rect 3810 18124 3852 18164
rect 3892 18124 3934 18164
rect 3974 18124 4016 18164
rect 4056 18124 4065 18164
rect 5644 18124 6316 18164
rect 6356 18124 6365 18164
rect 13603 18124 13612 18164
rect 13652 18124 13804 18164
rect 13844 18124 13853 18164
rect 14179 18124 14188 18164
rect 14228 18124 14380 18164
rect 14420 18124 14429 18164
rect 14755 18124 14764 18164
rect 14804 18124 18644 18164
rect 18799 18124 18808 18164
rect 18848 18124 18890 18164
rect 18930 18124 18972 18164
rect 19012 18124 19054 18164
rect 19094 18124 19136 18164
rect 19176 18124 19185 18164
rect 18604 18080 18644 18124
rect 2500 18040 11308 18080
rect 11348 18040 15244 18080
rect 15284 18040 15293 18080
rect 16771 18040 16780 18080
rect 16820 18040 18028 18080
rect 18068 18040 18077 18080
rect 18604 18040 19660 18080
rect 19700 18040 19709 18080
rect 0 17912 80 17932
rect 2500 17912 2540 18040
rect 3523 17996 3581 17997
rect 8899 17996 8957 17997
rect 14947 17996 15005 17997
rect 3427 17956 3436 17996
rect 3476 17956 3532 17996
rect 3572 17956 6412 17996
rect 6452 17956 8908 17996
rect 8948 17956 8957 17996
rect 13123 17956 13132 17996
rect 13172 17956 14708 17996
rect 3523 17955 3581 17956
rect 8899 17955 8957 17956
rect 14668 17912 14708 17956
rect 14947 17956 14956 17996
rect 14996 17956 15090 17996
rect 16483 17956 16492 17996
rect 16532 17956 16684 17996
rect 16724 17956 16733 17996
rect 14947 17955 15005 17956
rect 16780 17912 16820 18040
rect 18403 17996 18461 17997
rect 19180 17996 19220 18040
rect 17731 17956 17740 17996
rect 17780 17956 18412 17996
rect 18452 17956 18461 17996
rect 19171 17956 19180 17996
rect 19220 17956 19260 17996
rect 19459 17956 19468 17996
rect 19508 17956 20716 17996
rect 20756 17956 20765 17996
rect 18403 17955 18461 17956
rect 0 17872 2540 17912
rect 7747 17872 7756 17912
rect 7796 17872 7805 17912
rect 8035 17872 8044 17912
rect 8084 17872 8332 17912
rect 8372 17872 8381 17912
rect 8803 17872 8812 17912
rect 8852 17872 9292 17912
rect 9332 17872 9341 17912
rect 14371 17872 14380 17912
rect 14420 17872 14572 17912
rect 14612 17872 14621 17912
rect 14668 17872 16820 17912
rect 19459 17912 19517 17913
rect 21424 17912 21504 17932
rect 19459 17872 19468 17912
rect 19508 17872 21504 17912
rect 0 17852 80 17872
rect 7756 17828 7796 17872
rect 19459 17871 19517 17872
rect 21424 17852 21504 17872
rect 13603 17828 13661 17829
rect 15811 17828 15869 17829
rect 17251 17828 17309 17829
rect 1219 17788 1228 17828
rect 1268 17788 2284 17828
rect 2324 17788 2333 17828
rect 2467 17788 2476 17828
rect 2516 17788 7796 17828
rect 13518 17788 13612 17828
rect 13652 17788 13661 17828
rect 14755 17788 14764 17828
rect 14804 17788 15148 17828
rect 15188 17788 15197 17828
rect 15726 17788 15820 17828
rect 15860 17788 15869 17828
rect 17166 17788 17260 17828
rect 17300 17788 17309 17828
rect 13603 17787 13661 17788
rect 15811 17787 15869 17788
rect 17251 17787 17309 17788
rect 1603 17744 1661 17745
rect 4771 17744 4829 17745
rect 1507 17704 1516 17744
rect 1556 17704 1612 17744
rect 1652 17704 1661 17744
rect 1891 17704 1900 17744
rect 1940 17704 2668 17744
rect 2708 17704 3244 17744
rect 3284 17704 3293 17744
rect 4771 17704 4780 17744
rect 4820 17704 5932 17744
rect 5972 17704 6508 17744
rect 6548 17704 6557 17744
rect 7459 17704 7468 17744
rect 7508 17704 8332 17744
rect 8372 17704 8381 17744
rect 9379 17704 9388 17744
rect 9428 17704 10156 17744
rect 10196 17704 10205 17744
rect 12643 17704 12652 17744
rect 12692 17704 12701 17744
rect 13219 17704 13228 17744
rect 13268 17704 13516 17744
rect 13556 17704 13565 17744
rect 13699 17704 13708 17744
rect 13748 17704 18412 17744
rect 18452 17704 18461 17744
rect 1603 17703 1661 17704
rect 4771 17703 4829 17704
rect 163 17660 221 17661
rect 5347 17660 5405 17661
rect 7555 17660 7613 17661
rect 9475 17660 9533 17661
rect 12652 17660 12692 17704
rect 17827 17660 17885 17661
rect 163 17620 172 17660
rect 212 17620 2476 17660
rect 2516 17620 2525 17660
rect 5347 17620 5356 17660
rect 5396 17620 5780 17660
rect 6307 17620 6316 17660
rect 6356 17620 6892 17660
rect 6932 17620 6941 17660
rect 7470 17620 7564 17660
rect 7604 17620 7613 17660
rect 8899 17620 8908 17660
rect 8948 17620 9484 17660
rect 9524 17620 9676 17660
rect 9716 17620 9725 17660
rect 11587 17620 11596 17660
rect 11636 17620 12404 17660
rect 12652 17620 17780 17660
rect 163 17619 221 17620
rect 5347 17619 5405 17620
rect 0 17576 80 17596
rect 0 17536 3532 17576
rect 3572 17536 3581 17576
rect 0 17516 80 17536
rect 5539 17492 5597 17493
rect 5740 17492 5780 17620
rect 7555 17619 7613 17620
rect 9475 17619 9533 17620
rect 12364 17576 12404 17620
rect 17740 17576 17780 17620
rect 17827 17620 17836 17660
rect 17876 17620 18700 17660
rect 18740 17620 18749 17660
rect 17827 17619 17885 17620
rect 8803 17536 8812 17576
rect 8852 17536 9580 17576
rect 9620 17536 9629 17576
rect 12355 17536 12364 17576
rect 12404 17536 12413 17576
rect 12643 17536 12652 17576
rect 12692 17536 14860 17576
rect 14900 17536 14909 17576
rect 17731 17536 17740 17576
rect 17780 17536 17789 17576
rect 4579 17452 4588 17492
rect 4628 17452 5548 17492
rect 5588 17452 5597 17492
rect 5731 17452 5740 17492
rect 5780 17452 5789 17492
rect 5539 17451 5597 17452
rect 9763 17408 9821 17409
rect 21424 17408 21504 17428
rect 4919 17368 4928 17408
rect 4968 17368 5010 17408
rect 5050 17368 5092 17408
rect 5132 17368 5174 17408
rect 5214 17368 5256 17408
rect 5296 17368 5305 17408
rect 9678 17368 9772 17408
rect 9812 17368 9821 17408
rect 16963 17368 16972 17408
rect 17012 17368 17260 17408
rect 17300 17368 17309 17408
rect 20039 17368 20048 17408
rect 20088 17368 20130 17408
rect 20170 17368 20212 17408
rect 20252 17368 20294 17408
rect 20334 17368 20376 17408
rect 20416 17368 20425 17408
rect 21091 17368 21100 17408
rect 21140 17368 21504 17408
rect 9763 17367 9821 17368
rect 21424 17348 21504 17368
rect 1507 17324 1565 17325
rect 1315 17284 1324 17324
rect 1364 17284 1516 17324
rect 1556 17284 1565 17324
rect 2275 17284 2284 17324
rect 2324 17284 9964 17324
rect 10004 17284 10013 17324
rect 17347 17284 17356 17324
rect 17396 17284 17405 17324
rect 1507 17283 1565 17284
rect 0 17240 80 17260
rect 4771 17240 4829 17241
rect 17356 17240 17396 17284
rect 0 17200 4780 17240
rect 4820 17200 4829 17240
rect 5827 17200 5836 17240
rect 5876 17200 7276 17240
rect 7316 17200 7325 17240
rect 7843 17200 7852 17240
rect 7892 17200 8236 17240
rect 8276 17200 8285 17240
rect 9667 17200 9676 17240
rect 9716 17200 10828 17240
rect 10868 17200 10877 17240
rect 17068 17200 17396 17240
rect 0 17180 80 17200
rect 4771 17199 4829 17200
rect 13987 17156 14045 17157
rect 17068 17156 17108 17200
rect 1315 17116 1324 17156
rect 1364 17116 1612 17156
rect 1652 17116 1661 17156
rect 3907 17116 3916 17156
rect 3956 17116 5489 17156
rect 5529 17116 5538 17156
rect 12931 17116 12940 17156
rect 12980 17116 13996 17156
rect 14036 17116 14572 17156
rect 14612 17116 15860 17156
rect 17059 17116 17068 17156
rect 17108 17116 17117 17156
rect 17347 17116 17356 17156
rect 17396 17116 17836 17156
rect 17876 17116 17885 17156
rect 13987 17115 14045 17116
rect 2083 17072 2141 17073
rect 15820 17072 15860 17116
rect 20899 17072 20957 17073
rect 1795 17032 1804 17072
rect 1844 17032 2092 17072
rect 2132 17032 2141 17072
rect 2947 17032 2956 17072
rect 2996 17032 5164 17072
rect 5204 17032 5213 17072
rect 7171 17032 7180 17072
rect 7220 17032 9484 17072
rect 9524 17032 12268 17072
rect 12308 17032 12317 17072
rect 13987 17032 13996 17072
rect 14036 17032 14668 17072
rect 14708 17032 14717 17072
rect 15811 17032 15820 17072
rect 15860 17032 16204 17072
rect 16244 17032 16253 17072
rect 16387 17032 16396 17072
rect 16436 17032 16972 17072
rect 17012 17032 17021 17072
rect 18691 17032 18700 17072
rect 18740 17032 19180 17072
rect 19220 17032 19372 17072
rect 19412 17032 19421 17072
rect 19747 17032 19756 17072
rect 19796 17032 20908 17072
rect 20948 17032 20957 17072
rect 2083 17031 2141 17032
rect 20899 17031 20957 17032
rect 4099 16948 4108 16988
rect 4148 16948 4972 16988
rect 5012 16948 5021 16988
rect 11971 16948 11980 16988
rect 12020 16948 18124 16988
rect 18164 16948 18173 16988
rect 0 16904 80 16924
rect 1219 16904 1277 16905
rect 0 16864 1228 16904
rect 1268 16864 1277 16904
rect 0 16844 80 16864
rect 1219 16863 1277 16864
rect 4195 16904 4253 16905
rect 16291 16904 16349 16905
rect 21424 16904 21504 16924
rect 4195 16864 4204 16904
rect 4244 16864 4684 16904
rect 4724 16864 10060 16904
rect 10100 16864 10109 16904
rect 14755 16864 14764 16904
rect 14804 16864 14956 16904
rect 14996 16864 15005 16904
rect 16291 16864 16300 16904
rect 16340 16864 21504 16904
rect 4195 16863 4253 16864
rect 16291 16863 16349 16864
rect 21424 16844 21504 16864
rect 19747 16820 19805 16821
rect 2755 16780 2764 16820
rect 2804 16780 3244 16820
rect 3284 16780 3293 16820
rect 3619 16780 3628 16820
rect 3668 16780 4108 16820
rect 4148 16780 4157 16820
rect 16291 16780 16300 16820
rect 16340 16780 17260 16820
rect 17300 16780 17309 16820
rect 19662 16780 19756 16820
rect 19796 16780 19805 16820
rect 19747 16779 19805 16780
rect 10339 16736 10397 16737
rect 12547 16736 12605 16737
rect 10339 16696 10348 16736
rect 10388 16696 12556 16736
rect 12596 16696 12605 16736
rect 10339 16695 10397 16696
rect 12547 16695 12605 16696
rect 10627 16652 10685 16653
rect 11683 16652 11741 16653
rect 3679 16612 3688 16652
rect 3728 16612 3770 16652
rect 3810 16612 3852 16652
rect 3892 16612 3934 16652
rect 3974 16612 4016 16652
rect 4056 16612 4065 16652
rect 5731 16612 5740 16652
rect 5780 16612 7084 16652
rect 7124 16612 7133 16652
rect 8227 16612 8236 16652
rect 8276 16612 8524 16652
rect 8564 16612 8573 16652
rect 10627 16612 10636 16652
rect 10676 16612 11116 16652
rect 11156 16612 11165 16652
rect 11598 16612 11692 16652
rect 11732 16612 11741 16652
rect 16771 16612 16780 16652
rect 16820 16612 17356 16652
rect 17396 16612 17405 16652
rect 18799 16612 18808 16652
rect 18848 16612 18890 16652
rect 18930 16612 18972 16652
rect 19012 16612 19054 16652
rect 19094 16612 19136 16652
rect 19176 16612 19185 16652
rect 10627 16611 10685 16612
rect 11683 16611 11741 16612
rect 0 16568 80 16588
rect 16867 16568 16925 16569
rect 0 16528 11404 16568
rect 11444 16528 11788 16568
rect 11828 16528 11837 16568
rect 16867 16528 16876 16568
rect 16916 16528 17010 16568
rect 0 16508 80 16528
rect 16867 16527 16925 16528
rect 1411 16444 1420 16484
rect 1460 16444 1469 16484
rect 2179 16444 2188 16484
rect 2228 16444 17644 16484
rect 17684 16444 17693 16484
rect 19075 16444 19084 16484
rect 19124 16444 19948 16484
rect 19988 16444 19997 16484
rect 1420 16400 1460 16444
rect 8803 16400 8861 16401
rect 21283 16400 21341 16401
rect 21424 16400 21504 16420
rect 1420 16360 3436 16400
rect 3476 16360 3485 16400
rect 3907 16360 3916 16400
rect 3956 16360 4204 16400
rect 4244 16360 4253 16400
rect 5635 16360 5644 16400
rect 5684 16360 7180 16400
rect 7220 16360 7229 16400
rect 7939 16360 7948 16400
rect 7988 16360 8812 16400
rect 8852 16360 8861 16400
rect 9379 16360 9388 16400
rect 9428 16360 9437 16400
rect 10051 16360 10060 16400
rect 10100 16360 10964 16400
rect 12739 16360 12748 16400
rect 12788 16360 13516 16400
rect 13556 16360 14516 16400
rect 14947 16360 14956 16400
rect 14996 16360 15724 16400
rect 15764 16360 15773 16400
rect 16003 16360 16012 16400
rect 16052 16360 16684 16400
rect 16724 16360 16733 16400
rect 16780 16360 19180 16400
rect 19220 16360 19229 16400
rect 21283 16360 21292 16400
rect 21332 16360 21504 16400
rect 3043 16316 3101 16317
rect 3043 16276 3052 16316
rect 3092 16276 3820 16316
rect 3860 16276 3869 16316
rect 5923 16276 5932 16316
rect 5972 16276 6220 16316
rect 6260 16276 6269 16316
rect 3043 16275 3101 16276
rect 0 16232 80 16252
rect 3427 16232 3485 16233
rect 6508 16232 6548 16360
rect 8803 16359 8861 16360
rect 9388 16316 9428 16360
rect 7555 16276 7564 16316
rect 7604 16276 9428 16316
rect 10243 16276 10252 16316
rect 10292 16276 10540 16316
rect 10580 16276 10589 16316
rect 0 16192 2708 16232
rect 0 16172 80 16192
rect 1795 16108 1804 16148
rect 1844 16108 2540 16148
rect 2500 16064 2540 16108
rect 2500 16024 2572 16064
rect 2612 16024 2621 16064
rect 2668 15980 2708 16192
rect 3427 16192 3436 16232
rect 3476 16192 3724 16232
rect 3764 16192 3773 16232
rect 4195 16192 4204 16232
rect 4244 16192 6316 16232
rect 6356 16192 6365 16232
rect 6499 16192 6508 16232
rect 6548 16192 6557 16232
rect 6883 16192 6892 16232
rect 6932 16192 7084 16232
rect 7124 16192 7133 16232
rect 9859 16192 9868 16232
rect 9908 16192 10444 16232
rect 10484 16192 10493 16232
rect 3427 16191 3485 16192
rect 2755 16148 2813 16149
rect 10924 16148 10964 16360
rect 11683 16316 11741 16317
rect 14476 16316 14516 16360
rect 16780 16316 16820 16360
rect 21283 16359 21341 16360
rect 21424 16340 21504 16360
rect 11107 16276 11116 16316
rect 11156 16276 11692 16316
rect 11732 16276 14380 16316
rect 14420 16276 14429 16316
rect 14476 16276 16820 16316
rect 17155 16276 17164 16316
rect 17204 16276 19468 16316
rect 19508 16276 19517 16316
rect 11683 16275 11741 16276
rect 11011 16192 11020 16232
rect 11060 16192 14188 16232
rect 14228 16192 14237 16232
rect 14563 16192 14572 16232
rect 14612 16192 16204 16232
rect 16244 16192 16253 16232
rect 18979 16192 18988 16232
rect 19028 16192 19660 16232
rect 19700 16192 19709 16232
rect 13027 16148 13085 16149
rect 2755 16108 2764 16148
rect 2804 16108 5260 16148
rect 5300 16108 5309 16148
rect 5356 16108 7564 16148
rect 7604 16108 7613 16148
rect 10924 16108 11404 16148
rect 11444 16108 11453 16148
rect 13027 16108 13036 16148
rect 13076 16108 13612 16148
rect 13652 16108 13661 16148
rect 2755 16107 2813 16108
rect 5356 16064 5396 16108
rect 13027 16107 13085 16108
rect 6883 16064 6941 16065
rect 4675 16024 4684 16064
rect 4724 16024 4972 16064
rect 5012 16024 5021 16064
rect 5155 16024 5164 16064
rect 5204 16024 5396 16064
rect 6798 16024 6892 16064
rect 6932 16024 6941 16064
rect 6883 16023 6941 16024
rect 7459 16064 7517 16065
rect 8899 16064 8957 16065
rect 9283 16064 9341 16065
rect 11683 16064 11741 16065
rect 19939 16064 19997 16065
rect 7459 16024 7468 16064
rect 7508 16024 7756 16064
rect 7796 16024 7805 16064
rect 8814 16024 8908 16064
rect 8948 16024 8957 16064
rect 9198 16024 9292 16064
rect 9332 16024 9341 16064
rect 11598 16024 11692 16064
rect 11732 16024 11741 16064
rect 11875 16024 11884 16064
rect 11924 16024 13900 16064
rect 13940 16024 14572 16064
rect 14612 16024 14621 16064
rect 15235 16024 15244 16064
rect 15284 16024 16300 16064
rect 16340 16024 16349 16064
rect 19267 16024 19276 16064
rect 19316 16024 19756 16064
rect 19796 16024 19805 16064
rect 19939 16024 19948 16064
rect 19988 16024 20044 16064
rect 20084 16024 20093 16064
rect 7459 16023 7517 16024
rect 8899 16023 8957 16024
rect 9283 16023 9341 16024
rect 11683 16023 11741 16024
rect 19939 16023 19997 16024
rect 15523 15980 15581 15981
rect 19363 15980 19421 15981
rect 1987 15940 1996 15980
rect 2036 15940 2540 15980
rect 2668 15940 8524 15980
rect 8564 15940 8573 15980
rect 10531 15940 10540 15980
rect 10580 15940 15532 15980
rect 15572 15940 15581 15980
rect 15715 15940 15724 15980
rect 15764 15940 17548 15980
rect 17588 15940 17597 15980
rect 19363 15940 19372 15980
rect 19412 15940 20620 15980
rect 20660 15940 20669 15980
rect 0 15896 80 15916
rect 2500 15896 2540 15940
rect 15523 15939 15581 15940
rect 19363 15939 19421 15940
rect 21424 15897 21504 15916
rect 3139 15896 3197 15897
rect 9187 15896 9245 15897
rect 9763 15896 9821 15897
rect 14563 15896 14621 15897
rect 18691 15896 18749 15897
rect 21379 15896 21504 15897
rect 0 15856 1516 15896
rect 1556 15856 1565 15896
rect 2500 15856 3148 15896
rect 3188 15856 3197 15896
rect 4919 15856 4928 15896
rect 4968 15856 5010 15896
rect 5050 15856 5092 15896
rect 5132 15856 5174 15896
rect 5214 15856 5256 15896
rect 5296 15856 5305 15896
rect 7267 15856 7276 15896
rect 7316 15856 7852 15896
rect 7892 15856 9196 15896
rect 9236 15856 9772 15896
rect 9812 15856 9821 15896
rect 10435 15856 10444 15896
rect 10484 15856 11116 15896
rect 11156 15856 11165 15896
rect 11320 15856 11884 15896
rect 11924 15856 12076 15896
rect 12116 15856 12125 15896
rect 14563 15856 14572 15896
rect 14612 15856 17204 15896
rect 18606 15856 18700 15896
rect 18740 15856 18749 15896
rect 20039 15856 20048 15896
rect 20088 15856 20130 15896
rect 20170 15856 20212 15896
rect 20252 15856 20294 15896
rect 20334 15856 20376 15896
rect 20416 15856 20425 15896
rect 21379 15856 21388 15896
rect 21428 15856 21504 15896
rect 0 15836 80 15856
rect 3139 15855 3197 15856
rect 9187 15855 9245 15856
rect 9763 15855 9821 15856
rect 2659 15812 2717 15813
rect 7075 15812 7133 15813
rect 11320 15812 11360 15856
rect 14563 15855 14621 15856
rect 17164 15812 17204 15856
rect 18691 15855 18749 15856
rect 21379 15855 21504 15856
rect 21424 15836 21504 15855
rect 20515 15812 20573 15813
rect 2659 15772 2668 15812
rect 2708 15772 3724 15812
rect 3764 15772 3773 15812
rect 6019 15772 6028 15812
rect 6068 15772 7084 15812
rect 7124 15772 11360 15812
rect 12355 15772 12364 15812
rect 12404 15772 15724 15812
rect 15764 15772 15773 15812
rect 17164 15772 20524 15812
rect 20564 15772 20573 15812
rect 2659 15771 2717 15772
rect 7075 15771 7133 15772
rect 20515 15771 20573 15772
rect 13795 15728 13853 15729
rect 4771 15688 4780 15728
rect 4820 15688 5164 15728
rect 5204 15688 5213 15728
rect 5827 15688 5836 15728
rect 5876 15688 8620 15728
rect 8660 15688 8669 15728
rect 13411 15688 13420 15728
rect 13460 15688 13804 15728
rect 13844 15688 13853 15728
rect 14179 15688 14188 15728
rect 14228 15688 16012 15728
rect 16052 15688 16061 15728
rect 18403 15688 18412 15728
rect 18452 15688 18700 15728
rect 18740 15688 19084 15728
rect 19124 15688 19133 15728
rect 19459 15688 19468 15728
rect 19508 15688 20044 15728
rect 20084 15688 20093 15728
rect 13795 15687 13853 15688
rect 9091 15644 9149 15645
rect 20995 15644 21053 15645
rect 3235 15604 3244 15644
rect 3284 15604 5932 15644
rect 5972 15604 5981 15644
rect 7555 15604 7564 15644
rect 7604 15604 9100 15644
rect 9140 15604 9149 15644
rect 10915 15604 10924 15644
rect 10964 15604 11212 15644
rect 11252 15604 11261 15644
rect 13219 15604 13228 15644
rect 13268 15604 14956 15644
rect 14996 15604 15005 15644
rect 17923 15604 17932 15644
rect 17972 15604 21004 15644
rect 21044 15604 21053 15644
rect 9091 15603 9149 15604
rect 0 15560 80 15580
rect 1699 15560 1757 15561
rect 2755 15560 2813 15561
rect 9187 15560 9245 15561
rect 11875 15560 11933 15561
rect 19468 15560 19508 15604
rect 20995 15603 21053 15604
rect 0 15520 1516 15560
rect 1556 15520 1565 15560
rect 1699 15520 1708 15560
rect 1748 15520 2764 15560
rect 2804 15520 2813 15560
rect 3043 15520 3052 15560
rect 3092 15520 4012 15560
rect 4052 15520 4061 15560
rect 8227 15520 8236 15560
rect 8276 15520 8620 15560
rect 8660 15520 8669 15560
rect 9187 15520 9196 15560
rect 9236 15520 9484 15560
rect 9524 15520 9533 15560
rect 10243 15520 10252 15560
rect 10292 15520 10444 15560
rect 10484 15520 10493 15560
rect 11491 15520 11500 15560
rect 11540 15520 11884 15560
rect 11924 15520 12268 15560
rect 12308 15520 12317 15560
rect 13603 15520 13612 15560
rect 13652 15520 17356 15560
rect 17396 15520 17405 15560
rect 17827 15520 17836 15560
rect 17876 15520 18988 15560
rect 19028 15520 19037 15560
rect 19459 15520 19468 15560
rect 19508 15520 19517 15560
rect 0 15500 80 15520
rect 1699 15519 1757 15520
rect 2755 15519 2813 15520
rect 9187 15519 9245 15520
rect 11875 15519 11933 15520
rect 16867 15476 16925 15477
rect 19363 15476 19421 15477
rect 1699 15436 1708 15476
rect 1748 15436 15532 15476
rect 15572 15436 15581 15476
rect 16771 15436 16780 15476
rect 16820 15436 16876 15476
rect 16916 15436 16925 15476
rect 18115 15436 18124 15476
rect 18164 15436 18173 15476
rect 18787 15436 18796 15476
rect 18836 15436 19372 15476
rect 19412 15436 19421 15476
rect 16867 15435 16925 15436
rect 13603 15392 13661 15393
rect 2659 15352 2668 15392
rect 2708 15352 5836 15392
rect 5876 15352 8044 15392
rect 8084 15352 8093 15392
rect 13315 15352 13324 15392
rect 13364 15352 13612 15392
rect 13652 15352 13661 15392
rect 18124 15392 18164 15436
rect 19363 15435 19421 15436
rect 21424 15392 21504 15412
rect 18124 15352 19988 15392
rect 21187 15352 21196 15392
rect 21236 15352 21504 15392
rect 13603 15351 13661 15352
rect 1603 15308 1661 15309
rect 16963 15308 17021 15309
rect 17635 15308 17693 15309
rect 19948 15308 19988 15352
rect 21424 15332 21504 15352
rect 1603 15268 1612 15308
rect 1652 15268 4396 15308
rect 4436 15268 4445 15308
rect 12739 15268 12748 15308
rect 12788 15268 13228 15308
rect 13268 15268 13277 15308
rect 13699 15268 13708 15308
rect 13748 15268 13900 15308
rect 13940 15268 13949 15308
rect 14947 15268 14956 15308
rect 14996 15268 15532 15308
rect 15572 15268 15581 15308
rect 16963 15268 16972 15308
rect 17012 15268 17164 15308
rect 17204 15268 17213 15308
rect 17635 15268 17644 15308
rect 17684 15268 17740 15308
rect 17780 15268 17789 15308
rect 18307 15268 18316 15308
rect 18356 15268 18700 15308
rect 18740 15268 18749 15308
rect 19075 15268 19084 15308
rect 19124 15268 19468 15308
rect 19508 15268 19517 15308
rect 19939 15268 19948 15308
rect 19988 15268 19997 15308
rect 1603 15267 1661 15268
rect 16963 15267 17021 15268
rect 17635 15267 17693 15268
rect 0 15224 80 15244
rect 14947 15224 15005 15225
rect 0 15184 14956 15224
rect 14996 15184 15005 15224
rect 16387 15184 16396 15224
rect 16436 15184 16588 15224
rect 16628 15184 16637 15224
rect 17059 15184 17068 15224
rect 17108 15184 19372 15224
rect 19412 15184 19421 15224
rect 19651 15184 19660 15224
rect 19700 15184 19852 15224
rect 19892 15184 19901 15224
rect 0 15164 80 15184
rect 14947 15183 15005 15184
rect 19660 15141 19700 15184
rect 4579 15140 4637 15141
rect 5635 15140 5693 15141
rect 12451 15140 12509 15141
rect 16387 15140 16445 15141
rect 17155 15140 17213 15141
rect 19651 15140 19709 15141
rect 3679 15100 3688 15140
rect 3728 15100 3770 15140
rect 3810 15100 3852 15140
rect 3892 15100 3934 15140
rect 3974 15100 4016 15140
rect 4056 15100 4065 15140
rect 4494 15100 4588 15140
rect 4628 15100 4637 15140
rect 5443 15100 5452 15140
rect 5492 15100 5644 15140
rect 5684 15100 5693 15140
rect 7651 15100 7660 15140
rect 7700 15100 9964 15140
rect 10004 15100 10013 15140
rect 12366 15100 12460 15140
rect 12500 15100 12509 15140
rect 13123 15100 13132 15140
rect 13172 15100 15052 15140
rect 15092 15100 15101 15140
rect 16387 15100 16396 15140
rect 16436 15100 17164 15140
rect 17204 15100 17213 15140
rect 17443 15100 17452 15140
rect 17492 15100 17740 15140
rect 17780 15100 17789 15140
rect 18799 15100 18808 15140
rect 18848 15100 18890 15140
rect 18930 15100 18972 15140
rect 19012 15100 19054 15140
rect 19094 15100 19136 15140
rect 19176 15100 19185 15140
rect 19372 15100 19660 15140
rect 19700 15100 19709 15140
rect 4579 15099 4637 15100
rect 5635 15099 5693 15100
rect 12451 15099 12509 15100
rect 67 15056 125 15057
rect 1411 15056 1469 15057
rect 67 15016 76 15056
rect 116 15016 1420 15056
rect 1460 15016 1469 15056
rect 67 15015 125 15016
rect 1411 15015 1469 15016
rect 2467 14972 2525 14973
rect 5827 14972 5885 14973
rect 13132 14972 13172 15100
rect 16387 15099 16445 15100
rect 17155 15099 17213 15100
rect 19372 15056 19412 15100
rect 19651 15099 19709 15100
rect 16675 15016 16684 15056
rect 16724 15016 17356 15056
rect 17396 15016 17405 15056
rect 18115 15016 18124 15056
rect 18164 15016 18508 15056
rect 18548 15016 18557 15056
rect 19363 15016 19372 15056
rect 19412 15016 19421 15056
rect 19651 15016 19660 15056
rect 19700 15016 20236 15056
rect 20276 15016 20285 15056
rect 1219 14932 1228 14972
rect 1268 14932 1277 14972
rect 2382 14932 2476 14972
rect 2516 14932 2525 14972
rect 2659 14932 2668 14972
rect 2708 14932 4300 14972
rect 4340 14932 4349 14972
rect 5827 14932 5836 14972
rect 5876 14932 6028 14972
rect 6068 14932 8140 14972
rect 8180 14932 8189 14972
rect 11320 14932 13172 14972
rect 16195 14932 16204 14972
rect 16244 14932 17836 14972
rect 17876 14932 19468 14972
rect 19508 14932 19517 14972
rect 0 14888 80 14908
rect 1228 14888 1268 14932
rect 2467 14931 2525 14932
rect 5827 14931 5885 14932
rect 3139 14888 3197 14889
rect 9955 14888 10013 14889
rect 0 14848 1268 14888
rect 1987 14848 1996 14888
rect 2036 14848 3148 14888
rect 3188 14848 3916 14888
rect 3956 14848 9964 14888
rect 10004 14848 10828 14888
rect 10868 14848 10877 14888
rect 0 14828 80 14848
rect 3139 14847 3197 14848
rect 9955 14847 10013 14848
rect 3043 14804 3101 14805
rect 4195 14804 4253 14805
rect 11320 14804 11360 14932
rect 21187 14888 21245 14889
rect 21424 14888 21504 14908
rect 12163 14848 12172 14888
rect 12212 14848 12940 14888
rect 12980 14848 16492 14888
rect 16532 14848 16541 14888
rect 16771 14848 16780 14888
rect 16820 14848 18892 14888
rect 18932 14848 18941 14888
rect 19555 14848 19564 14888
rect 19604 14848 20044 14888
rect 20084 14848 20093 14888
rect 21187 14848 21196 14888
rect 21236 14848 21504 14888
rect 21187 14847 21245 14848
rect 21424 14828 21504 14848
rect 12739 14804 12797 14805
rect 2958 14764 3052 14804
rect 3092 14764 3101 14804
rect 4003 14764 4012 14804
rect 4052 14764 4204 14804
rect 4244 14764 4253 14804
rect 5635 14764 5644 14804
rect 5684 14764 5693 14804
rect 6220 14764 11360 14804
rect 12547 14764 12556 14804
rect 12596 14764 12748 14804
rect 12788 14764 12797 14804
rect 3043 14763 3101 14764
rect 4195 14763 4253 14764
rect 3523 14720 3581 14721
rect 1219 14680 1228 14720
rect 1268 14680 1364 14720
rect 2467 14680 2476 14720
rect 2516 14680 2956 14720
rect 2996 14680 3005 14720
rect 3438 14680 3532 14720
rect 3572 14680 3581 14720
rect 1324 14636 1364 14680
rect 3523 14679 3581 14680
rect 4483 14720 4541 14721
rect 5644 14720 5684 14764
rect 6220 14721 6260 14764
rect 12739 14763 12797 14764
rect 13795 14804 13853 14805
rect 13795 14764 13804 14804
rect 13844 14764 16108 14804
rect 16148 14764 16157 14804
rect 18499 14764 18508 14804
rect 18548 14764 19084 14804
rect 19124 14764 19133 14804
rect 19372 14764 19852 14804
rect 19892 14764 19901 14804
rect 13795 14763 13853 14764
rect 4483 14680 4492 14720
rect 4532 14680 5684 14720
rect 5731 14720 5789 14721
rect 6211 14720 6269 14721
rect 10435 14720 10493 14721
rect 10915 14720 10973 14721
rect 15715 14720 15773 14721
rect 5731 14680 5740 14720
rect 5780 14680 5932 14720
rect 5972 14680 5981 14720
rect 6126 14680 6220 14720
rect 6260 14680 6269 14720
rect 7171 14680 7180 14720
rect 7220 14680 7468 14720
rect 7508 14680 7517 14720
rect 8995 14680 9004 14720
rect 9044 14680 9964 14720
rect 10004 14680 10156 14720
rect 10196 14680 10205 14720
rect 10339 14680 10348 14720
rect 10388 14680 10444 14720
rect 10484 14680 10924 14720
rect 10964 14680 10973 14720
rect 12739 14680 12748 14720
rect 12788 14680 15724 14720
rect 15764 14680 18220 14720
rect 18260 14680 18269 14720
rect 18595 14680 18604 14720
rect 18644 14680 19276 14720
rect 19316 14680 19325 14720
rect 4483 14679 4541 14680
rect 5731 14679 5789 14680
rect 6211 14679 6269 14680
rect 10435 14679 10493 14680
rect 10915 14679 10973 14680
rect 15715 14679 15773 14680
rect 1987 14636 2045 14637
rect 5923 14636 5981 14637
rect 6220 14636 6260 14679
rect 8899 14636 8957 14637
rect 9475 14636 9533 14637
rect 16387 14636 16445 14637
rect 19372 14636 19412 14764
rect 19843 14720 19901 14721
rect 19843 14680 19852 14720
rect 19892 14680 19948 14720
rect 19988 14680 19997 14720
rect 19843 14679 19901 14680
rect 1324 14596 1996 14636
rect 2036 14596 4108 14636
rect 4148 14596 5876 14636
rect 1987 14595 2045 14596
rect 0 14552 80 14572
rect 1891 14552 1949 14553
rect 0 14512 1228 14552
rect 1268 14512 1277 14552
rect 1806 14512 1900 14552
rect 1940 14512 1949 14552
rect 3139 14512 3148 14552
rect 3188 14512 4972 14552
rect 5012 14512 5021 14552
rect 0 14492 80 14512
rect 1891 14511 1949 14512
rect 4771 14428 4780 14468
rect 4820 14428 5740 14468
rect 5780 14428 5789 14468
rect 1708 14344 2380 14384
rect 2420 14344 2429 14384
rect 4919 14344 4928 14384
rect 4968 14344 5010 14384
rect 5050 14344 5092 14384
rect 5132 14344 5174 14384
rect 5214 14344 5256 14384
rect 5296 14344 5305 14384
rect 1708 14300 1748 14344
rect 5836 14300 5876 14596
rect 5923 14596 5932 14636
rect 5972 14596 6260 14636
rect 8515 14596 8524 14636
rect 8564 14596 8908 14636
rect 8948 14596 9484 14636
rect 9524 14596 9533 14636
rect 5923 14595 5981 14596
rect 8899 14595 8957 14596
rect 9475 14595 9533 14596
rect 9580 14596 10732 14636
rect 10772 14596 13996 14636
rect 14036 14596 14764 14636
rect 14804 14596 14813 14636
rect 16301 14596 16396 14636
rect 16436 14596 16684 14636
rect 16724 14596 16733 14636
rect 18403 14596 18412 14636
rect 18452 14596 19412 14636
rect 19651 14636 19709 14637
rect 19651 14596 19660 14636
rect 19700 14596 19756 14636
rect 19796 14596 19805 14636
rect 20035 14596 20044 14636
rect 20084 14596 20093 14636
rect 6499 14512 6508 14552
rect 6548 14512 8428 14552
rect 8468 14512 8812 14552
rect 8852 14512 8861 14552
rect 9580 14468 9620 14596
rect 16387 14595 16445 14596
rect 19651 14595 19709 14596
rect 16867 14552 16925 14553
rect 11779 14512 11788 14552
rect 11828 14512 11980 14552
rect 12020 14512 12029 14552
rect 15619 14512 15628 14552
rect 15668 14512 16204 14552
rect 16244 14512 16253 14552
rect 16579 14512 16588 14552
rect 16628 14512 16876 14552
rect 16916 14512 16925 14552
rect 17635 14512 17644 14552
rect 17684 14512 19564 14552
rect 19604 14512 19613 14552
rect 16867 14511 16925 14512
rect 18691 14468 18749 14469
rect 20044 14468 20084 14596
rect 7651 14428 7660 14468
rect 7700 14428 9620 14468
rect 18403 14428 18412 14468
rect 18452 14428 18700 14468
rect 18740 14428 19084 14468
rect 19124 14428 19133 14468
rect 19939 14428 19948 14468
rect 19988 14428 20084 14468
rect 18691 14427 18749 14428
rect 11203 14384 11261 14385
rect 17635 14384 17693 14385
rect 21424 14384 21504 14404
rect 8515 14344 8524 14384
rect 8564 14344 9676 14384
rect 9716 14344 9725 14384
rect 11118 14344 11212 14384
rect 11252 14344 11261 14384
rect 11683 14344 11692 14384
rect 11732 14344 11980 14384
rect 12020 14344 12029 14384
rect 17550 14344 17644 14384
rect 17684 14344 17693 14384
rect 20039 14344 20048 14384
rect 20088 14344 20130 14384
rect 20170 14344 20212 14384
rect 20252 14344 20294 14384
rect 20334 14344 20376 14384
rect 20416 14344 20425 14384
rect 21187 14344 21196 14384
rect 21236 14344 21504 14384
rect 11203 14343 11261 14344
rect 17635 14343 17693 14344
rect 21424 14324 21504 14344
rect 9091 14300 9149 14301
rect 1699 14260 1708 14300
rect 1748 14260 1757 14300
rect 4099 14260 4108 14300
rect 4148 14260 5356 14300
rect 5396 14260 5405 14300
rect 5836 14260 9100 14300
rect 9140 14260 9149 14300
rect 9475 14260 9484 14300
rect 9524 14260 9533 14300
rect 13123 14260 13132 14300
rect 13172 14260 13516 14300
rect 13556 14260 13565 14300
rect 15811 14260 15820 14300
rect 15860 14260 16396 14300
rect 16436 14260 16445 14300
rect 9091 14259 9149 14260
rect 0 14216 80 14236
rect 6115 14216 6173 14217
rect 9484 14216 9524 14260
rect 11299 14216 11357 14217
rect 16291 14216 16349 14217
rect 0 14176 212 14216
rect 2275 14176 2284 14216
rect 2324 14176 3052 14216
rect 3092 14176 3101 14216
rect 4963 14176 4972 14216
rect 5012 14176 5452 14216
rect 5492 14176 5501 14216
rect 5731 14176 5740 14216
rect 5780 14176 6124 14216
rect 6164 14176 7276 14216
rect 7316 14176 7756 14216
rect 7796 14176 7805 14216
rect 9187 14176 9196 14216
rect 9236 14176 9524 14216
rect 9571 14176 9580 14216
rect 9620 14176 9868 14216
rect 9908 14176 9917 14216
rect 11214 14176 11308 14216
rect 11348 14176 11357 14216
rect 11587 14176 11596 14216
rect 11636 14176 16300 14216
rect 16340 14176 16349 14216
rect 0 14156 80 14176
rect 172 14048 212 14176
rect 6115 14175 6173 14176
rect 11299 14175 11357 14176
rect 16291 14175 16349 14176
rect 6211 14132 6269 14133
rect 13603 14132 13661 14133
rect 259 14092 268 14132
rect 308 14092 2860 14132
rect 2900 14092 2909 14132
rect 4204 14092 6028 14132
rect 6068 14092 6077 14132
rect 6211 14092 6220 14132
rect 6260 14092 10100 14132
rect 3811 14048 3869 14049
rect 4204 14048 4244 14092
rect 6211 14091 6269 14092
rect 10060 14048 10100 14092
rect 13603 14092 13612 14132
rect 13652 14092 14380 14132
rect 14420 14092 14429 14132
rect 16003 14092 16012 14132
rect 16052 14092 17164 14132
rect 17204 14092 17213 14132
rect 19651 14092 19660 14132
rect 19700 14092 20140 14132
rect 20180 14092 20189 14132
rect 13603 14091 13661 14092
rect 19747 14048 19805 14049
rect 172 14008 1228 14048
rect 1268 14008 1277 14048
rect 1795 14008 1804 14048
rect 1844 14008 2092 14048
rect 2132 14008 2141 14048
rect 3726 14008 3820 14048
rect 3860 14008 3869 14048
rect 4195 14008 4204 14048
rect 4244 14008 4253 14048
rect 6220 14008 6796 14048
rect 6836 14008 6988 14048
rect 7028 14008 7037 14048
rect 8419 14008 8428 14048
rect 8468 14008 9580 14048
rect 9620 14008 9629 14048
rect 10051 14008 10060 14048
rect 10100 14008 10636 14048
rect 10676 14008 10685 14048
rect 11980 14008 15188 14048
rect 15235 14008 15244 14048
rect 15284 14008 16972 14048
rect 17012 14008 17836 14048
rect 17876 14008 17885 14048
rect 19747 14008 19756 14048
rect 19796 14008 19852 14048
rect 19892 14008 19901 14048
rect 3811 14007 3869 14008
rect 6220 13964 6260 14008
rect 9187 13964 9245 13965
rect 11980 13964 12020 14008
rect 12355 13964 12413 13965
rect 15148 13964 15188 14008
rect 19747 14007 19805 14008
rect 1411 13924 1420 13964
rect 1460 13924 2572 13964
rect 2612 13924 2621 13964
rect 6019 13924 6028 13964
rect 6068 13924 6260 13964
rect 6307 13924 6316 13964
rect 6356 13924 6700 13964
rect 6740 13924 6749 13964
rect 8995 13924 9004 13964
rect 9044 13924 9196 13964
rect 9236 13924 9245 13964
rect 9187 13923 9245 13924
rect 10060 13924 10540 13964
rect 10580 13924 10589 13964
rect 11971 13924 11980 13964
rect 12020 13924 12029 13964
rect 12270 13924 12364 13964
rect 12404 13924 12413 13964
rect 12835 13924 12844 13964
rect 12884 13924 13228 13964
rect 13268 13924 13277 13964
rect 15148 13924 17452 13964
rect 17492 13924 17501 13964
rect 17836 13924 20180 13964
rect 0 13880 80 13900
rect 5635 13880 5693 13881
rect 10060 13880 10100 13924
rect 12355 13923 12413 13924
rect 0 13840 460 13880
rect 500 13840 509 13880
rect 2179 13840 2188 13880
rect 2228 13840 2612 13880
rect 2755 13840 2764 13880
rect 2804 13840 4300 13880
rect 4340 13840 4349 13880
rect 5635 13840 5644 13880
rect 5684 13840 10100 13880
rect 10147 13880 10205 13881
rect 11779 13880 11837 13881
rect 12163 13880 12221 13881
rect 17836 13880 17876 13924
rect 19468 13880 19508 13924
rect 19939 13880 19997 13881
rect 10147 13840 10156 13880
rect 10196 13840 10205 13880
rect 11694 13840 11788 13880
rect 11828 13840 11837 13880
rect 12078 13840 12172 13880
rect 12212 13840 12221 13880
rect 12643 13840 12652 13880
rect 12692 13840 13804 13880
rect 13844 13840 13853 13880
rect 15523 13840 15532 13880
rect 15572 13840 17260 13880
rect 17300 13840 17876 13880
rect 17923 13840 17932 13880
rect 17972 13840 19276 13880
rect 19316 13840 19325 13880
rect 19459 13840 19468 13880
rect 19508 13840 19517 13880
rect 19854 13840 19948 13880
rect 19988 13840 19997 13880
rect 20140 13880 20180 13924
rect 21424 13880 21504 13900
rect 20140 13840 21504 13880
rect 0 13820 80 13840
rect 2572 13796 2612 13840
rect 5635 13839 5693 13840
rect 10147 13839 10205 13840
rect 11779 13839 11837 13840
rect 12163 13839 12221 13840
rect 19939 13839 19997 13840
rect 4483 13796 4541 13797
rect 2572 13756 3244 13796
rect 3284 13756 4492 13796
rect 4532 13756 4541 13796
rect 4483 13755 4541 13756
rect 4675 13796 4733 13797
rect 10156 13796 10196 13839
rect 21424 13820 21504 13840
rect 12451 13796 12509 13797
rect 4675 13756 4684 13796
rect 4724 13756 8140 13796
rect 8180 13756 8189 13796
rect 10156 13756 12460 13796
rect 12500 13756 12509 13796
rect 15715 13756 15724 13796
rect 15764 13756 16204 13796
rect 16244 13756 16253 13796
rect 16387 13756 16396 13796
rect 16436 13756 17068 13796
rect 17108 13756 17117 13796
rect 4675 13755 4733 13756
rect 12451 13755 12509 13756
rect 15811 13712 15869 13713
rect 18691 13712 18749 13713
rect 19267 13712 19325 13713
rect 1411 13672 1420 13712
rect 1460 13672 15436 13712
rect 15476 13672 15485 13712
rect 15811 13672 15820 13712
rect 15860 13672 16588 13712
rect 16628 13672 16637 13712
rect 18691 13672 18700 13712
rect 18740 13672 19276 13712
rect 19316 13672 19325 13712
rect 15811 13671 15869 13672
rect 18691 13671 18749 13672
rect 19267 13671 19325 13672
rect 2467 13628 2525 13629
rect 12259 13628 12317 13629
rect 13219 13628 13277 13629
rect 2371 13588 2380 13628
rect 2420 13588 2476 13628
rect 2516 13588 2525 13628
rect 3235 13588 3244 13628
rect 3284 13588 3532 13628
rect 3572 13588 3581 13628
rect 3679 13588 3688 13628
rect 3728 13588 3770 13628
rect 3810 13588 3852 13628
rect 3892 13588 3934 13628
rect 3974 13588 4016 13628
rect 4056 13588 4065 13628
rect 4291 13588 4300 13628
rect 4340 13588 7756 13628
rect 7796 13588 7805 13628
rect 12259 13588 12268 13628
rect 12308 13588 13228 13628
rect 13268 13588 13277 13628
rect 18799 13588 18808 13628
rect 18848 13588 18890 13628
rect 18930 13588 18972 13628
rect 19012 13588 19054 13628
rect 19094 13588 19136 13628
rect 19176 13588 19185 13628
rect 2467 13587 2525 13588
rect 12259 13587 12317 13588
rect 13219 13587 13277 13588
rect 0 13544 80 13564
rect 4579 13544 4637 13545
rect 7459 13544 7517 13545
rect 0 13504 4588 13544
rect 4628 13504 4637 13544
rect 6787 13504 6796 13544
rect 6836 13504 7468 13544
rect 7508 13504 11360 13544
rect 13219 13504 13228 13544
rect 13268 13504 15820 13544
rect 15860 13504 15869 13544
rect 0 13484 80 13504
rect 4579 13503 4637 13504
rect 7459 13503 7517 13504
rect 1027 13460 1085 13461
rect 10435 13460 10493 13461
rect 1027 13420 1036 13460
rect 1076 13420 2540 13460
rect 3331 13420 3340 13460
rect 3380 13420 4588 13460
rect 4628 13420 4637 13460
rect 5635 13420 5644 13460
rect 5684 13420 7564 13460
rect 7604 13420 7613 13460
rect 7660 13420 10444 13460
rect 10484 13420 10493 13460
rect 1027 13419 1085 13420
rect 2500 13292 2540 13420
rect 7660 13376 7700 13420
rect 10435 13419 10493 13420
rect 11320 13376 11360 13504
rect 13228 13460 13268 13504
rect 19363 13460 19421 13461
rect 11491 13420 11500 13460
rect 11540 13420 13268 13460
rect 13411 13420 13420 13460
rect 13460 13420 13612 13460
rect 13652 13420 13661 13460
rect 17731 13420 17740 13460
rect 17780 13420 18124 13460
rect 18164 13420 18604 13460
rect 18644 13420 18653 13460
rect 18883 13420 18892 13460
rect 18932 13420 19372 13460
rect 19412 13420 19421 13460
rect 18604 13376 18644 13420
rect 19363 13419 19421 13420
rect 19939 13376 19997 13377
rect 21424 13376 21504 13396
rect 2659 13336 2668 13376
rect 2708 13336 2860 13376
rect 2900 13336 2909 13376
rect 3619 13336 3628 13376
rect 3668 13336 7700 13376
rect 7843 13336 7852 13376
rect 7892 13336 9772 13376
rect 9812 13336 9821 13376
rect 11320 13336 15244 13376
rect 15284 13336 15293 13376
rect 18604 13336 18988 13376
rect 19028 13336 19180 13376
rect 19220 13336 19229 13376
rect 19843 13336 19852 13376
rect 19892 13336 19948 13376
rect 19988 13336 19997 13376
rect 19939 13335 19997 13336
rect 20140 13336 21504 13376
rect 8323 13292 8381 13293
rect 20140 13292 20180 13336
rect 21424 13316 21504 13336
rect 2500 13252 8332 13292
rect 8372 13252 8381 13292
rect 8323 13251 8381 13252
rect 11308 13252 11500 13292
rect 11540 13252 11549 13292
rect 11683 13252 11692 13292
rect 11732 13252 16780 13292
rect 16820 13252 16829 13292
rect 17731 13252 17740 13292
rect 17780 13252 20180 13292
rect 0 13208 80 13228
rect 2467 13208 2525 13209
rect 4099 13208 4157 13209
rect 4579 13208 4637 13209
rect 5347 13208 5405 13209
rect 6307 13208 6365 13209
rect 9763 13208 9821 13209
rect 11308 13208 11348 13252
rect 0 13168 940 13208
rect 980 13168 989 13208
rect 1699 13168 1708 13208
rect 1748 13168 2476 13208
rect 2516 13168 4108 13208
rect 4148 13168 4157 13208
rect 4494 13168 4588 13208
rect 4628 13168 4637 13208
rect 5251 13168 5260 13208
rect 5300 13168 5356 13208
rect 5396 13168 5405 13208
rect 5539 13168 5548 13208
rect 5588 13168 6028 13208
rect 6068 13168 6077 13208
rect 6307 13168 6316 13208
rect 6356 13168 9772 13208
rect 9812 13168 9868 13208
rect 9908 13168 9917 13208
rect 9964 13168 11116 13208
rect 11156 13168 11348 13208
rect 11395 13208 11453 13209
rect 19363 13208 19421 13209
rect 11395 13168 11404 13208
rect 11444 13168 11538 13208
rect 11779 13168 11788 13208
rect 11828 13168 12268 13208
rect 12308 13168 12317 13208
rect 13891 13168 13900 13208
rect 13940 13168 16492 13208
rect 16532 13168 16541 13208
rect 18211 13168 18220 13208
rect 18260 13168 19372 13208
rect 19412 13168 19468 13208
rect 19508 13168 19517 13208
rect 0 13148 80 13168
rect 2467 13167 2525 13168
rect 4099 13167 4157 13168
rect 4579 13167 4637 13168
rect 5347 13167 5405 13168
rect 6307 13167 6365 13168
rect 9763 13167 9821 13168
rect 2947 13124 3005 13125
rect 9964 13124 10004 13168
rect 11395 13167 11453 13168
rect 19363 13167 19421 13168
rect 2862 13084 2956 13124
rect 2996 13084 5300 13124
rect 8131 13084 8140 13124
rect 8180 13084 8428 13124
rect 8468 13084 8477 13124
rect 9379 13084 9388 13124
rect 9428 13084 10004 13124
rect 10051 13124 10109 13125
rect 19459 13124 19517 13125
rect 10051 13084 10060 13124
rect 10100 13084 10252 13124
rect 10292 13084 10301 13124
rect 13603 13084 13612 13124
rect 13652 13084 14188 13124
rect 14228 13084 14237 13124
rect 19459 13084 19468 13124
rect 19508 13084 20140 13124
rect 20180 13084 20189 13124
rect 2947 13083 3005 13084
rect 5260 13040 5300 13084
rect 10051 13083 10109 13084
rect 19459 13083 19517 13084
rect 11395 13040 11453 13041
rect 739 13000 748 13040
rect 788 13000 3340 13040
rect 3380 13000 3389 13040
rect 5260 13000 5396 13040
rect 7651 13000 7660 13040
rect 7700 13000 10828 13040
rect 10868 13000 10877 13040
rect 11395 13000 11404 13040
rect 11444 13000 11500 13040
rect 11540 13000 11549 13040
rect 14083 13000 14092 13040
rect 14132 13000 17740 13040
rect 17780 13000 17789 13040
rect 19843 13000 19852 13040
rect 19892 13000 20044 13040
rect 20084 13000 20093 13040
rect 0 12872 80 12892
rect 835 12872 893 12873
rect 3139 12872 3197 12873
rect 0 12832 212 12872
rect 0 12812 80 12832
rect 172 12704 212 12832
rect 835 12832 844 12872
rect 884 12832 3148 12872
rect 3188 12832 3197 12872
rect 835 12831 893 12832
rect 3139 12831 3197 12832
rect 4387 12872 4445 12873
rect 5356 12872 5396 13000
rect 11395 12999 11453 13000
rect 9955 12872 10013 12873
rect 21424 12872 21504 12892
rect 4387 12832 4396 12872
rect 4436 12832 4530 12872
rect 4919 12832 4928 12872
rect 4968 12832 5010 12872
rect 5050 12832 5092 12872
rect 5132 12832 5174 12872
rect 5214 12832 5256 12872
rect 5296 12832 5305 12872
rect 5356 12832 9388 12872
rect 9428 12832 9437 12872
rect 9763 12832 9772 12872
rect 9812 12832 9964 12872
rect 10004 12832 14228 12872
rect 20039 12832 20048 12872
rect 20088 12832 20130 12872
rect 20170 12832 20212 12872
rect 20252 12832 20294 12872
rect 20334 12832 20376 12872
rect 20416 12832 20425 12872
rect 20812 12832 21504 12872
rect 4387 12831 4445 12832
rect 9955 12831 10013 12832
rect 4771 12788 4829 12789
rect 11971 12788 12029 12789
rect 643 12748 652 12788
rect 692 12748 3724 12788
rect 3764 12748 3773 12788
rect 4771 12748 4780 12788
rect 4820 12748 5932 12788
rect 5972 12748 5981 12788
rect 11320 12748 11980 12788
rect 12020 12748 12029 12788
rect 14188 12788 14228 12832
rect 20812 12788 20852 12832
rect 21424 12812 21504 12832
rect 14188 12748 20852 12788
rect 4771 12747 4829 12748
rect 11320 12704 11360 12748
rect 11971 12747 12029 12748
rect 172 12664 11360 12704
rect 14284 12664 17164 12704
rect 17204 12664 17213 12704
rect 17443 12664 17452 12704
rect 17492 12664 17501 12704
rect 18979 12664 18988 12704
rect 19028 12664 19852 12704
rect 19892 12664 19901 12704
rect 355 12620 413 12621
rect 4195 12620 4253 12621
rect 8611 12620 8669 12621
rect 14284 12620 14324 12664
rect 270 12580 364 12620
rect 404 12580 413 12620
rect 1699 12580 1708 12620
rect 1748 12580 2860 12620
rect 2900 12580 2909 12620
rect 4003 12580 4012 12620
rect 4052 12580 4204 12620
rect 4244 12580 6700 12620
rect 6740 12580 6749 12620
rect 7747 12580 7756 12620
rect 7796 12580 8236 12620
rect 8276 12580 8285 12620
rect 8611 12580 8620 12620
rect 8660 12580 8716 12620
rect 8756 12580 8765 12620
rect 9091 12580 9100 12620
rect 9140 12580 10100 12620
rect 355 12579 413 12580
rect 4195 12579 4253 12580
rect 8611 12579 8669 12580
rect 0 12536 80 12556
rect 3523 12536 3581 12537
rect 5155 12536 5213 12537
rect 7075 12536 7133 12537
rect 10060 12536 10100 12580
rect 11320 12580 14324 12620
rect 15427 12580 15436 12620
rect 15476 12580 17260 12620
rect 17300 12580 17309 12620
rect 11320 12536 11360 12580
rect 17452 12536 17492 12664
rect 18019 12580 18028 12620
rect 18068 12580 19084 12620
rect 19124 12580 19133 12620
rect 0 12496 172 12536
rect 212 12496 221 12536
rect 3438 12496 3532 12536
rect 3572 12496 4532 12536
rect 4579 12496 4588 12536
rect 4628 12496 4972 12536
rect 5012 12496 5021 12536
rect 5070 12496 5164 12536
rect 5204 12496 5213 12536
rect 0 12476 80 12496
rect 3523 12495 3581 12496
rect 355 12452 413 12453
rect 1507 12452 1565 12453
rect 4492 12452 4532 12496
rect 5155 12495 5213 12496
rect 5260 12496 5876 12536
rect 6211 12496 6220 12536
rect 6260 12496 6796 12536
rect 6836 12496 7084 12536
rect 7124 12496 7133 12536
rect 7843 12496 7852 12536
rect 7892 12496 9484 12536
rect 9524 12496 9533 12536
rect 10051 12496 10060 12536
rect 10100 12496 10109 12536
rect 10339 12496 10348 12536
rect 10388 12496 11116 12536
rect 11156 12496 11308 12536
rect 11348 12496 11360 12536
rect 11683 12496 11692 12536
rect 11732 12496 12364 12536
rect 12404 12496 13036 12536
rect 13076 12496 13900 12536
rect 13940 12496 13949 12536
rect 14083 12496 14092 12536
rect 14132 12496 15476 12536
rect 16579 12496 16588 12536
rect 16628 12496 17396 12536
rect 17452 12496 19276 12536
rect 19316 12496 19325 12536
rect 5260 12452 5300 12496
rect 355 12412 364 12452
rect 404 12412 1516 12452
rect 1556 12412 1565 12452
rect 2467 12412 2476 12452
rect 2516 12412 2540 12452
rect 4492 12412 5300 12452
rect 355 12411 413 12412
rect 1507 12411 1565 12412
rect 2500 12368 2540 12412
rect 2947 12368 3005 12369
rect 5836 12368 5876 12496
rect 7075 12495 7133 12496
rect 15436 12452 15476 12496
rect 17356 12452 17396 12496
rect 5923 12412 5932 12452
rect 5972 12412 6412 12452
rect 6452 12412 6461 12452
rect 7459 12412 7468 12452
rect 7508 12412 8840 12452
rect 9283 12412 9292 12452
rect 9332 12412 15340 12452
rect 15380 12412 15389 12452
rect 15436 12412 17164 12452
rect 17204 12412 17213 12452
rect 17347 12412 17356 12452
rect 17396 12412 19756 12452
rect 19796 12412 19805 12452
rect 2500 12328 2956 12368
rect 2996 12328 3005 12368
rect 2947 12327 3005 12328
rect 3724 12328 4780 12368
rect 4820 12328 4829 12368
rect 5836 12328 6316 12368
rect 6356 12328 6365 12368
rect 3724 12284 3764 12328
rect 6115 12284 6173 12285
rect 2275 12244 2284 12284
rect 2324 12244 3764 12284
rect 3907 12244 3916 12284
rect 3956 12244 4204 12284
rect 4244 12244 4253 12284
rect 5347 12244 5356 12284
rect 5396 12244 5644 12284
rect 5684 12244 6124 12284
rect 6164 12244 6173 12284
rect 8800 12284 8840 12412
rect 11320 12368 11360 12412
rect 9379 12328 9388 12368
rect 9428 12328 11060 12368
rect 11107 12328 11116 12368
rect 11156 12328 11360 12368
rect 12259 12368 12317 12369
rect 21424 12368 21504 12388
rect 12259 12328 12268 12368
rect 12308 12328 21504 12368
rect 8800 12244 9004 12284
rect 9044 12244 9292 12284
rect 9332 12244 9341 12284
rect 10147 12244 10156 12284
rect 10196 12244 10444 12284
rect 10484 12244 10493 12284
rect 6115 12243 6173 12244
rect 0 12200 80 12220
rect 3427 12200 3485 12201
rect 11020 12200 11060 12328
rect 12259 12327 12317 12328
rect 21424 12308 21504 12328
rect 14467 12284 14525 12285
rect 20035 12284 20093 12285
rect 11971 12244 11980 12284
rect 12020 12244 12364 12284
rect 12404 12244 12413 12284
rect 13699 12244 13708 12284
rect 13748 12244 14188 12284
rect 14228 12244 14237 12284
rect 14467 12244 14476 12284
rect 14516 12244 14860 12284
rect 14900 12244 14909 12284
rect 19267 12244 19276 12284
rect 19316 12244 19852 12284
rect 19892 12244 19901 12284
rect 19950 12244 20044 12284
rect 20084 12244 20093 12284
rect 14467 12243 14525 12244
rect 20035 12243 20093 12244
rect 0 12160 2092 12200
rect 2132 12160 2141 12200
rect 3427 12160 3436 12200
rect 3476 12160 6452 12200
rect 6691 12160 6700 12200
rect 6740 12160 9868 12200
rect 9908 12160 9917 12200
rect 11020 12160 12748 12200
rect 12788 12160 12797 12200
rect 13507 12160 13516 12200
rect 13556 12160 13996 12200
rect 14036 12160 15916 12200
rect 15956 12160 20524 12200
rect 20564 12160 20573 12200
rect 0 12140 80 12160
rect 3427 12159 3485 12160
rect 6307 12116 6365 12117
rect 3679 12076 3688 12116
rect 3728 12076 3770 12116
rect 3810 12076 3852 12116
rect 3892 12076 3934 12116
rect 3974 12076 4016 12116
rect 4056 12076 4065 12116
rect 4675 12076 4684 12116
rect 4724 12076 5068 12116
rect 5108 12076 5117 12116
rect 5356 12076 6316 12116
rect 6356 12076 6365 12116
rect 5356 12032 5396 12076
rect 6307 12075 6365 12076
rect 1315 11992 1324 12032
rect 1364 11992 5396 12032
rect 5539 12032 5597 12033
rect 5539 11992 5548 12032
rect 5588 11992 5836 12032
rect 5876 11992 5885 12032
rect 5539 11991 5597 11992
rect 2083 11948 2141 11949
rect 4771 11948 4829 11949
rect 6412 11948 6452 12160
rect 6595 12116 6653 12117
rect 10147 12116 10205 12117
rect 6595 12076 6604 12116
rect 6644 12076 10156 12116
rect 10196 12076 10205 12116
rect 6595 12075 6653 12076
rect 10147 12075 10205 12076
rect 12547 12116 12605 12117
rect 12547 12076 12556 12116
rect 12596 12076 14476 12116
rect 14516 12076 14525 12116
rect 18799 12076 18808 12116
rect 18848 12076 18890 12116
rect 18930 12076 18972 12116
rect 19012 12076 19054 12116
rect 19094 12076 19136 12116
rect 19176 12076 19185 12116
rect 12547 12075 12605 12076
rect 6883 11992 6892 12032
rect 6932 11992 7468 12032
rect 7508 11992 7517 12032
rect 7660 11992 8236 12032
rect 8276 11992 10636 12032
rect 10676 11992 10685 12032
rect 13411 11992 13420 12032
rect 13460 11992 14092 12032
rect 14132 11992 14141 12032
rect 14380 11992 18700 12032
rect 18740 11992 18749 12032
rect 7660 11948 7700 11992
rect 7843 11948 7901 11949
rect 9187 11948 9245 11949
rect 14380 11948 14420 11992
rect 2083 11908 2092 11948
rect 2132 11908 3148 11948
rect 3188 11908 4780 11948
rect 4820 11908 4829 11948
rect 5155 11908 5164 11948
rect 5204 11908 6124 11948
rect 6164 11908 6173 11948
rect 6412 11908 7604 11948
rect 7651 11908 7660 11948
rect 7700 11908 7709 11948
rect 7843 11908 7852 11948
rect 7892 11908 9196 11948
rect 9236 11908 9245 11948
rect 9763 11908 9772 11948
rect 9812 11908 10732 11948
rect 10772 11908 10781 11948
rect 11587 11908 11596 11948
rect 11636 11908 14420 11948
rect 14467 11908 14476 11948
rect 14516 11908 19468 11948
rect 19508 11908 19517 11948
rect 19939 11908 19948 11948
rect 19988 11908 20716 11948
rect 20756 11908 20765 11948
rect 2083 11907 2141 11908
rect 4771 11907 4829 11908
rect 0 11864 80 11884
rect 3427 11864 3485 11865
rect 5347 11864 5405 11865
rect 7564 11864 7604 11908
rect 7843 11907 7901 11908
rect 9187 11907 9245 11908
rect 8227 11864 8285 11865
rect 12643 11864 12701 11865
rect 13507 11864 13565 11865
rect 15139 11864 15197 11865
rect 16963 11864 17021 11865
rect 0 11824 556 11864
rect 596 11824 605 11864
rect 2764 11824 3436 11864
rect 3476 11824 3485 11864
rect 4675 11824 4684 11864
rect 4724 11824 5356 11864
rect 5396 11824 7276 11864
rect 7316 11824 7325 11864
rect 7564 11824 8236 11864
rect 8276 11824 8285 11864
rect 9859 11824 9868 11864
rect 9908 11824 9917 11864
rect 10435 11824 10444 11864
rect 10484 11824 11116 11864
rect 11156 11824 11165 11864
rect 12558 11824 12652 11864
rect 12692 11824 13516 11864
rect 13556 11824 13565 11864
rect 15043 11824 15052 11864
rect 15092 11824 15148 11864
rect 15188 11824 15197 11864
rect 15619 11824 15628 11864
rect 15668 11824 16972 11864
rect 17012 11824 17021 11864
rect 0 11804 80 11824
rect 2764 11696 2804 11824
rect 3427 11823 3485 11824
rect 5347 11823 5405 11824
rect 8227 11823 8285 11824
rect 5155 11780 5213 11781
rect 5635 11780 5693 11781
rect 6691 11780 6749 11781
rect 2947 11740 2956 11780
rect 2996 11740 5108 11780
rect 3715 11696 3773 11697
rect 1315 11656 1324 11696
rect 1364 11656 2804 11696
rect 2851 11656 2860 11696
rect 2900 11656 3724 11696
rect 3764 11656 3773 11696
rect 3715 11655 3773 11656
rect 1699 11612 1757 11613
rect 5068 11612 5108 11740
rect 5155 11740 5164 11780
rect 5204 11740 5644 11780
rect 5684 11740 5693 11780
rect 5923 11740 5932 11780
rect 5972 11740 6316 11780
rect 6356 11740 6508 11780
rect 6548 11740 6557 11780
rect 6691 11740 6700 11780
rect 6740 11740 6796 11780
rect 6836 11740 6845 11780
rect 5155 11739 5213 11740
rect 5635 11739 5693 11740
rect 6691 11739 6749 11740
rect 9667 11696 9725 11697
rect 5827 11656 5836 11696
rect 5876 11656 8524 11696
rect 8564 11656 8573 11696
rect 9091 11656 9100 11696
rect 9140 11656 9388 11696
rect 9428 11656 9437 11696
rect 9571 11656 9580 11696
rect 9620 11656 9676 11696
rect 9716 11656 9725 11696
rect 9868 11696 9908 11824
rect 12643 11823 12701 11824
rect 13507 11823 13565 11824
rect 15139 11823 15197 11824
rect 16963 11823 17021 11824
rect 18019 11864 18077 11865
rect 19747 11864 19805 11865
rect 21424 11864 21504 11884
rect 18019 11824 18028 11864
rect 18068 11824 19084 11864
rect 19124 11824 19133 11864
rect 19747 11824 19756 11864
rect 19796 11824 21504 11864
rect 18019 11823 18077 11824
rect 19747 11823 19805 11824
rect 21424 11804 21504 11824
rect 10435 11780 10493 11781
rect 10435 11740 10444 11780
rect 10484 11740 10732 11780
rect 10772 11740 10781 11780
rect 11116 11740 21004 11780
rect 21044 11740 21053 11780
rect 10435 11739 10493 11740
rect 11116 11696 11156 11740
rect 9868 11656 11156 11696
rect 11971 11696 12029 11697
rect 13027 11696 13085 11697
rect 13795 11696 13853 11697
rect 15811 11696 15869 11697
rect 11971 11656 11980 11696
rect 12020 11656 12268 11696
rect 12308 11656 13036 11696
rect 13076 11656 13085 11696
rect 13219 11656 13228 11696
rect 13268 11656 13804 11696
rect 13844 11656 13853 11696
rect 14275 11656 14284 11696
rect 14324 11656 14476 11696
rect 14516 11656 14525 11696
rect 15523 11656 15532 11696
rect 15572 11656 15820 11696
rect 15860 11656 15869 11696
rect 9667 11655 9725 11656
rect 11971 11655 12029 11656
rect 13027 11655 13085 11656
rect 13795 11655 13853 11656
rect 15811 11655 15869 11656
rect 16675 11696 16733 11697
rect 16963 11696 17021 11697
rect 16675 11656 16684 11696
rect 16724 11656 16780 11696
rect 16820 11656 16829 11696
rect 16963 11656 16972 11696
rect 17012 11656 19468 11696
rect 19508 11656 19517 11696
rect 16675 11655 16733 11656
rect 16963 11655 17021 11656
rect 6307 11612 6365 11613
rect 7267 11612 7325 11613
rect 1027 11572 1036 11612
rect 1076 11572 1708 11612
rect 1748 11572 1757 11612
rect 2755 11572 2764 11612
rect 2804 11572 4972 11612
rect 5012 11572 5021 11612
rect 5068 11572 6068 11612
rect 1699 11571 1757 11572
rect 0 11528 80 11548
rect 6028 11528 6068 11572
rect 6307 11572 6316 11612
rect 6356 11572 6796 11612
rect 6836 11572 6845 11612
rect 7267 11572 7276 11612
rect 7316 11572 11360 11612
rect 12931 11572 12940 11612
rect 12980 11572 13804 11612
rect 13844 11572 13853 11612
rect 13996 11572 17012 11612
rect 18787 11572 18796 11612
rect 18836 11572 19948 11612
rect 19988 11572 19997 11612
rect 6307 11571 6365 11572
rect 7267 11571 7325 11572
rect 7843 11528 7901 11529
rect 11320 11528 11360 11572
rect 13996 11528 14036 11572
rect 14179 11528 14237 11529
rect 16972 11528 17012 11572
rect 20035 11528 20093 11529
rect 0 11488 1900 11528
rect 1940 11488 1949 11528
rect 4483 11488 4492 11528
rect 4532 11488 5932 11528
rect 5972 11488 5981 11528
rect 6028 11488 7852 11528
rect 7892 11488 7901 11528
rect 9667 11488 9676 11528
rect 9716 11488 9964 11528
rect 10004 11488 10013 11528
rect 11320 11488 14036 11528
rect 14083 11488 14092 11528
rect 14132 11488 14188 11528
rect 14228 11488 14237 11528
rect 14563 11488 14572 11528
rect 14612 11488 14764 11528
rect 14804 11488 14813 11528
rect 16771 11488 16780 11528
rect 16820 11488 16829 11528
rect 16963 11488 16972 11528
rect 17012 11488 17021 11528
rect 17731 11488 17740 11528
rect 17780 11488 19372 11528
rect 19412 11488 19421 11528
rect 19950 11488 20044 11528
rect 20084 11488 20093 11528
rect 0 11468 80 11488
rect 7843 11487 7901 11488
rect 14179 11487 14237 11488
rect 15427 11444 15485 11445
rect 2467 11404 2476 11444
rect 2516 11404 2668 11444
rect 2708 11404 2717 11444
rect 3148 11404 3436 11444
rect 3476 11404 3485 11444
rect 5548 11404 7564 11444
rect 7604 11404 7613 11444
rect 7939 11404 7948 11444
rect 7988 11404 11308 11444
rect 11348 11404 11357 11444
rect 14476 11404 15436 11444
rect 15476 11404 15485 11444
rect 16780 11444 16820 11488
rect 20035 11487 20093 11488
rect 18883 11444 18941 11445
rect 19747 11444 19805 11445
rect 16780 11404 17012 11444
rect 3148 11276 3188 11404
rect 5548 11360 5588 11404
rect 7075 11360 7133 11361
rect 9475 11360 9533 11361
rect 13507 11360 13565 11361
rect 14476 11360 14516 11404
rect 15427 11403 15485 11404
rect 16972 11360 17012 11404
rect 18883 11404 18892 11444
rect 18932 11404 19756 11444
rect 19796 11404 19805 11444
rect 18883 11403 18941 11404
rect 19747 11403 19805 11404
rect 21091 11360 21149 11361
rect 21424 11360 21504 11380
rect 4919 11320 4928 11360
rect 4968 11320 5010 11360
rect 5050 11320 5092 11360
rect 5132 11320 5174 11360
rect 5214 11320 5256 11360
rect 5296 11320 5305 11360
rect 5508 11320 5548 11360
rect 5588 11320 5597 11360
rect 7075 11320 7084 11360
rect 7124 11320 7180 11360
rect 7220 11320 7229 11360
rect 9388 11320 9484 11360
rect 9524 11320 9868 11360
rect 9908 11320 9917 11360
rect 10339 11320 10348 11360
rect 10388 11320 10397 11360
rect 13315 11320 13324 11360
rect 13364 11320 13516 11360
rect 13556 11320 13565 11360
rect 14436 11320 14476 11360
rect 14516 11320 14525 11360
rect 16932 11320 16972 11360
rect 17012 11320 17021 11360
rect 19660 11320 19892 11360
rect 20039 11320 20048 11360
rect 20088 11320 20130 11360
rect 20170 11320 20212 11360
rect 20252 11320 20294 11360
rect 20334 11320 20376 11360
rect 20416 11320 20425 11360
rect 21091 11320 21100 11360
rect 21140 11320 21504 11360
rect 7075 11319 7133 11320
rect 2851 11236 2860 11276
rect 2900 11236 3188 11276
rect 4099 11276 4157 11277
rect 9388 11276 9428 11320
rect 9475 11319 9533 11320
rect 10348 11276 10388 11320
rect 13507 11319 13565 11320
rect 10435 11276 10493 11277
rect 14083 11276 14141 11277
rect 16387 11276 16445 11277
rect 18979 11276 19037 11277
rect 19660 11276 19700 11320
rect 19852 11276 19892 11320
rect 21091 11319 21149 11320
rect 21424 11300 21504 11320
rect 4099 11236 4108 11276
rect 4148 11236 4396 11276
rect 4436 11236 4445 11276
rect 5443 11236 5452 11276
rect 5492 11236 6220 11276
rect 6260 11236 6269 11276
rect 7843 11236 7852 11276
rect 7892 11236 8140 11276
rect 8180 11236 8189 11276
rect 9379 11236 9388 11276
rect 9428 11236 9437 11276
rect 10348 11236 10444 11276
rect 10484 11236 10493 11276
rect 13891 11236 13900 11276
rect 13940 11236 14092 11276
rect 14132 11236 14141 11276
rect 14563 11236 14572 11276
rect 14612 11236 16396 11276
rect 16436 11236 16445 11276
rect 18894 11236 18988 11276
rect 19028 11236 19037 11276
rect 19171 11236 19180 11276
rect 19220 11236 19700 11276
rect 19747 11236 19756 11276
rect 19796 11236 19805 11276
rect 19852 11236 20180 11276
rect 4099 11235 4157 11236
rect 10435 11235 10493 11236
rect 14083 11235 14141 11236
rect 16387 11235 16445 11236
rect 18979 11235 19037 11236
rect 0 11192 80 11212
rect 19756 11192 19796 11236
rect 20140 11192 20180 11236
rect 0 11152 940 11192
rect 980 11152 989 11192
rect 6019 11152 6028 11192
rect 6068 11152 10540 11192
rect 10580 11152 10589 11192
rect 11683 11152 11692 11192
rect 11732 11152 14380 11192
rect 14420 11152 14429 11192
rect 15811 11152 15820 11192
rect 15860 11152 16396 11192
rect 16436 11152 16445 11192
rect 17059 11152 17068 11192
rect 17108 11152 18412 11192
rect 18452 11152 18700 11192
rect 18740 11152 20044 11192
rect 20084 11152 20093 11192
rect 20140 11152 20236 11192
rect 20276 11152 20285 11192
rect 0 11132 80 11152
rect 4099 11108 4157 11109
rect 11491 11108 11549 11109
rect 16771 11108 16829 11109
rect 1603 11068 1612 11108
rect 1652 11068 1804 11108
rect 1844 11068 2764 11108
rect 2804 11068 2813 11108
rect 3427 11068 3436 11108
rect 3476 11068 4108 11108
rect 4148 11068 5068 11108
rect 5108 11068 6700 11108
rect 6740 11068 6749 11108
rect 6979 11068 6988 11108
rect 7028 11068 11020 11108
rect 11060 11068 11069 11108
rect 11395 11068 11404 11108
rect 11444 11068 11500 11108
rect 11540 11068 11549 11108
rect 12259 11068 12268 11108
rect 12308 11068 12556 11108
rect 12596 11068 12605 11108
rect 13123 11068 13132 11108
rect 13172 11068 15052 11108
rect 15092 11068 15101 11108
rect 16099 11068 16108 11108
rect 16148 11068 16492 11108
rect 16532 11068 16541 11108
rect 16771 11068 16780 11108
rect 16820 11068 19180 11108
rect 19220 11068 19229 11108
rect 19651 11068 19660 11108
rect 19700 11068 20620 11108
rect 20660 11068 20669 11108
rect 4099 11067 4157 11068
rect 11491 11067 11549 11068
rect 16771 11067 16829 11068
rect 9571 11024 9629 11025
rect 16867 11024 16925 11025
rect 1315 10984 1324 11024
rect 1364 10984 2476 11024
rect 2516 10984 2525 11024
rect 3811 10984 3820 11024
rect 3860 10984 7372 11024
rect 7412 10984 9580 11024
rect 9620 10984 15244 11024
rect 15284 10984 15293 11024
rect 15907 10984 15916 11024
rect 15956 10984 16876 11024
rect 16916 10984 16925 11024
rect 18499 10984 18508 11024
rect 18548 10984 19564 11024
rect 19604 10984 19613 11024
rect 9571 10983 9629 10984
rect 16867 10983 16925 10984
rect 16675 10940 16733 10941
rect 1987 10900 1996 10940
rect 2036 10900 13324 10940
rect 13364 10900 13373 10940
rect 14275 10900 14284 10940
rect 14324 10900 14668 10940
rect 14708 10900 14717 10940
rect 16675 10900 16684 10940
rect 16724 10900 16876 10940
rect 16916 10900 16925 10940
rect 18595 10900 18604 10940
rect 18644 10900 19660 10940
rect 19700 10900 19709 10940
rect 16675 10899 16733 10900
rect 0 10856 80 10876
rect 547 10856 605 10857
rect 2851 10856 2909 10857
rect 10243 10856 10301 10857
rect 18307 10856 18365 10857
rect 0 10816 556 10856
rect 596 10816 605 10856
rect 1123 10816 1132 10856
rect 1172 10816 2860 10856
rect 2900 10816 2909 10856
rect 3235 10816 3244 10856
rect 3284 10816 4492 10856
rect 4532 10816 4541 10856
rect 5443 10816 5452 10856
rect 5492 10816 6028 10856
rect 6068 10816 6077 10856
rect 10243 10816 10252 10856
rect 10292 10816 11692 10856
rect 11732 10816 11741 10856
rect 14467 10816 14476 10856
rect 14516 10816 18316 10856
rect 18356 10816 18365 10856
rect 0 10796 80 10816
rect 547 10815 605 10816
rect 2851 10815 2909 10816
rect 10243 10815 10301 10816
rect 18307 10815 18365 10816
rect 18499 10856 18557 10857
rect 21424 10856 21504 10876
rect 18499 10816 18508 10856
rect 18548 10816 19084 10856
rect 19124 10816 19133 10856
rect 21091 10816 21100 10856
rect 21140 10816 21504 10856
rect 18499 10815 18557 10816
rect 21424 10796 21504 10816
rect 835 10772 893 10773
rect 2275 10772 2333 10773
rect 4771 10772 4829 10773
rect 9667 10772 9725 10773
rect 835 10732 844 10772
rect 884 10732 2284 10772
rect 2324 10732 2333 10772
rect 4291 10732 4300 10772
rect 4340 10732 4588 10772
rect 4628 10732 4637 10772
rect 4771 10732 4780 10772
rect 4820 10732 8140 10772
rect 8180 10732 8189 10772
rect 9667 10732 9676 10772
rect 9716 10732 10060 10772
rect 10100 10732 11980 10772
rect 12020 10732 12029 10772
rect 13027 10732 13036 10772
rect 13076 10732 14668 10772
rect 14708 10732 16588 10772
rect 16628 10732 17452 10772
rect 17492 10732 17501 10772
rect 18019 10732 18028 10772
rect 18068 10732 20140 10772
rect 20180 10732 20189 10772
rect 835 10731 893 10732
rect 2275 10731 2333 10732
rect 4771 10731 4829 10732
rect 9667 10731 9725 10732
rect 1795 10688 1853 10689
rect 5443 10688 5501 10689
rect 13708 10688 13748 10732
rect 1795 10648 1804 10688
rect 1844 10648 5452 10688
rect 5492 10648 5501 10688
rect 9667 10648 9676 10688
rect 9716 10648 12460 10688
rect 12500 10648 12509 10688
rect 13699 10648 13708 10688
rect 13748 10648 13788 10688
rect 14371 10648 14380 10688
rect 14420 10648 17644 10688
rect 17684 10648 17693 10688
rect 1795 10647 1853 10648
rect 5443 10647 5501 10648
rect 931 10604 989 10605
rect 3427 10604 3485 10605
rect 4291 10604 4349 10605
rect 9475 10604 9533 10605
rect 16099 10604 16157 10605
rect 931 10564 940 10604
rect 980 10564 3436 10604
rect 3476 10564 3485 10604
rect 3679 10564 3688 10604
rect 3728 10564 3770 10604
rect 3810 10564 3852 10604
rect 3892 10564 3934 10604
rect 3974 10564 4016 10604
rect 4056 10564 4065 10604
rect 4291 10564 4300 10604
rect 4340 10564 5836 10604
rect 5876 10564 5885 10604
rect 7843 10564 7852 10604
rect 7892 10564 8620 10604
rect 8660 10564 9484 10604
rect 9524 10564 10252 10604
rect 10292 10564 10301 10604
rect 11875 10564 11884 10604
rect 11924 10564 12940 10604
rect 12980 10564 12989 10604
rect 16099 10564 16108 10604
rect 16148 10564 17164 10604
rect 17204 10564 17213 10604
rect 18799 10564 18808 10604
rect 18848 10564 18890 10604
rect 18930 10564 18972 10604
rect 19012 10564 19054 10604
rect 19094 10564 19136 10604
rect 19176 10564 19185 10604
rect 931 10563 989 10564
rect 3427 10563 3485 10564
rect 4291 10563 4349 10564
rect 9475 10563 9533 10564
rect 16099 10563 16157 10564
rect 0 10520 80 10540
rect 4771 10520 4829 10521
rect 0 10480 4300 10520
rect 4340 10480 4349 10520
rect 4771 10480 4780 10520
rect 4820 10480 7084 10520
rect 7124 10480 7133 10520
rect 8131 10480 8140 10520
rect 8180 10480 16972 10520
rect 17012 10480 17021 10520
rect 19747 10480 19756 10520
rect 19796 10480 20044 10520
rect 20084 10480 20093 10520
rect 0 10460 80 10480
rect 4771 10479 4829 10480
rect 2755 10436 2813 10437
rect 2947 10436 3005 10437
rect 2179 10396 2188 10436
rect 2228 10396 2764 10436
rect 2804 10396 2956 10436
rect 2996 10396 3005 10436
rect 2755 10395 2813 10396
rect 2947 10395 3005 10396
rect 3235 10436 3293 10437
rect 20803 10436 20861 10437
rect 3235 10396 3244 10436
rect 3284 10396 6028 10436
rect 6068 10396 6077 10436
rect 8707 10396 8716 10436
rect 8756 10396 10348 10436
rect 10388 10396 10397 10436
rect 11011 10396 11020 10436
rect 11060 10396 13844 10436
rect 14083 10396 14092 10436
rect 14132 10396 15340 10436
rect 15380 10396 15389 10436
rect 15715 10396 15724 10436
rect 15764 10396 16588 10436
rect 16628 10396 16637 10436
rect 17251 10396 17260 10436
rect 17300 10396 18796 10436
rect 18836 10396 18845 10436
rect 19363 10396 19372 10436
rect 19412 10396 20812 10436
rect 20852 10396 20861 10436
rect 3235 10395 3293 10396
rect 5539 10352 5597 10353
rect 6307 10352 6365 10353
rect 8515 10352 8573 10353
rect 13804 10352 13844 10396
rect 20803 10395 20861 10396
rect 21424 10352 21504 10372
rect 355 10312 364 10352
rect 404 10312 2540 10352
rect 3523 10312 3532 10352
rect 3572 10312 4684 10352
rect 4724 10312 4733 10352
rect 4780 10312 5548 10352
rect 5588 10312 5597 10352
rect 6192 10312 6220 10352
rect 6260 10312 6316 10352
rect 6356 10312 7180 10352
rect 7220 10312 7229 10352
rect 8323 10312 8332 10352
rect 8372 10312 8524 10352
rect 8564 10312 8573 10352
rect 10243 10312 10252 10352
rect 10292 10312 11596 10352
rect 11636 10312 11645 10352
rect 13804 10312 21504 10352
rect 2083 10268 2141 10269
rect 2500 10268 2540 10312
rect 4780 10268 4820 10312
rect 5539 10311 5597 10312
rect 6307 10311 6365 10312
rect 8515 10311 8573 10312
rect 21424 10292 21504 10312
rect 20707 10268 20765 10269
rect 2083 10228 2092 10268
rect 2132 10228 2188 10268
rect 2228 10228 2237 10268
rect 2500 10228 4820 10268
rect 5251 10228 5260 10268
rect 5300 10228 6892 10268
rect 6932 10228 6941 10268
rect 7459 10228 7468 10268
rect 7508 10228 9868 10268
rect 9908 10228 9917 10268
rect 10051 10228 10060 10268
rect 10100 10228 10828 10268
rect 10868 10228 10877 10268
rect 16003 10228 16012 10268
rect 16052 10228 19468 10268
rect 19508 10228 19517 10268
rect 20227 10228 20236 10268
rect 20276 10228 20716 10268
rect 20756 10228 20765 10268
rect 2083 10227 2141 10228
rect 20707 10227 20765 10228
rect 0 10184 80 10204
rect 1507 10184 1565 10185
rect 2275 10184 2333 10185
rect 5443 10184 5501 10185
rect 5923 10184 5981 10185
rect 7555 10184 7613 10185
rect 9955 10184 10013 10185
rect 15811 10184 15869 10185
rect 20611 10184 20669 10185
rect 0 10144 172 10184
rect 212 10144 221 10184
rect 1411 10144 1420 10184
rect 1460 10144 1516 10184
rect 1556 10144 2284 10184
rect 2324 10144 2333 10184
rect 2563 10144 2572 10184
rect 2612 10144 4684 10184
rect 4724 10144 4733 10184
rect 5358 10144 5452 10184
rect 5492 10144 5501 10184
rect 0 10124 80 10144
rect 1507 10143 1565 10144
rect 2275 10143 2333 10144
rect 5443 10143 5501 10144
rect 5548 10144 5932 10184
rect 5972 10144 7564 10184
rect 7604 10144 7613 10184
rect 7939 10144 7948 10184
rect 7988 10144 9772 10184
rect 9812 10144 9821 10184
rect 9955 10144 9964 10184
rect 10004 10144 10098 10184
rect 10243 10144 10252 10184
rect 10292 10144 12364 10184
rect 12404 10144 12413 10184
rect 13123 10144 13132 10184
rect 13172 10144 15052 10184
rect 15092 10144 15101 10184
rect 15811 10144 15820 10184
rect 15860 10144 16724 10184
rect 17059 10144 17068 10184
rect 17108 10144 18028 10184
rect 18068 10144 18077 10184
rect 19075 10144 19084 10184
rect 19124 10144 20620 10184
rect 20660 10144 20669 10184
rect 5548 10100 5588 10144
rect 5923 10143 5981 10144
rect 7555 10143 7613 10144
rect 9955 10143 10013 10144
rect 15811 10143 15869 10144
rect 14755 10100 14813 10101
rect 15235 10100 15293 10101
rect 16003 10100 16061 10101
rect 16579 10100 16637 10101
rect 4483 10060 4492 10100
rect 4532 10060 5588 10100
rect 6211 10060 6220 10100
rect 6260 10060 6604 10100
rect 6644 10060 6653 10100
rect 7267 10060 7276 10100
rect 7316 10060 8812 10100
rect 8852 10060 9004 10100
rect 9044 10060 9053 10100
rect 11587 10060 11596 10100
rect 11636 10060 12748 10100
rect 12788 10060 12797 10100
rect 14668 10060 14764 10100
rect 14804 10060 14813 10100
rect 15139 10060 15148 10100
rect 15188 10060 15244 10100
rect 15284 10060 15293 10100
rect 5827 10016 5885 10017
rect 5635 9976 5644 10016
rect 5684 9976 5836 10016
rect 5876 9976 5885 10016
rect 5827 9975 5885 9976
rect 7459 10016 7517 10017
rect 13603 10016 13661 10017
rect 14668 10016 14708 10060
rect 14755 10059 14813 10060
rect 15235 10059 15293 10060
rect 15340 10060 16012 10100
rect 16052 10060 16061 10100
rect 16483 10060 16492 10100
rect 16532 10060 16588 10100
rect 16628 10060 16637 10100
rect 16684 10100 16724 10144
rect 20611 10143 20669 10144
rect 20995 10100 21053 10101
rect 16684 10060 18220 10100
rect 18260 10060 18269 10100
rect 20035 10060 20044 10100
rect 20084 10060 21004 10100
rect 21044 10060 21053 10100
rect 15340 10016 15380 10060
rect 16003 10059 16061 10060
rect 16579 10059 16637 10060
rect 20995 10059 21053 10060
rect 7459 9976 7468 10016
rect 7508 9976 11404 10016
rect 11444 9976 11453 10016
rect 12067 9976 12076 10016
rect 12116 9976 13228 10016
rect 13268 9976 13277 10016
rect 13518 9976 13612 10016
rect 13652 9976 13661 10016
rect 14659 9976 14668 10016
rect 14708 9976 14717 10016
rect 15331 9976 15340 10016
rect 15380 9976 15389 10016
rect 17260 9976 17452 10016
rect 17492 9976 17501 10016
rect 7459 9975 7517 9976
rect 13603 9975 13661 9976
rect 5731 9932 5789 9933
rect 5923 9932 5981 9933
rect 8707 9932 8765 9933
rect 17155 9932 17213 9933
rect 17260 9932 17300 9976
rect 2275 9892 2284 9932
rect 2324 9892 5684 9932
rect 0 9848 80 9868
rect 5644 9848 5684 9892
rect 5731 9892 5740 9932
rect 5780 9892 5932 9932
rect 5972 9892 5981 9932
rect 8323 9892 8332 9932
rect 8372 9892 8716 9932
rect 8756 9892 8765 9932
rect 10339 9892 10348 9932
rect 10388 9892 14092 9932
rect 14132 9892 14141 9932
rect 15235 9892 15244 9932
rect 15284 9892 17164 9932
rect 17204 9892 17300 9932
rect 5731 9891 5789 9892
rect 5923 9891 5981 9892
rect 8707 9891 8765 9892
rect 17155 9891 17213 9892
rect 11203 9848 11261 9849
rect 13987 9848 14045 9849
rect 21424 9848 21504 9868
rect 0 9808 1996 9848
rect 2036 9808 2045 9848
rect 2371 9808 2380 9848
rect 2420 9808 3052 9848
rect 3092 9808 3101 9848
rect 4919 9808 4928 9848
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 5296 9808 5305 9848
rect 5644 9808 11212 9848
rect 11252 9808 11261 9848
rect 11395 9808 11404 9848
rect 11444 9808 12076 9848
rect 12116 9808 12125 9848
rect 13987 9808 13996 9848
rect 14036 9808 15820 9848
rect 15860 9808 15869 9848
rect 20039 9808 20048 9848
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20416 9808 20425 9848
rect 20812 9808 21504 9848
rect 0 9788 80 9808
rect 11203 9807 11261 9808
rect 13987 9807 14045 9808
rect 8707 9764 8765 9765
rect 9379 9764 9437 9765
rect 11875 9764 11933 9765
rect 20812 9764 20852 9808
rect 21424 9788 21504 9808
rect 1603 9724 1612 9764
rect 1652 9724 8044 9764
rect 8084 9724 8093 9764
rect 8707 9724 8716 9764
rect 8756 9724 8908 9764
rect 8948 9724 8957 9764
rect 9379 9724 9388 9764
rect 9428 9724 11348 9764
rect 11779 9724 11788 9764
rect 11828 9724 11884 9764
rect 11924 9724 11933 9764
rect 14947 9724 14956 9764
rect 14996 9724 15005 9764
rect 16099 9724 16108 9764
rect 16148 9724 20852 9764
rect 8707 9723 8765 9724
rect 9379 9723 9437 9724
rect 2947 9680 3005 9681
rect 7075 9680 7133 9681
rect 2947 9640 2956 9680
rect 2996 9640 7084 9680
rect 7124 9640 7133 9680
rect 11308 9680 11348 9724
rect 11875 9723 11933 9724
rect 11308 9640 11500 9680
rect 11540 9640 11549 9680
rect 2947 9639 3005 9640
rect 7075 9639 7133 9640
rect 14956 9596 14996 9724
rect 16579 9680 16637 9681
rect 20035 9680 20093 9681
rect 15523 9640 15532 9680
rect 15572 9640 15916 9680
rect 15956 9640 15965 9680
rect 16494 9640 16588 9680
rect 16628 9640 16637 9680
rect 16771 9640 16780 9680
rect 16820 9640 17447 9680
rect 17487 9640 17496 9680
rect 17539 9640 17548 9680
rect 17588 9640 17932 9680
rect 17972 9640 17981 9680
rect 19939 9640 19948 9680
rect 19988 9640 20044 9680
rect 20084 9640 20093 9680
rect 16579 9639 16637 9640
rect 20035 9639 20093 9640
rect 2947 9556 2956 9596
rect 2996 9556 3340 9596
rect 3380 9556 3389 9596
rect 4771 9556 4780 9596
rect 4820 9556 12268 9596
rect 12308 9556 12317 9596
rect 14956 9556 20812 9596
rect 20852 9556 20861 9596
rect 0 9512 80 9532
rect 9091 9512 9149 9513
rect 11203 9512 11261 9513
rect 15523 9512 15581 9513
rect 18307 9512 18365 9513
rect 19555 9512 19613 9513
rect 19939 9512 19997 9513
rect 0 9472 844 9512
rect 884 9472 893 9512
rect 1219 9472 1228 9512
rect 1268 9472 2380 9512
rect 2420 9472 2429 9512
rect 2659 9472 2668 9512
rect 2708 9472 4972 9512
rect 5012 9472 5021 9512
rect 5539 9472 5548 9512
rect 5588 9472 5932 9512
rect 5972 9472 5981 9512
rect 7075 9472 7084 9512
rect 7124 9472 8044 9512
rect 8084 9472 8093 9512
rect 9091 9472 9100 9512
rect 9140 9472 9196 9512
rect 9236 9472 9245 9512
rect 9379 9472 9388 9512
rect 9428 9472 10444 9512
rect 10484 9472 10493 9512
rect 11107 9472 11116 9512
rect 11156 9472 11212 9512
rect 11252 9472 11261 9512
rect 13315 9472 13324 9512
rect 13364 9472 13516 9512
rect 13556 9472 13708 9512
rect 13748 9472 13757 9512
rect 14371 9472 14380 9512
rect 14420 9472 14764 9512
rect 14804 9472 14813 9512
rect 15139 9472 15148 9512
rect 15188 9472 15532 9512
rect 15572 9472 15581 9512
rect 16675 9472 16684 9512
rect 16724 9472 17164 9512
rect 17204 9472 17644 9512
rect 17684 9472 17693 9512
rect 18222 9472 18316 9512
rect 18356 9472 18365 9512
rect 18691 9472 18700 9512
rect 18740 9472 19564 9512
rect 19604 9472 19613 9512
rect 19854 9472 19948 9512
rect 19988 9472 19997 9512
rect 20227 9472 20236 9512
rect 20276 9472 20716 9512
rect 20756 9472 20765 9512
rect 0 9452 80 9472
rect 9091 9471 9149 9472
rect 11203 9471 11261 9472
rect 15523 9471 15581 9472
rect 18307 9471 18365 9472
rect 19555 9471 19613 9472
rect 19939 9471 19997 9472
rect 7555 9428 7613 9429
rect 19747 9428 19805 9429
rect 4003 9388 4012 9428
rect 4052 9388 4396 9428
rect 4436 9388 6412 9428
rect 6452 9388 6604 9428
rect 6644 9388 6653 9428
rect 7555 9388 7564 9428
rect 7604 9388 7660 9428
rect 7700 9388 7709 9428
rect 8995 9388 9004 9428
rect 9044 9388 11020 9428
rect 11060 9388 11069 9428
rect 15043 9388 15052 9428
rect 15092 9388 16972 9428
rect 17012 9388 17021 9428
rect 19662 9388 19756 9428
rect 19796 9388 19805 9428
rect 7555 9387 7613 9388
rect 19747 9387 19805 9388
rect 2467 9344 2525 9345
rect 4675 9344 4733 9345
rect 11107 9344 11165 9345
rect 17155 9344 17213 9345
rect 21424 9344 21504 9364
rect 1603 9304 1612 9344
rect 1652 9304 1900 9344
rect 1940 9304 1949 9344
rect 2467 9304 2476 9344
rect 2516 9304 2860 9344
rect 2900 9304 2909 9344
rect 4099 9304 4108 9344
rect 4148 9304 4684 9344
rect 4724 9304 6316 9344
rect 6356 9304 8524 9344
rect 8564 9304 9676 9344
rect 9716 9304 9725 9344
rect 11022 9304 11116 9344
rect 11156 9304 11165 9344
rect 2467 9303 2525 9304
rect 4675 9303 4733 9304
rect 11107 9303 11165 9304
rect 11212 9304 15244 9344
rect 15284 9304 15293 9344
rect 15532 9304 17164 9344
rect 17204 9304 21504 9344
rect 5923 9260 5981 9261
rect 6691 9260 6749 9261
rect 9091 9260 9149 9261
rect 11212 9260 11252 9304
rect 15532 9260 15572 9304
rect 17155 9303 17213 9304
rect 21424 9284 21504 9304
rect 1411 9220 1420 9260
rect 1460 9220 3436 9260
rect 3476 9220 3485 9260
rect 3907 9220 3916 9260
rect 3956 9220 5932 9260
rect 5972 9220 6412 9260
rect 6452 9220 6461 9260
rect 6691 9220 6700 9260
rect 6740 9220 6988 9260
rect 7028 9220 7037 9260
rect 9091 9220 9100 9260
rect 9140 9220 11252 9260
rect 13795 9220 13804 9260
rect 13844 9220 15532 9260
rect 15572 9220 15581 9260
rect 15715 9220 15724 9260
rect 15764 9220 17452 9260
rect 17492 9220 17501 9260
rect 20227 9220 20236 9260
rect 20276 9220 20620 9260
rect 20660 9220 20669 9260
rect 5923 9219 5981 9220
rect 6691 9219 6749 9220
rect 9091 9219 9149 9220
rect 0 9176 80 9196
rect 10051 9176 10109 9177
rect 0 9136 10060 9176
rect 10100 9136 10109 9176
rect 0 9116 80 9136
rect 10051 9135 10109 9136
rect 10435 9176 10493 9177
rect 14467 9176 14525 9177
rect 10435 9136 10444 9176
rect 10484 9136 11020 9176
rect 11060 9136 11069 9176
rect 13699 9136 13708 9176
rect 13748 9136 14476 9176
rect 14516 9136 14525 9176
rect 10435 9135 10493 9136
rect 14467 9135 14525 9136
rect 15139 9176 15197 9177
rect 19267 9176 19325 9177
rect 15139 9136 15148 9176
rect 15188 9136 19276 9176
rect 19316 9136 19325 9176
rect 19459 9136 19468 9176
rect 19508 9136 20140 9176
rect 20180 9136 20189 9176
rect 15139 9135 15197 9136
rect 19267 9135 19325 9136
rect 4963 9092 5021 9093
rect 1795 9052 1804 9092
rect 1844 9052 1853 9092
rect 3679 9052 3688 9092
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 4056 9052 4065 9092
rect 4483 9052 4492 9092
rect 4532 9052 4972 9092
rect 5012 9052 5021 9092
rect 6307 9052 6316 9092
rect 6356 9052 6604 9092
rect 6644 9052 6653 9092
rect 6700 9052 8852 9092
rect 8899 9052 8908 9092
rect 8948 9052 13036 9092
rect 13076 9052 13085 9092
rect 18799 9052 18808 9092
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 19176 9052 19185 9092
rect 1804 9008 1844 9052
rect 4963 9051 5021 9052
rect 4291 9008 4349 9009
rect 6700 9008 6740 9052
rect 172 8968 1844 9008
rect 3331 8968 3340 9008
rect 3380 8968 4300 9008
rect 4340 8968 4349 9008
rect 6499 8968 6508 9008
rect 6548 8968 6740 9008
rect 6787 8968 6796 9008
rect 6836 8968 7468 9008
rect 7508 8968 7517 9008
rect 8707 8968 8716 9008
rect 8756 8968 8765 9008
rect 0 8840 80 8860
rect 172 8840 212 8968
rect 4291 8967 4349 8968
rect 1507 8924 1565 8925
rect 1507 8884 1516 8924
rect 1556 8884 3244 8924
rect 3284 8884 3293 8924
rect 1507 8883 1565 8884
rect 0 8800 212 8840
rect 451 8800 460 8840
rect 500 8800 1228 8840
rect 1268 8800 1277 8840
rect 1322 8800 1331 8840
rect 1371 8800 2284 8840
rect 2324 8800 2333 8840
rect 2500 8800 4780 8840
rect 4820 8800 4829 8840
rect 0 8780 80 8800
rect 1795 8756 1853 8757
rect 1411 8716 1420 8756
rect 1460 8716 1469 8756
rect 1710 8716 1804 8756
rect 1844 8716 1853 8756
rect 1420 8672 1460 8716
rect 1795 8715 1853 8716
rect 2500 8672 2540 8800
rect 8716 8756 8756 8968
rect 8812 8924 8852 9052
rect 10627 9008 10685 9009
rect 12547 9008 12605 9009
rect 9283 8968 9292 9008
rect 9332 8968 9580 9008
rect 9620 8968 9629 9008
rect 10627 8968 10636 9008
rect 10676 8968 11308 9008
rect 11348 8968 11357 9008
rect 12462 8968 12556 9008
rect 12596 8968 12605 9008
rect 10627 8967 10685 8968
rect 12547 8967 12605 8968
rect 12739 9008 12797 9009
rect 12739 8968 12748 9008
rect 12788 8968 13516 9008
rect 13556 8968 13565 9008
rect 19747 8968 19756 9008
rect 19796 8968 20127 9008
rect 20167 8968 20176 9008
rect 12739 8967 12797 8968
rect 8812 8884 12172 8924
rect 12212 8884 20180 8924
rect 10339 8840 10397 8841
rect 14947 8840 15005 8841
rect 16387 8840 16445 8841
rect 19747 8840 19805 8841
rect 10254 8800 10348 8840
rect 10388 8800 10397 8840
rect 11107 8800 11116 8840
rect 11156 8800 13036 8840
rect 13076 8800 13085 8840
rect 14947 8800 14956 8840
rect 14996 8800 15092 8840
rect 15619 8800 15628 8840
rect 15668 8800 16396 8840
rect 16436 8800 16445 8840
rect 17059 8800 17068 8840
rect 17108 8800 17117 8840
rect 17251 8800 17260 8840
rect 17300 8800 17836 8840
rect 17876 8800 17885 8840
rect 18019 8800 18028 8840
rect 18068 8800 19180 8840
rect 19220 8800 19468 8840
rect 19508 8800 19517 8840
rect 19662 8800 19756 8840
rect 19796 8800 19805 8840
rect 20140 8840 20180 8884
rect 21424 8840 21504 8860
rect 20140 8800 21504 8840
rect 10339 8799 10397 8800
rect 14947 8799 15005 8800
rect 15052 8756 15092 8800
rect 16387 8799 16445 8800
rect 16963 8756 17021 8757
rect 17068 8756 17108 8800
rect 19747 8799 19805 8800
rect 21424 8780 21504 8800
rect 3811 8716 3820 8756
rect 3860 8716 8756 8756
rect 9484 8716 10580 8756
rect 10627 8716 10636 8756
rect 10676 8716 10828 8756
rect 10868 8716 10877 8756
rect 11500 8716 11884 8756
rect 11924 8716 11933 8756
rect 13411 8716 13420 8756
rect 13460 8716 13469 8756
rect 14563 8716 14572 8756
rect 14612 8716 14860 8756
rect 14900 8716 14909 8756
rect 15043 8716 15052 8756
rect 15092 8716 15101 8756
rect 15907 8716 15916 8756
rect 15956 8716 16108 8756
rect 16148 8716 16157 8756
rect 16963 8716 16972 8756
rect 17012 8716 17108 8756
rect 17443 8716 17452 8756
rect 17492 8716 19852 8756
rect 19892 8716 19901 8756
rect 9484 8672 9524 8716
rect 1420 8632 2540 8672
rect 3139 8632 3148 8672
rect 3188 8632 5068 8672
rect 5108 8632 5117 8672
rect 5347 8632 5356 8672
rect 5396 8632 6124 8672
rect 6164 8632 6173 8672
rect 6691 8632 6700 8672
rect 6740 8632 7180 8672
rect 7220 8632 7229 8672
rect 8812 8657 9524 8672
rect 5068 8588 5108 8632
rect 8803 8617 8812 8657
rect 8852 8632 9524 8657
rect 9571 8672 9629 8673
rect 10540 8672 10580 8716
rect 11500 8672 11540 8716
rect 13420 8672 13460 8716
rect 16963 8715 17021 8716
rect 19459 8672 19517 8673
rect 19747 8672 19805 8673
rect 9571 8632 9580 8672
rect 9620 8632 9868 8672
rect 9908 8632 9917 8672
rect 10540 8632 11540 8672
rect 11587 8632 11596 8672
rect 11636 8632 13132 8672
rect 13172 8632 13181 8672
rect 13420 8632 16300 8672
rect 16340 8632 16349 8672
rect 16396 8632 16820 8672
rect 16867 8632 16876 8672
rect 16916 8632 17356 8672
rect 17396 8632 17405 8672
rect 18307 8632 18316 8672
rect 18356 8632 18604 8672
rect 18644 8632 18653 8672
rect 19374 8632 19468 8672
rect 19508 8632 19517 8672
rect 19651 8632 19660 8672
rect 19700 8632 19756 8672
rect 19796 8632 19805 8672
rect 8852 8617 8861 8632
rect 9571 8631 9629 8632
rect 12259 8588 12317 8589
rect 13891 8588 13949 8589
rect 16396 8588 16436 8632
rect 16579 8588 16637 8589
rect 2563 8548 2572 8588
rect 2612 8548 3244 8588
rect 3284 8548 3293 8588
rect 5068 8548 8716 8588
rect 8756 8548 8765 8588
rect 10531 8548 10540 8588
rect 10580 8548 11348 8588
rect 12174 8548 12268 8588
rect 12308 8548 12317 8588
rect 12547 8548 12556 8588
rect 12596 8548 12748 8588
rect 12788 8548 12797 8588
rect 13891 8548 13900 8588
rect 13940 8548 15436 8588
rect 15476 8548 15485 8588
rect 15820 8548 16436 8588
rect 16483 8548 16492 8588
rect 16532 8548 16588 8588
rect 16628 8548 16637 8588
rect 16780 8588 16820 8632
rect 19459 8631 19517 8632
rect 19747 8631 19805 8632
rect 18499 8588 18557 8589
rect 16780 8548 16972 8588
rect 17012 8548 18508 8588
rect 18548 8548 18557 8588
rect 0 8504 80 8524
rect 11308 8504 11348 8548
rect 12259 8547 12317 8548
rect 13891 8547 13949 8548
rect 13795 8504 13853 8505
rect 15820 8504 15860 8548
rect 16579 8547 16637 8548
rect 18499 8547 18557 8548
rect 0 8464 1516 8504
rect 1556 8464 1565 8504
rect 2947 8464 2956 8504
rect 2996 8464 10252 8504
rect 10292 8464 11020 8504
rect 11060 8464 11069 8504
rect 11299 8464 11308 8504
rect 11348 8464 11357 8504
rect 13219 8464 13228 8504
rect 13268 8464 13277 8504
rect 13795 8464 13804 8504
rect 13844 8464 15860 8504
rect 15907 8464 15916 8504
rect 15956 8464 17932 8504
rect 17972 8464 17981 8504
rect 19363 8464 19372 8504
rect 19412 8464 20127 8504
rect 20167 8464 20176 8504
rect 20227 8464 20236 8504
rect 20276 8464 20716 8504
rect 20756 8464 20765 8504
rect 0 8444 80 8464
rect 5923 8420 5981 8421
rect 3523 8380 3532 8420
rect 3572 8380 5932 8420
rect 5972 8380 5981 8420
rect 5923 8379 5981 8380
rect 6115 8420 6173 8421
rect 13228 8420 13268 8464
rect 13795 8463 13853 8464
rect 20899 8420 20957 8421
rect 6115 8380 6124 8420
rect 6164 8380 13268 8420
rect 15619 8380 15628 8420
rect 15668 8380 16012 8420
rect 16052 8380 17836 8420
rect 17876 8380 17885 8420
rect 19564 8380 20908 8420
rect 20948 8380 20957 8420
rect 6115 8379 6173 8380
rect 2755 8336 2813 8337
rect 4195 8336 4253 8337
rect 7555 8336 7613 8337
rect 12355 8336 12413 8337
rect 2755 8296 2764 8336
rect 2804 8296 2860 8336
rect 2900 8296 2909 8336
rect 3043 8296 3052 8336
rect 3092 8296 4204 8336
rect 4244 8296 4300 8336
rect 4340 8296 4349 8336
rect 4919 8296 4928 8336
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 5296 8296 5305 8336
rect 7555 8296 7564 8336
rect 7604 8296 12364 8336
rect 12404 8296 12413 8336
rect 2755 8295 2813 8296
rect 4195 8295 4253 8296
rect 7555 8295 7613 8296
rect 12355 8295 12413 8296
rect 16387 8336 16445 8337
rect 17635 8336 17693 8337
rect 19564 8336 19604 8380
rect 20899 8379 20957 8380
rect 21424 8336 21504 8356
rect 16387 8296 16396 8336
rect 16436 8296 16492 8336
rect 16532 8296 16541 8336
rect 17251 8296 17260 8336
rect 17300 8296 17452 8336
rect 17492 8296 17501 8336
rect 17550 8296 17644 8336
rect 17684 8296 17693 8336
rect 19267 8296 19276 8336
rect 19316 8296 19604 8336
rect 20039 8296 20048 8336
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20416 8296 20425 8336
rect 20995 8296 21004 8336
rect 21044 8296 21504 8336
rect 16387 8295 16445 8296
rect 17635 8295 17693 8296
rect 21424 8276 21504 8296
rect 5923 8252 5981 8253
rect 5443 8212 5452 8252
rect 5492 8212 5740 8252
rect 5780 8212 5789 8252
rect 5923 8212 5932 8252
rect 5972 8212 9676 8252
rect 9716 8212 9725 8252
rect 13132 8212 13324 8252
rect 13364 8212 13373 8252
rect 16003 8212 16012 8252
rect 16052 8212 18220 8252
rect 18260 8212 18269 8252
rect 5923 8211 5981 8212
rect 0 8168 80 8188
rect 7843 8168 7901 8169
rect 9475 8168 9533 8169
rect 0 8128 1996 8168
rect 2036 8128 2045 8168
rect 2755 8128 2764 8168
rect 2804 8128 3052 8168
rect 3092 8128 3101 8168
rect 3907 8128 3916 8168
rect 3956 8128 4204 8168
rect 4244 8128 4253 8168
rect 5251 8128 5260 8168
rect 5300 8128 5548 8168
rect 5588 8128 6604 8168
rect 6644 8128 6653 8168
rect 7843 8128 7852 8168
rect 7892 8128 8428 8168
rect 8468 8128 9484 8168
rect 9524 8128 9533 8168
rect 0 8108 80 8128
rect 7843 8127 7901 8128
rect 9475 8127 9533 8128
rect 9667 8168 9725 8169
rect 9667 8128 9676 8168
rect 9716 8128 9964 8168
rect 10004 8128 10013 8168
rect 10915 8128 10924 8168
rect 10964 8128 12556 8168
rect 12596 8128 12605 8168
rect 9667 8127 9725 8128
rect 12259 8084 12317 8085
rect 13132 8084 13172 8212
rect 13795 8168 13853 8169
rect 13219 8128 13228 8168
rect 13268 8128 13804 8168
rect 13844 8128 13853 8168
rect 13795 8127 13853 8128
rect 16963 8168 17021 8169
rect 19939 8168 19997 8169
rect 16963 8128 16972 8168
rect 17012 8128 17164 8168
rect 17204 8128 17213 8168
rect 17539 8128 17548 8168
rect 17588 8128 18028 8168
rect 18068 8128 18077 8168
rect 18883 8128 18892 8168
rect 18932 8128 19276 8168
rect 19316 8128 19325 8168
rect 19939 8128 19948 8168
rect 19988 8128 20140 8168
rect 20180 8128 20189 8168
rect 16963 8127 17021 8128
rect 19939 8127 19997 8128
rect 17827 8084 17885 8085
rect 2500 8044 11884 8084
rect 11924 8044 11933 8084
rect 12163 8044 12172 8084
rect 12212 8044 12268 8084
rect 12308 8044 13172 8084
rect 14755 8044 14764 8084
rect 14804 8044 16684 8084
rect 16724 8044 16733 8084
rect 16780 8044 16972 8084
rect 17012 8044 17836 8084
rect 17876 8044 17885 8084
rect 1603 8000 1661 8001
rect 1518 7960 1612 8000
rect 1652 7960 1661 8000
rect 1603 7959 1661 7960
rect 2500 7916 2540 8044
rect 12259 8043 12317 8044
rect 4675 8000 4733 8001
rect 5443 8000 5501 8001
rect 10339 8000 10397 8001
rect 13219 8000 13277 8001
rect 16780 8000 16820 8044
rect 17827 8043 17885 8044
rect 18595 8084 18653 8085
rect 18595 8044 18604 8084
rect 18644 8044 18796 8084
rect 18836 8044 19852 8084
rect 19892 8044 19901 8084
rect 18595 8043 18653 8044
rect 19459 8000 19517 8001
rect 2947 7960 2956 8000
rect 2996 7960 4684 8000
rect 4724 7960 5068 8000
rect 5108 7960 5117 8000
rect 5358 7960 5452 8000
rect 5492 7960 5501 8000
rect 7171 7960 7180 8000
rect 7220 7960 9100 8000
rect 9140 7960 9149 8000
rect 10339 7960 10348 8000
rect 10388 7960 10444 8000
rect 10484 7960 10493 8000
rect 11395 7960 11404 8000
rect 11444 7960 12844 8000
rect 12884 7960 12893 8000
rect 13219 7960 13228 8000
rect 13268 7960 13324 8000
rect 13364 7960 13373 8000
rect 16195 7960 16204 8000
rect 16244 7960 16820 8000
rect 16867 7960 16876 8000
rect 16916 7960 17068 8000
rect 17108 7960 17644 8000
rect 17684 7960 17693 8000
rect 17923 7960 17932 8000
rect 17972 7960 18604 8000
rect 18644 7960 18653 8000
rect 19374 7960 19468 8000
rect 19508 7960 19517 8000
rect 4675 7959 4733 7960
rect 5068 7916 5108 7960
rect 5443 7959 5501 7960
rect 10339 7959 10397 7960
rect 13219 7959 13277 7960
rect 19459 7959 19517 7960
rect 8707 7916 8765 7917
rect 9475 7916 9533 7917
rect 10915 7916 10973 7917
rect 11683 7916 11741 7917
rect 14755 7916 14813 7917
rect 2179 7876 2188 7916
rect 2228 7876 2540 7916
rect 2755 7876 2764 7916
rect 2804 7876 4012 7916
rect 4052 7876 4061 7916
rect 5068 7876 5836 7916
rect 5876 7876 6700 7916
rect 6740 7876 6749 7916
rect 6883 7876 6892 7916
rect 6932 7876 7220 7916
rect 0 7832 80 7852
rect 163 7832 221 7833
rect 7180 7832 7220 7876
rect 8707 7876 8716 7916
rect 8756 7876 9196 7916
rect 9236 7876 9245 7916
rect 9390 7876 9484 7916
rect 9524 7876 9533 7916
rect 10830 7876 10924 7916
rect 10964 7876 11692 7916
rect 11732 7876 11741 7916
rect 12259 7876 12268 7916
rect 12308 7876 12556 7916
rect 12596 7876 12605 7916
rect 14659 7876 14668 7916
rect 14708 7876 14764 7916
rect 14804 7876 14813 7916
rect 8707 7875 8765 7876
rect 9196 7832 9236 7876
rect 9475 7875 9533 7876
rect 10915 7875 10973 7876
rect 11683 7875 11741 7876
rect 14755 7875 14813 7876
rect 21424 7832 21504 7852
rect 0 7792 172 7832
rect 212 7792 221 7832
rect 7171 7792 7180 7832
rect 7220 7792 7229 7832
rect 9196 7792 11060 7832
rect 13603 7792 13612 7832
rect 13652 7792 15340 7832
rect 15380 7792 15389 7832
rect 21004 7792 21504 7832
rect 0 7772 80 7792
rect 163 7791 221 7792
rect 8803 7748 8861 7749
rect 11020 7748 11060 7792
rect 16579 7748 16637 7749
rect 6115 7708 6124 7748
rect 6164 7708 8812 7748
rect 8852 7708 8861 7748
rect 8995 7708 9004 7748
rect 9044 7708 9772 7748
rect 9812 7708 9821 7748
rect 10147 7708 10156 7748
rect 10196 7708 10636 7748
rect 10676 7708 10685 7748
rect 11020 7708 11156 7748
rect 14563 7708 14572 7748
rect 14612 7708 14956 7748
rect 14996 7708 16588 7748
rect 16628 7708 16637 7748
rect 17635 7708 17644 7748
rect 17684 7708 20908 7748
rect 20948 7708 20957 7748
rect 8803 7707 8861 7708
rect 11116 7664 11156 7708
rect 16579 7707 16637 7708
rect 21004 7664 21044 7792
rect 21424 7772 21504 7792
rect 3523 7624 3532 7664
rect 3572 7624 11020 7664
rect 11060 7624 11069 7664
rect 11116 7624 18220 7664
rect 18260 7624 18269 7664
rect 18316 7624 21044 7664
rect 2371 7580 2429 7581
rect 4579 7580 4637 7581
rect 6691 7580 6749 7581
rect 7459 7580 7517 7581
rect 9379 7580 9437 7581
rect 547 7540 556 7580
rect 596 7540 2380 7580
rect 2420 7540 2429 7580
rect 3679 7540 3688 7580
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 4056 7540 4065 7580
rect 4579 7540 4588 7580
rect 4628 7540 5780 7580
rect 5827 7540 5836 7580
rect 5876 7540 6700 7580
rect 6740 7540 7468 7580
rect 7508 7540 7517 7580
rect 8803 7540 8812 7580
rect 8852 7540 9388 7580
rect 9428 7540 9437 7580
rect 2371 7539 2429 7540
rect 4579 7539 4637 7540
rect 0 7496 80 7516
rect 5635 7496 5693 7497
rect 0 7456 748 7496
rect 788 7456 797 7496
rect 1411 7456 1420 7496
rect 1460 7456 5644 7496
rect 5684 7456 5693 7496
rect 0 7436 80 7456
rect 5635 7455 5693 7456
rect 5740 7412 5780 7540
rect 6691 7539 6749 7540
rect 7459 7539 7517 7540
rect 9379 7539 9437 7540
rect 11011 7580 11069 7581
rect 11011 7540 11020 7580
rect 11060 7540 11500 7580
rect 11540 7540 11549 7580
rect 11779 7540 11788 7580
rect 11828 7540 15052 7580
rect 15092 7540 15101 7580
rect 16483 7540 16492 7580
rect 16532 7540 17068 7580
rect 17108 7540 18068 7580
rect 11011 7539 11069 7540
rect 8899 7496 8957 7497
rect 16483 7496 16541 7497
rect 16771 7496 16829 7497
rect 18028 7496 18068 7540
rect 18316 7496 18356 7624
rect 19843 7580 19901 7581
rect 18595 7540 18604 7580
rect 18644 7540 18740 7580
rect 18799 7540 18808 7580
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 19176 7540 19185 7580
rect 19651 7540 19660 7580
rect 19700 7540 19852 7580
rect 19892 7540 19901 7580
rect 6787 7456 6796 7496
rect 6836 7456 7276 7496
rect 7316 7456 7325 7496
rect 7372 7456 8852 7496
rect 7372 7412 7412 7456
rect 8812 7412 8852 7456
rect 8899 7456 8908 7496
rect 8948 7456 11980 7496
rect 12020 7456 12029 7496
rect 14083 7456 14092 7496
rect 14132 7456 14380 7496
rect 14420 7456 14429 7496
rect 14755 7456 14764 7496
rect 14804 7456 15148 7496
rect 15188 7456 15197 7496
rect 16483 7456 16492 7496
rect 16532 7456 16684 7496
rect 16724 7456 16780 7496
rect 16820 7456 16848 7496
rect 18028 7456 18356 7496
rect 8899 7455 8957 7456
rect 16483 7455 16541 7456
rect 16771 7455 16829 7456
rect 13795 7412 13853 7413
rect 14275 7412 14333 7413
rect 4099 7372 4108 7412
rect 4148 7372 5164 7412
rect 5204 7372 5213 7412
rect 5740 7372 7412 7412
rect 8131 7372 8140 7412
rect 8180 7372 8716 7412
rect 8756 7372 8765 7412
rect 8812 7372 10924 7412
rect 10964 7372 10973 7412
rect 11491 7372 11500 7412
rect 11540 7372 13804 7412
rect 13844 7372 13853 7412
rect 14190 7372 14284 7412
rect 14324 7372 14333 7412
rect 13795 7371 13853 7372
rect 14275 7371 14333 7372
rect 15811 7412 15869 7413
rect 16387 7412 16445 7413
rect 15811 7372 15820 7412
rect 15860 7372 16108 7412
rect 16148 7372 16157 7412
rect 16387 7372 16396 7412
rect 16436 7372 16588 7412
rect 16628 7372 16637 7412
rect 15811 7371 15869 7372
rect 16387 7371 16445 7372
rect 6115 7328 6173 7329
rect 6499 7328 6557 7329
rect 172 7288 6124 7328
rect 6164 7288 6173 7328
rect 6414 7288 6508 7328
rect 6548 7288 6557 7328
rect 6691 7288 6700 7328
rect 6740 7288 11212 7328
rect 11252 7288 11261 7328
rect 12739 7288 12748 7328
rect 12788 7288 13516 7328
rect 13556 7288 17932 7328
rect 17972 7288 17981 7328
rect 0 7160 80 7180
rect 172 7160 212 7288
rect 6115 7287 6173 7288
rect 6499 7287 6557 7288
rect 3043 7244 3101 7245
rect 17155 7244 17213 7245
rect 18700 7244 18740 7540
rect 19843 7539 19901 7540
rect 19459 7456 19468 7496
rect 19508 7456 19988 7496
rect 19948 7413 19988 7456
rect 18883 7412 18941 7413
rect 19939 7412 19997 7413
rect 18883 7372 18892 7412
rect 18932 7372 19660 7412
rect 19700 7372 19709 7412
rect 19939 7372 19948 7412
rect 19988 7372 20140 7412
rect 20180 7372 20189 7412
rect 18883 7371 18941 7372
rect 19939 7371 19997 7372
rect 20803 7328 20861 7329
rect 21424 7328 21504 7348
rect 18883 7288 18892 7328
rect 18932 7288 20812 7328
rect 20852 7288 20861 7328
rect 20803 7287 20861 7288
rect 21292 7288 21504 7328
rect 3043 7204 3052 7244
rect 3092 7204 3532 7244
rect 3572 7204 3581 7244
rect 5155 7204 5164 7244
rect 5204 7204 7852 7244
rect 7892 7204 7901 7244
rect 8236 7204 9676 7244
rect 9716 7204 9725 7244
rect 10339 7204 10348 7244
rect 10388 7204 10636 7244
rect 10676 7204 10685 7244
rect 14467 7204 14476 7244
rect 14516 7204 16108 7244
rect 16148 7204 16157 7244
rect 17155 7204 17164 7244
rect 17204 7204 17548 7244
rect 17588 7204 17597 7244
rect 18700 7204 18988 7244
rect 19028 7204 19037 7244
rect 3043 7203 3101 7204
rect 8236 7160 8276 7204
rect 17155 7203 17213 7204
rect 8707 7160 8765 7161
rect 21292 7160 21332 7288
rect 21424 7268 21504 7288
rect 0 7120 212 7160
rect 1315 7120 1324 7160
rect 1364 7120 2092 7160
rect 2132 7120 2141 7160
rect 4963 7120 4972 7160
rect 5012 7120 5356 7160
rect 5396 7120 5405 7160
rect 5923 7120 5932 7160
rect 5972 7120 6700 7160
rect 6740 7120 6749 7160
rect 6796 7120 7468 7160
rect 7508 7120 7517 7160
rect 7651 7120 7660 7160
rect 7700 7120 8276 7160
rect 8622 7120 8716 7160
rect 8756 7120 8765 7160
rect 14275 7120 14284 7160
rect 14324 7120 18604 7160
rect 18644 7120 18653 7160
rect 19075 7120 19084 7160
rect 19124 7120 19948 7160
rect 19988 7120 19997 7160
rect 20227 7120 20236 7160
rect 20276 7120 20812 7160
rect 20852 7120 20861 7160
rect 21292 7120 21484 7160
rect 0 7100 80 7120
rect 6115 7076 6173 7077
rect 6796 7076 6836 7120
rect 8707 7119 8765 7120
rect 12643 7076 12701 7077
rect 172 7036 5644 7076
rect 5684 7036 5693 7076
rect 6019 7036 6028 7076
rect 6068 7036 6124 7076
rect 6164 7036 6173 7076
rect 6307 7036 6316 7076
rect 6356 7036 6836 7076
rect 7363 7036 7372 7076
rect 7412 7036 9292 7076
rect 9332 7036 9580 7076
rect 9620 7036 9629 7076
rect 12643 7036 12652 7076
rect 12692 7036 13996 7076
rect 14036 7036 14045 7076
rect 14476 7036 19564 7076
rect 19604 7036 19613 7076
rect 0 6824 80 6844
rect 0 6764 116 6824
rect 76 6740 116 6764
rect 172 6740 212 7036
rect 6115 7035 6173 7036
rect 12643 7035 12701 7036
rect 739 6992 797 6993
rect 5443 6992 5501 6993
rect 739 6952 748 6992
rect 788 6952 844 6992
rect 884 6952 893 6992
rect 1315 6952 1324 6992
rect 1364 6952 1900 6992
rect 1940 6952 1949 6992
rect 2563 6952 2572 6992
rect 2612 6952 2860 6992
rect 2900 6952 2909 6992
rect 5358 6952 5452 6992
rect 5492 6952 5501 6992
rect 739 6951 797 6952
rect 5443 6951 5501 6952
rect 5827 6992 5885 6993
rect 9379 6992 9437 6993
rect 14083 6992 14141 6993
rect 14476 6992 14516 7036
rect 19363 6992 19421 6993
rect 21444 6992 21484 7120
rect 5827 6952 5836 6992
rect 5876 6952 8428 6992
rect 8468 6952 8477 6992
rect 8707 6952 8716 6992
rect 8756 6952 9004 6992
rect 9044 6952 9053 6992
rect 9294 6952 9388 6992
rect 9428 6952 9437 6992
rect 13998 6952 14092 6992
rect 14132 6952 14141 6992
rect 14467 6952 14476 6992
rect 14516 6952 14525 6992
rect 16291 6952 16300 6992
rect 16340 6952 16349 6992
rect 16963 6952 16972 6992
rect 17012 6952 19372 6992
rect 19412 6952 21484 6992
rect 5827 6951 5885 6952
rect 9379 6951 9437 6952
rect 14083 6951 14141 6952
rect 6211 6908 6269 6909
rect 1795 6868 1804 6908
rect 1844 6868 6220 6908
rect 6260 6868 6269 6908
rect 6211 6867 6269 6868
rect 6691 6908 6749 6909
rect 7651 6908 7709 6909
rect 16300 6908 16340 6952
rect 19363 6951 19421 6952
rect 6691 6868 6700 6908
rect 6740 6868 7660 6908
rect 7700 6868 7709 6908
rect 9091 6868 9100 6908
rect 9140 6868 11500 6908
rect 11540 6868 11549 6908
rect 16300 6868 19468 6908
rect 19508 6868 19517 6908
rect 19651 6868 19660 6908
rect 19700 6868 20908 6908
rect 20948 6868 20957 6908
rect 6691 6867 6749 6868
rect 7651 6867 7709 6868
rect 6307 6824 6365 6825
rect 15715 6824 15773 6825
rect 19843 6824 19901 6825
rect 21424 6824 21504 6844
rect 1891 6784 1900 6824
rect 1940 6784 4780 6824
rect 4820 6784 4829 6824
rect 4919 6784 4928 6824
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 5296 6784 5305 6824
rect 5539 6784 5548 6824
rect 5588 6784 6316 6824
rect 6356 6784 6365 6824
rect 6499 6784 6508 6824
rect 6548 6784 7084 6824
rect 7124 6784 7133 6824
rect 7459 6784 7468 6824
rect 7508 6784 9004 6824
rect 9044 6784 15724 6824
rect 15764 6784 15773 6824
rect 16099 6784 16108 6824
rect 16148 6784 19852 6824
rect 19892 6784 19901 6824
rect 20039 6784 20048 6824
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20416 6784 20425 6824
rect 21004 6784 21504 6824
rect 6307 6783 6365 6784
rect 15715 6783 15773 6784
rect 19843 6783 19901 6784
rect 6499 6740 6557 6741
rect 12355 6740 12413 6741
rect 16675 6740 16733 6741
rect 18403 6740 18461 6741
rect 76 6700 212 6740
rect 1708 6700 1996 6740
rect 2036 6700 2045 6740
rect 5635 6700 5644 6740
rect 5684 6700 6316 6740
rect 6356 6700 6365 6740
rect 6499 6700 6508 6740
rect 6548 6700 7372 6740
rect 7412 6700 7421 6740
rect 7555 6700 7564 6740
rect 7604 6700 8140 6740
rect 8180 6700 8189 6740
rect 8323 6700 8332 6740
rect 8372 6700 10348 6740
rect 10388 6700 10397 6740
rect 12355 6700 12364 6740
rect 12404 6700 16684 6740
rect 16724 6700 16733 6740
rect 17539 6700 17548 6740
rect 17588 6700 17597 6740
rect 18318 6700 18412 6740
rect 18452 6700 18461 6740
rect 0 6488 80 6508
rect 1507 6488 1565 6489
rect 0 6448 652 6488
rect 692 6448 701 6488
rect 1422 6448 1516 6488
rect 1556 6448 1565 6488
rect 0 6428 80 6448
rect 1507 6447 1565 6448
rect 1708 6320 1748 6700
rect 6499 6699 6557 6700
rect 12355 6699 12413 6700
rect 16675 6699 16733 6700
rect 2179 6656 2237 6657
rect 2755 6656 2813 6657
rect 3139 6656 3197 6657
rect 9475 6656 9533 6657
rect 2083 6616 2092 6656
rect 2132 6616 2188 6656
rect 2228 6616 2237 6656
rect 2670 6616 2764 6656
rect 2804 6616 3148 6656
rect 3188 6616 3197 6656
rect 4195 6616 4204 6656
rect 4244 6616 4588 6656
rect 4628 6616 4637 6656
rect 5059 6616 5068 6656
rect 5108 6616 5836 6656
rect 5876 6616 5885 6656
rect 6403 6616 6412 6656
rect 6452 6616 7028 6656
rect 7267 6616 7276 6656
rect 7316 6616 8236 6656
rect 8276 6616 8285 6656
rect 9283 6616 9292 6656
rect 9332 6616 9484 6656
rect 9524 6616 9533 6656
rect 2179 6615 2237 6616
rect 2755 6615 2813 6616
rect 3139 6615 3197 6616
rect 6988 6572 7028 6616
rect 9475 6615 9533 6616
rect 10051 6656 10109 6657
rect 17548 6656 17588 6700
rect 18403 6699 18461 6700
rect 18883 6740 18941 6741
rect 21004 6740 21044 6784
rect 21424 6764 21504 6784
rect 18883 6700 18892 6740
rect 18932 6700 21044 6740
rect 18883 6699 18941 6700
rect 10051 6616 10060 6656
rect 10100 6616 12076 6656
rect 12116 6616 12125 6656
rect 12835 6616 12844 6656
rect 12884 6616 16204 6656
rect 16244 6616 16253 6656
rect 17548 6616 18452 6656
rect 18499 6616 18508 6656
rect 18548 6616 20236 6656
rect 20276 6616 20285 6656
rect 10051 6615 10109 6616
rect 11683 6572 11741 6573
rect 18412 6572 18452 6616
rect 2500 6532 4396 6572
rect 4436 6532 4445 6572
rect 4675 6532 4684 6572
rect 4724 6532 6892 6572
rect 6932 6532 6941 6572
rect 6988 6532 7412 6572
rect 7459 6532 7468 6572
rect 7508 6532 7948 6572
rect 7988 6532 7997 6572
rect 8803 6532 8812 6572
rect 8852 6532 9100 6572
rect 9140 6532 9149 6572
rect 11683 6532 11692 6572
rect 11732 6532 14132 6572
rect 16579 6532 16588 6572
rect 16628 6532 17548 6572
rect 17588 6532 18028 6572
rect 18068 6532 18077 6572
rect 18412 6532 19468 6572
rect 19508 6532 19517 6572
rect 2500 6488 2540 6532
rect 4099 6488 4157 6489
rect 6019 6488 6077 6489
rect 2371 6448 2380 6488
rect 2420 6448 2540 6488
rect 2851 6448 2860 6488
rect 2900 6448 4012 6488
rect 4052 6448 4108 6488
rect 4148 6448 4176 6488
rect 4291 6448 4300 6488
rect 4340 6448 5548 6488
rect 5588 6448 5597 6488
rect 5934 6448 6028 6488
rect 6068 6448 6077 6488
rect 4099 6447 4157 6448
rect 6019 6447 6077 6448
rect 5827 6404 5885 6405
rect 5742 6364 5836 6404
rect 5876 6364 5885 6404
rect 5827 6363 5885 6364
rect 7372 6320 7412 6532
rect 11683 6531 11741 6532
rect 7843 6488 7901 6489
rect 8707 6488 8765 6489
rect 10339 6488 10397 6489
rect 12259 6488 12317 6489
rect 14092 6488 14132 6532
rect 18307 6488 18365 6489
rect 19651 6488 19709 6489
rect 7843 6448 7852 6488
rect 7892 6448 8332 6488
rect 8372 6448 8381 6488
rect 8622 6448 8716 6488
rect 8756 6448 8765 6488
rect 7843 6447 7901 6448
rect 8707 6447 8765 6448
rect 9964 6448 10292 6488
rect 9964 6404 10004 6448
rect 7459 6364 7468 6404
rect 7508 6364 10004 6404
rect 10051 6404 10109 6405
rect 10252 6404 10292 6448
rect 10339 6448 10348 6488
rect 10388 6448 11692 6488
rect 11732 6448 12268 6488
rect 12308 6448 13708 6488
rect 13748 6448 13757 6488
rect 14083 6448 14092 6488
rect 14132 6448 14141 6488
rect 15811 6448 15820 6488
rect 15860 6448 16108 6488
rect 16148 6448 16157 6488
rect 16675 6448 16684 6488
rect 16724 6448 17260 6488
rect 17300 6448 17309 6488
rect 17443 6448 17452 6488
rect 17492 6448 17836 6488
rect 17876 6448 17885 6488
rect 18307 6448 18316 6488
rect 18356 6448 19564 6488
rect 19604 6448 19660 6488
rect 19700 6448 19709 6488
rect 10339 6447 10397 6448
rect 12259 6447 12317 6448
rect 18307 6447 18365 6448
rect 19651 6447 19709 6448
rect 10051 6364 10060 6404
rect 10100 6364 10194 6404
rect 10252 6364 10484 6404
rect 16387 6364 16396 6404
rect 16436 6364 17660 6404
rect 10051 6363 10109 6364
rect 7555 6320 7613 6321
rect 10243 6320 10301 6321
rect 10444 6320 10484 6364
rect 17620 6320 17660 6364
rect 19939 6320 19997 6321
rect 1699 6280 1708 6320
rect 1748 6280 1757 6320
rect 2179 6280 2188 6320
rect 2228 6280 2380 6320
rect 2420 6280 2429 6320
rect 2563 6280 2572 6320
rect 2612 6280 3436 6320
rect 3476 6280 3485 6320
rect 5731 6280 5740 6320
rect 5780 6280 6740 6320
rect 7363 6280 7372 6320
rect 7412 6280 7421 6320
rect 7555 6280 7564 6320
rect 7604 6280 7698 6320
rect 7843 6280 7852 6320
rect 7892 6280 9580 6320
rect 9620 6280 9629 6320
rect 10158 6280 10252 6320
rect 10292 6280 10301 6320
rect 10435 6280 10444 6320
rect 10484 6280 10493 6320
rect 10915 6280 10924 6320
rect 10964 6280 16588 6320
rect 16628 6280 16637 6320
rect 17620 6280 19180 6320
rect 19220 6280 19229 6320
rect 19843 6280 19852 6320
rect 19892 6280 19948 6320
rect 19988 6280 19997 6320
rect 643 6236 701 6237
rect 558 6196 652 6236
rect 692 6196 701 6236
rect 5635 6196 5644 6236
rect 5684 6196 6124 6236
rect 6164 6196 6173 6236
rect 643 6195 701 6196
rect 0 6152 80 6172
rect 1891 6152 1949 6153
rect 4771 6152 4829 6153
rect 5443 6152 5501 6153
rect 6700 6152 6740 6280
rect 7555 6279 7613 6280
rect 10243 6279 10301 6280
rect 19939 6279 19997 6280
rect 20803 6320 20861 6321
rect 21424 6320 21504 6340
rect 20803 6280 20812 6320
rect 20852 6280 21504 6320
rect 20803 6279 20861 6280
rect 21424 6260 21504 6280
rect 7075 6236 7133 6237
rect 11971 6236 12029 6237
rect 6892 6196 7084 6236
rect 7124 6196 10196 6236
rect 11875 6196 11884 6236
rect 11924 6196 11980 6236
rect 12020 6196 12029 6236
rect 6892 6152 6932 6196
rect 7075 6195 7133 6196
rect 10051 6152 10109 6153
rect 0 6112 1900 6152
rect 1940 6112 1949 6152
rect 4195 6112 4204 6152
rect 4244 6112 4780 6152
rect 4820 6112 4829 6152
rect 5251 6112 5260 6152
rect 5300 6112 5452 6152
rect 5492 6112 5501 6152
rect 6691 6112 6700 6152
rect 6740 6112 6749 6152
rect 6883 6112 6892 6152
rect 6932 6112 6941 6152
rect 7651 6112 7660 6152
rect 7700 6112 8332 6152
rect 8372 6112 8716 6152
rect 8756 6112 8765 6152
rect 9868 6112 10060 6152
rect 10100 6112 10109 6152
rect 10156 6152 10196 6196
rect 11971 6195 12029 6196
rect 13411 6236 13469 6237
rect 19267 6236 19325 6237
rect 13411 6196 13420 6236
rect 13460 6196 14284 6236
rect 14324 6196 14333 6236
rect 15043 6196 15052 6236
rect 15092 6196 15532 6236
rect 15572 6196 15581 6236
rect 16195 6196 16204 6236
rect 16244 6196 19084 6236
rect 19124 6196 19133 6236
rect 19267 6196 19276 6236
rect 19316 6196 20044 6236
rect 20084 6196 20093 6236
rect 13411 6195 13469 6196
rect 19267 6195 19325 6196
rect 16579 6152 16637 6153
rect 10156 6112 16396 6152
rect 16436 6112 16445 6152
rect 16579 6112 16588 6152
rect 16628 6112 17644 6152
rect 17684 6112 17693 6152
rect 18019 6112 18028 6152
rect 18068 6112 18412 6152
rect 18452 6112 18461 6152
rect 0 6092 80 6112
rect 1891 6111 1949 6112
rect 4771 6111 4829 6112
rect 5443 6111 5501 6112
rect 9868 6068 9908 6112
rect 10051 6111 10109 6112
rect 16579 6111 16637 6112
rect 13987 6068 14045 6069
rect 14467 6068 14525 6069
rect 18307 6068 18365 6069
rect 3679 6028 3688 6068
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 4056 6028 4065 6068
rect 4396 6028 6796 6068
rect 6836 6028 6845 6068
rect 7276 6028 9908 6068
rect 10339 6028 10348 6068
rect 10388 6028 13996 6068
rect 14036 6028 14476 6068
rect 14516 6028 14525 6068
rect 17155 6028 17164 6068
rect 17204 6028 18316 6068
rect 18356 6028 18365 6068
rect 18799 6028 18808 6068
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 19176 6028 19185 6068
rect 4396 5984 4436 6028
rect 7276 5984 7316 6028
rect 13987 6027 14045 6028
rect 14467 6027 14525 6028
rect 18307 6027 18365 6028
rect 7459 5984 7517 5985
rect 14275 5984 14333 5985
rect 19555 5984 19613 5985
rect 3148 5944 4436 5984
rect 4483 5944 4492 5984
rect 4532 5944 6508 5984
rect 6548 5944 7276 5984
rect 7316 5944 7325 5984
rect 7374 5944 7468 5984
rect 7508 5944 7517 5984
rect 8323 5944 8332 5984
rect 8372 5944 12940 5984
rect 12980 5944 12989 5984
rect 14275 5944 14284 5984
rect 14324 5944 19564 5984
rect 19604 5944 19613 5984
rect 3148 5900 3188 5944
rect 7459 5943 7517 5944
rect 14275 5943 14333 5944
rect 19555 5943 19613 5944
rect 3139 5860 3148 5900
rect 3188 5860 3197 5900
rect 4387 5860 4396 5900
rect 4436 5860 8620 5900
rect 8660 5860 8669 5900
rect 8803 5860 8812 5900
rect 8852 5860 12268 5900
rect 12308 5860 12317 5900
rect 14563 5860 14572 5900
rect 14612 5860 20140 5900
rect 20180 5860 20189 5900
rect 0 5816 80 5836
rect 11395 5816 11453 5817
rect 21424 5816 21504 5836
rect 0 5776 268 5816
rect 308 5776 317 5816
rect 2764 5776 2860 5816
rect 2900 5776 2909 5816
rect 3811 5776 3820 5816
rect 3860 5776 10348 5816
rect 10388 5776 10397 5816
rect 11395 5776 11404 5816
rect 11444 5776 13612 5816
rect 13652 5776 13661 5816
rect 14179 5776 14188 5816
rect 14228 5776 15436 5816
rect 15476 5776 15485 5816
rect 16099 5776 16108 5816
rect 16148 5776 16300 5816
rect 16340 5776 16349 5816
rect 17923 5776 17932 5816
rect 17972 5776 18220 5816
rect 18260 5776 18269 5816
rect 20803 5776 20812 5816
rect 20852 5776 21004 5816
rect 21044 5776 21504 5816
rect 0 5756 80 5776
rect 1987 5648 2045 5649
rect 2764 5648 2804 5776
rect 11395 5775 11453 5776
rect 21424 5756 21504 5776
rect 19267 5732 19325 5733
rect 3436 5692 5780 5732
rect 5827 5692 5836 5732
rect 5876 5692 11360 5732
rect 12355 5692 12364 5732
rect 12404 5692 14612 5732
rect 17827 5692 17836 5732
rect 17876 5692 19276 5732
rect 19316 5692 19325 5732
rect 1219 5608 1228 5648
rect 1268 5608 1996 5648
rect 2036 5608 2045 5648
rect 2467 5608 2476 5648
rect 2516 5608 2804 5648
rect 3043 5608 3052 5648
rect 3092 5608 3101 5648
rect 3331 5608 3340 5648
rect 3380 5608 3389 5648
rect 1987 5607 2045 5608
rect 3052 5564 3092 5608
rect 2659 5524 2668 5564
rect 2708 5524 3092 5564
rect 0 5480 80 5500
rect 3340 5480 3380 5608
rect 0 5440 3380 5480
rect 0 5420 80 5440
rect 1027 5396 1085 5397
rect 3436 5396 3476 5692
rect 4675 5648 4733 5649
rect 5740 5648 5780 5692
rect 11320 5648 11360 5692
rect 14572 5648 14612 5692
rect 19267 5691 19325 5692
rect 18499 5648 18557 5649
rect 3523 5608 3532 5648
rect 3572 5608 3581 5648
rect 3907 5608 3916 5648
rect 3956 5608 4492 5648
rect 4532 5608 4541 5648
rect 4675 5608 4684 5648
rect 4724 5608 5068 5648
rect 5108 5608 5117 5648
rect 5740 5608 9620 5648
rect 9667 5608 9676 5648
rect 9716 5608 11212 5648
rect 11252 5608 11261 5648
rect 11320 5608 11788 5648
rect 11828 5608 12460 5648
rect 12500 5608 12509 5648
rect 14563 5608 14572 5648
rect 14612 5608 14621 5648
rect 15235 5608 15244 5648
rect 15284 5608 15820 5648
rect 15860 5608 15869 5648
rect 18115 5608 18124 5648
rect 18164 5608 18508 5648
rect 18548 5608 18557 5648
rect 3532 5564 3572 5608
rect 4675 5607 4733 5608
rect 9580 5564 9620 5608
rect 10435 5564 10493 5565
rect 3532 5524 6740 5564
rect 7171 5524 7180 5564
rect 7220 5524 8140 5564
rect 8180 5524 8189 5564
rect 8515 5524 8524 5564
rect 8564 5524 9004 5564
rect 9044 5524 9053 5564
rect 9580 5524 10444 5564
rect 10484 5524 10493 5564
rect 14572 5564 14612 5608
rect 18499 5607 18557 5608
rect 19459 5648 19517 5649
rect 19459 5608 19468 5648
rect 19508 5608 19756 5648
rect 19796 5608 19805 5648
rect 19459 5607 19517 5608
rect 15523 5564 15581 5565
rect 14572 5524 15532 5564
rect 15572 5524 19508 5564
rect 19939 5524 19948 5564
rect 19988 5524 20236 5564
rect 20276 5524 20620 5564
rect 20660 5524 20669 5564
rect 5827 5480 5885 5481
rect 6499 5480 6557 5481
rect 6700 5480 6740 5524
rect 8140 5480 8180 5524
rect 10435 5523 10493 5524
rect 15523 5523 15581 5524
rect 12931 5480 12989 5481
rect 19363 5480 19421 5481
rect 3523 5440 3532 5480
rect 3572 5440 5548 5480
rect 5588 5440 5597 5480
rect 5827 5440 5836 5480
rect 5876 5440 5932 5480
rect 5972 5440 5981 5480
rect 6403 5440 6412 5480
rect 6452 5440 6508 5480
rect 6548 5440 6557 5480
rect 6691 5440 6700 5480
rect 6740 5440 6749 5480
rect 8140 5440 11404 5480
rect 11444 5440 12940 5480
rect 12980 5440 13036 5480
rect 13076 5440 13085 5480
rect 14083 5440 14092 5480
rect 14132 5440 16588 5480
rect 16628 5440 16637 5480
rect 17827 5440 17836 5480
rect 17876 5440 19372 5480
rect 19412 5440 19421 5480
rect 5827 5439 5885 5440
rect 5932 5396 5972 5440
rect 6499 5439 6557 5440
rect 12931 5439 12989 5440
rect 14092 5396 14132 5440
rect 19363 5439 19421 5440
rect 18595 5396 18653 5397
rect 942 5356 1036 5396
rect 1076 5356 1085 5396
rect 1027 5355 1085 5356
rect 2500 5356 3476 5396
rect 3619 5356 3628 5396
rect 3668 5356 4588 5396
rect 4628 5356 5740 5396
rect 5780 5356 5789 5396
rect 5932 5356 7660 5396
rect 7700 5356 7709 5396
rect 10723 5356 10732 5396
rect 10772 5356 14132 5396
rect 15523 5356 15532 5396
rect 15572 5356 16108 5396
rect 16148 5356 16157 5396
rect 18115 5356 18124 5396
rect 18164 5356 18604 5396
rect 18644 5356 18653 5396
rect 0 5144 80 5164
rect 2500 5144 2540 5356
rect 4291 5312 4349 5313
rect 6307 5312 6365 5313
rect 10732 5312 10772 5356
rect 18595 5355 18653 5356
rect 3139 5272 3148 5312
rect 3188 5272 4300 5312
rect 4340 5272 4349 5312
rect 4919 5272 4928 5312
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 5296 5272 5305 5312
rect 6307 5272 6316 5312
rect 6356 5272 10772 5312
rect 13987 5312 14045 5313
rect 17059 5312 17117 5313
rect 13987 5272 13996 5312
rect 14036 5272 17068 5312
rect 17108 5272 17117 5312
rect 4291 5271 4349 5272
rect 6307 5271 6365 5272
rect 13987 5271 14045 5272
rect 17059 5271 17117 5272
rect 5443 5228 5501 5229
rect 8707 5228 8765 5229
rect 10819 5228 10877 5229
rect 11107 5228 11165 5229
rect 14467 5228 14525 5229
rect 19468 5228 19508 5524
rect 21424 5312 21504 5332
rect 20039 5272 20048 5312
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20416 5272 20425 5312
rect 20812 5272 21504 5312
rect 20812 5228 20852 5272
rect 21424 5252 21504 5272
rect 2851 5188 2860 5228
rect 2900 5188 3724 5228
rect 3764 5188 5452 5228
rect 5492 5188 5501 5228
rect 6595 5188 6604 5228
rect 6644 5188 6796 5228
rect 6836 5188 6845 5228
rect 8131 5188 8140 5228
rect 8180 5188 8332 5228
rect 8372 5188 8716 5228
rect 8756 5188 8765 5228
rect 10627 5188 10636 5228
rect 10676 5188 10828 5228
rect 10868 5188 10877 5228
rect 11022 5188 11116 5228
rect 11156 5188 11165 5228
rect 11395 5188 11404 5228
rect 11444 5188 11596 5228
rect 11636 5188 11884 5228
rect 11924 5188 11933 5228
rect 14467 5188 14476 5228
rect 14516 5188 18508 5228
rect 18548 5188 18557 5228
rect 19084 5188 19372 5228
rect 19412 5188 19421 5228
rect 19468 5188 20812 5228
rect 20852 5188 20861 5228
rect 5443 5187 5501 5188
rect 8707 5187 8765 5188
rect 10819 5187 10877 5188
rect 11107 5187 11165 5188
rect 14467 5187 14525 5188
rect 9667 5144 9725 5145
rect 10627 5144 10685 5145
rect 19084 5144 19124 5188
rect 19747 5144 19805 5145
rect 0 5104 2540 5144
rect 3427 5104 3436 5144
rect 3476 5104 4492 5144
rect 4532 5104 4541 5144
rect 9667 5104 9676 5144
rect 9716 5104 10100 5144
rect 0 5084 80 5104
rect 9667 5103 9725 5104
rect 8803 5060 8861 5061
rect 9571 5060 9629 5061
rect 10060 5060 10100 5104
rect 10627 5104 10636 5144
rect 10676 5104 11308 5144
rect 11348 5104 11357 5144
rect 11779 5104 11788 5144
rect 11828 5104 16916 5144
rect 16963 5104 16972 5144
rect 17012 5104 17356 5144
rect 17396 5104 17405 5144
rect 17827 5104 17836 5144
rect 17876 5104 18220 5144
rect 18260 5104 18269 5144
rect 18403 5104 18412 5144
rect 18452 5104 19124 5144
rect 19180 5104 19756 5144
rect 19796 5104 19805 5144
rect 10627 5103 10685 5104
rect 16876 5060 16916 5104
rect 19180 5060 19220 5104
rect 19747 5103 19805 5104
rect 2563 5020 2572 5060
rect 2612 5020 6124 5060
rect 6164 5020 6173 5060
rect 8803 5020 8812 5060
rect 8852 5020 9196 5060
rect 9236 5020 9245 5060
rect 9571 5020 9580 5060
rect 9620 5020 9812 5060
rect 10060 5020 11360 5060
rect 13987 5020 13996 5060
rect 14036 5020 14045 5060
rect 15043 5020 15052 5060
rect 15092 5020 15436 5060
rect 15476 5020 15485 5060
rect 16876 5020 19220 5060
rect 8803 5019 8861 5020
rect 9571 5019 9629 5020
rect 2659 4976 2717 4977
rect 9379 4976 9437 4977
rect 9772 4976 9812 5020
rect 10243 4976 10301 4977
rect 2659 4936 2668 4976
rect 2708 4936 3628 4976
rect 3668 4936 3677 4976
rect 4291 4936 4300 4976
rect 4340 4936 8812 4976
rect 8852 4936 8861 4976
rect 9379 4936 9388 4976
rect 9428 4936 9676 4976
rect 9716 4936 9725 4976
rect 9772 4936 10156 4976
rect 10196 4936 10252 4976
rect 10292 4936 10301 4976
rect 2659 4935 2717 4936
rect 9379 4935 9437 4936
rect 10243 4935 10301 4936
rect 10924 4936 11116 4976
rect 11156 4936 11165 4976
rect 1315 4892 1373 4893
rect 5347 4892 5405 4893
rect 8227 4892 8285 4893
rect 10924 4892 10964 4936
rect 1315 4852 1324 4892
rect 1364 4852 2092 4892
rect 2132 4852 2141 4892
rect 5347 4852 5356 4892
rect 5396 4852 6892 4892
rect 6932 4852 6941 4892
rect 7555 4852 7564 4892
rect 7604 4852 8236 4892
rect 8276 4852 8852 4892
rect 10243 4852 10252 4892
rect 10292 4852 10964 4892
rect 11320 4892 11360 5020
rect 13996 4976 14036 5020
rect 17827 4976 17885 4977
rect 18019 4976 18077 4977
rect 18403 4976 18461 4977
rect 11971 4936 11980 4976
rect 12020 4936 12556 4976
rect 12596 4936 12748 4976
rect 12788 4936 12797 4976
rect 13507 4936 13516 4976
rect 13556 4936 13900 4976
rect 13940 4936 13949 4976
rect 13996 4936 17164 4976
rect 17204 4936 17213 4976
rect 17731 4936 17740 4976
rect 17780 4936 17836 4976
rect 17876 4936 17885 4976
rect 17934 4936 18028 4976
rect 18068 4936 18077 4976
rect 18211 4936 18220 4976
rect 18260 4936 18412 4976
rect 18452 4936 18461 4976
rect 17827 4935 17885 4936
rect 18019 4935 18077 4936
rect 18403 4935 18461 4936
rect 18595 4976 18653 4977
rect 18595 4936 18604 4976
rect 18644 4936 18738 4976
rect 18595 4935 18653 4936
rect 16291 4892 16349 4893
rect 11320 4852 12460 4892
rect 12500 4852 14476 4892
rect 14516 4852 14525 4892
rect 16291 4852 16300 4892
rect 16340 4852 21196 4892
rect 21236 4852 21245 4892
rect 1315 4851 1373 4852
rect 5347 4851 5405 4852
rect 8227 4851 8285 4852
rect 0 4808 80 4828
rect 1219 4808 1277 4809
rect 8812 4808 8852 4852
rect 16291 4851 16349 4852
rect 16300 4808 16340 4851
rect 21424 4808 21504 4828
rect 0 4768 1228 4808
rect 1268 4768 1277 4808
rect 6307 4768 6316 4808
rect 6356 4768 7084 4808
rect 7124 4768 7988 4808
rect 8803 4768 8812 4808
rect 8852 4768 12748 4808
rect 12788 4768 12797 4808
rect 12931 4768 12940 4808
rect 12980 4768 16340 4808
rect 18307 4768 18316 4808
rect 18356 4768 18700 4808
rect 18740 4768 18749 4808
rect 20419 4768 20428 4808
rect 20468 4768 21504 4808
rect 0 4748 80 4768
rect 1219 4767 1277 4768
rect 7555 4724 7613 4725
rect 7948 4724 7988 4768
rect 21424 4748 21504 4768
rect 10339 4724 10397 4725
rect 15331 4724 15389 4725
rect 20611 4724 20669 4725
rect 2275 4684 2284 4724
rect 2324 4684 7564 4724
rect 7604 4684 7613 4724
rect 7939 4684 7948 4724
rect 7988 4684 9004 4724
rect 9044 4684 10348 4724
rect 10388 4684 10397 4724
rect 13411 4684 13420 4724
rect 13460 4684 13708 4724
rect 13748 4684 13757 4724
rect 15331 4684 15340 4724
rect 15380 4684 17660 4724
rect 7555 4683 7613 4684
rect 10339 4683 10397 4684
rect 15331 4683 15389 4684
rect 16483 4640 16541 4641
rect 2371 4600 2380 4640
rect 2420 4600 3148 4640
rect 3188 4600 5684 4640
rect 6979 4600 6988 4640
rect 7028 4600 8428 4640
rect 8468 4600 12460 4640
rect 12500 4600 12509 4640
rect 15811 4600 15820 4640
rect 15860 4600 16492 4640
rect 16532 4600 16541 4640
rect 17620 4640 17660 4684
rect 18604 4684 20620 4724
rect 20660 4684 20669 4724
rect 18499 4640 18557 4641
rect 17620 4600 18508 4640
rect 18548 4600 18557 4640
rect 5644 4556 5684 4600
rect 16483 4599 16541 4600
rect 18499 4599 18557 4600
rect 18604 4556 18644 4684
rect 20611 4683 20669 4684
rect 18691 4600 18700 4640
rect 18740 4600 20716 4640
rect 20756 4600 20765 4640
rect 21091 4556 21149 4557
rect 3679 4516 3688 4556
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 4056 4516 4065 4556
rect 5644 4516 12364 4556
rect 12404 4516 14380 4556
rect 14420 4516 14429 4556
rect 18019 4516 18028 4556
rect 18068 4516 18644 4556
rect 18799 4516 18808 4556
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 19176 4516 19185 4556
rect 19276 4516 21100 4556
rect 21140 4516 21149 4556
rect 0 4472 80 4492
rect 1411 4472 1469 4473
rect 0 4432 1420 4472
rect 1460 4432 1469 4472
rect 0 4412 80 4432
rect 1411 4431 1469 4432
rect 4291 4472 4349 4473
rect 6019 4472 6077 4473
rect 8515 4472 8573 4473
rect 17347 4472 17405 4473
rect 18403 4472 18461 4473
rect 4291 4432 4300 4472
rect 4340 4432 4396 4472
rect 4436 4432 5644 4472
rect 5684 4432 5693 4472
rect 6019 4432 6028 4472
rect 6068 4432 8524 4472
rect 8564 4432 11500 4472
rect 11540 4432 11549 4472
rect 12547 4432 12556 4472
rect 12596 4432 17300 4472
rect 4291 4431 4349 4432
rect 6019 4431 6077 4432
rect 8515 4431 8573 4432
rect 4771 4388 4829 4389
rect 6211 4388 6269 4389
rect 13315 4388 13373 4389
rect 14083 4388 14141 4389
rect 14755 4388 14813 4389
rect 2275 4348 2284 4388
rect 2324 4348 4780 4388
rect 4820 4348 4829 4388
rect 5827 4348 5836 4388
rect 5876 4348 6220 4388
rect 6260 4348 6269 4388
rect 6499 4348 6508 4388
rect 6548 4348 6796 4388
rect 6836 4348 6845 4388
rect 8707 4348 8716 4388
rect 8756 4348 10676 4388
rect 13230 4348 13324 4388
rect 13364 4348 13373 4388
rect 13507 4348 13516 4388
rect 13556 4348 13804 4388
rect 13844 4348 13853 4388
rect 13998 4348 14092 4388
rect 14132 4348 14141 4388
rect 14467 4348 14476 4388
rect 14516 4348 14764 4388
rect 14804 4348 14813 4388
rect 17260 4388 17300 4432
rect 17347 4432 17356 4472
rect 17396 4432 18412 4472
rect 18452 4432 18461 4472
rect 17347 4431 17405 4432
rect 18403 4431 18461 4432
rect 19276 4388 19316 4516
rect 21091 4515 21149 4516
rect 19651 4472 19709 4473
rect 19363 4432 19372 4472
rect 19412 4432 19660 4472
rect 19700 4432 19948 4472
rect 19988 4432 19997 4472
rect 19651 4431 19709 4432
rect 17260 4348 18700 4388
rect 18740 4348 19316 4388
rect 4771 4347 4829 4348
rect 6211 4347 6269 4348
rect 2755 4304 2813 4305
rect 10243 4304 10301 4305
rect 2755 4264 2764 4304
rect 2804 4264 10252 4304
rect 10292 4264 10301 4304
rect 2755 4263 2813 4264
rect 10243 4263 10301 4264
rect 10348 4264 10540 4304
rect 10580 4264 10589 4304
rect 2275 4220 2333 4221
rect 6595 4220 6653 4221
rect 10348 4220 10388 4264
rect 10636 4220 10676 4348
rect 13315 4347 13373 4348
rect 14083 4347 14141 4348
rect 14755 4347 14813 4348
rect 17635 4304 17693 4305
rect 21424 4304 21504 4324
rect 13891 4264 13900 4304
rect 13940 4264 14188 4304
rect 14228 4264 14237 4304
rect 14947 4264 14956 4304
rect 14996 4264 17644 4304
rect 17684 4264 18412 4304
rect 18452 4264 18461 4304
rect 20803 4264 20812 4304
rect 20852 4264 21504 4304
rect 17635 4263 17693 4264
rect 21424 4244 21504 4264
rect 1507 4180 1516 4220
rect 1556 4180 2284 4220
rect 2324 4180 2540 4220
rect 3043 4180 3052 4220
rect 3092 4180 3340 4220
rect 3380 4180 3389 4220
rect 4195 4180 4204 4220
rect 4244 4180 4684 4220
rect 4724 4180 5836 4220
rect 5876 4180 5885 4220
rect 6307 4180 6316 4220
rect 6356 4180 6604 4220
rect 6644 4180 7852 4220
rect 7892 4180 8716 4220
rect 8756 4180 8765 4220
rect 10051 4180 10060 4220
rect 10100 4180 10348 4220
rect 10388 4180 10397 4220
rect 10636 4180 11252 4220
rect 2275 4179 2333 4180
rect 0 4137 80 4156
rect 0 4136 125 4137
rect 1603 4136 1661 4137
rect 0 4096 76 4136
rect 116 4096 125 4136
rect 1315 4096 1324 4136
rect 1364 4096 1612 4136
rect 1652 4096 1661 4136
rect 2500 4136 2540 4180
rect 6595 4179 6653 4180
rect 7843 4136 7901 4137
rect 11212 4136 11252 4180
rect 11320 4180 11596 4220
rect 11636 4180 17740 4220
rect 17780 4180 17789 4220
rect 18316 4180 20180 4220
rect 2500 4096 4588 4136
rect 4628 4096 4637 4136
rect 5260 4096 6220 4136
rect 6260 4096 7852 4136
rect 7892 4096 7901 4136
rect 9091 4096 9100 4136
rect 9140 4096 10540 4136
rect 10580 4096 10589 4136
rect 11203 4096 11212 4136
rect 11252 4096 11261 4136
rect 0 4095 125 4096
rect 1603 4095 1661 4096
rect 0 4076 80 4095
rect 5260 4052 5300 4096
rect 7843 4095 7901 4096
rect 11320 4052 11360 4180
rect 16579 4136 16637 4137
rect 18316 4136 18356 4180
rect 18499 4136 18557 4137
rect 20140 4136 20180 4180
rect 12739 4096 12748 4136
rect 12788 4096 16396 4136
rect 16436 4096 16445 4136
rect 16579 4096 16588 4136
rect 16628 4096 18356 4136
rect 18414 4096 18508 4136
rect 18548 4096 18557 4136
rect 19171 4096 19180 4136
rect 19220 4096 19756 4136
rect 19796 4096 19805 4136
rect 20140 4096 21388 4136
rect 21428 4096 21437 4136
rect 16579 4095 16637 4096
rect 18499 4095 18557 4096
rect 4387 4012 4396 4052
rect 4436 4012 5300 4052
rect 5347 4012 5356 4052
rect 5396 4012 11360 4052
rect 12451 4012 12460 4052
rect 12500 4012 20428 4052
rect 20468 4012 20477 4052
rect 11971 3968 12029 3969
rect 2659 3928 2668 3968
rect 2708 3928 7372 3968
rect 7412 3928 7421 3968
rect 7651 3928 7660 3968
rect 7700 3928 8140 3968
rect 8180 3928 10636 3968
rect 10676 3928 10924 3968
rect 10964 3928 10973 3968
rect 11971 3928 11980 3968
rect 12020 3928 12308 3968
rect 14083 3928 14092 3968
rect 14132 3928 14668 3968
rect 14708 3928 14717 3968
rect 19363 3928 19372 3968
rect 19412 3928 19948 3968
rect 19988 3928 19997 3968
rect 11971 3927 12029 3928
rect 2755 3884 2813 3885
rect 10435 3884 10493 3885
rect 2755 3844 2764 3884
rect 2804 3844 3244 3884
rect 3284 3844 3293 3884
rect 4099 3844 4108 3884
rect 4148 3844 8948 3884
rect 10350 3844 10444 3884
rect 10484 3844 10493 3884
rect 2755 3843 2813 3844
rect 0 3800 80 3820
rect 355 3800 413 3801
rect 3139 3800 3197 3801
rect 0 3760 364 3800
rect 404 3760 413 3800
rect 2947 3760 2956 3800
rect 2996 3760 3148 3800
rect 3188 3760 3197 3800
rect 0 3740 80 3760
rect 355 3759 413 3760
rect 3139 3759 3197 3760
rect 3331 3800 3389 3801
rect 4099 3800 4157 3801
rect 4579 3800 4637 3801
rect 5827 3800 5885 3801
rect 6115 3800 6173 3801
rect 8908 3800 8948 3844
rect 10435 3843 10493 3844
rect 10627 3884 10685 3885
rect 12268 3884 12308 3928
rect 10627 3844 10636 3884
rect 10676 3844 11116 3884
rect 11156 3844 11165 3884
rect 11395 3844 11404 3884
rect 11444 3844 12172 3884
rect 12212 3844 12221 3884
rect 12268 3844 13505 3884
rect 13545 3844 13554 3884
rect 13987 3844 13996 3884
rect 14036 3844 15340 3884
rect 15380 3844 15389 3884
rect 15715 3844 15724 3884
rect 15764 3844 17164 3884
rect 17204 3844 17213 3884
rect 17731 3844 17740 3884
rect 17780 3844 18316 3884
rect 18356 3844 20812 3884
rect 20852 3844 20861 3884
rect 10627 3843 10685 3844
rect 11299 3800 11357 3801
rect 3331 3760 3340 3800
rect 3380 3760 3436 3800
rect 3476 3760 3485 3800
rect 3907 3760 3916 3800
rect 3956 3760 4108 3800
rect 4148 3760 4588 3800
rect 4628 3760 4637 3800
rect 4919 3760 4928 3800
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 5296 3760 5305 3800
rect 5731 3760 5740 3800
rect 5780 3760 5836 3800
rect 5876 3760 5885 3800
rect 6019 3760 6028 3800
rect 6068 3760 6124 3800
rect 6164 3760 6173 3800
rect 8899 3760 8908 3800
rect 8948 3760 8957 3800
rect 10147 3760 10156 3800
rect 10196 3760 11308 3800
rect 11348 3760 11357 3800
rect 3331 3759 3389 3760
rect 4099 3759 4157 3760
rect 4579 3759 4637 3760
rect 5827 3759 5885 3760
rect 6115 3759 6173 3760
rect 11299 3759 11357 3760
rect 12067 3800 12125 3801
rect 16771 3800 16829 3801
rect 21424 3800 21504 3820
rect 12067 3760 12076 3800
rect 12116 3760 14956 3800
rect 14996 3760 15005 3800
rect 16771 3760 16780 3800
rect 16820 3760 17356 3800
rect 17396 3760 17644 3800
rect 17684 3760 17693 3800
rect 17827 3760 17836 3800
rect 17876 3760 18028 3800
rect 18068 3760 18077 3800
rect 20039 3760 20048 3800
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20416 3760 20425 3800
rect 21379 3760 21388 3800
rect 21428 3760 21504 3800
rect 12067 3759 12125 3760
rect 16771 3759 16829 3760
rect 21424 3740 21504 3760
rect 7843 3716 7901 3717
rect 9283 3716 9341 3717
rect 4387 3676 4396 3716
rect 4436 3676 7660 3716
rect 7700 3676 7709 3716
rect 7843 3676 7852 3716
rect 7892 3676 9292 3716
rect 9332 3676 9341 3716
rect 10627 3676 10636 3716
rect 10676 3676 11020 3716
rect 11060 3676 11069 3716
rect 11116 3676 15340 3716
rect 15380 3676 18124 3716
rect 18164 3676 18173 3716
rect 7843 3675 7901 3676
rect 9283 3675 9341 3676
rect 1699 3632 1757 3633
rect 3043 3632 3101 3633
rect 11116 3632 11156 3676
rect 1699 3592 1708 3632
rect 1748 3592 1996 3632
rect 2036 3592 2045 3632
rect 2947 3592 2956 3632
rect 2996 3592 3052 3632
rect 3092 3592 3101 3632
rect 7939 3592 7948 3632
rect 7988 3592 11156 3632
rect 14083 3632 14141 3633
rect 14851 3632 14909 3633
rect 17827 3632 17885 3633
rect 14083 3592 14092 3632
rect 14132 3592 14860 3632
rect 14900 3592 17588 3632
rect 17635 3592 17644 3632
rect 17684 3592 17836 3632
rect 17876 3592 17885 3632
rect 19651 3592 19660 3632
rect 19700 3592 20044 3632
rect 20084 3592 20093 3632
rect 1699 3591 1757 3592
rect 3043 3591 3101 3592
rect 2659 3548 2717 3549
rect 5443 3548 5501 3549
rect 7948 3548 7988 3592
rect 14083 3591 14141 3592
rect 14851 3591 14909 3592
rect 11107 3548 11165 3549
rect 12931 3548 12989 3549
rect 15811 3548 15869 3549
rect 2574 3508 2668 3548
rect 2708 3508 2717 3548
rect 3715 3508 3724 3548
rect 3764 3508 4588 3548
rect 4628 3508 4637 3548
rect 5443 3508 5452 3548
rect 5492 3508 7988 3548
rect 8800 3508 10252 3548
rect 10292 3508 10540 3548
rect 10580 3508 10589 3548
rect 11107 3508 11116 3548
rect 11156 3508 12652 3548
rect 12692 3508 12701 3548
rect 12931 3508 12940 3548
rect 12980 3508 13036 3548
rect 13076 3508 13085 3548
rect 13315 3508 13324 3548
rect 13364 3508 13804 3548
rect 13844 3508 13853 3548
rect 15726 3508 15820 3548
rect 15860 3508 15869 3548
rect 17548 3548 17588 3592
rect 17827 3591 17885 3592
rect 19267 3548 19325 3549
rect 17548 3508 17836 3548
rect 17876 3508 17885 3548
rect 19267 3508 19276 3548
rect 19316 3508 19756 3548
rect 19796 3508 19805 3548
rect 2659 3507 2717 3508
rect 5443 3507 5501 3508
rect 0 3464 80 3484
rect 451 3464 509 3465
rect 0 3424 460 3464
rect 500 3424 509 3464
rect 2179 3424 2188 3464
rect 2228 3424 7756 3464
rect 7796 3424 7805 3464
rect 0 3404 80 3424
rect 451 3423 509 3424
rect 1507 3380 1565 3381
rect 7075 3380 7133 3381
rect 1422 3340 1516 3380
rect 1556 3340 1565 3380
rect 3619 3340 3628 3380
rect 3668 3340 5356 3380
rect 5396 3340 5405 3380
rect 5635 3340 5644 3380
rect 5684 3340 5932 3380
rect 5972 3340 6508 3380
rect 6548 3340 6557 3380
rect 6691 3340 6700 3380
rect 6740 3340 7084 3380
rect 7124 3340 7133 3380
rect 1507 3339 1565 3340
rect 7075 3339 7133 3340
rect 7651 3380 7709 3381
rect 8800 3380 8840 3508
rect 11107 3507 11165 3508
rect 12931 3507 12989 3508
rect 15811 3507 15869 3508
rect 19267 3507 19325 3508
rect 16291 3464 16349 3465
rect 16867 3464 16925 3465
rect 9667 3424 9676 3464
rect 9716 3424 11020 3464
rect 11060 3424 11069 3464
rect 11779 3424 11788 3464
rect 11828 3424 16108 3464
rect 16148 3424 16157 3464
rect 16291 3424 16300 3464
rect 16340 3424 16434 3464
rect 16867 3424 16876 3464
rect 16916 3424 18220 3464
rect 18260 3424 18269 3464
rect 18787 3424 18796 3464
rect 18836 3424 21004 3464
rect 21044 3424 21053 3464
rect 9571 3380 9629 3381
rect 7651 3340 7660 3380
rect 7700 3340 8840 3380
rect 8995 3340 9004 3380
rect 9044 3340 9580 3380
rect 9620 3340 9629 3380
rect 7651 3339 7709 3340
rect 9571 3339 9629 3340
rect 11788 3296 11828 3424
rect 16291 3423 16349 3424
rect 16867 3423 16925 3424
rect 13891 3380 13949 3381
rect 19363 3380 19421 3381
rect 13891 3340 13900 3380
rect 13940 3340 14380 3380
rect 14420 3340 14429 3380
rect 19363 3340 19372 3380
rect 19412 3340 19852 3380
rect 19892 3340 19901 3380
rect 19948 3340 20140 3380
rect 20180 3340 20189 3380
rect 13891 3339 13949 3340
rect 19363 3339 19421 3340
rect 16099 3296 16157 3297
rect 19948 3296 19988 3340
rect 21424 3296 21504 3316
rect 2659 3256 2668 3296
rect 2708 3256 4780 3296
rect 4820 3256 7084 3296
rect 7124 3256 7133 3296
rect 10531 3256 10540 3296
rect 10580 3256 11828 3296
rect 12835 3256 12844 3296
rect 12884 3256 13804 3296
rect 13844 3256 13853 3296
rect 14179 3256 14188 3296
rect 14228 3256 16108 3296
rect 16148 3256 16157 3296
rect 18019 3256 18028 3296
rect 18068 3256 19660 3296
rect 19700 3256 19709 3296
rect 19756 3256 19988 3296
rect 20140 3256 21504 3296
rect 16099 3255 16157 3256
rect 2851 3212 2909 3213
rect 17059 3212 17117 3213
rect 2755 3172 2764 3212
rect 2804 3172 2860 3212
rect 2900 3172 2909 3212
rect 3139 3172 3148 3212
rect 3188 3172 7468 3212
rect 7508 3172 7517 3212
rect 9475 3172 9484 3212
rect 9524 3172 11116 3212
rect 11156 3172 11165 3212
rect 11395 3172 11404 3212
rect 11444 3172 15436 3212
rect 15476 3172 15485 3212
rect 16974 3172 17068 3212
rect 17108 3172 17117 3212
rect 2851 3171 2909 3172
rect 17059 3171 17117 3172
rect 18691 3212 18749 3213
rect 19756 3212 19796 3256
rect 18691 3172 18700 3212
rect 18740 3172 19796 3212
rect 18691 3171 18749 3172
rect 0 3128 80 3148
rect 259 3128 317 3129
rect 19747 3128 19805 3129
rect 20140 3128 20180 3256
rect 21424 3236 21504 3256
rect 0 3088 268 3128
rect 308 3088 317 3128
rect 3331 3088 3340 3128
rect 3380 3088 6604 3128
rect 6644 3088 6653 3128
rect 7363 3088 7372 3128
rect 7412 3088 11788 3128
rect 11828 3088 11837 3128
rect 19747 3088 19756 3128
rect 19796 3088 20180 3128
rect 0 3068 80 3088
rect 259 3087 317 3088
rect 19747 3087 19805 3088
rect 14563 3044 14621 3045
rect 3679 3004 3688 3044
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 4056 3004 4065 3044
rect 4291 3004 4300 3044
rect 4340 3004 11308 3044
rect 11348 3004 11357 3044
rect 13507 3004 13516 3044
rect 13556 3004 14188 3044
rect 14228 3004 14237 3044
rect 14478 3004 14572 3044
rect 14612 3004 14621 3044
rect 14851 3004 14860 3044
rect 14900 3004 15052 3044
rect 15092 3004 15101 3044
rect 18799 3004 18808 3044
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 19176 3004 19185 3044
rect 14563 3003 14621 3004
rect 3523 2960 3581 2961
rect 7459 2960 7517 2961
rect 9091 2960 9149 2961
rect 3523 2920 3532 2960
rect 3572 2920 4396 2960
rect 4436 2920 7372 2960
rect 7412 2920 7468 2960
rect 7508 2920 7536 2960
rect 9091 2920 9100 2960
rect 9140 2920 14764 2960
rect 14804 2920 14813 2960
rect 15523 2920 15532 2960
rect 15572 2920 15916 2960
rect 15956 2920 15965 2960
rect 17923 2920 17932 2960
rect 17972 2920 19660 2960
rect 19700 2920 19709 2960
rect 3523 2919 3581 2920
rect 7459 2919 7517 2920
rect 9091 2919 9149 2920
rect 1795 2836 1804 2876
rect 1844 2836 4684 2876
rect 4724 2836 4733 2876
rect 9955 2836 9964 2876
rect 10004 2836 10013 2876
rect 10156 2836 14380 2876
rect 14420 2836 14429 2876
rect 16579 2836 16588 2876
rect 16628 2836 20180 2876
rect 20227 2836 20236 2876
rect 20276 2836 20716 2876
rect 20756 2836 20765 2876
rect 0 2792 80 2812
rect 835 2792 893 2793
rect 4771 2792 4829 2793
rect 9964 2792 10004 2836
rect 0 2752 844 2792
rect 884 2752 893 2792
rect 3235 2752 3244 2792
rect 3284 2752 3532 2792
rect 3572 2752 3581 2792
rect 3811 2752 3820 2792
rect 3860 2752 4780 2792
rect 4820 2752 4829 2792
rect 8707 2752 8716 2792
rect 8756 2752 10004 2792
rect 0 2732 80 2752
rect 835 2751 893 2752
rect 4771 2751 4829 2752
rect 3523 2708 3581 2709
rect 6883 2708 6941 2709
rect 7651 2708 7709 2709
rect 9379 2708 9437 2709
rect 10156 2708 10196 2836
rect 10819 2792 10877 2793
rect 20140 2792 20180 2836
rect 21424 2792 21504 2812
rect 10819 2752 10828 2792
rect 10868 2752 11884 2792
rect 11924 2752 11933 2792
rect 13027 2752 13036 2792
rect 13076 2752 13996 2792
rect 14036 2752 14045 2792
rect 16195 2752 16204 2792
rect 16244 2752 20044 2792
rect 20084 2752 20093 2792
rect 20140 2752 21504 2792
rect 10819 2751 10877 2752
rect 21424 2732 21504 2752
rect 10531 2708 10589 2709
rect 17251 2708 17309 2709
rect 2083 2668 2092 2708
rect 2132 2668 3148 2708
rect 3188 2668 3197 2708
rect 3523 2668 3532 2708
rect 3572 2668 3628 2708
rect 3668 2668 3677 2708
rect 3724 2668 6320 2708
rect 3523 2667 3581 2668
rect 547 2624 605 2625
rect 3724 2624 3764 2668
rect 5539 2624 5597 2625
rect 547 2584 556 2624
rect 596 2584 2708 2624
rect 2851 2584 2860 2624
rect 2900 2584 3764 2624
rect 5454 2584 5548 2624
rect 5588 2584 5597 2624
rect 547 2583 605 2584
rect 547 2500 556 2540
rect 596 2500 748 2540
rect 788 2500 797 2540
rect 0 2456 80 2476
rect 1219 2456 1277 2457
rect 0 2416 1228 2456
rect 1268 2416 1277 2456
rect 2668 2456 2708 2584
rect 5539 2583 5597 2584
rect 5923 2624 5981 2625
rect 5923 2584 5932 2624
rect 5972 2584 6124 2624
rect 6164 2584 6173 2624
rect 5923 2583 5981 2584
rect 2668 2416 4012 2456
rect 4052 2416 4061 2456
rect 0 2396 80 2416
rect 1219 2415 1277 2416
rect 6280 2372 6320 2668
rect 6883 2668 6892 2708
rect 6932 2668 6988 2708
rect 7028 2668 7037 2708
rect 7651 2668 7660 2708
rect 7700 2668 7756 2708
rect 7796 2668 7805 2708
rect 9294 2668 9388 2708
rect 9428 2668 9437 2708
rect 9763 2668 9772 2708
rect 9812 2668 10196 2708
rect 10446 2668 10540 2708
rect 10580 2668 10589 2708
rect 6883 2667 6941 2668
rect 7651 2667 7709 2668
rect 9379 2667 9437 2668
rect 10531 2667 10589 2668
rect 10732 2668 11116 2708
rect 11156 2668 11165 2708
rect 11692 2668 15052 2708
rect 15092 2668 15101 2708
rect 15811 2668 15820 2708
rect 15860 2668 17204 2708
rect 10732 2624 10772 2668
rect 11692 2624 11732 2668
rect 17164 2624 17204 2668
rect 17251 2668 17260 2708
rect 17300 2668 17452 2708
rect 17492 2668 17501 2708
rect 18115 2668 18124 2708
rect 18164 2668 21100 2708
rect 21140 2668 21149 2708
rect 17251 2667 17309 2668
rect 19651 2624 19709 2625
rect 6595 2584 6604 2624
rect 6644 2584 10772 2624
rect 10915 2584 10924 2624
rect 10964 2584 11732 2624
rect 11779 2584 11788 2624
rect 11828 2584 14900 2624
rect 9091 2540 9149 2541
rect 9955 2540 10013 2541
rect 10339 2540 10397 2541
rect 10627 2540 10685 2541
rect 6787 2500 6796 2540
rect 6836 2500 8044 2540
rect 8084 2500 8093 2540
rect 9091 2500 9100 2540
rect 9140 2500 9234 2540
rect 9955 2500 9964 2540
rect 10004 2500 10060 2540
rect 10100 2500 10109 2540
rect 10339 2500 10348 2540
rect 10388 2500 10397 2540
rect 10542 2500 10636 2540
rect 10676 2500 10685 2540
rect 9091 2499 9149 2500
rect 9955 2499 10013 2500
rect 10339 2499 10397 2500
rect 10627 2499 10685 2500
rect 10819 2540 10877 2541
rect 14860 2540 14900 2584
rect 15340 2584 16012 2624
rect 16052 2584 16061 2624
rect 17164 2584 19084 2624
rect 19124 2584 19133 2624
rect 19651 2584 19660 2624
rect 19700 2584 20140 2624
rect 20180 2584 20189 2624
rect 15235 2540 15293 2541
rect 15340 2540 15380 2584
rect 19651 2583 19709 2584
rect 10819 2500 10828 2540
rect 10868 2500 11020 2540
rect 11060 2500 11069 2540
rect 14860 2500 15244 2540
rect 15284 2500 15380 2540
rect 10819 2499 10877 2500
rect 15235 2499 15293 2500
rect 10348 2456 10388 2499
rect 20995 2456 21053 2457
rect 7171 2416 7180 2456
rect 7220 2416 7468 2456
rect 7508 2416 7517 2456
rect 8803 2416 8812 2456
rect 8852 2416 9004 2456
rect 9044 2416 10252 2456
rect 10292 2416 10301 2456
rect 10348 2416 10540 2456
rect 10580 2416 11404 2456
rect 11444 2416 11453 2456
rect 11587 2416 11596 2456
rect 11636 2416 16876 2456
rect 16916 2416 16925 2456
rect 20140 2416 21004 2456
rect 21044 2416 21053 2456
rect 14563 2372 14621 2373
rect 20140 2372 20180 2416
rect 20995 2415 21053 2416
rect 2371 2332 2380 2372
rect 2420 2332 6028 2372
rect 6068 2332 6077 2372
rect 6280 2332 9484 2372
rect 9524 2332 9533 2372
rect 9676 2332 11500 2372
rect 11540 2332 11549 2372
rect 14478 2332 14572 2372
rect 14612 2332 14621 2372
rect 14947 2332 14956 2372
rect 14996 2332 20180 2372
rect 20515 2332 20524 2372
rect 20564 2332 20573 2372
rect 4099 2288 4157 2289
rect 9676 2288 9716 2332
rect 14563 2331 14621 2332
rect 9859 2288 9917 2289
rect 10147 2288 10205 2289
rect 15331 2288 15389 2289
rect 4014 2248 4108 2288
rect 4148 2248 4157 2288
rect 4919 2248 4928 2288
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 5296 2248 5305 2288
rect 5635 2248 5644 2288
rect 5684 2248 7276 2288
rect 7316 2248 7325 2288
rect 9667 2248 9676 2288
rect 9716 2248 9725 2288
rect 9859 2248 9868 2288
rect 9908 2248 10002 2288
rect 10147 2248 10156 2288
rect 10196 2248 11692 2288
rect 11732 2248 11741 2288
rect 13411 2248 13420 2288
rect 13460 2248 15340 2288
rect 15380 2248 15389 2288
rect 20039 2248 20048 2288
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20416 2248 20425 2288
rect 4099 2247 4157 2248
rect 9859 2247 9917 2248
rect 10147 2247 10205 2248
rect 15331 2247 15389 2248
rect 8803 2204 8861 2205
rect 11203 2204 11261 2205
rect 13219 2204 13277 2205
rect 20524 2204 20564 2332
rect 1891 2164 1900 2204
rect 1940 2164 4396 2204
rect 4436 2164 4445 2204
rect 4675 2164 4684 2204
rect 4724 2164 8812 2204
rect 8852 2164 8861 2204
rect 8995 2164 9004 2204
rect 9044 2164 10828 2204
rect 10868 2164 10877 2204
rect 11203 2164 11212 2204
rect 11252 2164 11308 2204
rect 11348 2164 11357 2204
rect 13219 2164 13228 2204
rect 13268 2164 15724 2204
rect 15764 2164 15773 2204
rect 20140 2164 20564 2204
rect 8803 2163 8861 2164
rect 11203 2163 11261 2164
rect 13219 2163 13277 2164
rect 0 2120 80 2140
rect 9283 2120 9341 2121
rect 11875 2120 11933 2121
rect 19555 2120 19613 2121
rect 19843 2120 19901 2121
rect 0 2080 748 2120
rect 788 2080 797 2120
rect 2500 2080 7564 2120
rect 7604 2080 8908 2120
rect 8948 2080 8957 2120
rect 9198 2080 9292 2120
rect 9332 2080 9484 2120
rect 9524 2080 9533 2120
rect 9580 2080 11692 2120
rect 11732 2080 11741 2120
rect 11875 2080 11884 2120
rect 11924 2080 15436 2120
rect 15476 2080 15485 2120
rect 16579 2080 16588 2120
rect 16628 2080 17164 2120
rect 17204 2080 17213 2120
rect 19555 2080 19564 2120
rect 19604 2080 19660 2120
rect 19700 2080 19709 2120
rect 19843 2080 19852 2120
rect 19892 2080 20044 2120
rect 20084 2080 20093 2120
rect 0 2060 80 2080
rect 2500 2036 2540 2080
rect 9283 2079 9341 2080
rect 1507 1996 1516 2036
rect 1556 1996 2540 2036
rect 5539 2036 5597 2037
rect 5731 2036 5789 2037
rect 9580 2036 9620 2080
rect 11875 2079 11933 2080
rect 19555 2079 19613 2080
rect 19843 2079 19901 2080
rect 5539 1996 5548 2036
rect 5588 1996 5740 2036
rect 5780 1996 9620 2036
rect 10243 1996 10252 2036
rect 10292 1996 12172 2036
rect 12212 1996 16012 2036
rect 16052 1996 16061 2036
rect 5539 1995 5597 1996
rect 5731 1995 5789 1996
rect 3619 1952 3677 1953
rect 5923 1952 5981 1953
rect 9187 1952 9245 1953
rect 10051 1952 10109 1953
rect 11587 1952 11645 1953
rect 18115 1952 18173 1953
rect 2659 1912 2668 1952
rect 2708 1912 3628 1952
rect 3668 1912 3677 1952
rect 4003 1912 4012 1952
rect 4052 1912 5780 1952
rect 5838 1912 5932 1952
rect 5972 1912 5981 1952
rect 7651 1912 7660 1952
rect 7700 1912 8428 1952
rect 8468 1912 8477 1952
rect 8995 1912 9004 1952
rect 9044 1912 9196 1952
rect 9236 1912 9245 1952
rect 9379 1912 9388 1952
rect 9428 1912 10004 1952
rect 3619 1911 3677 1912
rect 1987 1868 2045 1869
rect 5635 1868 5693 1869
rect 835 1828 844 1868
rect 884 1828 1228 1868
rect 1268 1828 1277 1868
rect 1902 1828 1996 1868
rect 2036 1828 2045 1868
rect 5059 1828 5068 1868
rect 5108 1828 5644 1868
rect 5684 1828 5693 1868
rect 5740 1868 5780 1912
rect 5923 1911 5981 1912
rect 9187 1911 9245 1912
rect 9964 1868 10004 1912
rect 10051 1912 10060 1952
rect 10100 1912 11596 1952
rect 11636 1912 11645 1952
rect 14755 1912 14764 1952
rect 14804 1912 15052 1952
rect 15092 1912 16972 1952
rect 17012 1912 17021 1952
rect 17923 1912 17932 1952
rect 17972 1912 18124 1952
rect 18164 1912 18173 1952
rect 10051 1911 10109 1912
rect 11587 1911 11645 1912
rect 18115 1911 18173 1912
rect 19363 1952 19421 1953
rect 19939 1952 19997 1953
rect 19363 1912 19372 1952
rect 19412 1912 19756 1952
rect 19796 1912 19805 1952
rect 19854 1912 19948 1952
rect 19988 1912 19997 1952
rect 19363 1911 19421 1912
rect 19939 1911 19997 1912
rect 5740 1828 9676 1868
rect 9716 1828 9725 1868
rect 9964 1828 10060 1868
rect 10100 1828 10924 1868
rect 10964 1828 10973 1868
rect 11203 1828 11212 1868
rect 11252 1828 14860 1868
rect 14900 1828 14909 1868
rect 1987 1827 2045 1828
rect 5635 1827 5693 1828
rect 0 1784 80 1804
rect 2371 1784 2429 1785
rect 20140 1784 20180 2164
rect 0 1744 2380 1784
rect 2420 1744 2429 1784
rect 4867 1744 4876 1784
rect 4916 1744 12172 1784
rect 12212 1744 12221 1784
rect 13987 1744 13996 1784
rect 14036 1744 16492 1784
rect 16532 1744 16541 1784
rect 20035 1744 20044 1784
rect 20084 1744 20180 1784
rect 0 1724 80 1744
rect 2371 1743 2429 1744
rect 1411 1700 1469 1701
rect 1326 1660 1420 1700
rect 1460 1660 1469 1700
rect 2179 1660 2188 1700
rect 2228 1660 2237 1700
rect 4387 1660 4396 1700
rect 4436 1660 9388 1700
rect 9428 1660 9437 1700
rect 9667 1660 9676 1700
rect 9716 1660 11788 1700
rect 11828 1660 11837 1700
rect 11971 1660 11980 1700
rect 12020 1660 17356 1700
rect 17396 1660 17405 1700
rect 1411 1659 1469 1660
rect 2188 1616 2228 1660
rect 2188 1576 10444 1616
rect 10484 1576 10493 1616
rect 11320 1576 15628 1616
rect 15668 1576 17452 1616
rect 17492 1576 17501 1616
rect 9955 1532 10013 1533
rect 11203 1532 11261 1533
rect 3679 1492 3688 1532
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 4056 1492 4065 1532
rect 5731 1492 5740 1532
rect 5780 1492 9964 1532
rect 10004 1492 10540 1532
rect 10580 1492 11212 1532
rect 11252 1492 11261 1532
rect 9955 1491 10013 1492
rect 11203 1491 11261 1492
rect 0 1448 80 1468
rect 1027 1448 1085 1449
rect 11320 1448 11360 1576
rect 17539 1532 17597 1533
rect 13891 1492 13900 1532
rect 13940 1492 17548 1532
rect 17588 1492 17597 1532
rect 18799 1492 18808 1532
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 19176 1492 19185 1532
rect 17539 1491 17597 1492
rect 0 1408 1036 1448
rect 1076 1408 1085 1448
rect 1603 1408 1612 1448
rect 1652 1408 11360 1448
rect 12268 1408 17164 1448
rect 17204 1408 17213 1448
rect 0 1388 80 1408
rect 1027 1407 1085 1408
rect 12268 1364 12308 1408
rect 15907 1364 15965 1365
rect 1795 1324 1804 1364
rect 1844 1324 9044 1364
rect 9379 1324 9388 1364
rect 9428 1324 12308 1364
rect 12364 1324 13268 1364
rect 2563 1280 2621 1281
rect 3331 1280 3389 1281
rect 3715 1280 3773 1281
rect 6403 1280 6461 1281
rect 6787 1280 6845 1281
rect 6979 1280 7037 1281
rect 2563 1240 2572 1280
rect 2612 1240 2706 1280
rect 3139 1240 3148 1280
rect 3188 1240 3340 1280
rect 3380 1240 3389 1280
rect 3630 1240 3724 1280
rect 3764 1240 3773 1280
rect 4099 1240 4108 1280
rect 4148 1240 5836 1280
rect 5876 1240 5885 1280
rect 6318 1240 6412 1280
rect 6452 1240 6461 1280
rect 6702 1240 6796 1280
rect 6836 1240 6845 1280
rect 6894 1240 6988 1280
rect 7028 1240 7037 1280
rect 2563 1239 2621 1240
rect 3331 1239 3389 1240
rect 3715 1239 3773 1240
rect 6403 1239 6461 1240
rect 6787 1239 6845 1240
rect 6979 1239 7037 1240
rect 7171 1280 7229 1281
rect 8131 1280 8189 1281
rect 8323 1280 8381 1281
rect 8515 1280 8573 1281
rect 9004 1280 9044 1324
rect 12364 1280 12404 1324
rect 12547 1280 12605 1281
rect 7171 1240 7180 1280
rect 7220 1240 7314 1280
rect 7372 1240 7756 1280
rect 7796 1240 7805 1280
rect 8131 1240 8140 1280
rect 8180 1240 8274 1280
rect 8323 1240 8332 1280
rect 8372 1240 8466 1280
rect 8515 1240 8524 1280
rect 8564 1240 8658 1280
rect 9004 1240 10484 1280
rect 10531 1240 10540 1280
rect 10580 1240 11212 1280
rect 11252 1240 11261 1280
rect 11320 1240 12404 1280
rect 12462 1240 12556 1280
rect 12596 1240 12605 1280
rect 7171 1239 7229 1240
rect 931 1196 989 1197
rect 76 1156 940 1196
rect 980 1156 989 1196
rect 76 1132 116 1156
rect 931 1155 989 1156
rect 3427 1196 3485 1197
rect 5443 1196 5501 1197
rect 5635 1196 5693 1197
rect 7372 1196 7412 1240
rect 8131 1239 8189 1240
rect 8323 1239 8381 1240
rect 8515 1239 8573 1240
rect 10444 1196 10484 1240
rect 10915 1196 10973 1197
rect 3427 1156 3436 1196
rect 3476 1156 3532 1196
rect 3572 1156 3581 1196
rect 4012 1156 5452 1196
rect 5492 1156 5501 1196
rect 5550 1156 5644 1196
rect 5684 1156 5693 1196
rect 6115 1156 6124 1196
rect 6164 1156 7412 1196
rect 7468 1156 9484 1196
rect 9524 1156 9533 1196
rect 10444 1156 10924 1196
rect 10964 1156 10973 1196
rect 3427 1155 3485 1156
rect 0 1072 116 1132
rect 4012 1112 4052 1156
rect 5443 1155 5501 1156
rect 5635 1155 5693 1156
rect 460 1072 4052 1112
rect 4099 1112 4157 1113
rect 5059 1112 5117 1113
rect 7468 1112 7508 1156
rect 10915 1155 10973 1156
rect 11107 1196 11165 1197
rect 11320 1196 11360 1240
rect 12547 1239 12605 1240
rect 12739 1280 12797 1281
rect 13123 1280 13181 1281
rect 12739 1240 12748 1280
rect 12788 1240 12882 1280
rect 12931 1240 12940 1280
rect 12980 1240 13132 1280
rect 13172 1240 13181 1280
rect 12739 1239 12797 1240
rect 13123 1239 13181 1240
rect 13228 1196 13268 1324
rect 15907 1324 15916 1364
rect 15956 1324 18548 1364
rect 15907 1323 15965 1324
rect 13507 1280 13565 1281
rect 13422 1240 13516 1280
rect 13556 1240 13565 1280
rect 13507 1239 13565 1240
rect 13699 1280 13757 1281
rect 14659 1280 14717 1281
rect 15427 1280 15485 1281
rect 15619 1280 15677 1281
rect 13699 1240 13708 1280
rect 13748 1240 13842 1280
rect 14574 1240 14668 1280
rect 14708 1240 14717 1280
rect 15342 1240 15436 1280
rect 15476 1240 15485 1280
rect 15534 1240 15628 1280
rect 15668 1240 15677 1280
rect 13699 1239 13757 1240
rect 14659 1239 14717 1240
rect 15427 1239 15485 1240
rect 15619 1239 15677 1240
rect 17443 1280 17501 1281
rect 17731 1280 17789 1281
rect 17443 1240 17452 1280
rect 17492 1240 17548 1280
rect 17588 1240 17597 1280
rect 17646 1240 17740 1280
rect 17780 1240 17789 1280
rect 17443 1239 17501 1240
rect 17731 1239 17789 1240
rect 18211 1280 18269 1281
rect 18508 1280 18548 1324
rect 18211 1240 18220 1280
rect 18260 1240 18316 1280
rect 18356 1240 18365 1280
rect 18508 1240 18988 1280
rect 19028 1240 19037 1280
rect 18211 1239 18269 1240
rect 18403 1196 18461 1197
rect 11107 1156 11116 1196
rect 11156 1156 11360 1196
rect 11491 1156 11500 1196
rect 11540 1156 12844 1196
rect 12884 1156 12893 1196
rect 13228 1156 14284 1196
rect 14324 1156 15380 1196
rect 11107 1155 11165 1156
rect 8611 1112 8669 1113
rect 9571 1112 9629 1113
rect 15340 1112 15380 1156
rect 18403 1156 18412 1196
rect 18452 1156 18508 1196
rect 18548 1156 18557 1196
rect 18403 1155 18461 1156
rect 4099 1072 4108 1112
rect 4148 1072 4242 1112
rect 4780 1072 5068 1112
rect 5108 1072 5117 1112
rect 5251 1072 5260 1112
rect 5300 1072 7508 1112
rect 7555 1072 7564 1112
rect 7604 1072 8620 1112
rect 8660 1072 8669 1112
rect 9091 1072 9100 1112
rect 9140 1072 9388 1112
rect 9428 1072 9437 1112
rect 9571 1072 9580 1112
rect 9620 1072 11212 1112
rect 11252 1072 11261 1112
rect 12451 1072 12460 1112
rect 12500 1072 15244 1112
rect 15284 1072 15293 1112
rect 15340 1072 19084 1112
rect 19124 1072 19133 1112
rect 0 1052 80 1072
rect 460 1028 500 1072
rect 4099 1071 4157 1072
rect 4780 1028 4820 1072
rect 5059 1071 5117 1072
rect 8611 1071 8669 1072
rect 9571 1071 9629 1072
rect 8035 1028 8093 1029
rect 12460 1028 12500 1072
rect 13795 1028 13853 1029
rect 172 988 500 1028
rect 1987 988 1996 1028
rect 2036 988 4820 1028
rect 4867 988 4876 1028
rect 4916 988 5068 1028
rect 5108 988 8044 1028
rect 8084 988 8093 1028
rect 9187 988 9196 1028
rect 9236 988 9964 1028
rect 10004 988 10013 1028
rect 10060 988 12500 1028
rect 13315 988 13324 1028
rect 13364 988 13804 1028
rect 13844 988 13853 1028
rect 14179 988 14188 1028
rect 14228 988 17068 1028
rect 17108 988 17117 1028
rect 17827 988 17836 1028
rect 17876 988 19276 1028
rect 19316 988 19325 1028
rect 0 776 80 796
rect 172 776 212 988
rect 8035 987 8093 988
rect 4291 944 4349 945
rect 7363 944 7421 945
rect 7747 944 7805 945
rect 10060 944 10100 988
rect 13795 987 13853 988
rect 14275 944 14333 945
rect 17836 944 17876 988
rect 259 904 268 944
rect 308 904 2540 944
rect 4206 904 4300 944
rect 4340 904 4349 944
rect 5443 904 5452 944
rect 5492 904 5501 944
rect 7278 904 7372 944
rect 7412 904 7421 944
rect 7662 904 7756 944
rect 7796 904 7805 944
rect 8035 904 8044 944
rect 8084 904 8236 944
rect 8276 904 10100 944
rect 14190 904 14284 944
rect 14324 904 14333 944
rect 14563 904 14572 944
rect 14612 904 14956 944
rect 14996 904 15005 944
rect 16483 904 16492 944
rect 16532 904 16780 944
rect 16820 904 17876 944
rect 2500 860 2540 904
rect 4291 903 4349 904
rect 5452 860 5492 904
rect 7363 903 7421 904
rect 7747 903 7805 904
rect 14275 903 14333 904
rect 5923 860 5981 861
rect 10915 860 10973 861
rect 11107 860 11165 861
rect 18691 860 18749 861
rect 20515 860 20573 861
rect 2500 820 5492 860
rect 5827 820 5836 860
rect 5876 820 5932 860
rect 5972 820 5981 860
rect 7459 820 7468 860
rect 7508 820 10252 860
rect 10292 820 10301 860
rect 10830 820 10924 860
rect 10964 820 10973 860
rect 11022 820 11116 860
rect 11156 820 11165 860
rect 5923 819 5981 820
rect 10915 819 10973 820
rect 11107 819 11165 820
rect 11320 820 11404 860
rect 11444 820 11453 860
rect 18606 820 18700 860
rect 18740 820 18749 860
rect 18883 820 18892 860
rect 18932 820 20524 860
rect 20564 820 20573 860
rect 4675 776 4733 777
rect 11320 776 11360 820
rect 18691 819 18749 820
rect 20515 819 20573 820
rect 0 736 212 776
rect 4590 736 4684 776
rect 4724 736 4733 776
rect 4919 736 4928 776
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 5296 736 5305 776
rect 5347 736 5356 776
rect 5396 736 11360 776
rect 20039 736 20048 776
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20416 736 20425 776
rect 0 716 80 736
rect 4675 735 4733 736
rect 6211 692 6269 693
rect 7939 692 7997 693
rect 19267 692 19325 693
rect 4387 652 4396 692
rect 4436 652 6220 692
rect 6260 652 7276 692
rect 7316 652 7325 692
rect 7854 652 7948 692
rect 7988 652 7997 692
rect 8899 652 8908 692
rect 8948 652 16876 692
rect 16916 652 16925 692
rect 19182 652 19276 692
rect 19316 652 19325 692
rect 6211 651 6269 652
rect 7939 651 7997 652
rect 19267 651 19325 652
rect 4483 608 4541 609
rect 5347 608 5405 609
rect 3907 568 3916 608
rect 3956 568 4492 608
rect 4532 568 4541 608
rect 5059 568 5068 608
rect 5108 568 5356 608
rect 5396 568 5405 608
rect 7651 568 7660 608
rect 7700 568 11212 608
rect 11252 568 11261 608
rect 11320 568 15244 608
rect 15284 568 15293 608
rect 4483 567 4541 568
rect 5347 567 5405 568
rect 9763 524 9821 525
rect 5539 484 5548 524
rect 5588 484 9388 524
rect 9428 484 9437 524
rect 9763 484 9772 524
rect 9812 484 11116 524
rect 11156 484 11165 524
rect 9763 483 9821 484
rect 0 440 80 460
rect 6019 440 6077 441
rect 11320 440 11360 568
rect 15043 524 15101 525
rect 12355 484 12364 524
rect 12404 484 14764 524
rect 14804 484 14813 524
rect 15043 484 15052 524
rect 15092 484 19468 524
rect 19508 484 19517 524
rect 15043 483 15101 484
rect 0 400 652 440
rect 692 400 701 440
rect 2371 400 2380 440
rect 2420 400 6028 440
rect 6068 400 6077 440
rect 0 380 80 400
rect 6019 399 6077 400
rect 6124 400 11360 440
rect 13603 440 13661 441
rect 13603 400 13612 440
rect 13652 400 17932 440
rect 17972 400 17981 440
rect 6124 356 6164 400
rect 13603 399 13661 400
rect 6595 356 6653 357
rect 1027 316 1036 356
rect 1076 316 4876 356
rect 4916 316 4925 356
rect 4972 316 6164 356
rect 6510 316 6604 356
rect 6644 316 6653 356
rect 1123 272 1181 273
rect 4771 272 4829 273
rect 4972 272 5012 316
rect 6595 315 6653 316
rect 6883 356 6941 357
rect 6883 316 6892 356
rect 6932 316 9004 356
rect 9044 316 13036 356
rect 13076 316 15820 356
rect 15860 316 15869 356
rect 6883 315 6941 316
rect 5827 272 5885 273
rect 11299 272 11357 273
rect 16291 272 16349 273
rect 1123 232 1132 272
rect 1172 232 4492 272
rect 4532 232 4541 272
rect 4771 232 4780 272
rect 4820 232 5012 272
rect 5443 232 5452 272
rect 5492 232 5836 272
rect 5876 232 5885 272
rect 7267 232 7276 272
rect 7316 232 11252 272
rect 1123 231 1181 232
rect 4771 231 4829 232
rect 5827 231 5885 232
rect 5251 188 5309 189
rect 9763 188 9821 189
rect 3043 148 3052 188
rect 3092 148 3101 188
rect 5166 148 5260 188
rect 5300 148 5309 188
rect 0 104 80 124
rect 259 104 317 105
rect 0 64 268 104
rect 308 64 317 104
rect 3052 104 3092 148
rect 5251 147 5309 148
rect 5836 148 9772 188
rect 9812 148 9821 188
rect 5836 104 5876 148
rect 9763 147 9821 148
rect 6019 104 6077 105
rect 3052 64 5876 104
rect 5934 64 6028 104
rect 6068 64 6077 104
rect 11212 104 11252 232
rect 11299 232 11308 272
rect 11348 232 16108 272
rect 16148 232 16157 272
rect 16291 232 16300 272
rect 16340 232 18124 272
rect 18164 232 18173 272
rect 11299 231 11357 232
rect 16291 231 16349 232
rect 11299 148 11308 188
rect 11348 148 16588 188
rect 16628 148 16637 188
rect 16771 104 16829 105
rect 11212 64 16780 104
rect 16820 64 16829 104
rect 0 44 80 64
rect 259 63 317 64
rect 6019 63 6077 64
rect 16771 63 16829 64
<< via3 >>
rect 1228 42820 1268 42860
rect 4780 42652 4820 42692
rect 18508 42652 18548 42692
rect 10252 42316 10292 42356
rect 2860 42232 2900 42272
rect 4684 42148 4724 42188
rect 10156 42148 10196 42188
rect 15052 42232 15092 42272
rect 17548 41980 17588 42020
rect 17740 41980 17780 42020
rect 4204 41896 4244 41936
rect 2956 41812 2996 41852
rect 7852 41812 7892 41852
rect 15628 41812 15668 41852
rect 17836 41728 17876 41768
rect 12172 41644 12212 41684
rect 4928 41560 4968 41600
rect 5010 41560 5050 41600
rect 5092 41560 5132 41600
rect 5174 41560 5214 41600
rect 5256 41560 5296 41600
rect 12556 41560 12596 41600
rect 16780 41560 16820 41600
rect 1612 41392 1652 41432
rect 2572 41392 2612 41432
rect 9388 41392 9428 41432
rect 16972 41560 17012 41600
rect 18124 41560 18164 41600
rect 20048 41560 20088 41600
rect 20130 41560 20170 41600
rect 20212 41560 20252 41600
rect 20294 41560 20334 41600
rect 20376 41560 20416 41600
rect 2380 41308 2420 41348
rect 13900 41392 13940 41432
rect 3340 41224 3380 41264
rect 4108 41224 4148 41264
rect 1324 41140 1364 41180
rect 15244 41392 15284 41432
rect 17548 41308 17588 41348
rect 18028 41308 18068 41348
rect 12364 41224 12404 41264
rect 15340 41224 15380 41264
rect 14764 41056 14804 41096
rect 3532 40972 3572 41012
rect 4876 40972 4916 41012
rect 17164 40972 17204 41012
rect 17548 40972 17588 41012
rect 17932 40972 17972 41012
rect 18316 40972 18356 41012
rect 18700 40972 18740 41012
rect 3688 40804 3728 40844
rect 3770 40804 3810 40844
rect 3852 40804 3892 40844
rect 3934 40804 3974 40844
rect 4016 40804 4056 40844
rect 17644 40888 17684 40928
rect 17260 40804 17300 40844
rect 18808 40804 18848 40844
rect 18890 40804 18930 40844
rect 18972 40804 19012 40844
rect 19054 40804 19094 40844
rect 19136 40804 19176 40844
rect 14572 40720 14612 40760
rect 14380 40636 14420 40676
rect 14764 40552 14804 40592
rect 1420 40468 1460 40508
rect 5644 40468 5684 40508
rect 17068 40552 17108 40592
rect 17548 40552 17588 40592
rect 17932 40552 17972 40592
rect 10732 40468 10772 40508
rect 18604 40468 18644 40508
rect 1804 40384 1844 40424
rect 10444 40398 10483 40424
rect 10483 40398 10484 40424
rect 10444 40384 10484 40398
rect 16396 40384 16436 40424
rect 18892 40384 18932 40424
rect 19756 40384 19796 40424
rect 1036 40300 1076 40340
rect 7276 40300 7316 40340
rect 11596 40300 11636 40340
rect 1900 40216 1940 40256
rect 3436 40216 3476 40256
rect 4876 40216 4916 40256
rect 20620 40300 20660 40340
rect 19468 40216 19508 40256
rect 1420 40132 1460 40172
rect 7372 40132 7412 40172
rect 10060 40132 10100 40172
rect 3436 40048 3476 40088
rect 4300 40048 4340 40088
rect 4928 40048 4968 40088
rect 5010 40048 5050 40088
rect 5092 40048 5132 40088
rect 5174 40048 5214 40088
rect 5256 40048 5296 40088
rect 8332 40048 8372 40088
rect 10924 40048 10964 40088
rect 14284 40048 14324 40088
rect 16684 40048 16724 40088
rect 18508 40048 18548 40088
rect 20048 40048 20088 40088
rect 20130 40048 20170 40088
rect 20212 40048 20252 40088
rect 20294 40048 20334 40088
rect 20376 40048 20416 40088
rect 12460 39964 12500 40004
rect 16588 39880 16628 39920
rect 3628 39796 3668 39836
rect 11596 39796 11636 39836
rect 17836 39796 17876 39836
rect 1708 39712 1748 39752
rect 6220 39712 6260 39752
rect 12940 39712 12980 39752
rect 15916 39712 15956 39752
rect 16876 39712 16916 39752
rect 18508 39712 18548 39752
rect 3148 39628 3188 39668
rect 4492 39628 4532 39668
rect 4684 39628 4724 39668
rect 5740 39628 5780 39668
rect 6124 39628 6164 39668
rect 13900 39628 13940 39668
rect 16588 39628 16628 39668
rect 18220 39628 18260 39668
rect 14764 39544 14804 39584
rect 9868 39460 9908 39500
rect 14572 39460 14612 39500
rect 16108 39460 16148 39500
rect 18412 39460 18452 39500
rect 19372 39460 19412 39500
rect 7180 39376 7220 39416
rect 1996 39292 2036 39332
rect 3688 39292 3728 39332
rect 3770 39292 3810 39332
rect 3852 39292 3892 39332
rect 3934 39292 3974 39332
rect 4016 39292 4056 39332
rect 1708 39208 1748 39248
rect 6028 39208 6068 39248
rect 10636 39208 10676 39248
rect 1900 39124 1940 39164
rect 2764 39124 2804 39164
rect 3052 39124 3092 39164
rect 4012 39124 4052 39164
rect 11116 39208 11156 39248
rect 11500 39292 11540 39332
rect 18808 39292 18848 39332
rect 18890 39292 18930 39332
rect 18972 39292 19012 39332
rect 19054 39292 19094 39332
rect 19136 39292 19176 39332
rect 19276 39292 19316 39332
rect 12844 39208 12884 39248
rect 18124 39208 18164 39248
rect 18412 39208 18452 39248
rect 2092 39040 2132 39080
rect 3340 39040 3380 39080
rect 4300 39040 4340 39080
rect 7276 39040 7316 39080
rect 15820 39040 15860 39080
rect 17932 39040 17972 39080
rect 19276 39040 19316 39080
rect 19564 39040 19604 39080
rect 556 38956 596 38996
rect 2380 38956 2420 38996
rect 4108 38956 4148 38996
rect 6700 38956 6740 38996
rect 8044 38956 8084 38996
rect 21004 39040 21044 39080
rect 8236 38956 8276 38996
rect 10252 38956 10292 38996
rect 11020 38956 11060 38996
rect 11212 38956 11252 38996
rect 14860 38956 14900 38996
rect 17260 38956 17300 38996
rect 6412 38872 6452 38912
rect 8620 38872 8660 38912
rect 4012 38788 4052 38828
rect 13996 38788 14036 38828
rect 1132 38704 1172 38744
rect 7084 38704 7124 38744
rect 8236 38704 8276 38744
rect 10252 38704 10292 38744
rect 21292 38788 21332 38828
rect 18028 38704 18068 38744
rect 21388 38704 21428 38744
rect 2092 38536 2132 38576
rect 2956 38536 2996 38576
rect 11212 38620 11252 38660
rect 20908 38620 20948 38660
rect 4204 38536 4244 38576
rect 4928 38536 4968 38576
rect 5010 38536 5050 38576
rect 5092 38536 5132 38576
rect 5174 38536 5214 38576
rect 5256 38536 5296 38576
rect 8716 38536 8756 38576
rect 10060 38536 10100 38576
rect 12652 38536 12692 38576
rect 20048 38536 20088 38576
rect 20130 38536 20170 38576
rect 20212 38536 20252 38576
rect 20294 38536 20334 38576
rect 20376 38536 20416 38576
rect 15244 38452 15284 38492
rect 2188 38284 2228 38324
rect 7372 38284 7412 38324
rect 16876 38452 16916 38492
rect 19660 38452 19700 38492
rect 19852 38452 19892 38492
rect 16012 38368 16052 38408
rect 8044 38284 8084 38324
rect 9772 38284 9812 38324
rect 4588 38200 4628 38240
rect 5548 38200 5588 38240
rect 7660 38200 7700 38240
rect 8716 38200 8756 38240
rect 17644 38200 17684 38240
rect 19276 38200 19316 38240
rect 19948 38200 19988 38240
rect 2380 38116 2420 38156
rect 2572 38116 2612 38156
rect 3340 38116 3380 38156
rect 9964 38116 10004 38156
rect 13420 38116 13460 38156
rect 4876 38032 4916 38072
rect 8812 38032 8852 38072
rect 11500 38032 11540 38072
rect 16300 38116 16340 38156
rect 19852 38116 19892 38156
rect 19372 38032 19412 38072
rect 1516 37948 1556 37988
rect 2956 37864 2996 37904
rect 2764 37780 2804 37820
rect 940 37696 980 37736
rect 3688 37780 3728 37820
rect 3770 37780 3810 37820
rect 3852 37780 3892 37820
rect 3934 37780 3974 37820
rect 4016 37780 4056 37820
rect 9484 37780 9524 37820
rect 11116 37780 11156 37820
rect 3052 37696 3092 37736
rect 12844 37864 12884 37904
rect 15724 37864 15764 37904
rect 17452 37864 17492 37904
rect 13036 37780 13076 37820
rect 14188 37780 14228 37820
rect 16492 37780 16532 37820
rect 18808 37780 18848 37820
rect 18890 37780 18930 37820
rect 18972 37780 19012 37820
rect 19054 37780 19094 37820
rect 19136 37780 19176 37820
rect 11308 37696 11348 37736
rect 2572 37612 2612 37652
rect 9772 37612 9812 37652
rect 12652 37612 12692 37652
rect 15436 37612 15476 37652
rect 16492 37696 16532 37736
rect 16876 37696 16916 37736
rect 3724 37528 3764 37568
rect 11308 37528 11348 37568
rect 13324 37528 13364 37568
rect 19276 37528 19316 37568
rect 21196 37528 21236 37568
rect 1324 37444 1364 37484
rect 4108 37444 4148 37484
rect 4492 37444 4532 37484
rect 5644 37444 5684 37484
rect 8716 37444 8756 37484
rect 12364 37444 12404 37484
rect 15244 37444 15284 37484
rect 19372 37444 19412 37484
rect 2764 37360 2804 37400
rect 3244 37360 3284 37400
rect 9484 37360 9524 37400
rect 11692 37360 11732 37400
rect 17452 37360 17492 37400
rect 5644 37276 5684 37316
rect 5932 37276 5972 37316
rect 8908 37276 8948 37316
rect 15532 37276 15572 37316
rect 16492 37276 16532 37316
rect 17356 37276 17396 37316
rect 1132 37192 1172 37232
rect 5836 37108 5876 37148
rect 6028 37108 6068 37148
rect 4928 37024 4968 37064
rect 5010 37024 5050 37064
rect 5092 37024 5132 37064
rect 5174 37024 5214 37064
rect 5256 37024 5296 37064
rect 16204 37024 16244 37064
rect 16876 37192 16916 37232
rect 20048 37024 20088 37064
rect 20130 37024 20170 37064
rect 20212 37024 20252 37064
rect 20294 37024 20334 37064
rect 20376 37024 20416 37064
rect 20812 37024 20852 37064
rect 19948 36940 19988 36980
rect 2284 36856 2324 36896
rect 2956 36856 2996 36896
rect 8140 36856 8180 36896
rect 15628 36856 15668 36896
rect 16300 36772 16340 36812
rect 5836 36688 5876 36728
rect 7468 36688 7508 36728
rect 8044 36688 8084 36728
rect 8620 36688 8660 36728
rect 9100 36688 9140 36728
rect 16492 36772 16532 36812
rect 15436 36688 15476 36728
rect 16876 36688 16916 36728
rect 5452 36604 5492 36644
rect 14860 36604 14900 36644
rect 17452 36772 17492 36812
rect 19276 36604 19316 36644
rect 1324 36520 1364 36560
rect 5260 36520 5300 36560
rect 9292 36520 9332 36560
rect 10828 36520 10868 36560
rect 11884 36520 11924 36560
rect 15244 36520 15284 36560
rect 20620 36520 20660 36560
rect 1900 36436 1940 36476
rect 10924 36436 10964 36476
rect 16876 36436 16916 36476
rect 5740 36352 5780 36392
rect 17356 36352 17396 36392
rect 19468 36352 19508 36392
rect 3688 36268 3728 36308
rect 3770 36268 3810 36308
rect 3852 36268 3892 36308
rect 3934 36268 3974 36308
rect 4016 36268 4056 36308
rect 17644 36268 17684 36308
rect 18808 36268 18848 36308
rect 18890 36268 18930 36308
rect 18972 36268 19012 36308
rect 19054 36268 19094 36308
rect 19136 36268 19176 36308
rect 8236 36184 8276 36224
rect 1516 36016 1556 36056
rect 2860 36100 2900 36140
rect 4780 36100 4820 36140
rect 8332 36100 8372 36140
rect 7564 36016 7604 36056
rect 4780 35932 4820 35972
rect 10156 35932 10196 35972
rect 17452 35932 17492 35972
rect 7372 35848 7412 35888
rect 13132 35848 13172 35888
rect 19276 35848 19316 35888
rect 19564 35848 19604 35888
rect 844 35764 884 35804
rect 13228 35764 13268 35804
rect 14764 35764 14804 35804
rect 18700 35764 18740 35804
rect 460 35680 500 35720
rect 9964 35680 10004 35720
rect 1324 35596 1364 35636
rect 4396 35596 4436 35636
rect 8236 35596 8276 35636
rect 13324 35596 13364 35636
rect 16012 35596 16052 35636
rect 17836 35596 17876 35636
rect 18124 35596 18164 35636
rect 19852 35596 19892 35636
rect 3436 35512 3476 35552
rect 4928 35512 4968 35552
rect 5010 35512 5050 35552
rect 5092 35512 5132 35552
rect 5174 35512 5214 35552
rect 5256 35512 5296 35552
rect 20048 35512 20088 35552
rect 20130 35512 20170 35552
rect 20212 35512 20252 35552
rect 20294 35512 20334 35552
rect 20376 35512 20416 35552
rect 1804 35428 1844 35468
rect 2092 35428 2132 35468
rect 3052 35428 3092 35468
rect 15052 35428 15092 35468
rect 3340 35344 3380 35384
rect 1804 35260 1844 35300
rect 2476 35260 2516 35300
rect 18028 35428 18068 35468
rect 3628 35344 3668 35384
rect 16300 35344 16340 35384
rect 17356 35344 17396 35384
rect 5356 35260 5396 35300
rect 15148 35260 15188 35300
rect 15628 35260 15668 35300
rect 18412 35260 18452 35300
rect 2380 35176 2420 35216
rect 6316 35176 6356 35216
rect 6508 35176 6548 35216
rect 9676 35176 9716 35216
rect 11212 35176 11252 35216
rect 11692 35176 11732 35216
rect 13516 35176 13556 35216
rect 14092 35176 14132 35216
rect 18220 35176 18260 35216
rect 4108 35092 4148 35132
rect 14572 35092 14612 35132
rect 13228 35008 13268 35048
rect 18124 35008 18164 35048
rect 6124 34924 6164 34964
rect 16684 34924 16724 34964
rect 18508 34924 18548 34964
rect 76 34840 116 34880
rect 6316 34840 6356 34880
rect 19468 34840 19508 34880
rect 3688 34756 3728 34796
rect 3770 34756 3810 34796
rect 3852 34756 3892 34796
rect 3934 34756 3974 34796
rect 4016 34756 4056 34796
rect 18508 34756 18548 34796
rect 18808 34756 18848 34796
rect 18890 34756 18930 34796
rect 18972 34756 19012 34796
rect 19054 34756 19094 34796
rect 19136 34756 19176 34796
rect 6604 34672 6644 34712
rect 15436 34672 15476 34712
rect 4012 34588 4052 34628
rect 4492 34588 4532 34628
rect 16588 34588 16628 34628
rect 19564 34588 19604 34628
rect 1708 34504 1748 34544
rect 6508 34504 6548 34544
rect 8908 34420 8948 34460
rect 19756 34420 19796 34460
rect 1612 34336 1652 34376
rect 4108 34336 4148 34376
rect 6892 34336 6932 34376
rect 7372 34336 7412 34376
rect 7660 34336 7700 34376
rect 9196 34336 9236 34376
rect 12364 34336 12404 34376
rect 13516 34336 13556 34376
rect 14476 34336 14516 34376
rect 15628 34336 15668 34376
rect 18220 34336 18260 34376
rect 5356 34252 5396 34292
rect 18412 34252 18452 34292
rect 10060 34168 10100 34208
rect 13324 34168 13364 34208
rect 14188 34084 14228 34124
rect 4928 34000 4968 34040
rect 5010 34000 5050 34040
rect 5092 34000 5132 34040
rect 5174 34000 5214 34040
rect 5256 34000 5296 34040
rect 7276 34000 7316 34040
rect 2956 33916 2996 33956
rect 15052 34000 15092 34040
rect 15436 34000 15476 34040
rect 16012 34084 16052 34124
rect 17836 34084 17876 34124
rect 16492 34000 16532 34040
rect 17644 34000 17684 34040
rect 20048 34000 20088 34040
rect 20130 34000 20170 34040
rect 20212 34000 20252 34040
rect 20294 34000 20334 34040
rect 20376 34000 20416 34040
rect 11116 33916 11156 33956
rect 18508 33916 18548 33956
rect 1420 33832 1460 33872
rect 2764 33748 2804 33788
rect 8716 33748 8756 33788
rect 1228 33664 1268 33704
rect 9964 33664 10004 33704
rect 11788 33664 11828 33704
rect 14284 33664 14324 33704
rect 15244 33664 15284 33704
rect 16012 33664 16052 33704
rect 18124 33664 18164 33704
rect 2764 33580 2804 33620
rect 5548 33580 5588 33620
rect 3628 33496 3668 33536
rect 13900 33580 13940 33620
rect 16300 33580 16340 33620
rect 19852 33580 19892 33620
rect 7180 33496 7220 33536
rect 19468 33496 19508 33536
rect 2956 33412 2996 33452
rect 11308 33412 11348 33452
rect 3436 33328 3476 33368
rect 3688 33244 3728 33284
rect 3770 33244 3810 33284
rect 3852 33244 3892 33284
rect 3934 33244 3974 33284
rect 4016 33244 4056 33284
rect 13132 33244 13172 33284
rect 14476 33244 14516 33284
rect 20812 33496 20852 33536
rect 20620 33412 20660 33452
rect 18220 33244 18260 33284
rect 18808 33244 18848 33284
rect 18890 33244 18930 33284
rect 18972 33244 19012 33284
rect 19054 33244 19094 33284
rect 19136 33244 19176 33284
rect 1228 33160 1268 33200
rect 10636 33160 10676 33200
rect 15916 33076 15956 33116
rect 19276 33076 19316 33116
rect 3340 32992 3380 33032
rect 4204 32992 4244 33032
rect 17644 32992 17684 33032
rect 3916 32908 3956 32948
rect 20716 32992 20756 33032
rect 4108 32908 4148 32948
rect 15148 32908 15188 32948
rect 16684 32908 16724 32948
rect 940 32824 980 32864
rect 4780 32824 4820 32864
rect 7564 32824 7604 32864
rect 9196 32824 9236 32864
rect 19564 32824 19604 32864
rect 4300 32740 4340 32780
rect 10924 32740 10964 32780
rect 12364 32740 12404 32780
rect 13036 32740 13076 32780
rect 2956 32656 2996 32696
rect 11788 32656 11828 32696
rect 15436 32656 15476 32696
rect 16300 32656 16340 32696
rect 10060 32572 10100 32612
rect 15628 32572 15668 32612
rect 18028 32572 18068 32612
rect 4300 32488 4340 32528
rect 4928 32488 4968 32528
rect 5010 32488 5050 32528
rect 5092 32488 5132 32528
rect 5174 32488 5214 32528
rect 5256 32488 5296 32528
rect 15820 32488 15860 32528
rect 19564 32488 19604 32528
rect 20048 32488 20088 32528
rect 20130 32488 20170 32528
rect 20212 32488 20252 32528
rect 20294 32488 20334 32528
rect 20376 32488 20416 32528
rect 21004 32488 21044 32528
rect 1132 32404 1172 32444
rect 8428 32404 8468 32444
rect 8716 32404 8756 32444
rect 2092 32320 2132 32360
rect 3916 32320 3956 32360
rect 12652 32320 12692 32360
rect 12940 32320 12980 32360
rect 14956 32320 14996 32360
rect 15436 32320 15476 32360
rect 15916 32320 15956 32360
rect 18508 32320 18548 32360
rect 12268 32236 12308 32276
rect 2092 32152 2132 32192
rect 8332 32152 8372 32192
rect 9580 32152 9620 32192
rect 14476 32152 14516 32192
rect 15532 32152 15572 32192
rect 18700 32152 18740 32192
rect 1516 32068 1556 32108
rect 10924 32068 10964 32108
rect 18220 32068 18260 32108
rect 748 31984 788 32024
rect 4108 31984 4148 32024
rect 14956 31984 14996 32024
rect 15148 31984 15188 32024
rect 15340 31984 15380 32024
rect 19660 31984 19700 32024
rect 6988 31900 7028 31940
rect 19948 31900 19988 31940
rect 2668 31816 2708 31856
rect 9100 31816 9140 31856
rect 10060 31816 10100 31856
rect 12652 31816 12692 31856
rect 3688 31732 3728 31772
rect 3770 31732 3810 31772
rect 3852 31732 3892 31772
rect 3934 31732 3974 31772
rect 4016 31732 4056 31772
rect 9964 31732 10004 31772
rect 14956 31732 14996 31772
rect 18808 31732 18848 31772
rect 18890 31732 18930 31772
rect 18972 31732 19012 31772
rect 19054 31732 19094 31772
rect 19136 31732 19176 31772
rect 3532 31648 3572 31688
rect 12940 31648 12980 31688
rect 2380 31564 2420 31604
rect 3052 31564 3092 31604
rect 3628 31564 3668 31604
rect 12076 31564 12116 31604
rect 15148 31564 15188 31604
rect 9292 31480 9332 31520
rect 16876 31480 16916 31520
rect 20908 31480 20948 31520
rect 2860 31228 2900 31268
rect 4012 31228 4052 31268
rect 4588 31228 4628 31268
rect 9964 31228 10004 31268
rect 13228 31228 13268 31268
rect 17260 31312 17300 31352
rect 18220 31228 18260 31268
rect 1324 31144 1364 31184
rect 2764 31144 2804 31184
rect 3340 31144 3380 31184
rect 16396 31144 16436 31184
rect 18124 31144 18164 31184
rect 1996 31060 2036 31100
rect 6988 31060 7028 31100
rect 11788 31060 11828 31100
rect 4928 30976 4968 31016
rect 5010 30976 5050 31016
rect 5092 30976 5132 31016
rect 5174 30976 5214 31016
rect 5256 30976 5296 31016
rect 12076 30976 12116 31016
rect 20048 30976 20088 31016
rect 20130 30976 20170 31016
rect 20212 30976 20252 31016
rect 20294 30976 20334 31016
rect 20376 30976 20416 31016
rect 21292 30976 21332 31016
rect 2668 30892 2708 30932
rect 4012 30892 4052 30932
rect 4396 30892 4436 30932
rect 19756 30892 19796 30932
rect 3052 30808 3092 30848
rect 7372 30808 7412 30848
rect 17452 30808 17492 30848
rect 18796 30808 18836 30848
rect 11116 30724 11156 30764
rect 14284 30724 14324 30764
rect 2764 30640 2804 30680
rect 4012 30640 4052 30680
rect 17260 30640 17300 30680
rect 18412 30640 18452 30680
rect 18700 30640 18740 30680
rect 4108 30556 4148 30596
rect 11500 30556 11540 30596
rect 17452 30556 17492 30596
rect 20524 30640 20564 30680
rect 17932 30472 17972 30512
rect 21388 30472 21428 30512
rect 15148 30388 15188 30428
rect 5356 30304 5396 30344
rect 7756 30304 7796 30344
rect 14092 30304 14132 30344
rect 3688 30220 3728 30260
rect 3770 30220 3810 30260
rect 3852 30220 3892 30260
rect 3934 30220 3974 30260
rect 4016 30220 4056 30260
rect 18808 30220 18848 30260
rect 18890 30220 18930 30260
rect 18972 30220 19012 30260
rect 19054 30220 19094 30260
rect 19136 30220 19176 30260
rect 7084 30136 7124 30176
rect 9580 30136 9620 30176
rect 14860 30136 14900 30176
rect 21388 30136 21428 30176
rect 3148 30052 3188 30092
rect 14092 30052 14132 30092
rect 20716 29968 20756 30008
rect 4204 29884 4244 29924
rect 9004 29884 9044 29924
rect 14476 29884 14516 29924
rect 2764 29800 2804 29840
rect 6604 29800 6644 29840
rect 7276 29800 7316 29840
rect 10636 29800 10676 29840
rect 13324 29716 13364 29756
rect 16300 29716 16340 29756
rect 76 29632 116 29672
rect 7084 29632 7124 29672
rect 10060 29632 10100 29672
rect 11116 29632 11156 29672
rect 3052 29464 3092 29504
rect 4928 29464 4968 29504
rect 5010 29464 5050 29504
rect 5092 29464 5132 29504
rect 5174 29464 5214 29504
rect 5256 29464 5296 29504
rect 6508 29464 6548 29504
rect 8428 29464 8468 29504
rect 13324 29464 13364 29504
rect 15436 29464 15476 29504
rect 20048 29464 20088 29504
rect 20130 29464 20170 29504
rect 20212 29464 20252 29504
rect 20294 29464 20334 29504
rect 20376 29464 20416 29504
rect 20620 29464 20660 29504
rect 16876 29380 16916 29420
rect 940 29296 980 29336
rect 5740 29296 5780 29336
rect 6028 29296 6068 29336
rect 14284 29212 14324 29252
rect 1996 29128 2036 29168
rect 11212 29128 11252 29168
rect 12844 29128 12884 29168
rect 460 29044 500 29084
rect 13132 29128 13172 29168
rect 15820 29128 15860 29168
rect 16588 29128 16628 29168
rect 844 28960 884 29000
rect 9964 28960 10004 29000
rect 10828 28960 10868 29000
rect 15436 28960 15476 29000
rect 19948 29044 19988 29084
rect 19852 28960 19892 29000
rect 1804 28876 1844 28916
rect 6988 28792 7028 28832
rect 10636 28792 10676 28832
rect 3436 28708 3476 28748
rect 3688 28708 3728 28748
rect 3770 28708 3810 28748
rect 3852 28708 3892 28748
rect 3934 28708 3974 28748
rect 4016 28708 4056 28748
rect 18808 28708 18848 28748
rect 18890 28708 18930 28748
rect 18972 28708 19012 28748
rect 19054 28708 19094 28748
rect 19136 28708 19176 28748
rect 7948 28624 7988 28664
rect 8428 28624 8468 28664
rect 15436 28540 15476 28580
rect 9676 28372 9716 28412
rect 13612 28372 13652 28412
rect 19564 28372 19604 28412
rect 9484 28288 9524 28328
rect 6700 28204 6740 28244
rect 13996 28204 14036 28244
rect 1228 28120 1268 28160
rect 14956 28036 14996 28076
rect 3244 27952 3284 27992
rect 4928 27952 4968 27992
rect 5010 27952 5050 27992
rect 5092 27952 5132 27992
rect 5174 27952 5214 27992
rect 5256 27952 5296 27992
rect 5644 27952 5684 27992
rect 9484 27952 9524 27992
rect 20048 27952 20088 27992
rect 20130 27952 20170 27992
rect 20212 27952 20252 27992
rect 20294 27952 20334 27992
rect 20376 27952 20416 27992
rect 2668 27868 2708 27908
rect 17260 27868 17300 27908
rect 4492 27784 4532 27824
rect 4780 27784 4820 27824
rect 5548 27784 5588 27824
rect 13900 27784 13940 27824
rect 1900 27700 1940 27740
rect 9772 27700 9812 27740
rect 13612 27700 13652 27740
rect 2476 27616 2516 27656
rect 15340 27700 15380 27740
rect 12652 27616 12692 27656
rect 14092 27616 14132 27656
rect 9004 27532 9044 27572
rect 9580 27532 9620 27572
rect 15628 27700 15668 27740
rect 17452 27616 17492 27656
rect 7276 27448 7316 27488
rect 7756 27448 7796 27488
rect 14860 27448 14900 27488
rect 15724 27448 15764 27488
rect 16300 27448 16340 27488
rect 9388 27364 9428 27404
rect 9676 27364 9716 27404
rect 19372 27280 19412 27320
rect 3688 27196 3728 27236
rect 3770 27196 3810 27236
rect 3852 27196 3892 27236
rect 3934 27196 3974 27236
rect 4016 27196 4056 27236
rect 13420 27196 13460 27236
rect 16684 27196 16724 27236
rect 18808 27196 18848 27236
rect 18890 27196 18930 27236
rect 18972 27196 19012 27236
rect 19054 27196 19094 27236
rect 19136 27196 19176 27236
rect 7948 27112 7988 27152
rect 3628 27028 3668 27068
rect 6316 27028 6356 27068
rect 14092 27028 14132 27068
rect 17740 27028 17780 27068
rect 18700 27028 18740 27068
rect 3052 26944 3092 26984
rect 4300 26860 4340 26900
rect 6412 26860 6452 26900
rect 6508 26776 6548 26816
rect 9292 26776 9332 26816
rect 9676 26776 9716 26816
rect 9964 26776 10004 26816
rect 2764 26692 2804 26732
rect 6316 26692 6356 26732
rect 11980 26692 12020 26732
rect 4300 26608 4340 26648
rect 7180 26608 7220 26648
rect 9580 26608 9620 26648
rect 12940 26608 12980 26648
rect 13420 26608 13460 26648
rect 16780 26860 16820 26900
rect 17356 26860 17396 26900
rect 18028 26860 18068 26900
rect 19564 26860 19604 26900
rect 17452 26776 17492 26816
rect 19948 26692 19988 26732
rect 16684 26608 16724 26648
rect 17260 26608 17300 26648
rect 1324 26440 1364 26480
rect 4928 26440 4968 26480
rect 5010 26440 5050 26480
rect 5092 26440 5132 26480
rect 5174 26440 5214 26480
rect 5256 26440 5296 26480
rect 5644 26440 5684 26480
rect 6508 26440 6548 26480
rect 7276 26440 7316 26480
rect 19660 26440 19700 26480
rect 20048 26440 20088 26480
rect 20130 26440 20170 26480
rect 20212 26440 20252 26480
rect 20294 26440 20334 26480
rect 20376 26440 20416 26480
rect 2476 26356 2516 26396
rect 2956 26356 2996 26396
rect 3340 26356 3380 26396
rect 3724 26356 3764 26396
rect 7756 26356 7796 26396
rect 8620 26356 8660 26396
rect 18700 26356 18740 26396
rect 3436 26272 3476 26312
rect 6412 26272 6452 26312
rect 10060 26272 10100 26312
rect 11116 26272 11156 26312
rect 11884 26272 11924 26312
rect 10252 26188 10292 26228
rect 15148 26188 15188 26228
rect 16780 26188 16820 26228
rect 2476 26104 2516 26144
rect 4492 26104 4532 26144
rect 8428 26104 8468 26144
rect 8620 26104 8660 26144
rect 16684 26104 16724 26144
rect 17740 26104 17780 26144
rect 18412 26104 18452 26144
rect 6508 26020 6548 26060
rect 4204 25936 4244 25976
rect 13036 25936 13076 25976
rect 6220 25852 6260 25892
rect 6316 25768 6356 25808
rect 3688 25684 3728 25724
rect 3770 25684 3810 25724
rect 3852 25684 3892 25724
rect 3934 25684 3974 25724
rect 4016 25684 4056 25724
rect 7180 25684 7220 25724
rect 10060 25684 10100 25724
rect 16780 25684 16820 25724
rect 18808 25684 18848 25724
rect 18890 25684 18930 25724
rect 18972 25684 19012 25724
rect 19054 25684 19094 25724
rect 19136 25684 19176 25724
rect 3340 25516 3380 25556
rect 4684 25516 4724 25556
rect 14092 25516 14132 25556
rect 18028 25516 18068 25556
rect 16204 25432 16244 25472
rect 16780 25432 16820 25472
rect 2284 25348 2324 25388
rect 5452 25348 5492 25388
rect 5740 25348 5780 25388
rect 11596 25348 11636 25388
rect 13132 25348 13172 25388
rect 13612 25348 13652 25388
rect 15532 25348 15572 25388
rect 18508 25348 18548 25388
rect 19948 25348 19988 25388
rect 6988 25264 7028 25304
rect 12844 25264 12884 25304
rect 15820 25264 15860 25304
rect 17740 25264 17780 25304
rect 5932 25180 5972 25220
rect 8236 25180 8276 25220
rect 14092 25180 14132 25220
rect 15148 25180 15188 25220
rect 16204 25180 16244 25220
rect 16588 25180 16628 25220
rect 17068 25180 17108 25220
rect 3244 25096 3284 25136
rect 10444 25096 10484 25136
rect 12172 25096 12212 25136
rect 15436 25096 15476 25136
rect 19372 25096 19412 25136
rect 8620 25012 8660 25052
rect 11980 25012 12020 25052
rect 172 24928 212 24968
rect 4928 24928 4968 24968
rect 5010 24928 5050 24968
rect 5092 24928 5132 24968
rect 5174 24928 5214 24968
rect 5256 24928 5296 24968
rect 14092 24928 14132 24968
rect 20048 24928 20088 24968
rect 20130 24928 20170 24968
rect 20212 24928 20252 24968
rect 20294 24928 20334 24968
rect 20376 24928 20416 24968
rect 9772 24844 9812 24884
rect 5452 24760 5492 24800
rect 10828 24760 10868 24800
rect 14956 24760 14996 24800
rect 4588 24676 4628 24716
rect 1228 24592 1268 24632
rect 11884 24676 11924 24716
rect 18604 24676 18644 24716
rect 1420 24592 1460 24632
rect 13036 24592 13076 24632
rect 2476 24508 2516 24548
rect 8428 24508 8468 24548
rect 17740 24508 17780 24548
rect 2380 24424 2420 24464
rect 3688 24172 3728 24212
rect 3770 24172 3810 24212
rect 3852 24172 3892 24212
rect 3934 24172 3974 24212
rect 4016 24172 4056 24212
rect 4780 24172 4820 24212
rect 10636 24172 10676 24212
rect 18808 24172 18848 24212
rect 18890 24172 18930 24212
rect 18972 24172 19012 24212
rect 19054 24172 19094 24212
rect 19136 24172 19176 24212
rect 13516 24004 13556 24044
rect 10540 23920 10580 23960
rect 1612 23836 1652 23876
rect 10828 23920 10868 23960
rect 4300 23836 4340 23876
rect 1900 23752 1940 23792
rect 3052 23752 3092 23792
rect 7084 23752 7124 23792
rect 10540 23752 10580 23792
rect 12268 23752 12308 23792
rect 17932 23920 17972 23960
rect 18412 23920 18452 23960
rect 19372 23920 19412 23960
rect 20524 23920 20564 23960
rect 19852 23836 19892 23876
rect 16300 23752 16340 23792
rect 19372 23752 19412 23792
rect 11788 23668 11828 23708
rect 15340 23668 15380 23708
rect 16588 23668 16628 23708
rect 18508 23668 18548 23708
rect 3724 23584 3764 23624
rect 9772 23584 9812 23624
rect 4108 23500 4148 23540
rect 2764 23416 2804 23456
rect 4928 23416 4968 23456
rect 5010 23416 5050 23456
rect 5092 23416 5132 23456
rect 5174 23416 5214 23456
rect 5256 23416 5296 23456
rect 8620 23416 8660 23456
rect 10540 23416 10580 23456
rect 20048 23416 20088 23456
rect 20130 23416 20170 23456
rect 20212 23416 20252 23456
rect 20294 23416 20334 23456
rect 20376 23416 20416 23456
rect 3052 23332 3092 23372
rect 11788 23248 11828 23288
rect 12652 23248 12692 23288
rect 2764 23080 2804 23120
rect 6700 23080 6740 23120
rect 9100 23080 9140 23120
rect 10060 23164 10100 23204
rect 9580 23080 9620 23120
rect 15340 23080 15380 23120
rect 4300 22996 4340 23036
rect 10828 22996 10868 23036
rect 19372 22996 19412 23036
rect 3436 22912 3476 22952
rect 8716 22912 8756 22952
rect 4108 22828 4148 22868
rect 12844 22828 12884 22868
rect 10540 22744 10580 22784
rect 2284 22660 2324 22700
rect 3688 22660 3728 22700
rect 3770 22660 3810 22700
rect 3852 22660 3892 22700
rect 3934 22660 3974 22700
rect 4016 22660 4056 22700
rect 16492 22660 16532 22700
rect 17836 22660 17876 22700
rect 18700 22660 18740 22700
rect 18808 22660 18848 22700
rect 18890 22660 18930 22700
rect 18972 22660 19012 22700
rect 19054 22660 19094 22700
rect 19136 22660 19176 22700
rect 19564 22660 19604 22700
rect 3244 22492 3284 22532
rect 6316 22492 6356 22532
rect 19372 22492 19412 22532
rect 3532 22408 3572 22448
rect 13324 22408 13364 22448
rect 7084 22324 7124 22364
rect 11308 22324 11348 22364
rect 1228 22240 1268 22280
rect 5356 22240 5396 22280
rect 16492 22240 16532 22280
rect 17164 22240 17204 22280
rect 13900 22156 13940 22196
rect 3340 22072 3380 22112
rect 8236 22072 8276 22112
rect 8428 22072 8468 22112
rect 8620 22072 8660 22112
rect 12268 22072 12308 22112
rect 11788 21988 11828 22028
rect 16492 21988 16532 22028
rect 3436 21904 3476 21944
rect 4928 21904 4968 21944
rect 5010 21904 5050 21944
rect 5092 21904 5132 21944
rect 5174 21904 5214 21944
rect 5256 21904 5296 21944
rect 6124 21904 6164 21944
rect 20048 21904 20088 21944
rect 20130 21904 20170 21944
rect 20212 21904 20252 21944
rect 20294 21904 20334 21944
rect 20376 21904 20416 21944
rect 4108 21736 4148 21776
rect 16876 21736 16916 21776
rect 18124 21736 18164 21776
rect 268 21568 308 21608
rect 1804 21568 1844 21608
rect 2188 21568 2228 21608
rect 4492 21568 4532 21608
rect 4684 21568 4724 21608
rect 7372 21568 7412 21608
rect 16876 21568 16916 21608
rect 3436 21484 3476 21524
rect 3916 21484 3956 21524
rect 6412 21484 6452 21524
rect 8716 21484 8756 21524
rect 11308 21484 11348 21524
rect 3340 21400 3380 21440
rect 6316 21400 6356 21440
rect 7372 21400 7412 21440
rect 8524 21400 8564 21440
rect 9292 21400 9332 21440
rect 11884 21400 11924 21440
rect 12268 21400 12308 21440
rect 2092 21316 2132 21356
rect 7756 21316 7796 21356
rect 8812 21316 8852 21356
rect 17740 21316 17780 21356
rect 1996 21232 2036 21272
rect 9292 21232 9332 21272
rect 10348 21232 10388 21272
rect 2764 21148 2804 21188
rect 3688 21148 3728 21188
rect 3770 21148 3810 21188
rect 3852 21148 3892 21188
rect 3934 21148 3974 21188
rect 4016 21148 4056 21188
rect 6892 21148 6932 21188
rect 18808 21148 18848 21188
rect 18890 21148 18930 21188
rect 18972 21148 19012 21188
rect 19054 21148 19094 21188
rect 19136 21148 19176 21188
rect 13900 21064 13940 21104
rect 16492 21064 16532 21104
rect 2860 20896 2900 20936
rect 6508 20896 6548 20936
rect 7084 20896 7124 20936
rect 6220 20812 6260 20852
rect 9388 20812 9428 20852
rect 1996 20728 2036 20768
rect 4684 20728 4724 20768
rect 6316 20728 6356 20768
rect 7276 20728 7316 20768
rect 10540 20728 10580 20768
rect 10828 20728 10868 20768
rect 11212 20728 11252 20768
rect 18412 20728 18452 20768
rect 19372 20728 19412 20768
rect 15724 20644 15764 20684
rect 3436 20560 3476 20600
rect 4492 20560 4532 20600
rect 10924 20560 10964 20600
rect 18700 20560 18740 20600
rect 19660 20560 19700 20600
rect 2668 20392 2708 20432
rect 4108 20392 4148 20432
rect 4928 20392 4968 20432
rect 5010 20392 5050 20432
rect 5092 20392 5132 20432
rect 5174 20392 5214 20432
rect 5256 20392 5296 20432
rect 5452 20392 5492 20432
rect 20048 20392 20088 20432
rect 20130 20392 20170 20432
rect 20212 20392 20252 20432
rect 20294 20392 20334 20432
rect 20376 20392 20416 20432
rect 18028 20308 18068 20348
rect 2956 20140 2996 20180
rect 11308 20140 11348 20180
rect 2476 20056 2516 20096
rect 4300 20056 4340 20096
rect 6508 20056 6548 20096
rect 9004 20056 9044 20096
rect 10444 20056 10484 20096
rect 2188 19972 2228 20012
rect 9676 19972 9716 20012
rect 13804 19972 13844 20012
rect 14860 19972 14900 20012
rect 15820 19972 15860 20012
rect 16588 19888 16628 19928
rect 2764 19804 2804 19844
rect 3532 19804 3572 19844
rect 4204 19804 4244 19844
rect 13996 19804 14036 19844
rect 17164 19804 17204 19844
rect 3688 19636 3728 19676
rect 3770 19636 3810 19676
rect 3852 19636 3892 19676
rect 3934 19636 3974 19676
rect 4016 19636 4056 19676
rect 17644 19636 17684 19676
rect 18808 19636 18848 19676
rect 18890 19636 18930 19676
rect 18972 19636 19012 19676
rect 19054 19636 19094 19676
rect 19136 19636 19176 19676
rect 19372 19636 19412 19676
rect 19660 19636 19700 19676
rect 10924 19552 10964 19592
rect 16780 19552 16820 19592
rect 2668 19468 2708 19508
rect 2764 19384 2804 19424
rect 14380 19384 14420 19424
rect 17260 19384 17300 19424
rect 6028 19300 6068 19340
rect 6220 19300 6260 19340
rect 9484 19300 9524 19340
rect 10636 19300 10676 19340
rect 16012 19300 16052 19340
rect 2092 19216 2132 19256
rect 4108 19216 4148 19256
rect 4780 19216 4820 19256
rect 6508 19216 6548 19256
rect 9676 19216 9716 19256
rect 17164 19216 17204 19256
rect 1708 19132 1748 19172
rect 8332 19132 8372 19172
rect 4300 19048 4340 19088
rect 10828 19048 10868 19088
rect 13804 19132 13844 19172
rect 14380 19132 14420 19172
rect 20812 19132 20852 19172
rect 14092 19048 14132 19088
rect 17164 19048 17204 19088
rect 9292 18964 9332 19004
rect 13804 18964 13844 19004
rect 16876 18964 16916 19004
rect 4928 18880 4968 18920
rect 5010 18880 5050 18920
rect 5092 18880 5132 18920
rect 5174 18880 5214 18920
rect 5256 18880 5296 18920
rect 6028 18880 6068 18920
rect 10924 18880 10964 18920
rect 17644 18880 17684 18920
rect 20048 18880 20088 18920
rect 20130 18880 20170 18920
rect 20212 18880 20252 18920
rect 20294 18880 20334 18920
rect 20376 18880 20416 18920
rect 5452 18796 5492 18836
rect 5356 18712 5396 18752
rect 10444 18628 10484 18668
rect 6124 18544 6164 18584
rect 1516 18460 1556 18500
rect 3148 18460 3188 18500
rect 13228 18376 13268 18416
rect 16684 18376 16724 18416
rect 2956 18292 2996 18332
rect 3148 18292 3188 18332
rect 10636 18292 10676 18332
rect 5740 18208 5780 18248
rect 13804 18208 13844 18248
rect 3688 18124 3728 18164
rect 3770 18124 3810 18164
rect 3852 18124 3892 18164
rect 3934 18124 3974 18164
rect 4016 18124 4056 18164
rect 18808 18124 18848 18164
rect 18890 18124 18930 18164
rect 18972 18124 19012 18164
rect 19054 18124 19094 18164
rect 19136 18124 19176 18164
rect 3532 17956 3572 17996
rect 8908 17956 8948 17996
rect 14956 17956 14996 17996
rect 18412 17956 18452 17996
rect 19468 17872 19508 17912
rect 13612 17788 13652 17828
rect 15820 17788 15860 17828
rect 17260 17788 17300 17828
rect 1612 17704 1652 17744
rect 4780 17704 4820 17744
rect 172 17620 212 17660
rect 5356 17620 5396 17660
rect 7564 17620 7604 17660
rect 9484 17620 9524 17660
rect 17836 17620 17876 17660
rect 5548 17452 5588 17492
rect 4928 17368 4968 17408
rect 5010 17368 5050 17408
rect 5092 17368 5132 17408
rect 5174 17368 5214 17408
rect 5256 17368 5296 17408
rect 9772 17368 9812 17408
rect 20048 17368 20088 17408
rect 20130 17368 20170 17408
rect 20212 17368 20252 17408
rect 20294 17368 20334 17408
rect 20376 17368 20416 17408
rect 1516 17284 1556 17324
rect 4780 17200 4820 17240
rect 13996 17116 14036 17156
rect 2092 17032 2132 17072
rect 20908 17032 20948 17072
rect 1228 16864 1268 16904
rect 4204 16864 4244 16904
rect 16300 16864 16340 16904
rect 19756 16780 19796 16820
rect 10348 16696 10388 16736
rect 12556 16696 12596 16736
rect 3688 16612 3728 16652
rect 3770 16612 3810 16652
rect 3852 16612 3892 16652
rect 3934 16612 3974 16652
rect 4016 16612 4056 16652
rect 10636 16612 10676 16652
rect 11692 16612 11732 16652
rect 18808 16612 18848 16652
rect 18890 16612 18930 16652
rect 18972 16612 19012 16652
rect 19054 16612 19094 16652
rect 19136 16612 19176 16652
rect 16876 16528 16916 16568
rect 8812 16360 8852 16400
rect 21292 16360 21332 16400
rect 3052 16276 3092 16316
rect 3436 16192 3476 16232
rect 11692 16276 11732 16316
rect 2764 16108 2804 16148
rect 13036 16108 13076 16148
rect 6892 16024 6932 16064
rect 7468 16024 7508 16064
rect 8908 16024 8948 16064
rect 9292 16024 9332 16064
rect 11692 16024 11732 16064
rect 19948 16024 19988 16064
rect 15532 15940 15572 15980
rect 19372 15940 19412 15980
rect 3148 15856 3188 15896
rect 4928 15856 4968 15896
rect 5010 15856 5050 15896
rect 5092 15856 5132 15896
rect 5174 15856 5214 15896
rect 5256 15856 5296 15896
rect 9196 15856 9236 15896
rect 9772 15856 9812 15896
rect 14572 15856 14612 15896
rect 18700 15856 18740 15896
rect 20048 15856 20088 15896
rect 20130 15856 20170 15896
rect 20212 15856 20252 15896
rect 20294 15856 20334 15896
rect 20376 15856 20416 15896
rect 21388 15856 21428 15896
rect 2668 15772 2708 15812
rect 7084 15772 7124 15812
rect 20524 15772 20564 15812
rect 13804 15688 13844 15728
rect 9100 15604 9140 15644
rect 21004 15604 21044 15644
rect 1708 15520 1748 15560
rect 2764 15520 2804 15560
rect 9196 15520 9236 15560
rect 11884 15520 11924 15560
rect 16876 15436 16916 15476
rect 19372 15436 19412 15476
rect 13612 15352 13652 15392
rect 1612 15268 1652 15308
rect 16972 15268 17012 15308
rect 17644 15268 17684 15308
rect 14956 15184 14996 15224
rect 3688 15100 3728 15140
rect 3770 15100 3810 15140
rect 3852 15100 3892 15140
rect 3934 15100 3974 15140
rect 4016 15100 4056 15140
rect 4588 15100 4628 15140
rect 5644 15100 5684 15140
rect 12460 15100 12500 15140
rect 16396 15100 16436 15140
rect 17164 15100 17204 15140
rect 18808 15100 18848 15140
rect 18890 15100 18930 15140
rect 18972 15100 19012 15140
rect 19054 15100 19094 15140
rect 19136 15100 19176 15140
rect 19660 15100 19700 15140
rect 76 15016 116 15056
rect 1420 15016 1460 15056
rect 2476 14932 2516 14972
rect 5836 14932 5876 14972
rect 3148 14848 3188 14888
rect 9964 14848 10004 14888
rect 21196 14848 21236 14888
rect 3052 14764 3092 14804
rect 4204 14764 4244 14804
rect 12748 14764 12788 14804
rect 3532 14680 3572 14720
rect 13804 14764 13844 14804
rect 4492 14680 4532 14720
rect 5740 14680 5780 14720
rect 6220 14680 6260 14720
rect 10444 14680 10484 14720
rect 10924 14680 10964 14720
rect 15724 14680 15764 14720
rect 19852 14680 19892 14720
rect 1996 14596 2036 14636
rect 1900 14512 1940 14552
rect 4928 14344 4968 14384
rect 5010 14344 5050 14384
rect 5092 14344 5132 14384
rect 5174 14344 5214 14384
rect 5256 14344 5296 14384
rect 5932 14596 5972 14636
rect 8908 14596 8948 14636
rect 9484 14596 9524 14636
rect 16396 14596 16436 14636
rect 19660 14596 19700 14636
rect 16876 14512 16916 14552
rect 18700 14428 18740 14468
rect 11212 14344 11252 14384
rect 17644 14344 17684 14384
rect 20048 14344 20088 14384
rect 20130 14344 20170 14384
rect 20212 14344 20252 14384
rect 20294 14344 20334 14384
rect 20376 14344 20416 14384
rect 9100 14260 9140 14300
rect 6124 14176 6164 14216
rect 11308 14176 11348 14216
rect 16300 14176 16340 14216
rect 6220 14092 6260 14132
rect 13612 14092 13652 14132
rect 3820 14008 3860 14048
rect 19756 14008 19796 14048
rect 9196 13924 9236 13964
rect 12364 13924 12404 13964
rect 5644 13840 5684 13880
rect 10156 13840 10196 13880
rect 11788 13840 11828 13880
rect 12172 13840 12212 13880
rect 19948 13840 19988 13880
rect 4492 13756 4532 13796
rect 4684 13756 4724 13796
rect 12460 13756 12500 13796
rect 15820 13672 15860 13712
rect 18700 13672 18740 13712
rect 19276 13672 19316 13712
rect 2476 13588 2516 13628
rect 3688 13588 3728 13628
rect 3770 13588 3810 13628
rect 3852 13588 3892 13628
rect 3934 13588 3974 13628
rect 4016 13588 4056 13628
rect 12268 13588 12308 13628
rect 13228 13588 13268 13628
rect 18808 13588 18848 13628
rect 18890 13588 18930 13628
rect 18972 13588 19012 13628
rect 19054 13588 19094 13628
rect 19136 13588 19176 13628
rect 4588 13504 4628 13544
rect 7468 13504 7508 13544
rect 1036 13420 1076 13460
rect 10444 13420 10484 13460
rect 19372 13420 19412 13460
rect 19948 13336 19988 13376
rect 8332 13252 8372 13292
rect 2476 13168 2516 13208
rect 4108 13168 4148 13208
rect 4588 13168 4628 13208
rect 5356 13168 5396 13208
rect 6316 13168 6356 13208
rect 9772 13168 9812 13208
rect 11404 13168 11444 13208
rect 19372 13168 19412 13208
rect 2956 13084 2996 13124
rect 10060 13084 10100 13124
rect 19468 13084 19508 13124
rect 11404 13000 11444 13040
rect 844 12832 884 12872
rect 3148 12832 3188 12872
rect 4396 12832 4436 12872
rect 4928 12832 4968 12872
rect 5010 12832 5050 12872
rect 5092 12832 5132 12872
rect 5174 12832 5214 12872
rect 5256 12832 5296 12872
rect 9964 12832 10004 12872
rect 20048 12832 20088 12872
rect 20130 12832 20170 12872
rect 20212 12832 20252 12872
rect 20294 12832 20334 12872
rect 20376 12832 20416 12872
rect 4780 12748 4820 12788
rect 11980 12748 12020 12788
rect 364 12580 404 12620
rect 4204 12580 4244 12620
rect 8620 12580 8660 12620
rect 3532 12496 3572 12536
rect 5164 12496 5204 12536
rect 7084 12496 7124 12536
rect 364 12412 404 12452
rect 1516 12412 1556 12452
rect 2956 12328 2996 12368
rect 6124 12244 6164 12284
rect 12268 12328 12308 12368
rect 14476 12244 14516 12284
rect 20044 12244 20084 12284
rect 3436 12160 3476 12200
rect 3688 12076 3728 12116
rect 3770 12076 3810 12116
rect 3852 12076 3892 12116
rect 3934 12076 3974 12116
rect 4016 12076 4056 12116
rect 6316 12076 6356 12116
rect 5548 11992 5588 12032
rect 6604 12076 6644 12116
rect 10156 12076 10196 12116
rect 12556 12076 12596 12116
rect 18808 12076 18848 12116
rect 18890 12076 18930 12116
rect 18972 12076 19012 12116
rect 19054 12076 19094 12116
rect 19136 12076 19176 12116
rect 2092 11908 2132 11948
rect 4780 11908 4820 11948
rect 7852 11908 7892 11948
rect 9196 11908 9236 11948
rect 3436 11824 3476 11864
rect 5356 11824 5396 11864
rect 8236 11824 8276 11864
rect 12652 11824 12692 11864
rect 13516 11824 13556 11864
rect 15148 11824 15188 11864
rect 16972 11824 17012 11864
rect 3724 11656 3764 11696
rect 5164 11740 5204 11780
rect 5644 11740 5684 11780
rect 6700 11740 6740 11780
rect 9676 11656 9716 11696
rect 18028 11824 18068 11864
rect 19756 11824 19796 11864
rect 10444 11740 10484 11780
rect 11980 11656 12020 11696
rect 13036 11656 13076 11696
rect 13804 11656 13844 11696
rect 15820 11656 15860 11696
rect 16684 11656 16724 11696
rect 16972 11656 17012 11696
rect 1708 11572 1748 11612
rect 6316 11572 6356 11612
rect 7276 11572 7316 11612
rect 7852 11488 7892 11528
rect 14188 11488 14228 11528
rect 20044 11488 20084 11528
rect 15436 11404 15476 11444
rect 18892 11404 18932 11444
rect 19756 11404 19796 11444
rect 4928 11320 4968 11360
rect 5010 11320 5050 11360
rect 5092 11320 5132 11360
rect 5174 11320 5214 11360
rect 5256 11320 5296 11360
rect 7084 11320 7124 11360
rect 9484 11320 9524 11360
rect 13516 11320 13556 11360
rect 20048 11320 20088 11360
rect 20130 11320 20170 11360
rect 20212 11320 20252 11360
rect 20294 11320 20334 11360
rect 20376 11320 20416 11360
rect 21100 11320 21140 11360
rect 4108 11236 4148 11276
rect 10444 11236 10484 11276
rect 14092 11236 14132 11276
rect 16396 11236 16436 11276
rect 18988 11236 19028 11276
rect 4108 11068 4148 11108
rect 11500 11068 11540 11108
rect 16780 11068 16820 11108
rect 9580 10984 9620 11024
rect 16876 10984 16916 11024
rect 16684 10900 16724 10940
rect 556 10816 596 10856
rect 2860 10816 2900 10856
rect 10252 10816 10292 10856
rect 18316 10816 18356 10856
rect 18508 10816 18548 10856
rect 844 10732 884 10772
rect 2284 10732 2324 10772
rect 4780 10732 4820 10772
rect 9676 10732 9716 10772
rect 1804 10648 1844 10688
rect 5452 10648 5492 10688
rect 940 10564 980 10604
rect 3436 10564 3476 10604
rect 3688 10564 3728 10604
rect 3770 10564 3810 10604
rect 3852 10564 3892 10604
rect 3934 10564 3974 10604
rect 4016 10564 4056 10604
rect 4300 10564 4340 10604
rect 9484 10564 9524 10604
rect 16108 10564 16148 10604
rect 18808 10564 18848 10604
rect 18890 10564 18930 10604
rect 18972 10564 19012 10604
rect 19054 10564 19094 10604
rect 19136 10564 19176 10604
rect 4780 10480 4820 10520
rect 2764 10396 2804 10436
rect 2956 10396 2996 10436
rect 3244 10396 3284 10436
rect 20812 10396 20852 10436
rect 5548 10312 5588 10352
rect 6316 10312 6356 10352
rect 8524 10312 8564 10352
rect 2092 10228 2132 10268
rect 20716 10228 20756 10268
rect 1516 10144 1556 10184
rect 2284 10144 2324 10184
rect 5452 10144 5492 10184
rect 5932 10144 5972 10184
rect 7564 10144 7604 10184
rect 9964 10144 10004 10184
rect 15820 10144 15860 10184
rect 20620 10144 20660 10184
rect 14764 10060 14804 10100
rect 15244 10060 15284 10100
rect 5836 9976 5876 10016
rect 16012 10060 16052 10100
rect 16588 10060 16628 10100
rect 21004 10060 21044 10100
rect 7468 9976 7508 10016
rect 13612 9976 13652 10016
rect 5740 9892 5780 9932
rect 5932 9892 5972 9932
rect 8716 9892 8756 9932
rect 17164 9892 17204 9932
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 11212 9808 11252 9848
rect 13996 9808 14036 9848
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 8716 9724 8756 9764
rect 9388 9724 9428 9764
rect 11884 9724 11924 9764
rect 2956 9640 2996 9680
rect 7084 9640 7124 9680
rect 16588 9640 16628 9680
rect 20044 9640 20084 9680
rect 9100 9472 9140 9512
rect 11212 9472 11252 9512
rect 15532 9472 15572 9512
rect 18316 9472 18356 9512
rect 19564 9472 19604 9512
rect 19948 9472 19988 9512
rect 7564 9388 7604 9428
rect 19756 9388 19796 9428
rect 2476 9304 2516 9344
rect 4684 9304 4724 9344
rect 11116 9304 11156 9344
rect 17164 9304 17204 9344
rect 5932 9220 5972 9260
rect 6700 9220 6740 9260
rect 9100 9220 9140 9260
rect 10060 9136 10100 9176
rect 10444 9136 10484 9176
rect 14476 9136 14516 9176
rect 15148 9136 15188 9176
rect 19276 9136 19316 9176
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 4972 9052 5012 9092
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 4300 8968 4340 9008
rect 1516 8884 1556 8924
rect 1804 8716 1844 8756
rect 10636 8968 10676 9008
rect 12556 8968 12596 9008
rect 12748 8968 12788 9008
rect 10348 8800 10388 8840
rect 14956 8800 14996 8840
rect 16396 8800 16436 8840
rect 19756 8800 19796 8840
rect 16972 8716 17012 8756
rect 9580 8632 9620 8672
rect 19468 8632 19508 8672
rect 19756 8632 19796 8672
rect 12268 8548 12308 8588
rect 13900 8548 13940 8588
rect 16588 8548 16628 8588
rect 18508 8548 18548 8588
rect 13804 8464 13844 8504
rect 5932 8380 5972 8420
rect 6124 8380 6164 8420
rect 20908 8380 20948 8420
rect 2764 8296 2804 8336
rect 4204 8296 4244 8336
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 7564 8296 7604 8336
rect 12364 8296 12404 8336
rect 16396 8296 16436 8336
rect 17644 8296 17684 8336
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 5932 8212 5972 8252
rect 7852 8128 7892 8168
rect 9484 8128 9524 8168
rect 9676 8128 9716 8168
rect 13804 8128 13844 8168
rect 16972 8128 17012 8168
rect 19948 8128 19988 8168
rect 12268 8044 12308 8084
rect 17836 8044 17876 8084
rect 1612 7960 1652 8000
rect 18604 8044 18644 8084
rect 4684 7960 4724 8000
rect 5452 7960 5492 8000
rect 10348 7960 10388 8000
rect 13228 7960 13268 8000
rect 19468 7960 19508 8000
rect 8716 7876 8756 7916
rect 9484 7876 9524 7916
rect 10924 7876 10964 7916
rect 11692 7876 11732 7916
rect 14764 7876 14804 7916
rect 172 7792 212 7832
rect 8812 7708 8852 7748
rect 16588 7708 16628 7748
rect 2380 7540 2420 7580
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 4588 7540 4628 7580
rect 6700 7540 6740 7580
rect 7468 7540 7508 7580
rect 9388 7540 9428 7580
rect 5644 7456 5684 7496
rect 11020 7540 11060 7580
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 19852 7540 19892 7580
rect 8908 7456 8948 7496
rect 16492 7456 16532 7496
rect 16780 7456 16820 7496
rect 13804 7372 13844 7412
rect 14284 7372 14324 7412
rect 15820 7372 15860 7412
rect 16396 7372 16436 7412
rect 6124 7288 6164 7328
rect 6508 7288 6548 7328
rect 18892 7372 18932 7412
rect 19948 7372 19988 7412
rect 20812 7288 20852 7328
rect 3052 7204 3092 7244
rect 17164 7204 17204 7244
rect 8716 7120 8756 7160
rect 6124 7036 6164 7076
rect 12652 7036 12692 7076
rect 748 6952 788 6992
rect 5452 6952 5492 6992
rect 5836 6952 5876 6992
rect 9388 6952 9428 6992
rect 14092 6952 14132 6992
rect 19372 6952 19412 6992
rect 6220 6868 6260 6908
rect 6700 6868 6740 6908
rect 7660 6868 7700 6908
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 6316 6784 6356 6824
rect 15724 6784 15764 6824
rect 19852 6784 19892 6824
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 6508 6700 6548 6740
rect 12364 6700 12404 6740
rect 16684 6700 16724 6740
rect 18412 6700 18452 6740
rect 1516 6448 1556 6488
rect 2188 6616 2228 6656
rect 2764 6616 2804 6656
rect 3148 6616 3188 6656
rect 9484 6616 9524 6656
rect 18892 6700 18932 6740
rect 10060 6616 10100 6656
rect 11692 6532 11732 6572
rect 4108 6448 4148 6488
rect 6028 6448 6068 6488
rect 5836 6364 5876 6404
rect 7852 6448 7892 6488
rect 8716 6448 8756 6488
rect 10348 6448 10388 6488
rect 12268 6448 12308 6488
rect 18316 6448 18356 6488
rect 19660 6448 19700 6488
rect 10060 6364 10100 6404
rect 7564 6280 7604 6320
rect 10252 6280 10292 6320
rect 19948 6280 19988 6320
rect 652 6196 692 6236
rect 20812 6280 20852 6320
rect 7084 6196 7124 6236
rect 11980 6196 12020 6236
rect 1900 6112 1940 6152
rect 4780 6112 4820 6152
rect 5452 6112 5492 6152
rect 10060 6112 10100 6152
rect 13420 6196 13460 6236
rect 19276 6196 19316 6236
rect 16588 6112 16628 6152
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 13996 6028 14036 6068
rect 14476 6028 14516 6068
rect 18316 6028 18356 6068
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 7468 5944 7508 5984
rect 14284 5944 14324 5984
rect 19564 5944 19604 5984
rect 11404 5776 11444 5816
rect 19276 5692 19316 5732
rect 1996 5608 2036 5648
rect 4684 5608 4724 5648
rect 18508 5608 18548 5648
rect 10444 5524 10484 5564
rect 19468 5608 19508 5648
rect 15532 5524 15572 5564
rect 5836 5440 5876 5480
rect 6508 5440 6548 5480
rect 12940 5440 12980 5480
rect 19372 5440 19412 5480
rect 1036 5356 1076 5396
rect 18604 5356 18644 5396
rect 4300 5272 4340 5312
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 6316 5272 6356 5312
rect 13996 5272 14036 5312
rect 17068 5272 17108 5312
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 5452 5188 5492 5228
rect 8716 5188 8756 5228
rect 10828 5188 10868 5228
rect 11116 5188 11156 5228
rect 14476 5188 14516 5228
rect 9676 5104 9716 5144
rect 10636 5104 10676 5144
rect 19756 5104 19796 5144
rect 8812 5020 8852 5060
rect 9580 5020 9620 5060
rect 2668 4936 2708 4976
rect 9388 4936 9428 4976
rect 10252 4936 10292 4976
rect 1324 4852 1364 4892
rect 5356 4852 5396 4892
rect 8236 4852 8276 4892
rect 17836 4936 17876 4976
rect 18028 4936 18068 4976
rect 18412 4936 18452 4976
rect 18604 4936 18644 4976
rect 16300 4852 16340 4892
rect 1228 4768 1268 4808
rect 7564 4684 7604 4724
rect 10348 4684 10388 4724
rect 15340 4684 15380 4724
rect 16492 4600 16532 4640
rect 20620 4684 20660 4724
rect 18508 4600 18548 4640
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 21100 4516 21140 4556
rect 1420 4432 1460 4472
rect 4300 4432 4340 4472
rect 6028 4432 6068 4472
rect 8524 4432 8564 4472
rect 4780 4348 4820 4388
rect 6220 4348 6260 4388
rect 13324 4348 13364 4388
rect 14092 4348 14132 4388
rect 14764 4348 14804 4388
rect 17356 4432 17396 4472
rect 18412 4432 18452 4472
rect 19660 4432 19700 4472
rect 2764 4264 2804 4304
rect 10252 4264 10292 4304
rect 17644 4264 17684 4304
rect 2284 4180 2324 4220
rect 6604 4180 6644 4220
rect 76 4096 116 4136
rect 1612 4096 1652 4136
rect 7852 4096 7892 4136
rect 16588 4096 16628 4136
rect 18508 4096 18548 4136
rect 11980 3928 12020 3968
rect 2764 3844 2804 3884
rect 10444 3844 10484 3884
rect 364 3760 404 3800
rect 3148 3760 3188 3800
rect 10636 3844 10676 3884
rect 3340 3760 3380 3800
rect 4108 3760 4148 3800
rect 4588 3760 4628 3800
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 5836 3760 5876 3800
rect 6124 3760 6164 3800
rect 11308 3760 11348 3800
rect 12076 3760 12116 3800
rect 16780 3760 16820 3800
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 7852 3676 7892 3716
rect 9292 3676 9332 3716
rect 1708 3592 1748 3632
rect 3052 3592 3092 3632
rect 14092 3592 14132 3632
rect 14860 3592 14900 3632
rect 17836 3592 17876 3632
rect 2668 3508 2708 3548
rect 5452 3508 5492 3548
rect 11116 3508 11156 3548
rect 12940 3508 12980 3548
rect 15820 3508 15860 3548
rect 19276 3508 19316 3548
rect 460 3424 500 3464
rect 1516 3340 1556 3380
rect 7084 3340 7124 3380
rect 16300 3424 16340 3464
rect 16876 3424 16916 3464
rect 7660 3340 7700 3380
rect 9580 3340 9620 3380
rect 13900 3340 13940 3380
rect 19372 3340 19412 3380
rect 16108 3256 16148 3296
rect 2860 3172 2900 3212
rect 17068 3172 17108 3212
rect 18700 3172 18740 3212
rect 268 3088 308 3128
rect 19756 3088 19796 3128
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 14572 3004 14612 3044
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 3532 2920 3572 2960
rect 7468 2920 7508 2960
rect 9100 2920 9140 2960
rect 844 2752 884 2792
rect 4780 2752 4820 2792
rect 10828 2752 10868 2792
rect 3532 2668 3572 2708
rect 556 2584 596 2624
rect 5548 2584 5588 2624
rect 1228 2416 1268 2456
rect 5932 2584 5972 2624
rect 6892 2668 6932 2708
rect 7660 2668 7700 2708
rect 9388 2668 9428 2708
rect 10540 2668 10580 2708
rect 17260 2668 17300 2708
rect 9100 2500 9140 2540
rect 9964 2500 10004 2540
rect 10348 2500 10388 2540
rect 10636 2500 10676 2540
rect 19660 2584 19700 2624
rect 10828 2500 10868 2540
rect 15244 2500 15284 2540
rect 21004 2416 21044 2456
rect 14572 2332 14612 2372
rect 4108 2248 4148 2288
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 9868 2248 9908 2288
rect 10156 2248 10196 2288
rect 15340 2248 15380 2288
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 8812 2164 8852 2204
rect 11212 2164 11252 2204
rect 13228 2164 13268 2204
rect 9292 2080 9332 2120
rect 11884 2080 11924 2120
rect 19564 2080 19604 2120
rect 19852 2080 19892 2120
rect 5548 1996 5588 2036
rect 5740 1996 5780 2036
rect 3628 1912 3668 1952
rect 5932 1912 5972 1952
rect 9196 1912 9236 1952
rect 1996 1828 2036 1868
rect 5644 1828 5684 1868
rect 10060 1912 10100 1952
rect 11596 1912 11636 1952
rect 18124 1912 18164 1952
rect 19372 1912 19412 1952
rect 19948 1912 19988 1952
rect 2380 1744 2420 1784
rect 1420 1660 1460 1700
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 9964 1492 10004 1532
rect 11212 1492 11252 1532
rect 17548 1492 17588 1532
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 1036 1408 1076 1448
rect 2572 1240 2612 1280
rect 3340 1240 3380 1280
rect 3724 1240 3764 1280
rect 6412 1240 6452 1280
rect 6796 1240 6836 1280
rect 6988 1240 7028 1280
rect 7180 1240 7220 1280
rect 8140 1240 8180 1280
rect 8332 1240 8372 1280
rect 8524 1240 8564 1280
rect 12556 1240 12596 1280
rect 940 1156 980 1196
rect 3436 1156 3476 1196
rect 5452 1156 5492 1196
rect 5644 1156 5684 1196
rect 10924 1156 10964 1196
rect 12748 1240 12788 1280
rect 13132 1240 13172 1280
rect 15916 1324 15956 1364
rect 13516 1240 13556 1280
rect 13708 1240 13748 1280
rect 14668 1240 14708 1280
rect 15436 1240 15476 1280
rect 15628 1240 15668 1280
rect 17452 1240 17492 1280
rect 17740 1240 17780 1280
rect 18220 1240 18260 1280
rect 11116 1156 11156 1196
rect 18412 1156 18452 1196
rect 4108 1072 4148 1112
rect 5068 1072 5108 1112
rect 8620 1072 8660 1112
rect 9580 1072 9620 1112
rect 8044 988 8084 1028
rect 13804 988 13844 1028
rect 4300 904 4340 944
rect 7372 904 7412 944
rect 7756 904 7796 944
rect 14284 904 14324 944
rect 5932 820 5972 860
rect 10924 820 10964 860
rect 11116 820 11156 860
rect 18700 820 18740 860
rect 20524 820 20564 860
rect 4684 736 4724 776
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 6220 652 6260 692
rect 7948 652 7988 692
rect 19276 652 19316 692
rect 4492 568 4532 608
rect 5356 568 5396 608
rect 9772 484 9812 524
rect 15052 484 15092 524
rect 6028 400 6068 440
rect 13612 400 13652 440
rect 6604 316 6644 356
rect 6892 316 6932 356
rect 1132 232 1172 272
rect 4780 232 4820 272
rect 5836 232 5876 272
rect 5260 148 5300 188
rect 268 64 308 104
rect 9772 148 9812 188
rect 6028 64 6068 104
rect 11308 232 11348 272
rect 16300 232 16340 272
rect 16780 64 16820 104
<< metal4 >>
rect 1228 42860 1268 42869
rect 1036 40340 1076 40349
rect 363 39164 405 39173
rect 363 39124 364 39164
rect 404 39124 405 39164
rect 363 39115 405 39124
rect 171 36560 213 36569
rect 171 36520 172 36560
rect 212 36520 213 36560
rect 171 36511 213 36520
rect 76 34880 116 34889
rect 76 29672 116 34840
rect 76 29623 116 29632
rect 172 29000 212 36511
rect 76 28960 212 29000
rect 76 21785 116 28960
rect 171 28328 213 28337
rect 171 28288 172 28328
rect 212 28288 213 28328
rect 171 28279 213 28288
rect 172 24968 212 28279
rect 172 24919 212 24928
rect 267 22196 309 22205
rect 267 22156 268 22196
rect 308 22156 309 22196
rect 267 22147 309 22156
rect 75 21776 117 21785
rect 75 21736 76 21776
rect 116 21736 117 21776
rect 75 21727 117 21736
rect 268 21608 308 22147
rect 268 21559 308 21568
rect 172 17660 212 17669
rect 76 15056 116 15065
rect 76 4136 116 15016
rect 172 7832 212 17620
rect 364 12620 404 39115
rect 556 38996 596 39005
rect 460 35720 500 35729
rect 460 29084 500 35680
rect 460 29035 500 29044
rect 556 21449 596 38956
rect 940 37736 980 37745
rect 844 35804 884 35813
rect 748 32024 788 32033
rect 651 29672 693 29681
rect 651 29632 652 29672
rect 692 29632 693 29672
rect 651 29623 693 29632
rect 555 21440 597 21449
rect 555 21400 556 21440
rect 596 21400 597 21440
rect 555 21391 597 21400
rect 652 20180 692 29623
rect 748 29093 788 31984
rect 844 29168 884 35764
rect 940 33041 980 37696
rect 939 33032 981 33041
rect 939 32992 940 33032
rect 980 32992 981 33032
rect 939 32983 981 32992
rect 940 32864 980 32873
rect 940 29336 980 32824
rect 940 29287 980 29296
rect 844 29128 980 29168
rect 747 29084 789 29093
rect 747 29044 748 29084
rect 788 29044 789 29084
rect 747 29035 789 29044
rect 844 29000 884 29009
rect 652 20140 788 20180
rect 364 12571 404 12580
rect 364 12452 404 12461
rect 267 12284 309 12293
rect 267 12244 268 12284
rect 308 12244 309 12284
rect 267 12235 309 12244
rect 172 7783 212 7792
rect 76 4087 116 4096
rect 268 3128 308 12235
rect 364 3800 404 12412
rect 459 11948 501 11957
rect 459 11908 460 11948
rect 500 11908 501 11948
rect 459 11899 501 11908
rect 364 3751 404 3760
rect 460 3464 500 11899
rect 460 3415 500 3424
rect 556 10856 596 10865
rect 268 3079 308 3088
rect 556 2624 596 10816
rect 748 6992 788 20140
rect 844 12872 884 28960
rect 844 12823 884 12832
rect 748 6943 788 6952
rect 844 10772 884 10781
rect 651 6236 693 6245
rect 651 6196 652 6236
rect 692 6196 693 6236
rect 651 6187 693 6196
rect 652 6102 692 6187
rect 844 2792 884 10732
rect 940 10604 980 29128
rect 1036 13460 1076 40300
rect 1132 38744 1172 38753
rect 1132 37232 1172 38704
rect 1132 37183 1172 37192
rect 1228 33956 1268 42820
rect 4780 42692 4820 42701
rect 2860 42272 2900 42281
rect 1612 41432 1652 41441
rect 1323 41180 1365 41189
rect 1323 41140 1324 41180
rect 1364 41140 1365 41180
rect 1323 41131 1365 41140
rect 1324 41046 1364 41131
rect 1420 40508 1460 40517
rect 1420 40349 1460 40468
rect 1419 40340 1461 40349
rect 1419 40300 1420 40340
rect 1460 40300 1461 40340
rect 1419 40291 1461 40300
rect 1420 40172 1460 40181
rect 1323 37484 1365 37493
rect 1323 37444 1324 37484
rect 1364 37444 1365 37484
rect 1323 37435 1365 37444
rect 1324 37350 1364 37435
rect 1132 33916 1268 33956
rect 1324 36560 1364 36569
rect 1324 35636 1364 36520
rect 1132 32444 1172 33916
rect 1227 33704 1269 33713
rect 1227 33664 1228 33704
rect 1268 33664 1269 33704
rect 1324 33704 1364 35596
rect 1420 33872 1460 40132
rect 1516 37988 1556 37997
rect 1516 36056 1556 37948
rect 1612 37661 1652 41392
rect 2572 41432 2612 41441
rect 2380 41348 2420 41357
rect 1804 40424 1844 40433
rect 1707 39752 1749 39761
rect 1707 39712 1708 39752
rect 1748 39712 1749 39752
rect 1707 39703 1749 39712
rect 1708 39618 1748 39703
rect 1708 39248 1748 39257
rect 1611 37652 1653 37661
rect 1611 37612 1612 37652
rect 1652 37612 1653 37652
rect 1611 37603 1653 37612
rect 1516 34385 1556 36016
rect 1515 34376 1557 34385
rect 1515 34336 1516 34376
rect 1556 34336 1557 34376
rect 1515 34327 1557 34336
rect 1612 34376 1652 37603
rect 1708 34544 1748 39208
rect 1804 35468 1844 40384
rect 1804 35419 1844 35428
rect 1900 40256 1940 40265
rect 1900 39164 1940 40216
rect 1900 36476 1940 39124
rect 1708 34495 1748 34504
rect 1804 35300 1844 35309
rect 1612 34327 1652 34336
rect 1804 34292 1844 35260
rect 1420 33823 1460 33832
rect 1708 34252 1844 34292
rect 1324 33664 1460 33704
rect 1227 33655 1269 33664
rect 1228 33570 1268 33655
rect 1132 32395 1172 32404
rect 1228 33200 1268 33209
rect 1228 31277 1268 33160
rect 1227 31268 1269 31277
rect 1227 31228 1228 31268
rect 1268 31228 1269 31268
rect 1227 31219 1269 31228
rect 1323 31184 1365 31193
rect 1323 31144 1324 31184
rect 1364 31144 1365 31184
rect 1323 31135 1365 31144
rect 1227 31100 1269 31109
rect 1227 31060 1228 31100
rect 1268 31060 1269 31100
rect 1227 31051 1269 31060
rect 1131 30092 1173 30101
rect 1131 30052 1132 30092
rect 1172 30052 1173 30092
rect 1131 30043 1173 30052
rect 1036 13411 1076 13420
rect 940 10555 980 10564
rect 939 5564 981 5573
rect 939 5524 940 5564
rect 980 5524 981 5564
rect 939 5515 981 5524
rect 844 2743 884 2752
rect 556 2575 596 2584
rect 940 1196 980 5515
rect 1035 5396 1077 5405
rect 1035 5356 1036 5396
rect 1076 5356 1077 5396
rect 1035 5347 1077 5356
rect 1036 5262 1076 5347
rect 1035 5144 1077 5153
rect 1035 5104 1036 5144
rect 1076 5104 1077 5144
rect 1035 5095 1077 5104
rect 1036 1448 1076 5095
rect 1036 1399 1076 1408
rect 940 1147 980 1156
rect 1132 272 1172 30043
rect 1228 28160 1268 31051
rect 1324 31050 1364 31135
rect 1420 30932 1460 33664
rect 1611 33032 1653 33041
rect 1611 32992 1612 33032
rect 1652 32992 1653 33032
rect 1611 32983 1653 32992
rect 1515 32108 1557 32117
rect 1515 32068 1516 32108
rect 1556 32068 1557 32108
rect 1515 32059 1557 32068
rect 1516 31974 1556 32059
rect 1515 31856 1557 31865
rect 1515 31816 1516 31856
rect 1556 31816 1557 31856
rect 1515 31807 1557 31816
rect 1228 28111 1268 28120
rect 1324 30892 1460 30932
rect 1324 26480 1364 30892
rect 1419 30764 1461 30773
rect 1419 30724 1420 30764
rect 1460 30724 1461 30764
rect 1419 30715 1461 30724
rect 1324 26431 1364 26440
rect 1227 24632 1269 24641
rect 1227 24592 1228 24632
rect 1268 24592 1269 24632
rect 1227 24583 1269 24592
rect 1420 24632 1460 30715
rect 1420 24583 1460 24592
rect 1228 24498 1268 24583
rect 1227 22448 1269 22457
rect 1227 22408 1228 22448
rect 1268 22408 1269 22448
rect 1227 22399 1269 22408
rect 1228 22280 1268 22399
rect 1228 22231 1268 22240
rect 1419 19844 1461 19853
rect 1419 19804 1420 19844
rect 1460 19804 1461 19844
rect 1419 19795 1461 19804
rect 1227 17828 1269 17837
rect 1227 17788 1228 17828
rect 1268 17788 1269 17828
rect 1227 17779 1269 17788
rect 1228 16904 1268 17779
rect 1323 17744 1365 17753
rect 1323 17704 1324 17744
rect 1364 17704 1365 17744
rect 1323 17695 1365 17704
rect 1228 16855 1268 16864
rect 1324 16736 1364 17695
rect 1228 16696 1364 16736
rect 1228 10100 1268 16696
rect 1323 16232 1365 16241
rect 1323 16192 1324 16232
rect 1364 16192 1365 16232
rect 1323 16183 1365 16192
rect 1324 10184 1364 16183
rect 1420 15056 1460 19795
rect 1516 18500 1556 31807
rect 1612 30773 1652 32983
rect 1611 30764 1653 30773
rect 1611 30724 1612 30764
rect 1652 30724 1653 30764
rect 1611 30715 1653 30724
rect 1611 30596 1653 30605
rect 1611 30556 1612 30596
rect 1652 30556 1653 30596
rect 1611 30547 1653 30556
rect 1612 29000 1652 30547
rect 1708 29756 1748 34252
rect 1803 34124 1845 34133
rect 1803 34084 1804 34124
rect 1844 34084 1845 34124
rect 1803 34075 1845 34084
rect 1804 30605 1844 34075
rect 1803 30596 1845 30605
rect 1803 30556 1804 30596
rect 1844 30556 1845 30596
rect 1803 30547 1845 30556
rect 1708 29716 1844 29756
rect 1612 28960 1748 29000
rect 1612 23876 1652 23885
rect 1612 20861 1652 23836
rect 1611 20852 1653 20861
rect 1611 20812 1612 20852
rect 1652 20812 1653 20852
rect 1611 20803 1653 20812
rect 1516 18451 1556 18460
rect 1708 19172 1748 28960
rect 1804 28916 1844 29716
rect 1804 28867 1844 28876
rect 1900 27740 1940 36436
rect 1996 39332 2036 39341
rect 1996 31100 2036 39292
rect 2092 39080 2132 39089
rect 2092 38576 2132 39040
rect 2380 38996 2420 41308
rect 2092 38527 2132 38536
rect 2188 38956 2380 38996
rect 2188 38324 2228 38956
rect 2380 38947 2420 38956
rect 2092 35468 2132 35477
rect 2092 34133 2132 35428
rect 2091 34124 2133 34133
rect 2091 34084 2092 34124
rect 2132 34084 2133 34124
rect 2091 34075 2133 34084
rect 2091 32948 2133 32957
rect 2091 32908 2092 32948
rect 2132 32908 2133 32948
rect 2091 32899 2133 32908
rect 2092 32360 2132 32899
rect 2092 32311 2132 32320
rect 1996 31051 2036 31060
rect 2092 32192 2132 32201
rect 1996 29168 2036 29177
rect 1996 29009 2036 29128
rect 1995 29000 2037 29009
rect 1995 28960 1996 29000
rect 2036 28960 2037 29000
rect 1995 28951 2037 28960
rect 1940 27700 2036 27740
rect 1900 27691 1940 27700
rect 1899 23792 1941 23801
rect 1899 23752 1900 23792
rect 1940 23752 1941 23792
rect 1899 23743 1941 23752
rect 1900 23658 1940 23743
rect 1612 17744 1652 17753
rect 1516 17324 1556 17333
rect 1516 16241 1556 17284
rect 1515 16232 1557 16241
rect 1515 16192 1516 16232
rect 1556 16192 1557 16232
rect 1515 16183 1557 16192
rect 1515 16064 1557 16073
rect 1515 16024 1516 16064
rect 1556 16024 1557 16064
rect 1515 16015 1557 16024
rect 1420 15007 1460 15016
rect 1419 14720 1461 14729
rect 1419 14680 1420 14720
rect 1460 14680 1461 14720
rect 1419 14671 1461 14680
rect 1420 11360 1460 14671
rect 1516 12452 1556 16015
rect 1516 12403 1556 12412
rect 1612 15308 1652 17704
rect 1708 15560 1748 19132
rect 1708 15511 1748 15520
rect 1804 21608 1844 21617
rect 1420 11320 1556 11360
rect 1516 10184 1556 11320
rect 1324 10144 1460 10184
rect 1228 10060 1364 10100
rect 1227 8168 1269 8177
rect 1227 8128 1228 8168
rect 1268 8128 1269 8168
rect 1227 8119 1269 8128
rect 1228 5237 1268 8119
rect 1227 5228 1269 5237
rect 1227 5188 1228 5228
rect 1268 5188 1269 5228
rect 1227 5179 1269 5188
rect 1324 4892 1364 10060
rect 1324 4843 1364 4852
rect 1228 4808 1268 4819
rect 1228 4733 1268 4768
rect 1227 4724 1269 4733
rect 1227 4684 1228 4724
rect 1268 4684 1269 4724
rect 1227 4675 1269 4684
rect 1420 4472 1460 10144
rect 1516 10135 1556 10144
rect 1516 8924 1556 8933
rect 1516 6488 1556 8884
rect 1612 8000 1652 15268
rect 1612 7085 1652 7960
rect 1708 11612 1748 11621
rect 1611 7076 1653 7085
rect 1611 7036 1612 7076
rect 1652 7036 1653 7076
rect 1611 7027 1653 7036
rect 1516 6439 1556 6448
rect 1515 5816 1557 5825
rect 1515 5776 1516 5816
rect 1556 5776 1557 5816
rect 1515 5767 1557 5776
rect 1420 4423 1460 4432
rect 1516 3380 1556 5767
rect 1612 4136 1652 7027
rect 1612 4087 1652 4096
rect 1708 3632 1748 11572
rect 1804 10688 1844 21568
rect 1996 21272 2036 27700
rect 1996 20768 2036 21232
rect 1996 20719 2036 20728
rect 2092 21356 2132 32152
rect 2188 26237 2228 38284
rect 2379 38324 2421 38333
rect 2379 38284 2380 38324
rect 2420 38284 2421 38324
rect 2379 38275 2421 38284
rect 2380 38156 2420 38275
rect 2380 38107 2420 38116
rect 2572 38156 2612 41392
rect 2572 38107 2612 38116
rect 2764 39164 2804 39173
rect 2764 37820 2804 39124
rect 2764 37771 2804 37780
rect 2572 37652 2612 37661
rect 2284 36896 2324 36905
rect 2187 26228 2229 26237
rect 2187 26188 2188 26228
rect 2228 26188 2229 26228
rect 2187 26179 2229 26188
rect 2188 21608 2228 26179
rect 2284 25397 2324 36856
rect 2476 35300 2516 35309
rect 2379 35216 2421 35225
rect 2379 35176 2380 35216
rect 2420 35176 2421 35216
rect 2379 35167 2421 35176
rect 2380 35082 2420 35167
rect 2379 34376 2421 34385
rect 2379 34336 2380 34376
rect 2420 34336 2421 34376
rect 2379 34327 2421 34336
rect 2380 31865 2420 34327
rect 2379 31856 2421 31865
rect 2379 31816 2380 31856
rect 2420 31816 2421 31856
rect 2379 31807 2421 31816
rect 2476 31697 2516 35260
rect 2475 31688 2517 31697
rect 2475 31648 2476 31688
rect 2516 31648 2517 31688
rect 2475 31639 2517 31648
rect 2380 31604 2420 31613
rect 2283 25388 2325 25397
rect 2283 25348 2284 25388
rect 2324 25348 2325 25388
rect 2283 25339 2325 25348
rect 2284 25253 2324 25339
rect 2380 24464 2420 31564
rect 2475 30848 2517 30857
rect 2475 30808 2476 30848
rect 2516 30808 2517 30848
rect 2475 30799 2517 30808
rect 2476 27656 2516 30799
rect 2476 27607 2516 27616
rect 2475 26396 2517 26405
rect 2475 26356 2476 26396
rect 2516 26356 2517 26396
rect 2475 26347 2517 26356
rect 2476 26262 2516 26347
rect 2380 24415 2420 24424
rect 2476 26144 2516 26153
rect 2476 24548 2516 26104
rect 2188 21559 2228 21568
rect 2284 22700 2324 22709
rect 2092 19256 2132 21316
rect 2092 19207 2132 19216
rect 2188 20012 2228 20021
rect 2092 17072 2132 17081
rect 1996 14636 2036 14645
rect 1804 10639 1844 10648
rect 1900 14552 1940 14561
rect 1803 8756 1845 8765
rect 1803 8716 1804 8756
rect 1844 8716 1845 8756
rect 1803 8707 1845 8716
rect 1804 8622 1844 8707
rect 1900 6152 1940 14512
rect 1900 6103 1940 6112
rect 1996 5648 2036 14596
rect 2092 11948 2132 17032
rect 2092 10268 2132 11908
rect 2092 10219 2132 10228
rect 2091 9428 2133 9437
rect 2091 9388 2092 9428
rect 2132 9388 2133 9428
rect 2091 9379 2133 9388
rect 1996 5599 2036 5608
rect 1708 3583 1748 3592
rect 1516 3331 1556 3340
rect 2092 2540 2132 9379
rect 2188 6656 2228 19972
rect 2284 10772 2324 22660
rect 2476 20096 2516 24508
rect 2476 20047 2516 20056
rect 2476 14972 2516 14981
rect 2379 13880 2421 13889
rect 2379 13840 2380 13880
rect 2420 13840 2421 13880
rect 2379 13831 2421 13840
rect 2284 10723 2324 10732
rect 2188 6607 2228 6616
rect 2284 10184 2324 10193
rect 2284 4220 2324 10144
rect 2380 7580 2420 13831
rect 2476 13628 2516 14932
rect 2476 13579 2516 13588
rect 2476 13208 2516 13217
rect 2476 9344 2516 13168
rect 2476 9295 2516 9304
rect 2380 7531 2420 7540
rect 2379 5732 2421 5741
rect 2379 5692 2380 5732
rect 2420 5692 2421 5732
rect 2379 5683 2421 5692
rect 2284 4171 2324 4180
rect 1996 2500 2132 2540
rect 1227 2456 1269 2465
rect 1227 2416 1228 2456
rect 1268 2416 1269 2456
rect 1227 2407 1269 2416
rect 1228 2322 1268 2407
rect 1996 1868 2036 2500
rect 1996 1819 2036 1828
rect 2380 1784 2420 5683
rect 2380 1735 2420 1744
rect 1419 1700 1461 1709
rect 1419 1660 1420 1700
rect 1460 1660 1461 1700
rect 1419 1651 1461 1660
rect 1420 1566 1460 1651
rect 2572 1280 2612 37612
rect 2764 37400 2804 37409
rect 2764 33956 2804 37360
rect 2860 36308 2900 42232
rect 4684 42188 4724 42197
rect 4204 41936 4244 41945
rect 2956 41852 2996 41861
rect 2956 38576 2996 41812
rect 3340 41264 3380 41273
rect 3148 39668 3188 39677
rect 2956 38527 2996 38536
rect 3052 39164 3092 39173
rect 2956 37904 2996 37913
rect 2956 36896 2996 37864
rect 3052 37736 3092 39124
rect 3052 37687 3092 37696
rect 2956 36847 2996 36856
rect 2860 36268 2996 36308
rect 2668 33916 2804 33956
rect 2860 36140 2900 36149
rect 2668 32453 2708 33916
rect 2764 33788 2804 33797
rect 2764 33620 2804 33748
rect 2764 33571 2804 33580
rect 2763 32528 2805 32537
rect 2763 32488 2764 32528
rect 2804 32488 2805 32528
rect 2763 32479 2805 32488
rect 2667 32444 2709 32453
rect 2667 32404 2668 32444
rect 2708 32404 2709 32444
rect 2667 32395 2709 32404
rect 2667 32108 2709 32117
rect 2667 32068 2668 32108
rect 2708 32068 2709 32108
rect 2667 32059 2709 32068
rect 2668 31856 2708 32059
rect 2668 31807 2708 31816
rect 2667 31688 2709 31697
rect 2667 31648 2668 31688
rect 2708 31648 2709 31688
rect 2667 31639 2709 31648
rect 2668 30932 2708 31639
rect 2764 31184 2804 32479
rect 2764 31135 2804 31144
rect 2860 31268 2900 36100
rect 2956 33956 2996 36268
rect 2956 33907 2996 33916
rect 3052 35468 3092 35477
rect 2956 33452 2996 33461
rect 2956 32696 2996 33412
rect 2956 32647 2996 32656
rect 2955 32444 2997 32453
rect 2955 32404 2956 32444
rect 2996 32404 2997 32444
rect 2955 32395 2997 32404
rect 2668 30883 2708 30892
rect 2764 30680 2804 30689
rect 2764 29840 2804 30640
rect 2667 29168 2709 29177
rect 2667 29128 2668 29168
rect 2708 29128 2709 29168
rect 2667 29119 2709 29128
rect 2668 29009 2708 29119
rect 2667 29000 2709 29009
rect 2667 28960 2668 29000
rect 2708 28960 2709 29000
rect 2667 28951 2709 28960
rect 2668 27908 2708 27917
rect 2668 23969 2708 27868
rect 2764 26732 2804 29800
rect 2764 26683 2804 26692
rect 2763 26564 2805 26573
rect 2763 26524 2764 26564
rect 2804 26524 2805 26564
rect 2763 26515 2805 26524
rect 2667 23960 2709 23969
rect 2667 23920 2668 23960
rect 2708 23920 2709 23960
rect 2667 23911 2709 23920
rect 2764 23456 2804 26515
rect 2764 23407 2804 23416
rect 2764 23120 2804 23129
rect 2764 21188 2804 23080
rect 2764 21139 2804 21148
rect 2860 20936 2900 31228
rect 2956 26396 2996 32395
rect 3052 31604 3092 35428
rect 3052 31555 3092 31564
rect 3052 30848 3092 30857
rect 3052 29504 3092 30808
rect 3148 30092 3188 39628
rect 3340 39080 3380 41224
rect 4108 41264 4148 41273
rect 3532 41012 3572 41021
rect 3340 39031 3380 39040
rect 3436 40256 3476 40265
rect 3436 40088 3476 40216
rect 3339 38156 3381 38165
rect 3339 38116 3340 38156
rect 3380 38116 3381 38156
rect 3339 38107 3381 38116
rect 3340 38022 3380 38107
rect 3148 30043 3188 30052
rect 3244 37400 3284 37409
rect 3052 29455 3092 29464
rect 3051 29084 3093 29093
rect 3051 29044 3052 29084
rect 3092 29044 3093 29084
rect 3051 29035 3093 29044
rect 3052 28925 3092 29035
rect 3244 29000 3284 37360
rect 3436 35720 3476 40048
rect 3532 36140 3572 40972
rect 3688 40844 4056 40853
rect 3728 40804 3770 40844
rect 3810 40804 3852 40844
rect 3892 40804 3934 40844
rect 3974 40804 4016 40844
rect 3688 40795 4056 40804
rect 3627 39836 3669 39845
rect 3627 39796 3628 39836
rect 3668 39796 3669 39836
rect 3627 39787 3669 39796
rect 3628 39702 3668 39787
rect 3688 39332 4056 39341
rect 3728 39292 3770 39332
rect 3810 39292 3852 39332
rect 3892 39292 3934 39332
rect 3974 39292 4016 39332
rect 3688 39283 4056 39292
rect 4012 39164 4052 39173
rect 4012 38828 4052 39124
rect 4108 38996 4148 41224
rect 4108 38947 4148 38956
rect 4012 38779 4052 38788
rect 4204 38576 4244 41896
rect 4300 40088 4340 40097
rect 4300 39509 4340 40048
rect 4395 39752 4437 39761
rect 4395 39712 4396 39752
rect 4436 39712 4437 39752
rect 4395 39703 4437 39712
rect 4299 39500 4341 39509
rect 4299 39460 4300 39500
rect 4340 39460 4341 39500
rect 4299 39451 4341 39460
rect 4204 38527 4244 38536
rect 4300 39080 4340 39089
rect 3688 37820 4056 37829
rect 3728 37780 3770 37820
rect 3810 37780 3852 37820
rect 3892 37780 3934 37820
rect 3974 37780 4016 37820
rect 3688 37771 4056 37780
rect 3723 37568 3765 37577
rect 3723 37528 3724 37568
rect 3764 37528 3765 37568
rect 3723 37519 3765 37528
rect 3724 37434 3764 37519
rect 4108 37484 4148 37493
rect 4108 36569 4148 37444
rect 4107 36560 4149 36569
rect 4107 36520 4108 36560
rect 4148 36520 4149 36560
rect 4107 36511 4149 36520
rect 3688 36308 4056 36317
rect 3728 36268 3770 36308
rect 3810 36268 3852 36308
rect 3892 36268 3934 36308
rect 3974 36268 4016 36308
rect 3688 36259 4056 36268
rect 3532 36100 3668 36140
rect 3436 35680 3572 35720
rect 3436 35552 3476 35561
rect 3339 35384 3381 35393
rect 3339 35344 3340 35384
rect 3380 35344 3381 35384
rect 3339 35335 3381 35344
rect 3340 35250 3380 35335
rect 3436 33368 3476 35512
rect 3340 33032 3380 33041
rect 3340 31361 3380 32992
rect 3339 31352 3381 31361
rect 3339 31312 3340 31352
rect 3380 31312 3381 31352
rect 3339 31303 3381 31312
rect 3148 28960 3284 29000
rect 3340 31184 3380 31193
rect 3051 28916 3093 28925
rect 3051 28876 3052 28916
rect 3092 28876 3093 28916
rect 3051 28867 3093 28876
rect 3052 26984 3092 28867
rect 3052 26935 3092 26944
rect 2956 26347 2996 26356
rect 3148 26060 3188 28960
rect 2668 20432 2708 20441
rect 2668 19508 2708 20392
rect 2668 19459 2708 19468
rect 2764 19844 2804 19853
rect 2764 19424 2804 19804
rect 2764 19375 2804 19384
rect 2764 16148 2804 16157
rect 2668 15812 2708 15821
rect 2668 6488 2708 15772
rect 2764 15560 2804 16108
rect 2764 10436 2804 15520
rect 2860 11033 2900 20896
rect 2956 26020 3188 26060
rect 3244 27992 3284 28001
rect 2956 20180 2996 26020
rect 3147 25892 3189 25901
rect 3147 25852 3148 25892
rect 3188 25852 3189 25892
rect 3147 25843 3189 25852
rect 2956 18332 2996 20140
rect 2956 18283 2996 18292
rect 3052 23792 3092 23801
rect 3052 23372 3092 23752
rect 3052 16316 3092 23332
rect 3148 18500 3188 25843
rect 3244 25136 3284 27952
rect 3340 26573 3380 31144
rect 3436 28748 3476 33328
rect 3532 32705 3572 35680
rect 3628 35384 3668 36100
rect 3628 35335 3668 35344
rect 4108 35132 4148 35141
rect 3688 34796 4056 34805
rect 3728 34756 3770 34796
rect 3810 34756 3852 34796
rect 3892 34756 3934 34796
rect 3974 34756 4016 34796
rect 3688 34747 4056 34756
rect 4012 34628 4052 34637
rect 4012 34208 4052 34588
rect 4108 34376 4148 35092
rect 4108 34327 4148 34336
rect 4012 34168 4148 34208
rect 3628 33545 3668 33630
rect 3627 33536 3669 33545
rect 3627 33496 3628 33536
rect 3668 33496 3669 33536
rect 3627 33487 3669 33496
rect 3688 33284 4056 33293
rect 3728 33244 3770 33284
rect 3810 33244 3852 33284
rect 3892 33244 3934 33284
rect 3974 33244 4016 33284
rect 3688 33235 4056 33244
rect 3916 32948 3956 32957
rect 3531 32696 3573 32705
rect 3531 32656 3532 32696
rect 3572 32656 3573 32696
rect 3531 32647 3573 32656
rect 3532 32537 3572 32647
rect 3531 32528 3573 32537
rect 3531 32488 3532 32528
rect 3572 32488 3573 32528
rect 3531 32479 3573 32488
rect 3531 32360 3573 32369
rect 3531 32320 3532 32360
rect 3572 32320 3573 32360
rect 3531 32311 3573 32320
rect 3916 32360 3956 32908
rect 3916 32311 3956 32320
rect 4108 32948 4148 34168
rect 4300 33200 4340 39040
rect 4396 35636 4436 39703
rect 4492 39668 4532 39677
rect 4492 37745 4532 39628
rect 4684 39668 4724 42148
rect 4684 39619 4724 39628
rect 4588 38240 4628 38249
rect 4491 37736 4533 37745
rect 4491 37696 4492 37736
rect 4532 37696 4533 37736
rect 4491 37687 4533 37696
rect 4396 35587 4436 35596
rect 4492 37484 4532 37493
rect 4492 34628 4532 37444
rect 4492 34579 4532 34588
rect 4300 33160 4436 33200
rect 3532 31688 3572 32311
rect 4108 32024 4148 32908
rect 3688 31772 4056 31781
rect 3728 31732 3770 31772
rect 3810 31732 3852 31772
rect 3892 31732 3934 31772
rect 3974 31732 4016 31772
rect 3688 31723 4056 31732
rect 3532 31639 3572 31648
rect 3628 31604 3668 31613
rect 3628 31520 3668 31564
rect 3436 28699 3476 28708
rect 3532 31480 3668 31520
rect 3435 28412 3477 28421
rect 3435 28372 3436 28412
rect 3476 28372 3477 28412
rect 3435 28363 3477 28372
rect 3339 26564 3381 26573
rect 3339 26524 3340 26564
rect 3380 26524 3381 26564
rect 3339 26515 3381 26524
rect 3340 26396 3380 26405
rect 3340 25556 3380 26356
rect 3436 26312 3476 28363
rect 3436 26263 3476 26272
rect 3340 25507 3380 25516
rect 3244 25087 3284 25096
rect 3532 23120 3572 31480
rect 4012 31268 4052 31277
rect 4012 30932 4052 31228
rect 4108 31109 4148 31984
rect 4204 33032 4244 33041
rect 4107 31100 4149 31109
rect 4107 31060 4108 31100
rect 4148 31060 4149 31100
rect 4107 31051 4149 31060
rect 4012 30680 4052 30892
rect 4012 30631 4052 30640
rect 4108 30596 4148 30605
rect 3688 30260 4056 30269
rect 3728 30220 3770 30260
rect 3810 30220 3852 30260
rect 3892 30220 3934 30260
rect 3974 30220 4016 30260
rect 3688 30211 4056 30220
rect 3688 28748 4056 28757
rect 3728 28708 3770 28748
rect 3810 28708 3852 28748
rect 3892 28708 3934 28748
rect 3974 28708 4016 28748
rect 3688 28699 4056 28708
rect 3688 27236 4056 27245
rect 3728 27196 3770 27236
rect 3810 27196 3852 27236
rect 3892 27196 3934 27236
rect 3974 27196 4016 27236
rect 3688 27187 4056 27196
rect 3628 27068 3668 27077
rect 3628 25901 3668 27028
rect 3724 26396 3764 26405
rect 3724 25985 3764 26356
rect 3723 25976 3765 25985
rect 3723 25936 3724 25976
rect 3764 25936 3765 25976
rect 3723 25927 3765 25936
rect 3627 25892 3669 25901
rect 3627 25852 3628 25892
rect 3668 25852 3669 25892
rect 3627 25843 3669 25852
rect 3688 25724 4056 25733
rect 3728 25684 3770 25724
rect 3810 25684 3852 25724
rect 3892 25684 3934 25724
rect 3974 25684 4016 25724
rect 3688 25675 4056 25684
rect 3688 24212 4056 24221
rect 3728 24172 3770 24212
rect 3810 24172 3852 24212
rect 3892 24172 3934 24212
rect 3974 24172 4016 24212
rect 3688 24163 4056 24172
rect 3723 23960 3765 23969
rect 3723 23920 3724 23960
rect 3764 23920 3765 23960
rect 3723 23911 3765 23920
rect 3724 23624 3764 23911
rect 3724 23575 3764 23584
rect 3340 23080 3572 23120
rect 4108 23540 4148 30556
rect 4204 29924 4244 32992
rect 4204 26825 4244 29884
rect 4300 32780 4340 32789
rect 4300 32528 4340 32740
rect 4300 26900 4340 32488
rect 4396 30932 4436 33160
rect 4491 32948 4533 32957
rect 4491 32908 4492 32948
rect 4532 32908 4533 32948
rect 4491 32899 4533 32908
rect 4396 30883 4436 30892
rect 4492 27824 4532 32899
rect 4588 31268 4628 38200
rect 4683 37736 4725 37745
rect 4683 37696 4684 37736
rect 4724 37696 4725 37736
rect 4683 37687 4725 37696
rect 4684 37493 4724 37687
rect 4683 37484 4725 37493
rect 4683 37444 4684 37484
rect 4724 37444 4725 37484
rect 4683 37435 4725 37444
rect 4780 36140 4820 42652
rect 18508 42692 18548 42701
rect 10252 42356 10292 42365
rect 10156 42188 10196 42197
rect 7852 41852 7892 41861
rect 4928 41600 5296 41609
rect 4968 41560 5010 41600
rect 5050 41560 5092 41600
rect 5132 41560 5174 41600
rect 5214 41560 5256 41600
rect 4928 41551 5296 41560
rect 6699 41180 6741 41189
rect 6699 41140 6700 41180
rect 6740 41140 6741 41180
rect 6699 41131 6741 41140
rect 4876 41012 4916 41021
rect 4876 40256 4916 40972
rect 5643 40508 5685 40517
rect 5643 40468 5644 40508
rect 5684 40468 5685 40508
rect 5643 40459 5685 40468
rect 5644 40374 5684 40459
rect 4876 40207 4916 40216
rect 4928 40088 5296 40097
rect 4968 40048 5010 40088
rect 5050 40048 5092 40088
rect 5132 40048 5174 40088
rect 5214 40048 5256 40088
rect 4928 40039 5296 40048
rect 6027 39836 6069 39845
rect 6027 39796 6028 39836
rect 6068 39796 6069 39836
rect 6027 39787 6069 39796
rect 5740 39668 5780 39677
rect 4928 38576 5296 38585
rect 4968 38536 5010 38576
rect 5050 38536 5092 38576
rect 5132 38536 5174 38576
rect 5214 38536 5256 38576
rect 4928 38527 5296 38536
rect 5548 38240 5588 38249
rect 4875 38072 4917 38081
rect 4875 38032 4876 38072
rect 4916 38032 4917 38072
rect 4875 38023 4917 38032
rect 4876 37938 4916 38023
rect 4928 37064 5296 37073
rect 4968 37024 5010 37064
rect 5050 37024 5092 37064
rect 5132 37024 5174 37064
rect 5214 37024 5256 37064
rect 4928 37015 5296 37024
rect 5452 36644 5492 36653
rect 5259 36560 5301 36569
rect 5259 36520 5260 36560
rect 5300 36520 5301 36560
rect 5259 36511 5301 36520
rect 5260 36426 5300 36511
rect 4780 36091 4820 36100
rect 4780 35972 4820 35981
rect 4683 35384 4725 35393
rect 4683 35344 4684 35384
rect 4724 35344 4725 35384
rect 4683 35335 4725 35344
rect 4588 31219 4628 31228
rect 4492 27775 4532 27784
rect 4203 26816 4245 26825
rect 4203 26776 4204 26816
rect 4244 26776 4245 26816
rect 4203 26767 4245 26776
rect 4204 26396 4244 26767
rect 4300 26648 4340 26860
rect 4300 26599 4340 26608
rect 4491 26396 4533 26405
rect 4204 26356 4436 26396
rect 4203 25976 4245 25985
rect 4203 25936 4204 25976
rect 4244 25936 4245 25976
rect 4203 25927 4245 25936
rect 4204 25842 4244 25927
rect 3148 18451 3188 18460
rect 3244 22532 3284 22541
rect 3052 16267 3092 16276
rect 3148 18332 3188 18341
rect 3148 15896 3188 18292
rect 3148 15728 3188 15856
rect 3244 15812 3284 22492
rect 3340 22112 3380 23080
rect 3340 21440 3380 22072
rect 3436 22952 3476 22961
rect 3436 21944 3476 22912
rect 4108 22868 4148 23500
rect 4108 22819 4148 22828
rect 4300 23876 4340 23885
rect 4300 23036 4340 23836
rect 3688 22700 4056 22709
rect 3728 22660 3770 22700
rect 3810 22660 3852 22700
rect 3892 22660 3934 22700
rect 3974 22660 4016 22700
rect 3688 22651 4056 22660
rect 3436 21895 3476 21904
rect 3532 22448 3572 22457
rect 3435 21524 3477 21533
rect 3435 21484 3436 21524
rect 3476 21484 3477 21524
rect 3435 21475 3477 21484
rect 3340 21391 3380 21400
rect 3436 21390 3476 21475
rect 3339 21272 3381 21281
rect 3339 21232 3340 21272
rect 3380 21232 3381 21272
rect 3339 21223 3381 21232
rect 3340 15896 3380 21223
rect 3532 20777 3572 22408
rect 4203 22364 4245 22373
rect 4203 22324 4204 22364
rect 4244 22324 4245 22364
rect 4203 22315 4245 22324
rect 4204 22205 4244 22315
rect 4203 22196 4245 22205
rect 4203 22156 4204 22196
rect 4244 22156 4245 22196
rect 4203 22147 4245 22156
rect 3915 21776 3957 21785
rect 3915 21736 3916 21776
rect 3956 21736 3957 21776
rect 3915 21727 3957 21736
rect 4108 21776 4148 21785
rect 3627 21608 3669 21617
rect 3627 21568 3628 21608
rect 3668 21568 3669 21608
rect 3627 21559 3669 21568
rect 3628 21365 3668 21559
rect 3916 21524 3956 21727
rect 3916 21475 3956 21484
rect 3627 21356 3669 21365
rect 3627 21316 3628 21356
rect 3668 21316 3669 21356
rect 3627 21307 3669 21316
rect 3688 21188 4056 21197
rect 3728 21148 3770 21188
rect 3810 21148 3852 21188
rect 3892 21148 3934 21188
rect 3974 21148 4016 21188
rect 3688 21139 4056 21148
rect 3531 20768 3573 20777
rect 3531 20728 3532 20768
rect 3572 20728 3573 20768
rect 3531 20719 3573 20728
rect 3436 20600 3476 20609
rect 3436 16232 3476 20560
rect 4108 20432 4148 21736
rect 4204 20441 4244 22147
rect 4108 20383 4148 20392
rect 4203 20432 4245 20441
rect 4203 20392 4204 20432
rect 4244 20392 4245 20432
rect 4203 20383 4245 20392
rect 4300 20096 4340 22996
rect 4396 20609 4436 26356
rect 4491 26356 4492 26396
rect 4532 26356 4533 26396
rect 4491 26347 4533 26356
rect 4492 26144 4532 26347
rect 4492 26095 4532 26104
rect 4684 25556 4724 35335
rect 4780 32864 4820 35932
rect 4928 35552 5296 35561
rect 4968 35512 5010 35552
rect 5050 35512 5092 35552
rect 5132 35512 5174 35552
rect 5214 35512 5256 35552
rect 4928 35503 5296 35512
rect 5356 35300 5396 35309
rect 5356 34292 5396 35260
rect 4928 34040 5296 34049
rect 4968 34000 5010 34040
rect 5050 34000 5092 34040
rect 5132 34000 5174 34040
rect 5214 34000 5256 34040
rect 4928 33991 5296 34000
rect 4780 32815 4820 32824
rect 4928 32528 5296 32537
rect 4968 32488 5010 32528
rect 5050 32488 5092 32528
rect 5132 32488 5174 32528
rect 5214 32488 5256 32528
rect 4928 32479 5296 32488
rect 4928 31016 5296 31025
rect 4968 30976 5010 31016
rect 5050 30976 5092 31016
rect 5132 30976 5174 31016
rect 5214 30976 5256 31016
rect 4928 30967 5296 30976
rect 5356 30344 5396 34252
rect 5356 30295 5396 30304
rect 5355 30176 5397 30185
rect 5355 30136 5356 30176
rect 5396 30136 5397 30176
rect 5355 30127 5397 30136
rect 4928 29504 5296 29513
rect 4968 29464 5010 29504
rect 5050 29464 5092 29504
rect 5132 29464 5174 29504
rect 5214 29464 5256 29504
rect 4928 29455 5296 29464
rect 4928 27992 5296 28001
rect 4968 27952 5010 27992
rect 5050 27952 5092 27992
rect 5132 27952 5174 27992
rect 5214 27952 5256 27992
rect 4928 27943 5296 27952
rect 4588 24716 4628 24725
rect 4491 21608 4533 21617
rect 4491 21568 4492 21608
rect 4532 21568 4533 21608
rect 4491 21559 4533 21568
rect 4492 21474 4532 21559
rect 4395 20600 4437 20609
rect 4395 20560 4396 20600
rect 4436 20560 4437 20600
rect 4395 20551 4437 20560
rect 4492 20600 4532 20609
rect 4588 20600 4628 24676
rect 4684 21608 4724 25516
rect 4684 21559 4724 21568
rect 4780 27824 4820 27833
rect 4780 24212 4820 27784
rect 4928 26480 5296 26489
rect 4968 26440 5010 26480
rect 5050 26440 5092 26480
rect 5132 26440 5174 26480
rect 5214 26440 5256 26480
rect 4928 26431 5296 26440
rect 5356 25733 5396 30127
rect 5355 25724 5397 25733
rect 5355 25684 5356 25724
rect 5396 25684 5397 25724
rect 5355 25675 5397 25684
rect 5452 25556 5492 36604
rect 5548 33797 5588 38200
rect 5644 37484 5684 37493
rect 5644 37316 5684 37444
rect 5547 33788 5589 33797
rect 5547 33748 5548 33788
rect 5588 33748 5589 33788
rect 5547 33739 5589 33748
rect 5548 33620 5588 33629
rect 5548 32789 5588 33580
rect 5547 32780 5589 32789
rect 5547 32740 5548 32780
rect 5588 32740 5589 32780
rect 5547 32731 5589 32740
rect 5548 30185 5588 32731
rect 5547 30176 5589 30185
rect 5547 30136 5548 30176
rect 5588 30136 5589 30176
rect 5547 30127 5589 30136
rect 5644 27992 5684 37276
rect 5740 37157 5780 39628
rect 6028 39257 6068 39787
rect 6220 39752 6260 39761
rect 6124 39668 6164 39677
rect 6027 39248 6069 39257
rect 6027 39208 6028 39248
rect 6068 39208 6069 39248
rect 6027 39199 6069 39208
rect 6028 39114 6068 39199
rect 6124 39173 6164 39628
rect 6123 39164 6165 39173
rect 6123 39124 6124 39164
rect 6164 39124 6165 39164
rect 6123 39115 6165 39124
rect 5932 37316 5972 37325
rect 5739 37148 5781 37157
rect 5739 37108 5740 37148
rect 5780 37108 5781 37148
rect 5739 37099 5781 37108
rect 5836 37148 5876 37176
rect 5932 37148 5972 37276
rect 5876 37108 5972 37148
rect 5836 37099 5876 37108
rect 5932 36821 5972 37108
rect 6028 37148 6068 37157
rect 5931 36812 5973 36821
rect 5931 36772 5932 36812
rect 5972 36772 5973 36812
rect 5931 36763 5973 36772
rect 5836 36728 5876 36737
rect 5740 36392 5780 36401
rect 5740 29336 5780 36352
rect 5740 29287 5780 29296
rect 5644 27943 5684 27952
rect 5356 25516 5492 25556
rect 5548 27824 5588 27833
rect 4928 24968 5296 24977
rect 4968 24928 5010 24968
rect 5050 24928 5092 24968
rect 5132 24928 5174 24968
rect 5214 24928 5256 24968
rect 4928 24919 5296 24928
rect 4532 20560 4628 20600
rect 4684 20768 4724 20777
rect 4780 20768 4820 24172
rect 5356 23801 5396 25516
rect 5452 25388 5492 25397
rect 5452 24800 5492 25348
rect 5355 23792 5397 23801
rect 5355 23752 5356 23792
rect 5396 23752 5397 23792
rect 5355 23743 5397 23752
rect 4928 23456 5296 23465
rect 4968 23416 5010 23456
rect 5050 23416 5092 23456
rect 5132 23416 5174 23456
rect 5214 23416 5256 23456
rect 4928 23407 5296 23416
rect 5356 22280 5396 22289
rect 4928 21944 5296 21953
rect 4968 21904 5010 21944
rect 5050 21904 5092 21944
rect 5132 21904 5174 21944
rect 5214 21904 5256 21944
rect 4928 21895 5296 21904
rect 4724 20728 4820 20768
rect 4492 20551 4532 20560
rect 4395 20432 4437 20441
rect 4395 20392 4396 20432
rect 4436 20392 4437 20432
rect 4395 20383 4437 20392
rect 3532 19844 3572 19853
rect 3532 17996 3572 19804
rect 4203 19844 4245 19853
rect 4203 19804 4204 19844
rect 4244 19804 4245 19844
rect 4203 19795 4245 19804
rect 4204 19710 4244 19795
rect 3688 19676 4056 19685
rect 3728 19636 3770 19676
rect 3810 19636 3852 19676
rect 3892 19636 3934 19676
rect 3974 19636 4016 19676
rect 3688 19627 4056 19636
rect 4108 19256 4148 19265
rect 3688 18164 4056 18173
rect 3728 18124 3770 18164
rect 3810 18124 3852 18164
rect 3892 18124 3934 18164
rect 3974 18124 4016 18164
rect 3688 18115 4056 18124
rect 3532 17947 3572 17956
rect 3688 16652 4056 16661
rect 3728 16612 3770 16652
rect 3810 16612 3852 16652
rect 3892 16612 3934 16652
rect 3974 16612 4016 16652
rect 3688 16603 4056 16612
rect 3436 16183 3476 16192
rect 3340 15856 3476 15896
rect 3244 15772 3380 15812
rect 3148 15688 3284 15728
rect 3148 14888 3188 14897
rect 3051 14804 3093 14813
rect 3051 14764 3052 14804
rect 3092 14764 3093 14804
rect 3051 14755 3093 14764
rect 3052 14670 3092 14755
rect 2956 13124 2996 13133
rect 3148 13124 3188 14848
rect 2956 12368 2996 13084
rect 2956 12319 2996 12328
rect 3052 13084 3188 13124
rect 2859 11024 2901 11033
rect 2859 10984 2860 11024
rect 2900 10984 2901 11024
rect 2859 10975 2901 10984
rect 2764 10387 2804 10396
rect 2860 10856 2900 10865
rect 2764 8336 2804 8345
rect 2764 6656 2804 8296
rect 2764 6607 2804 6616
rect 2668 6448 2804 6488
rect 2667 6320 2709 6329
rect 2667 6280 2668 6320
rect 2708 6280 2709 6320
rect 2667 6271 2709 6280
rect 2668 5573 2708 6271
rect 2667 5564 2709 5573
rect 2667 5524 2668 5564
rect 2708 5524 2709 5564
rect 2667 5515 2709 5524
rect 2668 4976 2708 4985
rect 2668 3548 2708 4936
rect 2764 4304 2804 6448
rect 2764 3884 2804 4264
rect 2764 3835 2804 3844
rect 2668 3499 2708 3508
rect 2860 3212 2900 10816
rect 2956 10436 2996 10445
rect 2956 9680 2996 10396
rect 2956 9631 2996 9640
rect 3052 7244 3092 13084
rect 3147 12872 3189 12881
rect 3147 12832 3148 12872
rect 3188 12832 3189 12872
rect 3147 12823 3189 12832
rect 3148 12738 3188 12823
rect 3147 12620 3189 12629
rect 3147 12580 3148 12620
rect 3188 12580 3189 12620
rect 3147 12571 3189 12580
rect 3052 7195 3092 7204
rect 3148 6824 3188 12571
rect 3244 10436 3284 15688
rect 3244 10387 3284 10396
rect 3052 6784 3188 6824
rect 3052 3632 3092 6784
rect 3148 6656 3188 6665
rect 3148 4145 3188 6616
rect 3147 4136 3189 4145
rect 3147 4096 3148 4136
rect 3188 4096 3189 4136
rect 3147 4087 3189 4096
rect 3148 3800 3188 4087
rect 3148 3751 3188 3760
rect 3340 3800 3380 15772
rect 3436 12200 3476 15856
rect 3688 15140 4056 15149
rect 3728 15100 3770 15140
rect 3810 15100 3852 15140
rect 3892 15100 3934 15140
rect 3974 15100 4016 15140
rect 3688 15091 4056 15100
rect 3532 14720 3572 14729
rect 3532 12536 3572 14680
rect 3819 14132 3861 14141
rect 3819 14092 3820 14132
rect 3860 14092 3861 14132
rect 3819 14083 3861 14092
rect 3820 14048 3860 14083
rect 3820 13997 3860 14008
rect 3688 13628 4056 13637
rect 3728 13588 3770 13628
rect 3810 13588 3852 13628
rect 3892 13588 3934 13628
rect 3974 13588 4016 13628
rect 3688 13579 4056 13588
rect 4108 13208 4148 19216
rect 4300 19088 4340 20056
rect 4300 19039 4340 19048
rect 4108 13159 4148 13168
rect 4204 16904 4244 16913
rect 4204 14804 4244 16864
rect 4204 12788 4244 14764
rect 4299 12872 4341 12881
rect 4299 12832 4300 12872
rect 4340 12832 4341 12872
rect 4299 12823 4341 12832
rect 4396 12872 4436 20383
rect 4588 15140 4628 15149
rect 4492 14720 4532 14729
rect 4492 13796 4532 14680
rect 4492 13376 4532 13756
rect 4588 13544 4628 15100
rect 4684 13796 4724 20728
rect 4779 20600 4821 20609
rect 4779 20560 4780 20600
rect 4820 20560 4821 20600
rect 4779 20551 4821 20560
rect 4780 19256 4820 20551
rect 4928 20432 5296 20441
rect 4968 20392 5010 20432
rect 5050 20392 5092 20432
rect 5132 20392 5174 20432
rect 5214 20392 5256 20432
rect 4928 20383 5296 20392
rect 4780 19207 4820 19216
rect 4928 18920 5296 18929
rect 4968 18880 5010 18920
rect 5050 18880 5092 18920
rect 5132 18880 5174 18920
rect 5214 18880 5256 18920
rect 4928 18871 5296 18880
rect 5356 18752 5396 22240
rect 5452 20432 5492 24760
rect 5452 20383 5492 20392
rect 4780 17744 4820 17753
rect 4780 17240 4820 17704
rect 5356 17660 5396 18712
rect 5356 17611 5396 17620
rect 5452 18836 5492 18845
rect 4928 17408 5296 17417
rect 4968 17368 5010 17408
rect 5050 17368 5092 17408
rect 5132 17368 5174 17408
rect 5214 17368 5256 17408
rect 4928 17359 5296 17368
rect 4780 17191 4820 17200
rect 4928 15896 5296 15905
rect 4968 15856 5010 15896
rect 5050 15856 5092 15896
rect 5132 15856 5174 15896
rect 5214 15856 5256 15896
rect 4928 15847 5296 15856
rect 4928 14384 5296 14393
rect 4968 14344 5010 14384
rect 5050 14344 5092 14384
rect 5132 14344 5174 14384
rect 5214 14344 5256 14384
rect 4928 14335 5296 14344
rect 4684 13747 4724 13756
rect 4588 13495 4628 13504
rect 4492 13336 4724 13376
rect 4396 12823 4436 12832
rect 4588 13208 4628 13217
rect 3532 12487 3572 12496
rect 4108 12748 4244 12788
rect 3436 11864 3476 12160
rect 3688 12116 4056 12125
rect 3728 12076 3770 12116
rect 3810 12076 3852 12116
rect 3892 12076 3934 12116
rect 3974 12076 4016 12116
rect 3688 12067 4056 12076
rect 3436 11815 3476 11824
rect 3723 11696 3765 11705
rect 3723 11656 3724 11696
rect 3764 11656 3765 11696
rect 3723 11647 3765 11656
rect 3724 11562 3764 11647
rect 4108 11276 4148 12748
rect 4108 11227 4148 11236
rect 4204 12620 4244 12629
rect 4108 11108 4148 11117
rect 3531 11024 3573 11033
rect 3531 10984 3532 11024
rect 3572 10984 3573 11024
rect 3531 10975 3573 10984
rect 3340 3751 3380 3760
rect 3436 10604 3476 10613
rect 3436 3632 3476 10564
rect 3052 3583 3092 3592
rect 3340 3592 3476 3632
rect 2860 3163 2900 3172
rect 2572 1231 2612 1240
rect 3340 1280 3380 3592
rect 3435 3464 3477 3473
rect 3435 3424 3436 3464
rect 3476 3424 3477 3464
rect 3435 3415 3477 3424
rect 3340 1231 3380 1240
rect 3436 1196 3476 3415
rect 3532 2960 3572 10975
rect 3688 10604 4056 10613
rect 3728 10564 3770 10604
rect 3810 10564 3852 10604
rect 3892 10564 3934 10604
rect 3974 10564 4016 10604
rect 3688 10555 4056 10564
rect 3688 9092 4056 9101
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 3688 9043 4056 9052
rect 3688 7580 4056 7589
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 3688 7531 4056 7540
rect 4108 6488 4148 11068
rect 4204 8336 4244 12580
rect 4300 12368 4340 12823
rect 4300 12328 4436 12368
rect 4300 10604 4340 10613
rect 4300 9008 4340 10564
rect 4300 8959 4340 8968
rect 4204 8287 4244 8296
rect 4108 6439 4148 6448
rect 3688 6068 4056 6077
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 3688 6019 4056 6028
rect 4300 5312 4340 5321
rect 3688 4556 4056 4565
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 3688 4507 4056 4516
rect 4300 4472 4340 5272
rect 4300 4423 4340 4432
rect 4108 3800 4148 3809
rect 3688 3044 4056 3053
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 3688 2995 4056 3004
rect 3532 2911 3572 2920
rect 3532 2708 3572 2717
rect 3532 1373 3572 2668
rect 4108 2288 4148 3760
rect 4396 2540 4436 12328
rect 4491 12116 4533 12125
rect 4491 12076 4492 12116
rect 4532 12076 4533 12116
rect 4491 12067 4533 12076
rect 4108 2239 4148 2248
rect 4300 2500 4436 2540
rect 4107 2120 4149 2129
rect 4107 2080 4108 2120
rect 4148 2080 4149 2120
rect 4107 2071 4149 2080
rect 3628 1952 3668 1963
rect 3628 1877 3668 1912
rect 3627 1868 3669 1877
rect 3627 1828 3628 1868
rect 3668 1828 3669 1868
rect 3627 1819 3669 1828
rect 3688 1532 4056 1541
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 3688 1483 4056 1492
rect 3531 1364 3573 1373
rect 3531 1324 3532 1364
rect 3572 1324 3573 1364
rect 3531 1315 3573 1324
rect 3723 1280 3765 1289
rect 3723 1240 3724 1280
rect 3764 1240 3765 1280
rect 3723 1231 3765 1240
rect 3436 1147 3476 1156
rect 3724 1146 3764 1231
rect 4108 1112 4148 2071
rect 4108 1063 4148 1072
rect 4300 944 4340 2500
rect 4300 895 4340 904
rect 4492 608 4532 12067
rect 4588 7580 4628 13168
rect 4684 9344 4724 13336
rect 5356 13208 5396 13217
rect 4928 12872 5296 12881
rect 4968 12832 5010 12872
rect 5050 12832 5092 12872
rect 5132 12832 5174 12872
rect 5214 12832 5256 12872
rect 4928 12823 5296 12832
rect 4780 12788 4820 12797
rect 4780 11948 4820 12748
rect 4780 10772 4820 11908
rect 5164 12536 5204 12545
rect 5164 11780 5204 12496
rect 5356 11864 5396 13168
rect 5356 11815 5396 11824
rect 5164 11731 5204 11740
rect 4928 11360 5296 11369
rect 5452 11360 5492 18796
rect 5548 17492 5588 27784
rect 5643 26732 5685 26741
rect 5643 26692 5644 26732
rect 5684 26692 5685 26732
rect 5643 26683 5685 26692
rect 5644 26480 5684 26683
rect 5644 26431 5684 26440
rect 5739 25892 5781 25901
rect 5739 25852 5740 25892
rect 5780 25852 5781 25892
rect 5739 25843 5781 25852
rect 5643 25724 5685 25733
rect 5643 25684 5644 25724
rect 5684 25684 5685 25724
rect 5643 25675 5685 25684
rect 5644 22457 5684 25675
rect 5740 25388 5780 25843
rect 5643 22448 5685 22457
rect 5643 22408 5644 22448
rect 5684 22408 5685 22448
rect 5643 22399 5685 22408
rect 5740 21365 5780 25348
rect 5739 21356 5781 21365
rect 5739 21316 5740 21356
rect 5780 21316 5781 21356
rect 5739 21307 5781 21316
rect 5836 20180 5876 36688
rect 6028 35309 6068 37108
rect 6027 35300 6069 35309
rect 6027 35260 6028 35300
rect 6068 35260 6069 35300
rect 6027 35251 6069 35260
rect 6123 35132 6165 35141
rect 6123 35092 6124 35132
rect 6164 35092 6165 35132
rect 6123 35083 6165 35092
rect 6124 34964 6164 35083
rect 6124 34915 6164 34924
rect 6220 32033 6260 39712
rect 6700 38996 6740 41131
rect 6987 40508 7029 40517
rect 6987 40468 6988 40508
rect 7028 40468 7029 40508
rect 6987 40459 7029 40468
rect 6700 38947 6740 38956
rect 6412 38912 6452 38921
rect 6316 35216 6356 35225
rect 6316 34880 6356 35176
rect 6219 32024 6261 32033
rect 6219 31984 6220 32024
rect 6260 31984 6261 32024
rect 6219 31975 6261 31984
rect 5931 31352 5973 31361
rect 5931 31312 5932 31352
rect 5972 31312 5973 31352
rect 5931 31303 5973 31312
rect 5932 25220 5972 31303
rect 5932 25171 5972 25180
rect 6028 29336 6068 29345
rect 5740 20140 5876 20180
rect 5740 18248 5780 20140
rect 6028 19340 6068 29296
rect 6316 27068 6356 34840
rect 6412 31193 6452 38872
rect 6795 38156 6837 38165
rect 6795 38116 6796 38156
rect 6836 38116 6837 38156
rect 6795 38107 6837 38116
rect 6508 35216 6548 35225
rect 6508 34973 6548 35176
rect 6699 35132 6741 35141
rect 6699 35092 6700 35132
rect 6740 35092 6741 35132
rect 6699 35083 6741 35092
rect 6507 34964 6549 34973
rect 6507 34924 6508 34964
rect 6548 34924 6549 34964
rect 6507 34915 6549 34924
rect 6508 34544 6548 34915
rect 6508 34495 6548 34504
rect 6604 34712 6644 34721
rect 6411 31184 6453 31193
rect 6411 31144 6412 31184
rect 6452 31144 6453 31184
rect 6411 31135 6453 31144
rect 6604 29840 6644 34672
rect 6604 29791 6644 29800
rect 6316 27019 6356 27028
rect 6508 29504 6548 29513
rect 6412 26900 6452 26909
rect 6315 26732 6357 26741
rect 6315 26692 6316 26732
rect 6356 26692 6357 26732
rect 6315 26683 6357 26692
rect 6316 26598 6356 26683
rect 6412 26312 6452 26860
rect 6508 26816 6548 29464
rect 6508 26480 6548 26776
rect 6508 26431 6548 26440
rect 6700 28244 6740 35083
rect 6412 26263 6452 26272
rect 6508 26060 6548 26069
rect 6220 25892 6260 25901
rect 6220 25397 6260 25852
rect 6316 25808 6356 25817
rect 6219 25388 6261 25397
rect 6219 25348 6220 25388
rect 6260 25348 6261 25388
rect 6219 25339 6261 25348
rect 6316 22532 6356 25768
rect 6316 22483 6356 22492
rect 6219 22448 6261 22457
rect 6219 22408 6220 22448
rect 6260 22408 6261 22448
rect 6219 22399 6261 22408
rect 6124 21944 6164 21953
rect 6124 21701 6164 21904
rect 6123 21692 6165 21701
rect 6123 21652 6124 21692
rect 6164 21652 6165 21692
rect 6123 21643 6165 21652
rect 6123 21356 6165 21365
rect 6123 21316 6124 21356
rect 6164 21316 6165 21356
rect 6123 21307 6165 21316
rect 6028 19291 6068 19300
rect 5740 17837 5780 18208
rect 6028 18920 6068 18929
rect 5739 17828 5781 17837
rect 5739 17788 5740 17828
rect 5780 17788 5781 17828
rect 5739 17779 5781 17788
rect 5548 12032 5588 17452
rect 5548 11983 5588 11992
rect 5644 15140 5684 15149
rect 5644 13880 5684 15100
rect 5836 14972 5876 14981
rect 4968 11320 5010 11360
rect 5050 11320 5092 11360
rect 5132 11320 5174 11360
rect 5214 11320 5256 11360
rect 4928 11311 5296 11320
rect 5356 11320 5492 11360
rect 5644 11780 5684 13840
rect 4780 10723 4820 10732
rect 4684 9295 4724 9304
rect 4780 10520 4820 10529
rect 4588 3800 4628 7540
rect 4684 8000 4724 8009
rect 4684 5648 4724 7960
rect 4780 6152 4820 10480
rect 4928 9848 5296 9857
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 4928 9799 5296 9808
rect 4972 9092 5012 9101
rect 4972 8681 5012 9052
rect 5356 9008 5396 11320
rect 5452 10688 5492 10697
rect 5452 10184 5492 10648
rect 5452 10025 5492 10144
rect 5548 10352 5588 10361
rect 5451 10016 5493 10025
rect 5451 9976 5452 10016
rect 5492 9976 5493 10016
rect 5451 9967 5493 9976
rect 5356 8968 5492 9008
rect 4971 8672 5013 8681
rect 4971 8632 4972 8672
rect 5012 8632 5013 8672
rect 4971 8623 5013 8632
rect 5355 8672 5397 8681
rect 5355 8632 5356 8672
rect 5396 8632 5397 8672
rect 5355 8623 5397 8632
rect 4928 8336 5296 8345
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 4928 8287 5296 8296
rect 4928 6824 5296 6833
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 4928 6775 5296 6784
rect 4780 6103 4820 6112
rect 4779 5900 4821 5909
rect 4779 5860 4780 5900
rect 4820 5860 4821 5900
rect 4779 5851 4821 5860
rect 4684 5599 4724 5608
rect 4780 4388 4820 5851
rect 4928 5312 5296 5321
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 4928 5263 5296 5272
rect 5356 4892 5396 8623
rect 5452 8000 5492 8968
rect 5452 7925 5492 7960
rect 5451 7916 5493 7925
rect 5451 7876 5452 7916
rect 5492 7876 5493 7916
rect 5451 7867 5493 7876
rect 5452 7836 5492 7867
rect 5452 6992 5492 7001
rect 5452 6152 5492 6952
rect 5452 6103 5492 6112
rect 5356 4843 5396 4852
rect 5452 5228 5492 5237
rect 5355 4640 5397 4649
rect 5355 4600 5356 4640
rect 5396 4600 5397 4640
rect 5355 4591 5397 4600
rect 4780 4339 4820 4348
rect 4588 3751 4628 3760
rect 4928 3800 5296 3809
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 4928 3751 5296 3760
rect 4780 2792 4820 2801
rect 4683 776 4725 785
rect 4683 736 4684 776
rect 4724 736 4725 776
rect 4683 727 4725 736
rect 4684 642 4724 727
rect 4492 559 4532 568
rect 1132 223 1172 232
rect 4780 272 4820 2752
rect 4928 2288 5296 2297
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 4928 2239 5296 2248
rect 5067 1364 5109 1373
rect 5067 1324 5068 1364
rect 5108 1324 5109 1364
rect 5067 1315 5109 1324
rect 5068 1112 5108 1315
rect 5068 1063 5108 1072
rect 4928 776 5296 785
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 4928 727 5296 736
rect 5356 608 5396 4591
rect 5452 3548 5492 5188
rect 5548 3641 5588 10312
rect 5644 9764 5684 11740
rect 5740 14720 5780 14729
rect 5740 9932 5780 14680
rect 5740 9883 5780 9892
rect 5836 10016 5876 14932
rect 5932 14636 5972 14645
rect 5932 10184 5972 14596
rect 5932 10135 5972 10144
rect 5644 9724 5780 9764
rect 5643 7496 5685 7505
rect 5643 7456 5644 7496
rect 5684 7456 5685 7496
rect 5643 7447 5685 7456
rect 5644 7362 5684 7447
rect 5547 3632 5589 3641
rect 5547 3592 5548 3632
rect 5588 3592 5589 3632
rect 5547 3583 5589 3592
rect 5452 3499 5492 3508
rect 5643 3548 5685 3557
rect 5643 3508 5644 3548
rect 5684 3508 5685 3548
rect 5643 3499 5685 3508
rect 5451 3128 5493 3137
rect 5451 3088 5452 3128
rect 5492 3088 5493 3128
rect 5451 3079 5493 3088
rect 5452 1196 5492 3079
rect 5548 2624 5588 2633
rect 5548 2036 5588 2584
rect 5548 1987 5588 1996
rect 5644 1868 5684 3499
rect 5740 2036 5780 9724
rect 5836 6992 5876 9976
rect 5932 9932 5972 9941
rect 5932 9260 5972 9892
rect 5932 9211 5972 9220
rect 5836 6404 5876 6952
rect 5836 6355 5876 6364
rect 5932 8420 5972 8429
rect 5932 8252 5972 8380
rect 5836 5480 5876 5489
rect 5836 3800 5876 5440
rect 5836 3751 5876 3760
rect 5835 3632 5877 3641
rect 5835 3592 5836 3632
rect 5876 3592 5877 3632
rect 5835 3583 5877 3592
rect 5740 1987 5780 1996
rect 5644 1819 5684 1828
rect 5452 1147 5492 1156
rect 5643 1196 5685 1205
rect 5643 1156 5644 1196
rect 5684 1156 5685 1196
rect 5643 1147 5685 1156
rect 5644 1062 5684 1147
rect 5356 559 5396 568
rect 4780 223 4820 232
rect 5836 272 5876 3583
rect 5932 2624 5972 8212
rect 6028 6488 6068 18880
rect 6124 18584 6164 21307
rect 6220 20852 6260 22399
rect 6412 21524 6452 21533
rect 6315 21440 6357 21449
rect 6315 21400 6316 21440
rect 6356 21400 6357 21440
rect 6315 21391 6357 21400
rect 6316 21306 6356 21391
rect 6220 20803 6260 20812
rect 6316 20768 6356 20777
rect 6124 14729 6164 18544
rect 6220 19340 6260 19349
rect 6123 14720 6165 14729
rect 6123 14680 6124 14720
rect 6164 14680 6165 14720
rect 6123 14671 6165 14680
rect 6220 14720 6260 19300
rect 6220 14671 6260 14680
rect 6124 14216 6164 14225
rect 6124 12284 6164 14176
rect 6219 14132 6261 14141
rect 6219 14092 6220 14132
rect 6260 14092 6261 14132
rect 6219 14083 6261 14092
rect 6220 13998 6260 14083
rect 6316 13208 6356 20728
rect 6316 13159 6356 13168
rect 6124 12235 6164 12244
rect 6316 12116 6356 12125
rect 6316 11612 6356 12076
rect 6316 11563 6356 11572
rect 6316 10352 6356 10361
rect 6124 8420 6164 8429
rect 6124 7328 6164 8380
rect 6124 7279 6164 7288
rect 6124 7076 6164 7087
rect 6124 7001 6164 7036
rect 6219 7076 6261 7085
rect 6219 7036 6220 7076
rect 6260 7036 6261 7076
rect 6219 7027 6261 7036
rect 6123 6992 6165 7001
rect 6123 6952 6124 6992
rect 6164 6952 6165 6992
rect 6123 6943 6165 6952
rect 6220 6908 6260 7027
rect 6220 6859 6260 6868
rect 6316 6824 6356 10312
rect 6123 6656 6165 6665
rect 6123 6616 6124 6656
rect 6164 6616 6165 6656
rect 6123 6607 6165 6616
rect 6028 6439 6068 6448
rect 5932 2575 5972 2584
rect 6028 4472 6068 4481
rect 5931 1952 5973 1961
rect 5931 1912 5932 1952
rect 5972 1912 5973 1952
rect 5931 1903 5973 1912
rect 5932 1818 5972 1903
rect 5931 860 5973 869
rect 5931 820 5932 860
rect 5972 820 5973 860
rect 5931 811 5973 820
rect 5932 726 5972 811
rect 6028 440 6068 4432
rect 6124 3800 6164 6607
rect 6316 5312 6356 6784
rect 6316 5263 6356 5272
rect 6124 3751 6164 3760
rect 6220 4388 6260 4397
rect 6220 692 6260 4348
rect 6315 2288 6357 2297
rect 6315 2248 6316 2288
rect 6356 2248 6357 2288
rect 6315 2239 6357 2248
rect 6316 1373 6356 2239
rect 6315 1364 6357 1373
rect 6315 1324 6316 1364
rect 6356 1324 6357 1364
rect 6315 1315 6357 1324
rect 6412 1280 6452 21484
rect 6508 20936 6548 26020
rect 6508 20887 6548 20896
rect 6700 23120 6740 28204
rect 6508 20096 6548 20105
rect 6508 19256 6548 20056
rect 6508 11360 6548 19216
rect 6603 12116 6645 12125
rect 6603 12076 6604 12116
rect 6644 12076 6645 12116
rect 6603 12067 6645 12076
rect 6604 11982 6644 12067
rect 6700 11780 6740 23080
rect 6700 11731 6740 11740
rect 6508 11320 6644 11360
rect 6508 7328 6548 7337
rect 6508 6917 6548 7288
rect 6507 6908 6549 6917
rect 6507 6868 6508 6908
rect 6548 6868 6549 6908
rect 6507 6859 6549 6868
rect 6508 6740 6548 6749
rect 6508 5480 6548 6700
rect 6508 5431 6548 5440
rect 6604 4220 6644 11320
rect 6700 9260 6740 9269
rect 6700 7580 6740 9220
rect 6700 7531 6740 7540
rect 6604 4171 6644 4180
rect 6700 6908 6740 6917
rect 6700 1289 6740 6868
rect 6412 1231 6452 1240
rect 6699 1280 6741 1289
rect 6699 1240 6700 1280
rect 6740 1240 6741 1280
rect 6699 1231 6741 1240
rect 6796 1280 6836 38107
rect 6892 34376 6932 34385
rect 6892 27749 6932 34336
rect 6988 31940 7028 40459
rect 7276 40340 7316 40349
rect 7180 39416 7220 39425
rect 7084 38744 7124 38753
rect 7084 36149 7124 38704
rect 7083 36140 7125 36149
rect 7083 36100 7084 36140
rect 7124 36100 7125 36140
rect 7083 36091 7125 36100
rect 7180 35309 7220 39376
rect 7276 39080 7316 40300
rect 7372 40172 7412 40181
rect 7372 39761 7412 40132
rect 7371 39752 7413 39761
rect 7371 39712 7372 39752
rect 7412 39712 7413 39752
rect 7371 39703 7413 39712
rect 7276 39031 7316 39040
rect 7372 38324 7412 38333
rect 7275 36728 7317 36737
rect 7275 36688 7276 36728
rect 7316 36688 7317 36728
rect 7275 36679 7317 36688
rect 7179 35300 7221 35309
rect 7179 35260 7180 35300
rect 7220 35260 7221 35300
rect 7179 35251 7221 35260
rect 6988 31891 7028 31900
rect 7180 33536 7220 35251
rect 6988 31100 7028 31109
rect 6988 28832 7028 31060
rect 6891 27740 6933 27749
rect 6891 27700 6892 27740
rect 6932 27700 6933 27740
rect 6891 27691 6933 27700
rect 6891 26900 6933 26909
rect 6891 26860 6892 26900
rect 6932 26860 6933 26900
rect 6891 26851 6933 26860
rect 6892 21188 6932 26851
rect 6988 25304 7028 28792
rect 6988 25255 7028 25264
rect 7084 30176 7124 30185
rect 7084 29672 7124 30136
rect 7084 23792 7124 29632
rect 7180 26909 7220 33496
rect 7276 34040 7316 36679
rect 7372 36065 7412 38284
rect 7660 38240 7700 38249
rect 7468 36728 7508 36737
rect 7371 36056 7413 36065
rect 7371 36016 7372 36056
rect 7412 36016 7413 36056
rect 7371 36007 7413 36016
rect 7372 35888 7412 35897
rect 7372 34376 7412 35848
rect 7372 34327 7412 34336
rect 7276 30101 7316 34000
rect 7372 30848 7412 30857
rect 7275 30092 7317 30101
rect 7275 30052 7276 30092
rect 7316 30052 7317 30092
rect 7275 30043 7317 30052
rect 7276 29840 7316 29849
rect 7276 27488 7316 29800
rect 7179 26900 7221 26909
rect 7179 26860 7180 26900
rect 7220 26860 7221 26900
rect 7179 26851 7221 26860
rect 7180 26648 7220 26657
rect 7180 25724 7220 26608
rect 7276 26480 7316 27448
rect 7276 26431 7316 26440
rect 7220 25684 7316 25724
rect 7180 25675 7220 25684
rect 7084 23743 7124 23752
rect 7179 23792 7221 23801
rect 7179 23752 7180 23792
rect 7220 23752 7221 23792
rect 7179 23743 7221 23752
rect 6987 22700 7029 22709
rect 6987 22660 6988 22700
rect 7028 22660 7029 22700
rect 6987 22651 7029 22660
rect 6988 21533 7028 22651
rect 7083 22364 7125 22373
rect 7083 22324 7084 22364
rect 7124 22324 7125 22364
rect 7083 22315 7125 22324
rect 7084 22230 7124 22315
rect 6987 21524 7029 21533
rect 6987 21484 6988 21524
rect 7028 21484 7029 21524
rect 6987 21475 7029 21484
rect 6892 21139 6932 21148
rect 6892 16064 6932 16073
rect 6892 2708 6932 16024
rect 6892 2659 6932 2668
rect 6891 1868 6933 1877
rect 6891 1828 6892 1868
rect 6932 1828 6933 1868
rect 6891 1819 6933 1828
rect 6796 1231 6836 1240
rect 6220 643 6260 652
rect 6028 391 6068 400
rect 6603 356 6645 365
rect 6603 316 6604 356
rect 6644 316 6645 356
rect 6603 307 6645 316
rect 6892 356 6932 1819
rect 6988 1280 7028 21475
rect 7084 20936 7124 20945
rect 7084 15812 7124 20896
rect 7084 15763 7124 15772
rect 7084 12536 7124 12545
rect 7084 11360 7124 12496
rect 7084 11311 7124 11320
rect 7084 9680 7124 9689
rect 7084 6236 7124 9640
rect 7084 6187 7124 6196
rect 7083 3380 7125 3389
rect 7083 3340 7084 3380
rect 7124 3340 7125 3380
rect 7083 3331 7125 3340
rect 7084 3246 7124 3331
rect 6988 1231 7028 1240
rect 7180 1280 7220 23743
rect 7276 20768 7316 25684
rect 7372 21608 7412 30808
rect 7468 22709 7508 36688
rect 7564 36056 7604 36065
rect 7564 33545 7604 36016
rect 7660 34376 7700 38200
rect 7563 33536 7605 33545
rect 7563 33496 7564 33536
rect 7604 33496 7605 33536
rect 7563 33487 7605 33496
rect 7563 32948 7605 32957
rect 7563 32908 7564 32948
rect 7604 32908 7605 32948
rect 7563 32899 7605 32908
rect 7564 32864 7604 32899
rect 7564 32813 7604 32824
rect 7467 22700 7509 22709
rect 7467 22660 7468 22700
rect 7508 22660 7509 22700
rect 7467 22651 7509 22660
rect 7660 22289 7700 34336
rect 7756 30344 7796 30353
rect 7756 27488 7796 30304
rect 7756 27439 7796 27448
rect 7756 26396 7796 26405
rect 7659 22280 7701 22289
rect 7659 22240 7660 22280
rect 7700 22240 7701 22280
rect 7659 22231 7701 22240
rect 7660 21869 7700 22231
rect 7659 21860 7701 21869
rect 7659 21820 7660 21860
rect 7700 21820 7701 21860
rect 7659 21811 7701 21820
rect 7659 21692 7701 21701
rect 7756 21692 7796 26356
rect 7659 21652 7660 21692
rect 7700 21652 7796 21692
rect 7659 21643 7701 21652
rect 7372 21559 7412 21568
rect 7276 20719 7316 20728
rect 7372 21440 7412 21449
rect 7276 11612 7316 11621
rect 7276 6329 7316 11572
rect 7275 6320 7317 6329
rect 7275 6280 7276 6320
rect 7316 6280 7317 6320
rect 7275 6271 7317 6280
rect 7180 1231 7220 1240
rect 7372 944 7412 21400
rect 7563 17660 7605 17669
rect 7563 17620 7564 17660
rect 7604 17620 7605 17660
rect 7563 17611 7605 17620
rect 7564 17526 7604 17611
rect 7468 16064 7508 16073
rect 7468 13544 7508 16024
rect 7660 15896 7700 21643
rect 7468 13495 7508 13504
rect 7564 15856 7700 15896
rect 7756 21356 7796 21365
rect 7564 12629 7604 15856
rect 7659 15728 7701 15737
rect 7659 15688 7660 15728
rect 7700 15688 7701 15728
rect 7659 15679 7701 15688
rect 7563 12620 7605 12629
rect 7563 12580 7564 12620
rect 7604 12580 7605 12620
rect 7563 12571 7605 12580
rect 7467 11696 7509 11705
rect 7467 11656 7468 11696
rect 7508 11656 7509 11696
rect 7467 11647 7509 11656
rect 7468 10016 7508 11647
rect 7468 9967 7508 9976
rect 7564 10184 7604 10193
rect 7564 9428 7604 10144
rect 7564 9379 7604 9388
rect 7564 8336 7604 8345
rect 7468 7580 7508 7589
rect 7468 5984 7508 7540
rect 7564 6320 7604 8296
rect 7660 6908 7700 15679
rect 7660 6859 7700 6868
rect 7659 6740 7701 6749
rect 7659 6700 7660 6740
rect 7700 6700 7701 6740
rect 7659 6691 7701 6700
rect 7564 6271 7604 6280
rect 7468 5935 7508 5944
rect 7564 4724 7604 4733
rect 7564 3725 7604 4684
rect 7563 3716 7605 3725
rect 7563 3676 7564 3716
rect 7604 3676 7605 3716
rect 7563 3667 7605 3676
rect 7660 3380 7700 6691
rect 7468 2960 7508 2969
rect 7468 2717 7508 2920
rect 7467 2708 7509 2717
rect 7467 2668 7468 2708
rect 7508 2668 7509 2708
rect 7467 2659 7509 2668
rect 7660 2708 7700 3340
rect 7660 2659 7700 2668
rect 7372 895 7412 904
rect 7756 944 7796 21316
rect 7852 11948 7892 41812
rect 9388 41432 9428 41441
rect 8235 40340 8277 40349
rect 8235 40300 8236 40340
rect 8276 40300 8277 40340
rect 8235 40291 8277 40300
rect 8044 38996 8084 39005
rect 8044 38324 8084 38956
rect 8236 38996 8276 40291
rect 8236 38744 8276 38956
rect 8236 38695 8276 38704
rect 8332 40088 8372 40097
rect 8332 38576 8372 40048
rect 8619 38912 8661 38921
rect 8619 38872 8620 38912
rect 8660 38872 8661 38912
rect 8619 38863 8661 38872
rect 8620 38778 8660 38863
rect 7947 37736 7989 37745
rect 7947 37696 7948 37736
rect 7988 37696 7989 37736
rect 7947 37687 7989 37696
rect 7948 32621 7988 37687
rect 8044 36728 8084 38284
rect 8236 38536 8372 38576
rect 8716 38576 8756 38585
rect 8044 36679 8084 36688
rect 8140 36896 8180 36905
rect 8140 36560 8180 36856
rect 8236 36653 8276 38536
rect 8716 38240 8756 38536
rect 8716 38191 8756 38200
rect 8715 38072 8757 38081
rect 8715 38032 8716 38072
rect 8756 38032 8757 38072
rect 8715 38023 8757 38032
rect 8812 38072 8852 38081
rect 8716 37484 8756 38023
rect 8427 37148 8469 37157
rect 8427 37108 8428 37148
rect 8468 37108 8469 37148
rect 8427 37099 8469 37108
rect 8235 36644 8277 36653
rect 8235 36604 8236 36644
rect 8276 36604 8277 36644
rect 8235 36595 8277 36604
rect 8044 36520 8180 36560
rect 8331 36560 8373 36569
rect 8331 36520 8332 36560
rect 8372 36520 8373 36560
rect 7947 32612 7989 32621
rect 7947 32572 7948 32612
rect 7988 32572 7989 32612
rect 7947 32563 7989 32572
rect 7947 28664 7989 28673
rect 7947 28624 7948 28664
rect 7988 28624 7989 28664
rect 7947 28615 7989 28624
rect 7948 28530 7988 28615
rect 7852 11528 7892 11908
rect 7852 11479 7892 11488
rect 7948 27152 7988 27161
rect 7852 8168 7892 8177
rect 7852 6665 7892 8128
rect 7851 6656 7893 6665
rect 7851 6616 7852 6656
rect 7892 6616 7893 6656
rect 7851 6607 7893 6616
rect 7852 6488 7892 6497
rect 7852 4136 7892 6448
rect 7852 4087 7892 4096
rect 7852 3716 7892 3725
rect 7852 2465 7892 3676
rect 7851 2456 7893 2465
rect 7851 2416 7852 2456
rect 7892 2416 7893 2456
rect 7851 2407 7893 2416
rect 7756 895 7796 904
rect 7948 692 7988 27112
rect 8044 1028 8084 36520
rect 8331 36511 8373 36520
rect 8236 36224 8276 36233
rect 8236 35636 8276 36184
rect 8332 36140 8372 36511
rect 8332 36091 8372 36100
rect 8139 32612 8181 32621
rect 8139 32572 8140 32612
rect 8180 32572 8181 32612
rect 8139 32563 8181 32572
rect 8140 1280 8180 32563
rect 8236 25220 8276 35596
rect 8428 32444 8468 37099
rect 8620 36728 8660 36737
rect 8523 36644 8565 36653
rect 8523 36604 8524 36644
rect 8564 36604 8565 36644
rect 8523 36595 8565 36604
rect 8428 32395 8468 32404
rect 8236 25171 8276 25180
rect 8332 32192 8372 32201
rect 8235 22112 8277 22121
rect 8235 22072 8236 22112
rect 8276 22072 8277 22112
rect 8235 22063 8277 22072
rect 8236 21978 8276 22063
rect 8235 21860 8277 21869
rect 8235 21820 8236 21860
rect 8276 21820 8277 21860
rect 8235 21811 8277 21820
rect 8236 15737 8276 21811
rect 8332 19172 8372 32152
rect 8428 29504 8468 29513
rect 8428 28664 8468 29464
rect 8428 28615 8468 28624
rect 8428 26144 8468 26153
rect 8428 24548 8468 26104
rect 8428 24499 8468 24508
rect 8332 19123 8372 19132
rect 8428 22112 8468 22121
rect 8235 15728 8277 15737
rect 8235 15688 8236 15728
rect 8276 15688 8277 15728
rect 8235 15679 8277 15688
rect 8332 13292 8372 13301
rect 8236 11864 8276 11873
rect 8236 4892 8276 11824
rect 8236 4843 8276 4852
rect 8140 1231 8180 1240
rect 8332 1280 8372 13252
rect 8428 3473 8468 22072
rect 8524 21440 8564 36595
rect 8620 26396 8660 36688
rect 8716 36569 8756 37444
rect 8715 36560 8757 36569
rect 8715 36520 8716 36560
rect 8756 36520 8757 36560
rect 8715 36511 8757 36520
rect 8715 33788 8757 33797
rect 8715 33748 8716 33788
rect 8756 33748 8757 33788
rect 8715 33739 8757 33748
rect 8716 33654 8756 33739
rect 8620 26347 8660 26356
rect 8716 32444 8756 32453
rect 8619 26228 8661 26237
rect 8619 26188 8620 26228
rect 8660 26188 8661 26228
rect 8619 26179 8661 26188
rect 8620 26144 8660 26179
rect 8620 26093 8660 26104
rect 8620 25052 8660 25061
rect 8620 23456 8660 25012
rect 8620 23407 8660 23416
rect 8716 23120 8756 32404
rect 8620 23080 8756 23120
rect 8620 22112 8660 23080
rect 8715 22952 8757 22961
rect 8715 22912 8716 22952
rect 8756 22912 8757 22952
rect 8715 22903 8757 22912
rect 8716 22818 8756 22903
rect 8620 22063 8660 22072
rect 8715 21524 8757 21533
rect 8715 21484 8716 21524
rect 8756 21484 8757 21524
rect 8715 21475 8757 21484
rect 8524 21391 8564 21400
rect 8716 21390 8756 21475
rect 8812 21356 8852 38032
rect 8907 37736 8949 37745
rect 8907 37696 8908 37736
rect 8948 37696 8949 37736
rect 8907 37687 8949 37696
rect 8908 37316 8948 37687
rect 8908 37267 8948 37276
rect 9388 36821 9428 41392
rect 10060 40172 10100 40181
rect 9868 39500 9908 39509
rect 9772 38324 9812 38333
rect 9484 37820 9524 37829
rect 9484 37400 9524 37780
rect 9772 37652 9812 38284
rect 9772 37603 9812 37612
rect 9484 37351 9524 37360
rect 9387 36812 9429 36821
rect 9387 36772 9388 36812
rect 9428 36772 9429 36812
rect 9387 36763 9429 36772
rect 9099 36728 9141 36737
rect 9099 36688 9100 36728
rect 9140 36688 9141 36728
rect 9099 36679 9141 36688
rect 9100 36594 9140 36679
rect 9292 36560 9332 36569
rect 8812 21307 8852 21316
rect 8908 34460 8948 34469
rect 8908 17996 8948 34420
rect 9195 34376 9237 34385
rect 9195 34336 9196 34376
rect 9236 34336 9237 34376
rect 9195 34327 9237 34336
rect 9196 34049 9236 34327
rect 9195 34040 9237 34049
rect 9195 34000 9196 34040
rect 9236 34000 9237 34040
rect 9195 33991 9237 34000
rect 9195 33032 9237 33041
rect 9195 32992 9196 33032
rect 9236 32992 9237 33032
rect 9195 32983 9237 32992
rect 9196 32864 9236 32983
rect 9196 32815 9236 32824
rect 9292 32117 9332 36520
rect 9388 36317 9428 36763
rect 9771 36560 9813 36569
rect 9771 36520 9772 36560
rect 9812 36520 9813 36560
rect 9771 36511 9813 36520
rect 9387 36308 9429 36317
rect 9387 36268 9388 36308
rect 9428 36268 9429 36308
rect 9387 36259 9429 36268
rect 9675 35216 9717 35225
rect 9675 35176 9676 35216
rect 9716 35176 9717 35216
rect 9675 35167 9717 35176
rect 9579 32696 9621 32705
rect 9579 32656 9580 32696
rect 9620 32656 9621 32696
rect 9579 32647 9621 32656
rect 9580 32192 9620 32647
rect 9580 32143 9620 32152
rect 9291 32108 9333 32117
rect 9291 32068 9292 32108
rect 9332 32068 9333 32108
rect 9291 32059 9333 32068
rect 9100 31856 9140 31865
rect 9004 29924 9044 29933
rect 9004 27572 9044 29884
rect 9004 27523 9044 27532
rect 9100 23120 9140 31816
rect 9292 31520 9332 31529
rect 9292 26816 9332 31480
rect 9580 30176 9620 30185
rect 9484 28328 9524 28337
rect 9484 27992 9524 28288
rect 9292 26767 9332 26776
rect 9388 27404 9428 27413
rect 8908 17947 8948 17956
rect 9004 20096 9044 20105
rect 8812 16400 8852 16409
rect 8620 12620 8660 12629
rect 8524 10352 8564 10361
rect 8524 4472 8564 10312
rect 8524 4423 8564 4432
rect 8427 3464 8469 3473
rect 8427 3424 8428 3464
rect 8468 3424 8469 3464
rect 8427 3415 8469 3424
rect 8332 1231 8372 1240
rect 8523 1280 8565 1289
rect 8523 1240 8524 1280
rect 8564 1240 8565 1280
rect 8523 1231 8565 1240
rect 8524 1146 8564 1231
rect 8620 1112 8660 12580
rect 8716 9932 8756 9941
rect 8812 9932 8852 16360
rect 8907 16064 8949 16073
rect 8907 16024 8908 16064
rect 8948 16024 8949 16064
rect 8907 16015 8949 16024
rect 8908 15930 8948 16015
rect 8756 9892 8852 9932
rect 8908 14636 8948 14645
rect 8716 9883 8756 9892
rect 8716 9764 8756 9773
rect 8716 8429 8756 9724
rect 8811 9764 8853 9773
rect 8811 9724 8812 9764
rect 8852 9724 8853 9764
rect 8811 9715 8853 9724
rect 8812 8681 8852 9715
rect 8811 8672 8853 8681
rect 8811 8632 8812 8672
rect 8852 8632 8853 8672
rect 8811 8623 8853 8632
rect 8811 8504 8853 8513
rect 8811 8464 8812 8504
rect 8852 8464 8853 8504
rect 8811 8455 8853 8464
rect 8715 8420 8757 8429
rect 8715 8380 8716 8420
rect 8756 8380 8757 8420
rect 8715 8371 8757 8380
rect 8715 7916 8757 7925
rect 8715 7876 8716 7916
rect 8756 7876 8757 7916
rect 8715 7867 8757 7876
rect 8716 7782 8756 7867
rect 8812 7748 8852 8455
rect 8715 7160 8757 7169
rect 8715 7120 8716 7160
rect 8756 7120 8757 7160
rect 8715 7111 8757 7120
rect 8716 7026 8756 7111
rect 8716 6488 8756 6497
rect 8716 5228 8756 6448
rect 8716 5179 8756 5188
rect 8812 5060 8852 7708
rect 8908 7496 8948 14596
rect 8908 7447 8948 7456
rect 8812 5011 8852 5020
rect 8811 3800 8853 3809
rect 8811 3760 8812 3800
rect 8852 3760 8853 3800
rect 8811 3751 8853 3760
rect 8812 2204 8852 3751
rect 9004 3557 9044 20056
rect 9100 16232 9140 23080
rect 9292 21440 9332 21449
rect 9292 21272 9332 21400
rect 9292 19004 9332 21232
rect 9388 20852 9428 27364
rect 9388 20803 9428 20812
rect 9484 19340 9524 27952
rect 9580 27572 9620 30136
rect 9580 27523 9620 27532
rect 9676 28412 9716 35167
rect 9676 27404 9716 28372
rect 9772 27740 9812 36511
rect 9772 27691 9812 27700
rect 9676 27355 9716 27364
rect 9676 26816 9716 26825
rect 9580 26648 9620 26657
rect 9580 25733 9620 26608
rect 9579 25724 9621 25733
rect 9579 25684 9580 25724
rect 9620 25684 9621 25724
rect 9579 25675 9621 25684
rect 9484 19291 9524 19300
rect 9580 23120 9620 23129
rect 9292 18955 9332 18964
rect 9484 17660 9524 17669
rect 9100 16192 9428 16232
rect 9292 16064 9332 16073
rect 9196 15896 9236 15905
rect 9100 15644 9140 15653
rect 9100 14477 9140 15604
rect 9196 15560 9236 15856
rect 9099 14468 9141 14477
rect 9099 14428 9100 14468
rect 9140 14428 9141 14468
rect 9099 14419 9141 14428
rect 9100 14300 9140 14309
rect 9100 9512 9140 14260
rect 9196 13964 9236 15520
rect 9196 13915 9236 13924
rect 9100 9260 9140 9472
rect 9100 9211 9140 9220
rect 9196 11948 9236 11957
rect 9196 8840 9236 11908
rect 9100 8800 9236 8840
rect 9100 8681 9140 8800
rect 9099 8672 9141 8681
rect 9099 8632 9100 8672
rect 9140 8632 9141 8672
rect 9099 8623 9141 8632
rect 9195 8420 9237 8429
rect 9195 8380 9196 8420
rect 9236 8380 9237 8420
rect 9195 8371 9237 8380
rect 9003 3548 9045 3557
rect 9003 3508 9004 3548
rect 9044 3508 9045 3548
rect 9003 3499 9045 3508
rect 9100 2960 9140 2969
rect 9100 2540 9140 2920
rect 9100 2491 9140 2500
rect 8812 2155 8852 2164
rect 9196 1952 9236 8371
rect 9292 3716 9332 16024
rect 9388 9764 9428 16192
rect 9484 14636 9524 17620
rect 9484 14587 9524 14596
rect 9483 14468 9525 14477
rect 9483 14428 9484 14468
rect 9524 14428 9525 14468
rect 9483 14419 9525 14428
rect 9484 11360 9524 14419
rect 9484 11311 9524 11320
rect 9580 11024 9620 23080
rect 9676 20012 9716 26776
rect 9772 24884 9812 24893
rect 9772 23624 9812 24844
rect 9772 23575 9812 23584
rect 9676 19256 9716 19972
rect 9676 19207 9716 19216
rect 9772 17408 9812 17417
rect 9772 15896 9812 17368
rect 9772 15847 9812 15856
rect 9772 13208 9812 13217
rect 9580 10975 9620 10984
rect 9676 11696 9716 11705
rect 9676 10772 9716 11656
rect 9676 10723 9716 10732
rect 9484 10604 9524 10613
rect 9484 9773 9524 10564
rect 9388 8840 9428 9724
rect 9483 9764 9525 9773
rect 9483 9724 9484 9764
rect 9524 9724 9525 9764
rect 9483 9715 9525 9724
rect 9388 8800 9524 8840
rect 9387 8588 9429 8597
rect 9387 8548 9388 8588
rect 9428 8548 9429 8588
rect 9387 8539 9429 8548
rect 9388 7580 9428 8539
rect 9484 8513 9524 8800
rect 9579 8672 9621 8681
rect 9579 8632 9580 8672
rect 9620 8632 9621 8672
rect 9579 8623 9621 8632
rect 9483 8504 9525 8513
rect 9483 8464 9484 8504
rect 9524 8464 9525 8504
rect 9483 8455 9525 8464
rect 9483 8336 9525 8345
rect 9483 8296 9484 8336
rect 9524 8296 9525 8336
rect 9483 8287 9525 8296
rect 9484 8168 9524 8287
rect 9484 8119 9524 8128
rect 9388 7531 9428 7540
rect 9484 7916 9524 7925
rect 9292 3667 9332 3676
rect 9388 6992 9428 7001
rect 9388 4976 9428 6952
rect 9484 6656 9524 7876
rect 9484 6607 9524 6616
rect 9580 5060 9620 8623
rect 9676 8168 9716 8177
rect 9676 7001 9716 8128
rect 9675 6992 9717 7001
rect 9675 6952 9676 6992
rect 9716 6952 9717 6992
rect 9675 6943 9717 6952
rect 9676 5144 9716 6943
rect 9676 5095 9716 5104
rect 9580 5011 9620 5020
rect 9388 2708 9428 4936
rect 9388 2659 9428 2668
rect 9580 3380 9620 3389
rect 9291 2120 9333 2129
rect 9291 2080 9292 2120
rect 9332 2080 9333 2120
rect 9291 2071 9333 2080
rect 9292 1986 9332 2071
rect 9196 1903 9236 1912
rect 8620 1063 8660 1072
rect 9580 1112 9620 3340
rect 9580 1063 9620 1072
rect 8044 979 8084 988
rect 7948 643 7988 652
rect 6892 307 6932 316
rect 9772 524 9812 13168
rect 9868 3809 9908 39460
rect 10060 38576 10100 40132
rect 10060 38527 10100 38536
rect 9964 38156 10004 38165
rect 9964 35720 10004 38116
rect 9964 35671 10004 35680
rect 10156 35972 10196 42148
rect 10252 38996 10292 42316
rect 15052 42272 15092 42281
rect 12172 41684 12212 41693
rect 10732 40508 10772 40517
rect 10252 38947 10292 38956
rect 10444 40424 10484 40433
rect 10347 38912 10389 38921
rect 10347 38872 10348 38912
rect 10388 38872 10389 38912
rect 10347 38863 10389 38872
rect 10059 34208 10101 34217
rect 10059 34168 10060 34208
rect 10100 34168 10101 34208
rect 10059 34159 10101 34168
rect 10060 34074 10100 34159
rect 9964 33704 10004 33713
rect 9964 31772 10004 33664
rect 10060 32612 10100 32621
rect 10060 31856 10100 32572
rect 10060 31807 10100 31816
rect 9964 31723 10004 31732
rect 9964 31268 10004 31277
rect 9964 29261 10004 31228
rect 10059 29672 10101 29681
rect 10059 29632 10060 29672
rect 10100 29632 10101 29672
rect 10059 29623 10101 29632
rect 10060 29538 10100 29623
rect 9963 29252 10005 29261
rect 9963 29212 9964 29252
rect 10004 29212 10005 29252
rect 9963 29203 10005 29212
rect 9964 29000 10004 29203
rect 9964 28951 10004 28960
rect 9963 26816 10005 26825
rect 9963 26776 9964 26816
rect 10004 26776 10005 26816
rect 9963 26767 10005 26776
rect 9964 26682 10004 26767
rect 10060 26312 10100 26321
rect 10060 25724 10100 26272
rect 10060 23204 10100 25684
rect 10060 23155 10100 23164
rect 9964 14888 10004 14897
rect 9964 13217 10004 14848
rect 10156 13880 10196 35932
rect 10252 38744 10292 38753
rect 10252 26228 10292 38704
rect 10252 26179 10292 26188
rect 10251 24548 10293 24557
rect 10251 24508 10252 24548
rect 10292 24508 10293 24548
rect 10251 24499 10293 24508
rect 10156 13831 10196 13840
rect 9963 13208 10005 13217
rect 9963 13168 9964 13208
rect 10004 13168 10005 13208
rect 9963 13159 10005 13168
rect 10060 13124 10100 13133
rect 9964 12872 10004 12881
rect 9964 10184 10004 12832
rect 10060 11360 10100 13084
rect 10252 12788 10292 24499
rect 10348 21272 10388 38863
rect 10444 26489 10484 40384
rect 10732 39257 10772 40468
rect 11596 40340 11636 40349
rect 10924 40088 10964 40097
rect 10636 39248 10676 39257
rect 10636 33200 10676 39208
rect 10731 39248 10773 39257
rect 10731 39208 10732 39248
rect 10772 39208 10773 39248
rect 10731 39199 10773 39208
rect 10636 33151 10676 33160
rect 10539 32024 10581 32033
rect 10539 31984 10540 32024
rect 10580 31984 10581 32024
rect 10539 31975 10581 31984
rect 10443 26480 10485 26489
rect 10443 26440 10444 26480
rect 10484 26440 10485 26480
rect 10443 26431 10485 26440
rect 10348 21223 10388 21232
rect 10444 25136 10484 25145
rect 10444 20096 10484 25096
rect 10540 24557 10580 31975
rect 10636 29840 10676 29849
rect 10636 28832 10676 29800
rect 10636 28783 10676 28792
rect 10539 24548 10581 24557
rect 10539 24508 10540 24548
rect 10580 24508 10581 24548
rect 10539 24499 10581 24508
rect 10636 24212 10676 24221
rect 10540 23960 10580 23969
rect 10540 23792 10580 23920
rect 10540 23743 10580 23752
rect 10540 23456 10580 23465
rect 10540 22784 10580 23416
rect 10540 22735 10580 22744
rect 10636 22280 10676 24172
rect 10540 22240 10676 22280
rect 10540 20768 10580 22240
rect 10635 22112 10677 22121
rect 10635 22072 10636 22112
rect 10676 22072 10677 22112
rect 10635 22063 10677 22072
rect 10540 20719 10580 20728
rect 10636 20180 10676 22063
rect 10444 20047 10484 20056
rect 10540 20140 10676 20180
rect 10444 18668 10484 18677
rect 10156 12748 10292 12788
rect 10348 16736 10388 16745
rect 10156 12116 10196 12748
rect 10156 12067 10196 12076
rect 10060 11320 10196 11360
rect 9964 10135 10004 10144
rect 9963 9932 10005 9941
rect 9963 9892 9964 9932
rect 10004 9892 10005 9932
rect 9963 9883 10005 9892
rect 9867 3800 9909 3809
rect 9867 3760 9868 3800
rect 9908 3760 9909 3800
rect 9867 3751 9909 3760
rect 9964 3632 10004 9883
rect 10060 9176 10100 9185
rect 10060 6656 10100 9136
rect 10060 6607 10100 6616
rect 10060 6404 10100 6413
rect 10060 6152 10100 6364
rect 10060 6103 10100 6112
rect 10156 4649 10196 11320
rect 10252 10856 10292 10865
rect 10252 6320 10292 10816
rect 10348 8840 10388 16696
rect 10444 14720 10484 18628
rect 10444 14671 10484 14680
rect 10443 13460 10485 13469
rect 10443 13420 10444 13460
rect 10484 13420 10485 13460
rect 10443 13411 10485 13420
rect 10444 13326 10484 13411
rect 10443 13208 10485 13217
rect 10443 13168 10444 13208
rect 10484 13168 10485 13208
rect 10443 13159 10485 13168
rect 10444 11780 10484 13159
rect 10444 11731 10484 11740
rect 10444 11276 10484 11285
rect 10444 9176 10484 11236
rect 10444 9127 10484 9136
rect 10348 8791 10388 8800
rect 10252 6271 10292 6280
rect 10348 8000 10388 8009
rect 10348 6488 10388 7960
rect 10252 4976 10292 4985
rect 10155 4640 10197 4649
rect 10155 4600 10156 4640
rect 10196 4600 10197 4640
rect 10155 4591 10197 4600
rect 10252 4556 10292 4936
rect 10348 4724 10388 6448
rect 10348 4675 10388 4684
rect 10444 5564 10484 5573
rect 10252 4516 10388 4556
rect 10251 4304 10293 4313
rect 10251 4264 10252 4304
rect 10292 4264 10293 4304
rect 10251 4255 10293 4264
rect 10252 4170 10292 4255
rect 9868 3592 10004 3632
rect 9868 2288 9908 3592
rect 9868 2239 9908 2248
rect 9964 2540 10004 2549
rect 9964 1532 10004 2500
rect 10348 2540 10388 4516
rect 10444 3884 10484 5524
rect 10444 3835 10484 3844
rect 10540 2708 10580 20140
rect 10636 19340 10676 19349
rect 10636 18332 10676 19300
rect 10636 18283 10676 18292
rect 10636 16652 10676 16661
rect 10636 9008 10676 16612
rect 10636 8959 10676 8968
rect 10636 5144 10676 5153
rect 10636 4313 10676 5104
rect 10635 4304 10677 4313
rect 10635 4264 10636 4304
rect 10676 4264 10677 4304
rect 10635 4255 10677 4264
rect 10636 3884 10676 4255
rect 10636 3835 10676 3844
rect 10635 3716 10677 3725
rect 10635 3676 10636 3716
rect 10676 3676 10677 3716
rect 10635 3667 10677 3676
rect 10540 2659 10580 2668
rect 10348 2491 10388 2500
rect 10636 2540 10676 3667
rect 10636 2491 10676 2500
rect 10732 2381 10772 39199
rect 10827 36560 10869 36569
rect 10827 36520 10828 36560
rect 10868 36520 10869 36560
rect 10827 36511 10869 36520
rect 10828 36426 10868 36511
rect 10924 36476 10964 40048
rect 11596 39836 11636 40300
rect 11596 39787 11636 39796
rect 11500 39332 11540 39341
rect 11116 39248 11156 39257
rect 10924 36427 10964 36436
rect 11020 38996 11060 39005
rect 10923 32780 10965 32789
rect 10923 32740 10924 32780
rect 10964 32740 10965 32780
rect 10923 32731 10965 32740
rect 10924 32646 10964 32731
rect 10924 32108 10964 32117
rect 10827 29000 10869 29009
rect 10827 28960 10828 29000
rect 10868 28960 10869 29000
rect 10827 28951 10869 28960
rect 10828 28866 10868 28951
rect 10828 24800 10868 24809
rect 10828 23960 10868 24760
rect 10828 23036 10868 23920
rect 10828 22987 10868 22996
rect 10828 20768 10868 20777
rect 10828 19256 10868 20728
rect 10924 20600 10964 32068
rect 10924 19592 10964 20560
rect 10924 19543 10964 19552
rect 10828 19216 10964 19256
rect 10828 19088 10868 19097
rect 10828 12125 10868 19048
rect 10924 18920 10964 19216
rect 10924 18871 10964 18880
rect 10924 14720 10964 14729
rect 10827 12116 10869 12125
rect 10827 12076 10828 12116
rect 10868 12076 10869 12116
rect 10827 12067 10869 12076
rect 10924 7916 10964 14680
rect 10924 7867 10964 7876
rect 11020 7580 11060 38956
rect 11116 37820 11156 39208
rect 11212 38996 11252 39005
rect 11212 38660 11252 38956
rect 11212 38611 11252 38620
rect 11500 38072 11540 39292
rect 11500 38023 11540 38032
rect 11116 37771 11156 37780
rect 11308 37736 11348 37745
rect 11308 37568 11348 37696
rect 11308 37519 11348 37528
rect 11692 37400 11732 37409
rect 11212 35216 11252 35227
rect 11212 35141 11252 35176
rect 11692 35216 11732 37360
rect 11211 35132 11253 35141
rect 11211 35092 11212 35132
rect 11252 35092 11253 35132
rect 11211 35083 11253 35092
rect 11116 33956 11156 33965
rect 11116 30764 11156 33916
rect 11116 29672 11156 30724
rect 11116 29623 11156 29632
rect 11308 33452 11348 33461
rect 11115 29252 11157 29261
rect 11115 29212 11116 29252
rect 11156 29212 11157 29252
rect 11115 29203 11157 29212
rect 11116 26312 11156 29203
rect 11116 26263 11156 26272
rect 11212 29168 11252 29177
rect 11115 20852 11157 20861
rect 11115 20812 11116 20852
rect 11156 20812 11157 20852
rect 11115 20803 11157 20812
rect 11116 9344 11156 20803
rect 11212 20768 11252 29128
rect 11308 28673 11348 33412
rect 11500 30596 11540 30605
rect 11307 28664 11349 28673
rect 11307 28624 11308 28664
rect 11348 28624 11349 28664
rect 11307 28615 11349 28624
rect 11403 26480 11445 26489
rect 11403 26440 11404 26480
rect 11444 26440 11445 26480
rect 11403 26431 11445 26440
rect 11212 20719 11252 20728
rect 11308 22364 11348 22373
rect 11308 21524 11348 22324
rect 11308 20180 11348 21484
rect 11308 20131 11348 20140
rect 11212 14384 11252 14393
rect 11212 9848 11252 14344
rect 11308 14216 11348 14225
rect 11308 12293 11348 14176
rect 11404 13208 11444 26431
rect 11404 13159 11444 13168
rect 11404 13040 11444 13049
rect 11307 12284 11349 12293
rect 11307 12244 11308 12284
rect 11348 12244 11349 12284
rect 11307 12235 11349 12244
rect 11307 12116 11349 12125
rect 11307 12076 11308 12116
rect 11348 12076 11349 12116
rect 11307 12067 11349 12076
rect 11212 9799 11252 9808
rect 11116 9295 11156 9304
rect 11212 9512 11252 9521
rect 11020 7531 11060 7540
rect 10828 5228 10868 5237
rect 10828 2792 10868 5188
rect 11116 5228 11156 5237
rect 11116 3548 11156 5188
rect 11116 3389 11156 3508
rect 11115 3380 11157 3389
rect 11115 3340 11116 3380
rect 11156 3340 11157 3380
rect 11115 3331 11157 3340
rect 10828 2540 10868 2752
rect 10828 2491 10868 2500
rect 10731 2372 10773 2381
rect 10731 2332 10732 2372
rect 10772 2332 10773 2372
rect 11212 2372 11252 9472
rect 11308 3800 11348 12067
rect 11404 11957 11444 13000
rect 11403 11948 11445 11957
rect 11403 11908 11404 11948
rect 11444 11908 11445 11948
rect 11403 11899 11445 11908
rect 11403 11780 11445 11789
rect 11403 11740 11404 11780
rect 11444 11740 11445 11780
rect 11403 11731 11445 11740
rect 11404 5909 11444 11731
rect 11500 11612 11540 30556
rect 11596 25388 11636 25397
rect 11596 25229 11636 25348
rect 11595 25220 11637 25229
rect 11595 25180 11596 25220
rect 11636 25180 11637 25220
rect 11595 25171 11637 25180
rect 11692 20180 11732 35176
rect 11884 36560 11924 36569
rect 11788 33704 11828 33713
rect 11788 32696 11828 33664
rect 11788 32647 11828 32656
rect 11788 31100 11828 31109
rect 11788 23708 11828 31060
rect 11884 26312 11924 36520
rect 12076 31604 12116 31613
rect 12076 31016 12116 31564
rect 12076 30967 12116 30976
rect 11884 26263 11924 26272
rect 11980 26732 12020 26741
rect 11980 26144 12020 26692
rect 11788 23659 11828 23668
rect 11884 26104 12020 26144
rect 11884 24716 11924 26104
rect 12172 25136 12212 41644
rect 12556 41600 12596 41609
rect 12364 41264 12404 41273
rect 12364 37484 12404 41224
rect 12364 37435 12404 37444
rect 12460 40004 12500 40013
rect 12364 34376 12404 34385
rect 12364 32780 12404 34336
rect 12268 32276 12308 32285
rect 12268 31529 12308 32236
rect 12267 31520 12309 31529
rect 12267 31480 12268 31520
rect 12308 31480 12309 31520
rect 12267 31471 12309 31480
rect 12172 25087 12212 25096
rect 11788 23288 11828 23297
rect 11788 22028 11828 23248
rect 11788 21979 11828 21988
rect 11884 21440 11924 24676
rect 11884 21391 11924 21400
rect 11980 25052 12020 25061
rect 11596 20140 11732 20180
rect 11596 11789 11636 20140
rect 11692 16652 11732 16661
rect 11692 16316 11732 16612
rect 11692 16267 11732 16276
rect 11692 16064 11732 16073
rect 11692 13628 11732 16024
rect 11884 15560 11924 15569
rect 11787 13880 11829 13889
rect 11787 13840 11788 13880
rect 11828 13840 11829 13880
rect 11787 13831 11829 13840
rect 11788 13746 11828 13831
rect 11692 13588 11828 13628
rect 11595 11780 11637 11789
rect 11595 11740 11596 11780
rect 11636 11740 11637 11780
rect 11595 11731 11637 11740
rect 11500 11572 11636 11612
rect 11500 11108 11540 11117
rect 11403 5900 11445 5909
rect 11403 5860 11404 5900
rect 11444 5860 11445 5900
rect 11403 5851 11445 5860
rect 11404 5816 11444 5851
rect 11404 5736 11444 5776
rect 11308 3751 11348 3760
rect 11212 2332 11348 2372
rect 10731 2323 10773 2332
rect 10156 2288 10196 2297
rect 9964 1483 10004 1492
rect 10060 1952 10100 1961
rect 5836 223 5876 232
rect 6604 222 6644 307
rect 267 188 309 197
rect 267 148 268 188
rect 308 148 309 188
rect 267 139 309 148
rect 5259 188 5301 197
rect 5259 148 5260 188
rect 5300 148 5301 188
rect 5259 139 5301 148
rect 268 104 308 139
rect 268 53 308 64
rect 5260 54 5300 139
rect 6028 113 6068 198
rect 9772 188 9812 484
rect 9772 139 9812 148
rect 10060 113 10100 1912
rect 10156 869 10196 2248
rect 11212 2204 11252 2213
rect 11212 1532 11252 2164
rect 11212 1483 11252 1492
rect 10924 1196 10964 1205
rect 10155 860 10197 869
rect 10155 820 10156 860
rect 10196 820 10197 860
rect 10155 811 10197 820
rect 10924 860 10964 1156
rect 10924 811 10964 820
rect 11116 1196 11156 1205
rect 11116 860 11156 1156
rect 11116 811 11156 820
rect 11308 272 11348 2332
rect 11308 223 11348 232
rect 11500 197 11540 11068
rect 11596 1952 11636 11572
rect 11788 9437 11828 13588
rect 11884 9764 11924 15520
rect 11980 12788 12020 25012
rect 12268 23792 12308 23801
rect 12268 22112 12308 23752
rect 12075 21524 12117 21533
rect 12075 21484 12076 21524
rect 12116 21484 12117 21524
rect 12075 21475 12117 21484
rect 11980 12739 12020 12748
rect 11884 9715 11924 9724
rect 11980 11696 12020 11705
rect 11787 9428 11829 9437
rect 11787 9388 11788 9428
rect 11828 9388 11829 9428
rect 11787 9379 11829 9388
rect 11692 7916 11732 7925
rect 11692 6572 11732 7876
rect 11692 6523 11732 6532
rect 11980 6236 12020 11656
rect 11980 6187 12020 6196
rect 11980 3968 12020 3977
rect 11980 3137 12020 3928
rect 12076 3800 12116 21475
rect 12268 21440 12308 22072
rect 12268 21391 12308 21400
rect 12364 20180 12404 32740
rect 12268 20140 12404 20180
rect 12172 13880 12212 13889
rect 12172 8177 12212 13840
rect 12268 13628 12308 20140
rect 12460 15140 12500 39964
rect 12556 16736 12596 41560
rect 13900 41432 13940 41441
rect 13707 40508 13749 40517
rect 13707 40468 13708 40508
rect 13748 40468 13749 40508
rect 13707 40459 13749 40468
rect 12940 39752 12980 39761
rect 12747 39500 12789 39509
rect 12747 39460 12748 39500
rect 12788 39460 12789 39500
rect 12747 39451 12789 39460
rect 12652 38576 12692 38585
rect 12652 37652 12692 38536
rect 12652 37603 12692 37612
rect 12748 37241 12788 39451
rect 12844 39248 12884 39257
rect 12844 37904 12884 39208
rect 12844 37855 12884 37864
rect 12747 37232 12789 37241
rect 12747 37192 12748 37232
rect 12788 37192 12789 37232
rect 12747 37183 12789 37192
rect 12652 32360 12692 32369
rect 12652 31856 12692 32320
rect 12940 32360 12980 39712
rect 13420 38156 13460 38165
rect 13036 37820 13076 37829
rect 13036 35477 13076 37780
rect 13131 37652 13173 37661
rect 13131 37612 13132 37652
rect 13172 37612 13173 37652
rect 13131 37603 13173 37612
rect 13132 37493 13172 37603
rect 13324 37568 13364 37577
rect 13131 37484 13173 37493
rect 13131 37444 13132 37484
rect 13172 37444 13173 37484
rect 13131 37435 13173 37444
rect 13132 35888 13172 35897
rect 13035 35468 13077 35477
rect 13035 35428 13036 35468
rect 13076 35428 13077 35468
rect 13035 35419 13077 35428
rect 13132 35300 13172 35848
rect 12940 32311 12980 32320
rect 13036 35260 13172 35300
rect 13228 35804 13268 35813
rect 13036 32780 13076 35260
rect 13228 35048 13268 35764
rect 13324 35636 13364 37528
rect 13324 35587 13364 35596
rect 12652 27665 12692 31816
rect 12940 31688 12980 31697
rect 12844 29168 12884 29177
rect 12651 27656 12693 27665
rect 12651 27616 12652 27656
rect 12692 27616 12693 27656
rect 12651 27607 12693 27616
rect 12652 23288 12692 27607
rect 12844 25304 12884 29128
rect 12940 26648 12980 31648
rect 12940 26599 12980 26608
rect 12844 25255 12884 25264
rect 13036 25976 13076 32740
rect 13036 24632 13076 25936
rect 13132 33284 13172 33293
rect 13132 29168 13172 33244
rect 13228 31436 13268 35008
rect 13324 34208 13364 34217
rect 13324 33629 13364 34168
rect 13323 33620 13365 33629
rect 13323 33580 13324 33620
rect 13364 33580 13365 33620
rect 13323 33571 13365 33580
rect 13420 32369 13460 38116
rect 13516 35216 13556 35225
rect 13516 35057 13556 35176
rect 13515 35048 13557 35057
rect 13515 35008 13516 35048
rect 13556 35008 13557 35048
rect 13515 34999 13557 35008
rect 13516 34376 13556 34999
rect 13516 34327 13556 34336
rect 13515 33620 13557 33629
rect 13515 33580 13516 33620
rect 13556 33580 13557 33620
rect 13515 33571 13557 33580
rect 13419 32360 13461 32369
rect 13419 32320 13420 32360
rect 13460 32320 13461 32360
rect 13419 32311 13461 32320
rect 13228 31396 13460 31436
rect 13227 31268 13269 31277
rect 13227 31228 13228 31268
rect 13268 31228 13269 31268
rect 13227 31219 13269 31228
rect 13228 31134 13268 31219
rect 13323 31184 13365 31193
rect 13323 31144 13324 31184
rect 13364 31144 13365 31184
rect 13323 31135 13365 31144
rect 13324 29756 13364 31135
rect 13324 29707 13364 29716
rect 13132 25388 13172 29128
rect 13132 25339 13172 25348
rect 13324 29504 13364 29513
rect 13036 24583 13076 24592
rect 12652 23239 12692 23248
rect 12556 16687 12596 16696
rect 12844 22868 12884 22877
rect 12460 15091 12500 15100
rect 12748 14804 12788 14813
rect 12268 13579 12308 13588
rect 12364 13964 12404 13973
rect 12268 12368 12308 12377
rect 12268 8588 12308 12328
rect 12268 8539 12308 8548
rect 12364 8336 12404 13924
rect 12364 8287 12404 8296
rect 12460 13796 12500 13805
rect 12171 8168 12213 8177
rect 12171 8128 12172 8168
rect 12212 8128 12213 8168
rect 12171 8119 12213 8128
rect 12268 8084 12308 8093
rect 12268 6488 12308 8044
rect 12268 6439 12308 6448
rect 12364 6740 12404 6749
rect 12076 3751 12116 3760
rect 11979 3128 12021 3137
rect 11979 3088 11980 3128
rect 12020 3088 12021 3128
rect 11979 3079 12021 3088
rect 11883 2708 11925 2717
rect 11883 2668 11884 2708
rect 11924 2668 11925 2708
rect 11883 2659 11925 2668
rect 11884 2120 11924 2659
rect 11884 2071 11924 2080
rect 11596 1903 11636 1912
rect 12364 1121 12404 6700
rect 12460 3221 12500 13756
rect 12556 12116 12596 12125
rect 12556 9941 12596 12076
rect 12652 11864 12692 11873
rect 12652 11285 12692 11824
rect 12651 11276 12693 11285
rect 12651 11236 12652 11276
rect 12692 11236 12693 11276
rect 12651 11227 12693 11236
rect 12555 9932 12597 9941
rect 12555 9892 12556 9932
rect 12596 9892 12597 9932
rect 12555 9883 12597 9892
rect 12556 9008 12596 9017
rect 12459 3212 12501 3221
rect 12459 3172 12460 3212
rect 12500 3172 12501 3212
rect 12459 3163 12501 3172
rect 12556 1280 12596 8968
rect 12748 9008 12788 14764
rect 12748 8959 12788 8968
rect 12651 7076 12693 7085
rect 12651 7036 12652 7076
rect 12692 7036 12693 7076
rect 12651 7027 12693 7036
rect 12652 6942 12692 7027
rect 12844 5069 12884 22828
rect 13324 22448 13364 29464
rect 13420 27236 13460 31396
rect 13420 27187 13460 27196
rect 13324 22399 13364 22408
rect 13420 26648 13460 26657
rect 13228 18416 13268 18425
rect 13036 16148 13076 16157
rect 13036 11696 13076 16108
rect 13228 15476 13268 18376
rect 13228 15436 13364 15476
rect 13036 11647 13076 11656
rect 13228 13628 13268 13637
rect 13131 10184 13173 10193
rect 13131 10144 13132 10184
rect 13172 10144 13173 10184
rect 13131 10135 13173 10144
rect 13035 6320 13077 6329
rect 13035 6280 13036 6320
rect 13076 6280 13077 6320
rect 13035 6271 13077 6280
rect 12940 5480 12980 5489
rect 12843 5060 12885 5069
rect 12843 5020 12844 5060
rect 12884 5020 12885 5060
rect 12843 5011 12885 5020
rect 12940 3548 12980 5440
rect 12940 3499 12980 3508
rect 13036 2540 13076 6271
rect 13132 5825 13172 10135
rect 13228 8177 13268 13588
rect 13227 8168 13269 8177
rect 13227 8128 13228 8168
rect 13268 8128 13269 8168
rect 13227 8119 13269 8128
rect 13228 8000 13268 8009
rect 13324 8000 13364 15436
rect 13268 7960 13364 8000
rect 13131 5816 13173 5825
rect 13131 5776 13132 5816
rect 13172 5776 13173 5816
rect 13131 5767 13173 5776
rect 13036 2500 13172 2540
rect 12556 1231 12596 1240
rect 12747 1280 12789 1289
rect 12747 1240 12748 1280
rect 12788 1240 12789 1280
rect 12747 1231 12789 1240
rect 13132 1280 13172 2500
rect 13228 2204 13268 7960
rect 13420 6236 13460 26608
rect 13516 24044 13556 33571
rect 13611 28664 13653 28673
rect 13611 28624 13612 28664
rect 13652 28624 13653 28664
rect 13611 28615 13653 28624
rect 13612 28412 13652 28615
rect 13612 27740 13652 28372
rect 13612 27691 13652 27700
rect 13516 23995 13556 24004
rect 13612 25388 13652 25397
rect 13612 17828 13652 25348
rect 13516 17788 13612 17828
rect 13516 11864 13556 17788
rect 13612 17779 13652 17788
rect 13611 15392 13653 15401
rect 13611 15352 13612 15392
rect 13652 15352 13653 15392
rect 13611 15343 13653 15352
rect 13612 15258 13652 15343
rect 13611 15140 13653 15149
rect 13611 15100 13612 15140
rect 13652 15100 13653 15140
rect 13611 15091 13653 15100
rect 13612 14729 13652 15091
rect 13611 14720 13653 14729
rect 13611 14680 13612 14720
rect 13652 14680 13653 14720
rect 13611 14671 13653 14680
rect 13516 11815 13556 11824
rect 13612 14132 13652 14141
rect 13420 6187 13460 6196
rect 13516 11360 13556 11369
rect 13323 4724 13365 4733
rect 13323 4684 13324 4724
rect 13364 4684 13365 4724
rect 13323 4675 13365 4684
rect 13324 4388 13364 4675
rect 13324 4339 13364 4348
rect 13228 2045 13268 2164
rect 13227 2036 13269 2045
rect 13227 1996 13228 2036
rect 13268 1996 13269 2036
rect 13227 1987 13269 1996
rect 13132 1231 13172 1240
rect 13516 1280 13556 11320
rect 13612 10193 13652 14092
rect 13611 10184 13653 10193
rect 13611 10144 13612 10184
rect 13652 10144 13653 10184
rect 13611 10135 13653 10144
rect 13611 10016 13653 10025
rect 13611 9976 13612 10016
rect 13652 9976 13653 10016
rect 13611 9967 13653 9976
rect 13612 9882 13652 9967
rect 13611 8168 13653 8177
rect 13611 8128 13612 8168
rect 13652 8128 13653 8168
rect 13611 8119 13653 8128
rect 13516 1231 13556 1240
rect 12748 1146 12788 1231
rect 12363 1112 12405 1121
rect 12363 1072 12364 1112
rect 12404 1072 12405 1112
rect 12363 1063 12405 1072
rect 13612 440 13652 8119
rect 13708 1280 13748 40459
rect 13900 39668 13940 41392
rect 14764 41096 14804 41105
rect 14572 40760 14612 40769
rect 14380 40676 14420 40685
rect 13900 39619 13940 39628
rect 14284 40088 14324 40097
rect 13996 38828 14036 38837
rect 13996 37493 14036 38788
rect 14188 37820 14228 37829
rect 13995 37484 14037 37493
rect 13995 37444 13996 37484
rect 14036 37444 14037 37484
rect 13995 37435 14037 37444
rect 13803 35132 13845 35141
rect 13803 35092 13804 35132
rect 13844 35092 13845 35132
rect 13803 35083 13845 35092
rect 13804 32453 13844 35083
rect 13900 33620 13940 33629
rect 13803 32444 13845 32453
rect 13803 32404 13804 32444
rect 13844 32404 13845 32444
rect 13803 32395 13845 32404
rect 13804 20012 13844 32395
rect 13900 27824 13940 33580
rect 13900 27775 13940 27784
rect 13996 28244 14036 37435
rect 14188 35225 14228 37780
rect 14092 35216 14132 35225
rect 14092 30344 14132 35176
rect 14187 35216 14229 35225
rect 14187 35176 14188 35216
rect 14228 35176 14229 35216
rect 14187 35167 14229 35176
rect 14092 30295 14132 30304
rect 14188 34124 14228 34133
rect 13804 19172 13844 19972
rect 13804 19123 13844 19132
rect 13900 22196 13940 22205
rect 13996 22196 14036 28204
rect 14092 30092 14132 30101
rect 14092 27656 14132 30052
rect 14188 29000 14228 34084
rect 14284 33704 14324 40048
rect 14380 39761 14420 40636
rect 14379 39752 14421 39761
rect 14379 39712 14380 39752
rect 14420 39712 14421 39752
rect 14379 39703 14421 39712
rect 14284 33655 14324 33664
rect 14284 30764 14324 30773
rect 14284 29252 14324 30724
rect 14284 29203 14324 29212
rect 14188 28960 14324 29000
rect 14092 27607 14132 27616
rect 14092 27068 14132 27077
rect 14092 25556 14132 27028
rect 14092 25507 14132 25516
rect 13940 22156 14036 22196
rect 14092 25220 14132 25229
rect 14092 24968 14132 25180
rect 13900 21104 13940 22156
rect 13804 19004 13844 19013
rect 13804 18248 13844 18964
rect 13804 18199 13844 18208
rect 13804 15728 13844 15737
rect 13804 14804 13844 15688
rect 13804 11696 13844 14764
rect 13804 8504 13844 11656
rect 13900 8924 13940 21064
rect 13996 19844 14036 19853
rect 13996 17156 14036 19804
rect 14092 19088 14132 24928
rect 14092 19039 14132 19048
rect 13996 17107 14036 17116
rect 13995 14888 14037 14897
rect 13995 14848 13996 14888
rect 14036 14848 14037 14888
rect 13995 14839 14037 14848
rect 13996 9848 14036 14839
rect 14188 11528 14228 11537
rect 13996 9799 14036 9808
rect 14092 11276 14132 11285
rect 13900 8884 14036 8924
rect 13899 8756 13941 8765
rect 13899 8716 13900 8756
rect 13940 8716 13941 8756
rect 13899 8707 13941 8716
rect 13900 8588 13940 8707
rect 13900 8539 13940 8548
rect 13804 8168 13844 8464
rect 13804 8119 13844 8128
rect 13804 7412 13844 7421
rect 13804 4985 13844 7372
rect 13996 6068 14036 8884
rect 14092 7505 14132 11236
rect 14091 7496 14133 7505
rect 14091 7456 14092 7496
rect 14132 7456 14133 7496
rect 14091 7447 14133 7456
rect 13996 6019 14036 6028
rect 14092 6992 14132 7001
rect 13996 5312 14036 5321
rect 13899 5060 13941 5069
rect 13899 5020 13900 5060
rect 13940 5020 13941 5060
rect 13899 5011 13941 5020
rect 13803 4976 13845 4985
rect 13803 4936 13804 4976
rect 13844 4936 13845 4976
rect 13803 4927 13845 4936
rect 13900 3380 13940 5011
rect 13900 3331 13940 3340
rect 13996 3212 14036 5272
rect 14092 4388 14132 6952
rect 14188 5741 14228 11488
rect 14284 11360 14324 28960
rect 14380 19424 14420 39703
rect 14572 39500 14612 40720
rect 14764 40592 14804 41056
rect 14764 39584 14804 40552
rect 14764 39535 14804 39544
rect 14572 39451 14612 39460
rect 14667 39500 14709 39509
rect 14667 39460 14668 39500
rect 14708 39460 14709 39500
rect 14667 39451 14709 39460
rect 14572 35132 14612 35141
rect 14476 34376 14516 34385
rect 14476 33284 14516 34336
rect 14476 33235 14516 33244
rect 14476 32192 14516 32201
rect 14476 29924 14516 32152
rect 14476 29875 14516 29884
rect 14380 19172 14420 19384
rect 14380 19123 14420 19132
rect 14572 15896 14612 35092
rect 14572 15847 14612 15856
rect 14476 12284 14516 12293
rect 14284 11320 14420 11360
rect 14284 7412 14324 7421
rect 14284 5984 14324 7372
rect 14284 5935 14324 5944
rect 14187 5732 14229 5741
rect 14187 5692 14188 5732
rect 14228 5692 14229 5732
rect 14187 5683 14229 5692
rect 14092 4339 14132 4348
rect 13708 1231 13748 1240
rect 13900 3172 14036 3212
rect 14092 3632 14132 3641
rect 13804 1028 13844 1037
rect 13900 1028 13940 3172
rect 14092 2540 14132 3592
rect 13996 2500 14132 2540
rect 13996 2297 14036 2500
rect 13995 2288 14037 2297
rect 13995 2248 13996 2288
rect 14036 2248 14037 2288
rect 13995 2239 14037 2248
rect 13844 988 13940 1028
rect 13804 979 13844 988
rect 14283 944 14325 953
rect 14283 904 14284 944
rect 14324 904 14325 944
rect 14283 895 14325 904
rect 14284 810 14324 895
rect 14380 701 14420 11320
rect 14476 9176 14516 12244
rect 14571 11528 14613 11537
rect 14571 11488 14572 11528
rect 14612 11488 14613 11528
rect 14571 11479 14613 11488
rect 14476 9127 14516 9136
rect 14572 6161 14612 11479
rect 14571 6152 14613 6161
rect 14571 6112 14572 6152
rect 14612 6112 14613 6152
rect 14571 6103 14613 6112
rect 14476 6068 14516 6077
rect 14476 5228 14516 6028
rect 14476 5179 14516 5188
rect 14571 3044 14613 3053
rect 14571 3004 14572 3044
rect 14612 3004 14613 3044
rect 14571 2995 14613 3004
rect 14572 2910 14612 2995
rect 14571 2372 14613 2381
rect 14571 2332 14572 2372
rect 14612 2332 14613 2372
rect 14571 2323 14613 2332
rect 14572 2238 14612 2323
rect 14668 1280 14708 39451
rect 14860 38996 14900 39005
rect 14860 36644 14900 38956
rect 14764 35804 14804 35813
rect 14764 10100 14804 35764
rect 14860 30176 14900 36604
rect 15052 35468 15092 42232
rect 17548 42020 17588 42029
rect 15628 41852 15668 41861
rect 15244 41432 15284 41441
rect 15147 40760 15189 40769
rect 15147 40720 15148 40760
rect 15188 40720 15189 40760
rect 15147 40711 15189 40720
rect 15148 39425 15188 40711
rect 15147 39416 15189 39425
rect 15147 39376 15148 39416
rect 15188 39376 15189 39416
rect 15147 39367 15189 39376
rect 15244 38492 15284 41392
rect 15244 38443 15284 38452
rect 15340 41264 15380 41273
rect 15244 37484 15284 37493
rect 15147 36812 15189 36821
rect 15147 36772 15148 36812
rect 15188 36772 15189 36812
rect 15147 36763 15189 36772
rect 15052 35419 15092 35428
rect 15148 35300 15188 36763
rect 15244 36560 15284 37444
rect 15244 36511 15284 36520
rect 15340 35393 15380 41224
rect 15435 37652 15477 37661
rect 15435 37612 15436 37652
rect 15476 37612 15477 37652
rect 15435 37603 15477 37612
rect 15436 37518 15476 37603
rect 15532 37316 15572 37325
rect 15436 36728 15476 36737
rect 15339 35384 15381 35393
rect 15339 35344 15340 35384
rect 15380 35344 15381 35384
rect 15339 35335 15381 35344
rect 15148 35251 15188 35260
rect 15052 34040 15092 34049
rect 14956 32360 14996 32369
rect 14956 32024 14996 32320
rect 14956 31975 14996 31984
rect 14860 30127 14900 30136
rect 14956 31772 14996 31781
rect 14956 29000 14996 31732
rect 14860 28960 14996 29000
rect 14860 27488 14900 28960
rect 14860 27439 14900 27448
rect 14956 28076 14996 28085
rect 14956 24800 14996 28036
rect 14956 24751 14996 24760
rect 14764 10051 14804 10060
rect 14860 20012 14900 20021
rect 14764 7916 14804 7925
rect 14764 4388 14804 7876
rect 14764 4339 14804 4348
rect 14860 3632 14900 19972
rect 14956 17996 14996 18005
rect 14956 15224 14996 17956
rect 14956 15175 14996 15184
rect 14955 13460 14997 13469
rect 14955 13420 14956 13460
rect 14996 13420 14997 13460
rect 14955 13411 14997 13420
rect 14956 8840 14996 13411
rect 14956 8791 14996 8800
rect 14860 3583 14900 3592
rect 14668 1231 14708 1240
rect 14379 692 14421 701
rect 14379 652 14380 692
rect 14420 652 14421 692
rect 14379 643 14421 652
rect 15052 524 15092 34000
rect 15244 33704 15284 33713
rect 15148 32948 15188 32957
rect 15148 32024 15188 32908
rect 15148 31975 15188 31984
rect 15148 31604 15188 31613
rect 15148 30428 15188 31564
rect 15148 30379 15188 30388
rect 15244 28421 15284 33664
rect 15340 32024 15380 35335
rect 15436 34712 15476 36688
rect 15436 34663 15476 34672
rect 15436 34040 15476 34049
rect 15436 32696 15476 34000
rect 15436 32647 15476 32656
rect 15340 31975 15380 31984
rect 15436 32360 15476 32369
rect 15436 29672 15476 32320
rect 15340 29632 15476 29672
rect 15532 32192 15572 37276
rect 15628 36896 15668 41812
rect 16780 41600 16820 41609
rect 16587 40508 16629 40517
rect 16587 40468 16588 40508
rect 16628 40468 16629 40508
rect 16587 40459 16629 40468
rect 16396 40424 16436 40433
rect 15916 39752 15956 39761
rect 15820 39080 15860 39089
rect 15628 36847 15668 36856
rect 15724 37904 15764 37913
rect 15627 35300 15669 35309
rect 15627 35260 15628 35300
rect 15668 35260 15669 35300
rect 15627 35251 15669 35260
rect 15628 35166 15668 35251
rect 15724 35141 15764 37864
rect 15820 36485 15860 39040
rect 15819 36476 15861 36485
rect 15819 36436 15820 36476
rect 15860 36436 15861 36476
rect 15819 36427 15861 36436
rect 15723 35132 15765 35141
rect 15723 35092 15724 35132
rect 15764 35092 15765 35132
rect 15723 35083 15765 35092
rect 15628 34376 15668 34385
rect 15628 32612 15668 34336
rect 15723 34040 15765 34049
rect 15723 34000 15724 34040
rect 15764 34000 15765 34040
rect 15723 33991 15765 34000
rect 15628 32563 15668 32572
rect 15243 28412 15285 28421
rect 15243 28372 15244 28412
rect 15284 28372 15285 28412
rect 15243 28363 15285 28372
rect 15340 27740 15380 29632
rect 15436 29504 15476 29513
rect 15436 29000 15476 29464
rect 15436 28951 15476 28960
rect 15340 27691 15380 27700
rect 15436 28580 15476 28589
rect 15148 26228 15188 26237
rect 15148 25220 15188 26188
rect 15148 25171 15188 25180
rect 15436 25136 15476 28540
rect 15532 25388 15572 32152
rect 15532 25339 15572 25348
rect 15628 27740 15668 27749
rect 15436 25087 15476 25096
rect 15340 23708 15380 23717
rect 15340 23120 15380 23668
rect 15148 11864 15188 11873
rect 15148 9176 15188 11824
rect 15148 9127 15188 9136
rect 15244 10100 15284 10109
rect 15244 6497 15284 10060
rect 15340 8345 15380 23080
rect 15532 15980 15572 15989
rect 15436 11453 15476 11538
rect 15435 11444 15477 11453
rect 15435 11404 15436 11444
rect 15476 11404 15477 11444
rect 15435 11395 15477 11404
rect 15435 10940 15477 10949
rect 15435 10900 15436 10940
rect 15476 10900 15477 10940
rect 15435 10891 15477 10900
rect 15339 8336 15381 8345
rect 15339 8296 15340 8336
rect 15380 8296 15381 8336
rect 15339 8287 15381 8296
rect 15243 6488 15285 6497
rect 15243 6448 15244 6488
rect 15284 6448 15285 6488
rect 15243 6439 15285 6448
rect 15244 2540 15284 6439
rect 15244 2491 15284 2500
rect 15340 4724 15380 8287
rect 15436 5657 15476 10891
rect 15532 9512 15572 15940
rect 15532 9463 15572 9472
rect 15531 7328 15573 7337
rect 15531 7288 15532 7328
rect 15572 7288 15573 7328
rect 15531 7279 15573 7288
rect 15435 5648 15477 5657
rect 15435 5608 15436 5648
rect 15476 5608 15477 5648
rect 15435 5599 15477 5608
rect 15532 5564 15572 7279
rect 15532 5515 15572 5524
rect 15340 2288 15380 4684
rect 15340 2239 15380 2248
rect 15435 1700 15477 1709
rect 15435 1660 15436 1700
rect 15476 1660 15477 1700
rect 15435 1651 15477 1660
rect 15436 1280 15476 1651
rect 15436 1231 15476 1240
rect 15628 1280 15668 27700
rect 15724 27488 15764 33991
rect 15916 33116 15956 39712
rect 16108 39500 16148 39509
rect 16012 38408 16052 38417
rect 16012 35636 16052 38368
rect 16012 35587 16052 35596
rect 16012 34124 16052 34133
rect 16012 33704 16052 34084
rect 16012 33655 16052 33664
rect 15956 33076 16052 33116
rect 15916 33067 15956 33076
rect 15724 27439 15764 27448
rect 15820 32528 15860 32537
rect 15820 29168 15860 32488
rect 15915 32360 15957 32369
rect 15915 32320 15916 32360
rect 15956 32320 15957 32360
rect 15915 32311 15957 32320
rect 15723 25976 15765 25985
rect 15723 25936 15724 25976
rect 15764 25936 15765 25976
rect 15723 25927 15765 25936
rect 15724 20684 15764 25927
rect 15820 25304 15860 29128
rect 15820 25255 15860 25264
rect 15724 20635 15764 20644
rect 15820 20012 15860 20021
rect 15820 17828 15860 19972
rect 15820 17779 15860 17788
rect 15724 14720 15764 14729
rect 15724 7337 15764 14680
rect 15820 13712 15860 13721
rect 15820 11696 15860 13672
rect 15820 10184 15860 11656
rect 15820 10135 15860 10144
rect 15820 7412 15860 7421
rect 15723 7328 15765 7337
rect 15723 7288 15724 7328
rect 15764 7288 15765 7328
rect 15723 7279 15765 7288
rect 15724 6824 15764 6835
rect 15724 6749 15764 6784
rect 15723 6740 15765 6749
rect 15723 6700 15724 6740
rect 15764 6700 15765 6740
rect 15723 6691 15765 6700
rect 15820 3548 15860 7372
rect 15820 3499 15860 3508
rect 15916 1364 15956 32311
rect 16012 19340 16052 33076
rect 16012 19291 16052 19300
rect 16011 12284 16053 12293
rect 16011 12244 16012 12284
rect 16052 12244 16053 12284
rect 16011 12235 16053 12244
rect 16012 10949 16052 12235
rect 16011 10940 16053 10949
rect 16011 10900 16012 10940
rect 16052 10900 16053 10940
rect 16011 10891 16053 10900
rect 16108 10772 16148 39460
rect 16300 38156 16340 38165
rect 16204 37064 16244 37073
rect 16204 36644 16244 37024
rect 16300 36812 16340 38116
rect 16396 36821 16436 40384
rect 16588 39920 16628 40459
rect 16588 39871 16628 39880
rect 16684 40088 16724 40097
rect 16588 39668 16628 39677
rect 16492 37820 16532 37860
rect 16492 37736 16532 37780
rect 16492 37687 16532 37696
rect 16492 37316 16532 37325
rect 16300 36763 16340 36772
rect 16395 36812 16437 36821
rect 16395 36772 16396 36812
rect 16436 36772 16437 36812
rect 16395 36763 16437 36772
rect 16492 36812 16532 37276
rect 16492 36763 16532 36772
rect 16204 36604 16436 36644
rect 16203 36476 16245 36485
rect 16203 36436 16204 36476
rect 16244 36436 16245 36476
rect 16203 36427 16245 36436
rect 16204 35057 16244 36427
rect 16300 35384 16340 35395
rect 16300 35309 16340 35344
rect 16299 35300 16341 35309
rect 16299 35260 16300 35300
rect 16340 35260 16341 35300
rect 16299 35251 16341 35260
rect 16203 35048 16245 35057
rect 16203 35008 16204 35048
rect 16244 35008 16245 35048
rect 16203 34999 16245 35008
rect 16204 25472 16244 34999
rect 16299 34964 16341 34973
rect 16299 34924 16300 34964
rect 16340 34924 16341 34964
rect 16299 34915 16341 34924
rect 16300 33620 16340 34915
rect 16300 33571 16340 33580
rect 16300 32696 16340 32705
rect 16300 29756 16340 32656
rect 16300 29707 16340 29716
rect 16396 31184 16436 36604
rect 16588 34628 16628 39628
rect 16684 34964 16724 40048
rect 16684 34915 16724 34924
rect 16588 34579 16628 34588
rect 16492 34040 16532 34049
rect 16492 33965 16532 34000
rect 16491 33956 16533 33965
rect 16491 33916 16492 33956
rect 16532 33916 16533 33956
rect 16491 33907 16533 33916
rect 16492 33905 16532 33907
rect 16683 32948 16725 32957
rect 16683 32908 16684 32948
rect 16724 32908 16725 32948
rect 16683 32899 16725 32908
rect 16684 32814 16724 32899
rect 16780 31940 16820 41560
rect 16972 41600 17012 41609
rect 16875 39752 16917 39761
rect 16875 39712 16876 39752
rect 16916 39712 16917 39752
rect 16875 39703 16917 39712
rect 16876 39618 16916 39703
rect 16876 38492 16916 38501
rect 16876 37736 16916 38452
rect 16876 37687 16916 37696
rect 16876 37232 16916 37241
rect 16876 36728 16916 37192
rect 16876 36679 16916 36688
rect 16204 25423 16244 25432
rect 16300 27488 16340 27497
rect 16012 10732 16148 10772
rect 16204 25220 16244 25229
rect 16012 10100 16052 10732
rect 16012 10051 16052 10060
rect 16108 10604 16148 10613
rect 16108 3296 16148 10564
rect 16108 3247 16148 3256
rect 16204 2540 16244 25180
rect 16300 23792 16340 27448
rect 16300 23743 16340 23752
rect 16299 22952 16341 22961
rect 16299 22912 16300 22952
rect 16340 22912 16341 22952
rect 16299 22903 16341 22912
rect 16300 16904 16340 22903
rect 16300 16855 16340 16864
rect 16396 15140 16436 31144
rect 16492 31900 16820 31940
rect 16876 36476 16916 36485
rect 16492 22700 16532 31900
rect 16876 31520 16916 36436
rect 16780 31480 16876 31520
rect 16587 29252 16629 29261
rect 16587 29212 16588 29252
rect 16628 29212 16629 29252
rect 16780 29252 16820 31480
rect 16876 31471 16916 31480
rect 16875 31268 16917 31277
rect 16875 31228 16876 31268
rect 16916 31228 16917 31268
rect 16875 31219 16917 31228
rect 16876 29420 16916 31219
rect 16876 29371 16916 29380
rect 16780 29212 16916 29252
rect 16587 29203 16629 29212
rect 16588 29168 16628 29203
rect 16588 29117 16628 29128
rect 16684 27236 16724 27245
rect 16587 26732 16629 26741
rect 16587 26692 16588 26732
rect 16628 26692 16629 26732
rect 16587 26683 16629 26692
rect 16588 25220 16628 26683
rect 16684 26648 16724 27196
rect 16684 26599 16724 26608
rect 16780 26900 16820 26909
rect 16780 26396 16820 26860
rect 16684 26356 16820 26396
rect 16684 26144 16724 26356
rect 16684 26095 16724 26104
rect 16780 26228 16820 26237
rect 16683 25724 16725 25733
rect 16683 25684 16684 25724
rect 16724 25684 16725 25724
rect 16683 25675 16725 25684
rect 16780 25724 16820 26188
rect 16780 25675 16820 25684
rect 16588 25171 16628 25180
rect 16492 22651 16532 22660
rect 16588 23708 16628 23717
rect 16492 22280 16532 22289
rect 16492 22028 16532 22240
rect 16492 21104 16532 21988
rect 16492 21055 16532 21064
rect 16588 19928 16628 23668
rect 16491 15980 16533 15989
rect 16491 15940 16492 15980
rect 16532 15940 16533 15980
rect 16491 15931 16533 15940
rect 16492 15149 16532 15931
rect 16396 15091 16436 15100
rect 16491 15140 16533 15149
rect 16491 15100 16492 15140
rect 16532 15100 16533 15140
rect 16491 15091 16533 15100
rect 16588 14972 16628 19888
rect 16684 18416 16724 25675
rect 16780 25472 16820 25481
rect 16780 20441 16820 25432
rect 16876 24641 16916 29212
rect 16875 24632 16917 24641
rect 16875 24592 16876 24632
rect 16916 24592 16917 24632
rect 16875 24583 16917 24592
rect 16876 21776 16916 21785
rect 16876 21608 16916 21736
rect 16876 21559 16916 21568
rect 16972 20600 17012 41560
rect 17548 41348 17588 41980
rect 17548 41299 17588 41308
rect 17740 42020 17780 42029
rect 17164 41012 17204 41021
rect 17068 40592 17108 40601
rect 17068 25220 17108 40552
rect 17068 25171 17108 25180
rect 17164 24044 17204 40972
rect 17547 41012 17589 41021
rect 17547 40972 17548 41012
rect 17588 40972 17589 41012
rect 17547 40963 17589 40972
rect 17548 40878 17588 40963
rect 17644 40928 17684 40937
rect 17260 40844 17300 40853
rect 17260 38996 17300 40804
rect 17644 40685 17684 40888
rect 17643 40676 17685 40685
rect 17643 40636 17644 40676
rect 17684 40636 17685 40676
rect 17643 40627 17685 40636
rect 17260 38947 17300 38956
rect 17548 40592 17588 40601
rect 17452 37904 17492 37913
rect 17452 37400 17492 37864
rect 17452 37351 17492 37360
rect 17356 37316 17396 37325
rect 17356 36392 17396 37276
rect 17356 36343 17396 36352
rect 17452 36812 17492 36821
rect 17452 35972 17492 36772
rect 17452 35923 17492 35932
rect 17356 35384 17396 35393
rect 17259 35216 17301 35225
rect 17259 35176 17260 35216
rect 17300 35176 17301 35216
rect 17259 35167 17301 35176
rect 17260 31352 17300 35167
rect 17356 35141 17396 35344
rect 17355 35132 17397 35141
rect 17355 35092 17356 35132
rect 17396 35092 17397 35132
rect 17355 35083 17397 35092
rect 17260 31303 17300 31312
rect 17451 31268 17493 31277
rect 17451 31228 17452 31268
rect 17492 31228 17493 31268
rect 17451 31219 17493 31228
rect 17452 30848 17492 31219
rect 17452 30799 17492 30808
rect 17260 30680 17300 30689
rect 17260 27908 17300 30640
rect 17260 26648 17300 27868
rect 17452 30596 17492 30605
rect 17452 27656 17492 30556
rect 17452 27607 17492 27616
rect 17260 26599 17300 26608
rect 17356 26900 17396 26909
rect 17259 24632 17301 24641
rect 17259 24592 17260 24632
rect 17300 24592 17301 24632
rect 17259 24583 17301 24592
rect 16876 20560 17012 20600
rect 17068 24004 17204 24044
rect 16779 20432 16821 20441
rect 16779 20392 16780 20432
rect 16820 20392 16821 20432
rect 16779 20383 16821 20392
rect 16684 18367 16724 18376
rect 16780 19592 16820 19601
rect 16492 14932 16628 14972
rect 16396 14636 16436 14645
rect 16300 14216 16340 14225
rect 16300 7421 16340 14176
rect 16396 11276 16436 14596
rect 16396 11227 16436 11236
rect 16396 8840 16436 8849
rect 16396 8336 16436 8800
rect 16396 8287 16436 8296
rect 16492 8168 16532 14932
rect 16780 14888 16820 19552
rect 16876 19004 16916 20560
rect 16971 20432 17013 20441
rect 16971 20392 16972 20432
rect 17012 20392 17013 20432
rect 16971 20383 17013 20392
rect 16876 18955 16916 18964
rect 16876 16568 16916 16577
rect 16876 15644 16916 16528
rect 16972 15821 17012 20383
rect 17068 15989 17108 24004
rect 17163 22280 17205 22289
rect 17163 22240 17164 22280
rect 17204 22240 17205 22280
rect 17163 22231 17205 22240
rect 17164 22146 17204 22231
rect 17164 19844 17204 19853
rect 17164 19256 17204 19804
rect 17164 19207 17204 19216
rect 17260 19424 17300 24583
rect 17164 19088 17204 19097
rect 17067 15980 17109 15989
rect 17067 15940 17068 15980
rect 17108 15940 17109 15980
rect 17067 15931 17109 15940
rect 16971 15812 17013 15821
rect 16971 15772 16972 15812
rect 17012 15772 17013 15812
rect 16971 15763 17013 15772
rect 16876 15604 17108 15644
rect 16588 14848 16820 14888
rect 16876 15476 16916 15485
rect 16588 10100 16628 14848
rect 16876 14552 16916 15436
rect 16876 14503 16916 14512
rect 16972 15308 17012 15317
rect 16972 11864 17012 15268
rect 16684 11696 16724 11705
rect 16684 11276 16724 11656
rect 16972 11696 17012 11824
rect 16972 11647 17012 11656
rect 16684 11236 16820 11276
rect 16780 11108 16820 11236
rect 16588 10051 16628 10060
rect 16684 10940 16724 10949
rect 16396 8128 16532 8168
rect 16588 9680 16628 9689
rect 16588 8588 16628 9640
rect 16299 7412 16341 7421
rect 16299 7372 16300 7412
rect 16340 7372 16341 7412
rect 16299 7363 16341 7372
rect 16396 7412 16436 8128
rect 16588 7748 16628 8548
rect 16396 7363 16436 7372
rect 16492 7496 16532 7505
rect 16300 4892 16340 4901
rect 16300 3464 16340 4852
rect 16492 4640 16532 7456
rect 16588 6152 16628 7708
rect 16684 6740 16724 10900
rect 16780 7496 16820 11068
rect 16780 7447 16820 7456
rect 16876 11024 16916 11033
rect 16684 6691 16724 6700
rect 16588 6103 16628 6112
rect 16492 4136 16532 4600
rect 16588 4136 16628 4145
rect 16492 4096 16588 4136
rect 16588 4087 16628 4096
rect 16300 3415 16340 3424
rect 16780 3800 16820 3809
rect 16204 2500 16340 2540
rect 15916 1315 15956 1324
rect 15628 1231 15668 1240
rect 15052 475 15092 484
rect 13612 391 13652 400
rect 16300 272 16340 2500
rect 16300 223 16340 232
rect 11499 188 11541 197
rect 11499 148 11500 188
rect 11540 148 11541 188
rect 11499 139 11541 148
rect 6027 104 6069 113
rect 6027 64 6028 104
rect 6068 64 6069 104
rect 6027 55 6069 64
rect 10059 104 10101 113
rect 10059 64 10060 104
rect 10100 64 10101 104
rect 10059 55 10101 64
rect 16780 104 16820 3760
rect 16876 3464 16916 10984
rect 16972 8756 17012 8765
rect 16972 8168 17012 8716
rect 16972 8119 17012 8128
rect 17068 5312 17108 15604
rect 17164 15308 17204 19048
rect 17260 17828 17300 19384
rect 17260 17779 17300 17788
rect 17164 15268 17300 15308
rect 17164 15140 17204 15149
rect 17164 9932 17204 15100
rect 17164 9883 17204 9892
rect 17164 9344 17204 9353
rect 17164 7244 17204 9304
rect 17164 7195 17204 7204
rect 17068 5263 17108 5272
rect 16876 3415 16916 3424
rect 17067 3212 17109 3221
rect 17067 3172 17068 3212
rect 17108 3172 17109 3212
rect 17067 3163 17109 3172
rect 17068 3078 17108 3163
rect 17260 2708 17300 15268
rect 17356 4472 17396 26860
rect 17452 26816 17492 26827
rect 17452 26741 17492 26776
rect 17451 26732 17493 26741
rect 17451 26692 17452 26732
rect 17492 26692 17493 26732
rect 17451 26683 17493 26692
rect 17451 15812 17493 15821
rect 17451 15772 17452 15812
rect 17492 15772 17493 15812
rect 17451 15763 17493 15772
rect 17356 4423 17396 4432
rect 17260 2659 17300 2668
rect 17452 1280 17492 15763
rect 17548 1532 17588 40552
rect 17644 38240 17684 38249
rect 17644 36308 17684 38200
rect 17644 36259 17684 36268
rect 17644 34040 17684 34049
rect 17644 33965 17684 34000
rect 17643 33956 17685 33965
rect 17643 33916 17644 33956
rect 17684 33916 17685 33956
rect 17643 33907 17685 33916
rect 17644 33032 17684 33907
rect 17644 32983 17684 32992
rect 17740 27068 17780 41980
rect 17836 41768 17876 41777
rect 17836 39836 17876 41728
rect 18124 41600 18164 41609
rect 18028 41348 18068 41357
rect 17932 41012 17972 41021
rect 17932 40769 17972 40972
rect 17931 40760 17973 40769
rect 17931 40720 17932 40760
rect 17972 40720 17973 40760
rect 17931 40711 17973 40720
rect 17932 40592 17972 40601
rect 17932 40349 17972 40552
rect 17931 40340 17973 40349
rect 17931 40300 17932 40340
rect 17972 40300 17973 40340
rect 17931 40291 17973 40300
rect 17836 39787 17876 39796
rect 17932 39080 17972 39089
rect 17835 35636 17877 35645
rect 17835 35596 17836 35636
rect 17876 35596 17877 35636
rect 17835 35587 17877 35596
rect 17836 35502 17876 35587
rect 17740 27019 17780 27028
rect 17836 34124 17876 34133
rect 17740 26144 17780 26153
rect 17740 25304 17780 26104
rect 17740 25255 17780 25264
rect 17643 25220 17685 25229
rect 17643 25180 17644 25220
rect 17684 25180 17685 25220
rect 17643 25171 17685 25180
rect 17644 20180 17684 25171
rect 17740 24548 17780 24557
rect 17740 21356 17780 24508
rect 17836 22700 17876 34084
rect 17932 30512 17972 39040
rect 18028 38744 18068 41308
rect 18124 39248 18164 41560
rect 18316 41012 18356 41021
rect 18124 39199 18164 39208
rect 18220 39668 18260 39677
rect 18028 38695 18068 38704
rect 18220 35645 18260 39628
rect 18124 35636 18164 35645
rect 18028 35468 18068 35477
rect 18028 32612 18068 35428
rect 18124 35048 18164 35596
rect 18219 35636 18261 35645
rect 18219 35596 18220 35636
rect 18260 35596 18261 35636
rect 18219 35587 18261 35596
rect 18124 34999 18164 35008
rect 18220 35216 18260 35587
rect 18220 34376 18260 35176
rect 18220 34327 18260 34336
rect 18028 32563 18068 32572
rect 18124 33704 18164 33713
rect 17932 30463 17972 30472
rect 18124 31184 18164 33664
rect 18220 33284 18260 33293
rect 18220 32108 18260 33244
rect 18220 31268 18260 32068
rect 18220 31219 18260 31228
rect 18124 28337 18164 31144
rect 18123 28328 18165 28337
rect 18123 28288 18124 28328
rect 18164 28288 18165 28328
rect 18123 28279 18165 28288
rect 18027 27656 18069 27665
rect 18027 27616 18028 27656
rect 18068 27616 18069 27656
rect 18027 27607 18069 27616
rect 18028 26900 18068 27607
rect 18028 26851 18068 26860
rect 18028 25556 18068 25565
rect 17931 24716 17973 24725
rect 17931 24676 17932 24716
rect 17972 24676 17973 24716
rect 17931 24667 17973 24676
rect 17932 23960 17972 24667
rect 17932 23911 17972 23920
rect 17836 22651 17876 22660
rect 17740 21307 17780 21316
rect 18028 20348 18068 25516
rect 18219 23960 18261 23969
rect 18219 23920 18220 23960
rect 18260 23920 18261 23960
rect 18219 23911 18261 23920
rect 18028 20299 18068 20308
rect 18124 21776 18164 21785
rect 17644 20140 17780 20180
rect 17644 19676 17684 19685
rect 17644 18920 17684 19636
rect 17644 18871 17684 18880
rect 17644 15308 17684 15317
rect 17644 14384 17684 15268
rect 17644 14335 17684 14344
rect 17644 8336 17684 8345
rect 17644 4304 17684 8296
rect 17644 4255 17684 4264
rect 17548 1483 17588 1492
rect 17452 1231 17492 1240
rect 17740 1280 17780 20140
rect 17836 17660 17876 17669
rect 17836 8084 17876 17620
rect 17836 8035 17876 8044
rect 18028 11864 18068 11873
rect 17835 4976 17877 4985
rect 17835 4936 17836 4976
rect 17876 4936 17877 4976
rect 17835 4927 17877 4936
rect 18028 4976 18068 11824
rect 18028 4927 18068 4936
rect 17836 3632 17876 4927
rect 17836 3583 17876 3592
rect 18124 1952 18164 21736
rect 18124 1903 18164 1912
rect 17740 1231 17780 1240
rect 18220 1280 18260 23911
rect 18316 10856 18356 40972
rect 18508 40088 18548 42652
rect 20048 41600 20416 41609
rect 20088 41560 20130 41600
rect 20170 41560 20212 41600
rect 20252 41560 20294 41600
rect 20334 41560 20376 41600
rect 20048 41551 20416 41560
rect 18700 41012 18740 41021
rect 18508 40039 18548 40048
rect 18604 40508 18644 40517
rect 18508 39752 18548 39761
rect 18411 39500 18453 39509
rect 18411 39460 18412 39500
rect 18452 39460 18453 39500
rect 18411 39451 18453 39460
rect 18412 39366 18452 39451
rect 18412 39248 18452 39257
rect 18412 37745 18452 39208
rect 18411 37736 18453 37745
rect 18411 37696 18412 37736
rect 18452 37696 18453 37736
rect 18411 37687 18453 37696
rect 18412 35300 18452 35309
rect 18412 34292 18452 35260
rect 18508 34964 18548 39712
rect 18508 34915 18548 34924
rect 18412 30857 18452 34252
rect 18508 34796 18548 34805
rect 18508 33956 18548 34756
rect 18508 32360 18548 33916
rect 18508 32311 18548 32320
rect 18507 32108 18549 32117
rect 18507 32068 18508 32108
rect 18548 32068 18549 32108
rect 18507 32059 18549 32068
rect 18411 30848 18453 30857
rect 18411 30808 18412 30848
rect 18452 30808 18453 30848
rect 18411 30799 18453 30808
rect 18412 30680 18452 30689
rect 18412 26144 18452 30640
rect 18412 26095 18452 26104
rect 18508 25388 18548 32059
rect 18412 23960 18452 23969
rect 18412 20768 18452 23920
rect 18508 23708 18548 25348
rect 18604 25229 18644 40468
rect 18700 35804 18740 40972
rect 18808 40844 19176 40853
rect 18848 40804 18890 40844
rect 18930 40804 18972 40844
rect 19012 40804 19054 40844
rect 19094 40804 19136 40844
rect 18808 40795 19176 40804
rect 18891 40676 18933 40685
rect 18891 40636 18892 40676
rect 18932 40636 18933 40676
rect 18891 40627 18933 40636
rect 18892 40424 18932 40627
rect 18892 40375 18932 40384
rect 19756 40424 19796 40433
rect 19468 40256 19508 40265
rect 19372 39500 19412 39509
rect 18808 39332 19176 39341
rect 18848 39292 18890 39332
rect 18930 39292 18972 39332
rect 19012 39292 19054 39332
rect 19094 39292 19136 39332
rect 18808 39283 19176 39292
rect 19276 39332 19316 39341
rect 19276 39080 19316 39292
rect 19276 39031 19316 39040
rect 19276 38240 19316 38249
rect 18808 37820 19176 37829
rect 18848 37780 18890 37820
rect 18930 37780 18972 37820
rect 19012 37780 19054 37820
rect 19094 37780 19136 37820
rect 18808 37771 19176 37780
rect 19276 37568 19316 38200
rect 19372 38072 19412 39460
rect 19372 38023 19412 38032
rect 19276 36644 19316 37528
rect 19276 36595 19316 36604
rect 19372 37484 19412 37493
rect 18808 36308 19176 36317
rect 18848 36268 18890 36308
rect 18930 36268 18972 36308
rect 19012 36268 19054 36308
rect 19094 36268 19136 36308
rect 18808 36259 19176 36268
rect 18700 35755 18740 35764
rect 19276 35888 19316 35897
rect 18808 34796 19176 34805
rect 18848 34756 18890 34796
rect 18930 34756 18972 34796
rect 19012 34756 19054 34796
rect 19094 34756 19136 34796
rect 18808 34747 19176 34756
rect 18808 33284 19176 33293
rect 18848 33244 18890 33284
rect 18930 33244 18972 33284
rect 19012 33244 19054 33284
rect 19094 33244 19136 33284
rect 18808 33235 19176 33244
rect 19276 33116 19316 35848
rect 19276 33067 19316 33076
rect 18700 32192 18740 32201
rect 18700 30680 18740 32152
rect 18808 31772 19176 31781
rect 18848 31732 18890 31772
rect 18930 31732 18972 31772
rect 19012 31732 19054 31772
rect 19094 31732 19136 31772
rect 18808 31723 19176 31732
rect 18795 30848 18837 30857
rect 18795 30808 18796 30848
rect 18836 30808 18837 30848
rect 18795 30799 18837 30808
rect 18796 30714 18836 30799
rect 18700 30631 18740 30640
rect 18808 30260 19176 30269
rect 18848 30220 18890 30260
rect 18930 30220 18972 30260
rect 19012 30220 19054 30260
rect 19094 30220 19136 30260
rect 18808 30211 19176 30220
rect 19372 29000 19412 37444
rect 19468 36392 19508 40216
rect 19468 36343 19508 36352
rect 19564 39080 19604 39089
rect 19564 35888 19604 39040
rect 19468 34880 19508 34889
rect 19468 33704 19508 34840
rect 19564 34628 19604 35848
rect 19564 34579 19604 34588
rect 19660 38492 19700 38501
rect 19468 33664 19604 33704
rect 19276 28960 19412 29000
rect 19468 33536 19508 33545
rect 18808 28748 19176 28757
rect 18848 28708 18890 28748
rect 18930 28708 18972 28748
rect 19012 28708 19054 28748
rect 19094 28708 19136 28748
rect 18808 28699 19176 28708
rect 18808 27236 19176 27245
rect 18848 27196 18890 27236
rect 18930 27196 18972 27236
rect 19012 27196 19054 27236
rect 19094 27196 19136 27236
rect 18808 27187 19176 27196
rect 18700 27068 18740 27077
rect 18700 26396 18740 27028
rect 18700 26347 18740 26356
rect 18808 25724 19176 25733
rect 18848 25684 18890 25724
rect 18930 25684 18972 25724
rect 19012 25684 19054 25724
rect 19094 25684 19136 25724
rect 18808 25675 19176 25684
rect 18603 25220 18645 25229
rect 18603 25180 18604 25220
rect 18644 25180 18645 25220
rect 18603 25171 18645 25180
rect 18603 24716 18645 24725
rect 18603 24676 18604 24716
rect 18644 24676 18645 24716
rect 18603 24667 18645 24676
rect 18604 24582 18644 24667
rect 18808 24212 19176 24221
rect 18848 24172 18890 24212
rect 18930 24172 18972 24212
rect 19012 24172 19054 24212
rect 19094 24172 19136 24212
rect 18808 24163 19176 24172
rect 18508 23659 18548 23668
rect 18412 17996 18452 20728
rect 18700 22700 18740 22709
rect 18700 20600 18740 22660
rect 18808 22700 19176 22709
rect 18848 22660 18890 22700
rect 18930 22660 18972 22700
rect 19012 22660 19054 22700
rect 19094 22660 19136 22700
rect 18808 22651 19176 22660
rect 18808 21188 19176 21197
rect 18848 21148 18890 21188
rect 18930 21148 18972 21188
rect 19012 21148 19054 21188
rect 19094 21148 19136 21188
rect 18808 21139 19176 21148
rect 18700 20551 18740 20560
rect 18808 19676 19176 19685
rect 18848 19636 18890 19676
rect 18930 19636 18972 19676
rect 19012 19636 19054 19676
rect 19094 19636 19136 19676
rect 18808 19627 19176 19636
rect 18808 18164 19176 18173
rect 18848 18124 18890 18164
rect 18930 18124 18972 18164
rect 19012 18124 19054 18164
rect 19094 18124 19136 18164
rect 18808 18115 19176 18124
rect 18412 17947 18452 17956
rect 18808 16652 19176 16661
rect 18848 16612 18890 16652
rect 18930 16612 18972 16652
rect 19012 16612 19054 16652
rect 19094 16612 19136 16652
rect 18808 16603 19176 16612
rect 18700 15896 18740 15905
rect 18700 14468 18740 15856
rect 18808 15140 19176 15149
rect 18848 15100 18890 15140
rect 18930 15100 18972 15140
rect 19012 15100 19054 15140
rect 19094 15100 19136 15140
rect 18808 15091 19176 15100
rect 18700 14419 18740 14428
rect 18700 13712 18740 13721
rect 18316 10807 18356 10816
rect 18508 10856 18548 10865
rect 18315 10016 18357 10025
rect 18315 9976 18316 10016
rect 18356 9976 18357 10016
rect 18315 9967 18357 9976
rect 18316 9512 18356 9967
rect 18316 9463 18356 9472
rect 18508 8588 18548 10816
rect 18412 6740 18452 6749
rect 18316 6488 18356 6497
rect 18316 6068 18356 6448
rect 18316 6019 18356 6028
rect 18412 4976 18452 6700
rect 18508 5648 18548 8548
rect 18508 5599 18548 5608
rect 18604 8084 18644 8093
rect 18604 5396 18644 8044
rect 18604 5347 18644 5356
rect 18412 4927 18452 4936
rect 18604 4976 18644 4985
rect 18508 4640 18548 4649
rect 18604 4640 18644 4936
rect 18548 4600 18644 4640
rect 18508 4591 18548 4600
rect 18220 1231 18260 1240
rect 18412 4472 18452 4481
rect 18412 1196 18452 4432
rect 18507 4136 18549 4145
rect 18507 4096 18508 4136
rect 18548 4096 18549 4136
rect 18507 4087 18549 4096
rect 18508 4002 18548 4087
rect 18700 3212 18740 13672
rect 19276 13712 19316 28960
rect 19372 27320 19412 27329
rect 19372 25136 19412 27280
rect 19372 23960 19412 25096
rect 19372 23911 19412 23920
rect 19372 23792 19412 23801
rect 19372 23036 19412 23752
rect 19372 22532 19412 22996
rect 19372 22483 19412 22492
rect 19372 20768 19412 20777
rect 19372 19676 19412 20728
rect 19372 19627 19412 19636
rect 19468 17912 19508 33496
rect 19564 32864 19604 33664
rect 19564 32815 19604 32824
rect 19564 32528 19604 32537
rect 19564 28412 19604 32488
rect 19660 32024 19700 38452
rect 19756 34460 19796 40384
rect 20620 40340 20660 40349
rect 20048 40088 20416 40097
rect 20088 40048 20130 40088
rect 20170 40048 20212 40088
rect 20252 40048 20294 40088
rect 20334 40048 20376 40088
rect 20048 40039 20416 40048
rect 20048 38576 20416 38585
rect 20088 38536 20130 38576
rect 20170 38536 20212 38576
rect 20252 38536 20294 38576
rect 20334 38536 20376 38576
rect 20048 38527 20416 38536
rect 19852 38492 19892 38501
rect 19852 38156 19892 38452
rect 19852 38107 19892 38116
rect 19948 38240 19988 38249
rect 19948 36980 19988 38200
rect 20048 37064 20416 37073
rect 20088 37024 20130 37064
rect 20170 37024 20212 37064
rect 20252 37024 20294 37064
rect 20334 37024 20376 37064
rect 20048 37015 20416 37024
rect 19948 36931 19988 36940
rect 20620 36560 20660 40300
rect 21004 39080 21044 39089
rect 20908 38660 20948 38669
rect 20811 37232 20853 37241
rect 20811 37192 20812 37232
rect 20852 37192 20853 37232
rect 20811 37183 20853 37192
rect 20812 37064 20852 37183
rect 20812 37015 20852 37024
rect 20620 36511 20660 36520
rect 20715 36140 20757 36149
rect 20715 36100 20716 36140
rect 20756 36100 20757 36140
rect 20715 36091 20757 36100
rect 19756 34411 19796 34420
rect 19852 35636 19892 35645
rect 19852 34292 19892 35596
rect 20048 35552 20416 35561
rect 20088 35512 20130 35552
rect 20170 35512 20212 35552
rect 20252 35512 20294 35552
rect 20334 35512 20376 35552
rect 20048 35503 20416 35512
rect 19660 31975 19700 31984
rect 19756 34252 19892 34292
rect 19756 30932 19796 34252
rect 20048 34040 20416 34049
rect 20088 34000 20130 34040
rect 20170 34000 20212 34040
rect 20252 34000 20294 34040
rect 20334 34000 20376 34040
rect 20048 33991 20416 34000
rect 19851 33620 19893 33629
rect 19851 33580 19852 33620
rect 19892 33580 19893 33620
rect 19851 33571 19893 33580
rect 19852 33486 19892 33571
rect 20620 33452 20660 33461
rect 20048 32528 20416 32537
rect 20088 32488 20130 32528
rect 20170 32488 20212 32528
rect 20252 32488 20294 32528
rect 20334 32488 20376 32528
rect 20048 32479 20416 32488
rect 19756 30883 19796 30892
rect 19948 31940 19988 31949
rect 19948 29084 19988 31900
rect 20048 31016 20416 31025
rect 20088 30976 20130 31016
rect 20170 30976 20212 31016
rect 20252 30976 20294 31016
rect 20334 30976 20376 31016
rect 20048 30967 20416 30976
rect 20524 30680 20564 30689
rect 20048 29504 20416 29513
rect 20088 29464 20130 29504
rect 20170 29464 20212 29504
rect 20252 29464 20294 29504
rect 20334 29464 20376 29504
rect 20048 29455 20416 29464
rect 19948 29035 19988 29044
rect 19852 29000 19892 29009
rect 19604 28372 19700 28412
rect 19564 28363 19604 28372
rect 19564 26900 19604 26909
rect 19564 22700 19604 26860
rect 19660 26480 19700 28372
rect 19660 26431 19700 26440
rect 19852 23876 19892 28960
rect 20048 27992 20416 28001
rect 20088 27952 20130 27992
rect 20170 27952 20212 27992
rect 20252 27952 20294 27992
rect 20334 27952 20376 27992
rect 20048 27943 20416 27952
rect 19948 26732 19988 26741
rect 19948 25388 19988 26692
rect 20048 26480 20416 26489
rect 20088 26440 20130 26480
rect 20170 26440 20212 26480
rect 20252 26440 20294 26480
rect 20334 26440 20376 26480
rect 20048 26431 20416 26440
rect 19948 25339 19988 25348
rect 20048 24968 20416 24977
rect 20088 24928 20130 24968
rect 20170 24928 20212 24968
rect 20252 24928 20294 24968
rect 20334 24928 20376 24968
rect 20048 24919 20416 24928
rect 20524 23960 20564 30640
rect 20620 29504 20660 33412
rect 20716 33032 20756 36091
rect 20811 36056 20853 36065
rect 20811 36016 20812 36056
rect 20852 36016 20853 36056
rect 20811 36007 20853 36016
rect 20812 33536 20852 36007
rect 20812 33487 20852 33496
rect 20716 32983 20756 32992
rect 20908 31520 20948 38620
rect 21004 32528 21044 39040
rect 21292 38828 21332 38837
rect 21196 37568 21236 37577
rect 21196 36569 21236 37528
rect 21195 36560 21237 36569
rect 21195 36520 21196 36560
rect 21236 36520 21237 36560
rect 21195 36511 21237 36520
rect 21004 32479 21044 32488
rect 20908 31471 20948 31480
rect 21292 31016 21332 38788
rect 21292 30967 21332 30976
rect 21388 38744 21428 38753
rect 21388 30512 21428 38704
rect 21388 30463 21428 30472
rect 21388 30176 21428 30185
rect 20620 29455 20660 29464
rect 20716 30008 20756 30017
rect 20524 23911 20564 23920
rect 19852 23827 19892 23836
rect 20048 23456 20416 23465
rect 20088 23416 20130 23456
rect 20170 23416 20212 23456
rect 20252 23416 20294 23456
rect 20334 23416 20376 23456
rect 20048 23407 20416 23416
rect 19564 22651 19604 22660
rect 20048 21944 20416 21953
rect 20088 21904 20130 21944
rect 20170 21904 20212 21944
rect 20252 21904 20294 21944
rect 20334 21904 20376 21944
rect 20048 21895 20416 21904
rect 19660 20600 19700 20609
rect 19660 19676 19700 20560
rect 20048 20432 20416 20441
rect 20088 20392 20130 20432
rect 20170 20392 20212 20432
rect 20252 20392 20294 20432
rect 20334 20392 20376 20432
rect 20048 20383 20416 20392
rect 19660 19627 19700 19636
rect 20048 18920 20416 18929
rect 20088 18880 20130 18920
rect 20170 18880 20212 18920
rect 20252 18880 20294 18920
rect 20334 18880 20376 18920
rect 20048 18871 20416 18880
rect 19468 17863 19508 17872
rect 20048 17408 20416 17417
rect 20088 17368 20130 17408
rect 20170 17368 20212 17408
rect 20252 17368 20294 17408
rect 20334 17368 20376 17408
rect 20048 17359 20416 17368
rect 19756 16820 19796 16829
rect 19276 13663 19316 13672
rect 19372 15980 19412 15989
rect 19372 15476 19412 15940
rect 18808 13628 19176 13637
rect 18848 13588 18890 13628
rect 18930 13588 18972 13628
rect 19012 13588 19054 13628
rect 19094 13588 19136 13628
rect 18808 13579 19176 13588
rect 19372 13460 19412 15436
rect 19660 15140 19700 15149
rect 19660 14636 19700 15100
rect 19660 14587 19700 14596
rect 19756 14048 19796 16780
rect 19948 16064 19988 16073
rect 19756 13999 19796 14008
rect 19852 14720 19892 14729
rect 19372 13411 19412 13420
rect 19372 13208 19412 13217
rect 18808 12116 19176 12125
rect 18848 12076 18890 12116
rect 18930 12076 18972 12116
rect 19012 12076 19054 12116
rect 19094 12076 19136 12116
rect 18808 12067 19176 12076
rect 18892 11453 18932 11538
rect 18891 11444 18933 11453
rect 18891 11404 18892 11444
rect 18932 11404 18933 11444
rect 18891 11395 18933 11404
rect 18987 11276 19029 11285
rect 18987 11236 18988 11276
rect 19028 11236 19029 11276
rect 18987 11227 19029 11236
rect 18988 11142 19028 11227
rect 18808 10604 19176 10613
rect 18848 10564 18890 10604
rect 18930 10564 18972 10604
rect 19012 10564 19054 10604
rect 19094 10564 19136 10604
rect 18808 10555 19176 10564
rect 19276 9176 19316 9185
rect 18808 9092 19176 9101
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 18808 9043 19176 9052
rect 18808 7580 19176 7589
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 18808 7531 19176 7540
rect 18891 7412 18933 7421
rect 18891 7372 18892 7412
rect 18932 7372 18933 7412
rect 18891 7363 18933 7372
rect 18892 7278 18932 7363
rect 18891 6740 18933 6749
rect 18891 6700 18892 6740
rect 18932 6700 18933 6740
rect 18891 6691 18933 6700
rect 18892 6606 18932 6691
rect 19276 6236 19316 9136
rect 19372 6992 19412 13168
rect 19468 13124 19508 13133
rect 19468 8672 19508 13084
rect 19756 11864 19796 11873
rect 19756 11444 19796 11824
rect 19756 11360 19796 11404
rect 19660 11320 19796 11360
rect 19468 8623 19508 8632
rect 19564 9512 19604 9521
rect 19372 6943 19412 6952
rect 19468 8000 19508 8009
rect 19564 8000 19604 9472
rect 19508 7960 19604 8000
rect 19276 6187 19316 6196
rect 18808 6068 19176 6077
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 18808 6019 19176 6028
rect 19276 5732 19316 5741
rect 18808 4556 19176 4565
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 18808 4507 19176 4516
rect 19276 3548 19316 5692
rect 19468 5648 19508 7960
rect 19660 6488 19700 11320
rect 19756 9428 19796 9437
rect 19756 8840 19796 9388
rect 19756 8791 19796 8800
rect 19660 6439 19700 6448
rect 19756 8672 19796 8681
rect 19468 5599 19508 5608
rect 19564 5984 19604 5993
rect 19276 3499 19316 3508
rect 19372 5480 19412 5489
rect 18700 1457 18740 3172
rect 19372 3380 19412 5440
rect 18808 3044 19176 3053
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 18808 2995 19176 3004
rect 19372 1952 19412 3340
rect 19564 2120 19604 5944
rect 19756 5144 19796 8632
rect 19852 7748 19892 14680
rect 19948 13880 19988 16024
rect 20048 15896 20416 15905
rect 20088 15856 20130 15896
rect 20170 15856 20212 15896
rect 20252 15856 20294 15896
rect 20334 15856 20376 15896
rect 20048 15847 20416 15856
rect 20524 15812 20564 15821
rect 20048 14384 20416 14393
rect 20088 14344 20130 14384
rect 20170 14344 20212 14384
rect 20252 14344 20294 14384
rect 20334 14344 20376 14384
rect 20048 14335 20416 14344
rect 19948 13831 19988 13840
rect 19948 13376 19988 13385
rect 19948 9512 19988 13336
rect 20048 12872 20416 12881
rect 20088 12832 20130 12872
rect 20170 12832 20212 12872
rect 20252 12832 20294 12872
rect 20334 12832 20376 12872
rect 20048 12823 20416 12832
rect 20043 12284 20085 12293
rect 20043 12244 20044 12284
rect 20084 12244 20085 12284
rect 20043 12235 20085 12244
rect 20044 12150 20084 12235
rect 20044 11537 20084 11622
rect 20043 11528 20085 11537
rect 20043 11488 20044 11528
rect 20084 11488 20085 11528
rect 20043 11479 20085 11488
rect 20048 11360 20416 11369
rect 20088 11320 20130 11360
rect 20170 11320 20212 11360
rect 20252 11320 20294 11360
rect 20334 11320 20376 11360
rect 20048 11311 20416 11320
rect 20048 9848 20416 9857
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20048 9799 20416 9808
rect 19948 9463 19988 9472
rect 20044 9680 20084 9689
rect 20044 8504 20084 9640
rect 19948 8464 20084 8504
rect 19948 8168 19988 8464
rect 20048 8336 20416 8345
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20048 8287 20416 8296
rect 19948 8119 19988 8128
rect 19852 7708 19988 7748
rect 19660 4472 19700 4481
rect 19660 2624 19700 4432
rect 19756 3128 19796 5104
rect 19756 3079 19796 3088
rect 19852 7580 19892 7589
rect 19852 6824 19892 7540
rect 19948 7412 19988 7708
rect 19948 7363 19988 7372
rect 19660 2575 19700 2584
rect 19564 2071 19604 2080
rect 19852 2120 19892 6784
rect 20048 6824 20416 6833
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20048 6775 20416 6784
rect 19852 2071 19892 2080
rect 19948 6320 19988 6329
rect 19372 1903 19412 1912
rect 19948 1952 19988 6280
rect 20048 5312 20416 5321
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20048 5263 20416 5272
rect 20048 3800 20416 3809
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20048 3751 20416 3760
rect 20048 2288 20416 2297
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20048 2239 20416 2248
rect 19948 1903 19988 1912
rect 18808 1532 19176 1541
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 18808 1483 19176 1492
rect 18699 1448 18741 1457
rect 18699 1408 18700 1448
rect 18740 1408 18741 1448
rect 18699 1399 18741 1408
rect 18412 1147 18452 1156
rect 18699 860 18741 869
rect 18699 820 18700 860
rect 18740 820 18741 860
rect 18699 811 18741 820
rect 20524 860 20564 15772
rect 20716 10268 20756 29968
rect 21291 29084 21333 29093
rect 21291 29044 21292 29084
rect 21332 29044 21333 29084
rect 21291 29035 21333 29044
rect 21195 20768 21237 20777
rect 21195 20728 21196 20768
rect 21236 20728 21237 20768
rect 21195 20719 21237 20728
rect 20716 10219 20756 10228
rect 20812 19172 20852 19181
rect 20812 10436 20852 19132
rect 20620 10184 20660 10193
rect 20620 4724 20660 10144
rect 20812 7328 20852 10396
rect 20908 17072 20948 17081
rect 20908 8420 20948 17032
rect 21004 15644 21044 15653
rect 21004 11360 21044 15604
rect 21196 14888 21236 20719
rect 21292 16400 21332 29035
rect 21292 16351 21332 16360
rect 21388 15896 21428 30136
rect 21388 15847 21428 15856
rect 21196 14839 21236 14848
rect 21100 11360 21140 11369
rect 21004 11320 21100 11360
rect 20908 8371 20948 8380
rect 21004 10100 21044 10109
rect 20812 7279 20852 7288
rect 20811 6488 20853 6497
rect 20811 6448 20812 6488
rect 20852 6448 20853 6488
rect 20811 6439 20853 6448
rect 20812 6320 20852 6439
rect 20812 6271 20852 6280
rect 20620 4675 20660 4684
rect 21004 2456 21044 10060
rect 21100 4556 21140 11320
rect 21100 4507 21140 4516
rect 21004 2407 21044 2416
rect 20524 811 20564 820
rect 18700 726 18740 811
rect 20048 776 20416 785
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20048 727 20416 736
rect 19275 692 19317 701
rect 19275 652 19276 692
rect 19316 652 19317 692
rect 19275 643 19317 652
rect 19276 558 19316 643
rect 16780 55 16820 64
<< via4 >>
rect 364 39124 404 39164
rect 172 36520 212 36560
rect 172 28288 212 28328
rect 268 22156 308 22196
rect 76 21736 116 21776
rect 652 29632 692 29672
rect 556 21400 596 21440
rect 940 32992 980 33032
rect 748 29044 788 29084
rect 268 12244 308 12284
rect 460 11908 500 11948
rect 652 6196 692 6236
rect 1324 41140 1364 41180
rect 1420 40300 1460 40340
rect 1324 37444 1364 37484
rect 1228 33664 1268 33704
rect 1708 39712 1748 39752
rect 1612 37612 1652 37652
rect 1516 34336 1556 34376
rect 1228 31228 1268 31268
rect 1324 31144 1364 31184
rect 1228 31060 1268 31100
rect 1132 30052 1172 30092
rect 940 5524 980 5564
rect 1036 5356 1076 5396
rect 1036 5104 1076 5144
rect 1612 32992 1652 33032
rect 1516 32068 1556 32108
rect 1516 31816 1556 31856
rect 1420 30724 1460 30764
rect 1228 24592 1268 24632
rect 1228 22408 1268 22448
rect 1420 19804 1460 19844
rect 1228 17788 1268 17828
rect 1324 17704 1364 17744
rect 1324 16192 1364 16232
rect 1612 30724 1652 30764
rect 1612 30556 1652 30596
rect 1804 34084 1844 34124
rect 1804 30556 1844 30596
rect 1612 20812 1652 20852
rect 2092 34084 2132 34124
rect 2092 32908 2132 32948
rect 1996 28960 2036 29000
rect 1900 23752 1940 23792
rect 1516 16192 1556 16232
rect 1516 16024 1556 16064
rect 1420 14680 1460 14720
rect 1228 8128 1268 8168
rect 1228 5188 1268 5228
rect 1228 4684 1268 4724
rect 1612 7036 1652 7076
rect 1516 5776 1556 5816
rect 2380 38284 2420 38324
rect 2188 26188 2228 26228
rect 2380 35176 2420 35216
rect 2380 34336 2420 34376
rect 2380 31816 2420 31856
rect 2476 31648 2516 31688
rect 2284 25348 2324 25388
rect 2476 30808 2516 30848
rect 2476 26356 2516 26396
rect 1804 8716 1844 8756
rect 2092 9388 2132 9428
rect 2380 13840 2420 13880
rect 2380 5692 2420 5732
rect 1228 2416 1268 2456
rect 1420 1660 1460 1700
rect 2764 32488 2804 32528
rect 2668 32404 2708 32444
rect 2668 32068 2708 32108
rect 2668 31648 2708 31688
rect 2956 32404 2996 32444
rect 2668 29128 2708 29168
rect 2668 28960 2708 29000
rect 2764 26524 2804 26564
rect 2668 23920 2708 23960
rect 3340 38116 3380 38156
rect 3052 29044 3092 29084
rect 3688 40804 3728 40844
rect 3770 40804 3810 40844
rect 3852 40804 3892 40844
rect 3934 40804 3974 40844
rect 4016 40804 4056 40844
rect 3628 39796 3668 39836
rect 3688 39292 3728 39332
rect 3770 39292 3810 39332
rect 3852 39292 3892 39332
rect 3934 39292 3974 39332
rect 4016 39292 4056 39332
rect 4396 39712 4436 39752
rect 4300 39460 4340 39500
rect 3688 37780 3728 37820
rect 3770 37780 3810 37820
rect 3852 37780 3892 37820
rect 3934 37780 3974 37820
rect 4016 37780 4056 37820
rect 3724 37528 3764 37568
rect 4108 36520 4148 36560
rect 3688 36268 3728 36308
rect 3770 36268 3810 36308
rect 3852 36268 3892 36308
rect 3934 36268 3974 36308
rect 4016 36268 4056 36308
rect 3340 35344 3380 35384
rect 3340 31312 3380 31352
rect 3052 28876 3092 28916
rect 3148 25852 3188 25892
rect 3688 34756 3728 34796
rect 3770 34756 3810 34796
rect 3852 34756 3892 34796
rect 3934 34756 3974 34796
rect 4016 34756 4056 34796
rect 3628 33496 3668 33536
rect 3688 33244 3728 33284
rect 3770 33244 3810 33284
rect 3852 33244 3892 33284
rect 3934 33244 3974 33284
rect 4016 33244 4056 33284
rect 3532 32656 3572 32696
rect 3532 32488 3572 32528
rect 3532 32320 3572 32360
rect 4492 37696 4532 37736
rect 3688 31732 3728 31772
rect 3770 31732 3810 31772
rect 3852 31732 3892 31772
rect 3934 31732 3974 31772
rect 4016 31732 4056 31772
rect 3436 28372 3476 28412
rect 3340 26524 3380 26564
rect 4108 31060 4148 31100
rect 3688 30220 3728 30260
rect 3770 30220 3810 30260
rect 3852 30220 3892 30260
rect 3934 30220 3974 30260
rect 4016 30220 4056 30260
rect 3688 28708 3728 28748
rect 3770 28708 3810 28748
rect 3852 28708 3892 28748
rect 3934 28708 3974 28748
rect 4016 28708 4056 28748
rect 3688 27196 3728 27236
rect 3770 27196 3810 27236
rect 3852 27196 3892 27236
rect 3934 27196 3974 27236
rect 4016 27196 4056 27236
rect 3724 25936 3764 25976
rect 3628 25852 3668 25892
rect 3688 25684 3728 25724
rect 3770 25684 3810 25724
rect 3852 25684 3892 25724
rect 3934 25684 3974 25724
rect 4016 25684 4056 25724
rect 3688 24172 3728 24212
rect 3770 24172 3810 24212
rect 3852 24172 3892 24212
rect 3934 24172 3974 24212
rect 4016 24172 4056 24212
rect 3724 23920 3764 23960
rect 4492 32908 4532 32948
rect 4684 37696 4724 37736
rect 4684 37444 4724 37484
rect 4928 41560 4968 41600
rect 5010 41560 5050 41600
rect 5092 41560 5132 41600
rect 5174 41560 5214 41600
rect 5256 41560 5296 41600
rect 6700 41140 6740 41180
rect 5644 40468 5684 40508
rect 4928 40048 4968 40088
rect 5010 40048 5050 40088
rect 5092 40048 5132 40088
rect 5174 40048 5214 40088
rect 5256 40048 5296 40088
rect 6028 39796 6068 39836
rect 4928 38536 4968 38576
rect 5010 38536 5050 38576
rect 5092 38536 5132 38576
rect 5174 38536 5214 38576
rect 5256 38536 5296 38576
rect 4876 38032 4916 38072
rect 4928 37024 4968 37064
rect 5010 37024 5050 37064
rect 5092 37024 5132 37064
rect 5174 37024 5214 37064
rect 5256 37024 5296 37064
rect 5260 36520 5300 36560
rect 4684 35344 4724 35384
rect 4204 26776 4244 26816
rect 4204 25936 4244 25976
rect 3688 22660 3728 22700
rect 3770 22660 3810 22700
rect 3852 22660 3892 22700
rect 3934 22660 3974 22700
rect 4016 22660 4056 22700
rect 3436 21484 3476 21524
rect 3340 21232 3380 21272
rect 4204 22324 4244 22364
rect 4204 22156 4244 22196
rect 3916 21736 3956 21776
rect 3628 21568 3668 21608
rect 3628 21316 3668 21356
rect 3688 21148 3728 21188
rect 3770 21148 3810 21188
rect 3852 21148 3892 21188
rect 3934 21148 3974 21188
rect 4016 21148 4056 21188
rect 3532 20728 3572 20768
rect 4204 20392 4244 20432
rect 4492 26356 4532 26396
rect 4928 35512 4968 35552
rect 5010 35512 5050 35552
rect 5092 35512 5132 35552
rect 5174 35512 5214 35552
rect 5256 35512 5296 35552
rect 4928 34000 4968 34040
rect 5010 34000 5050 34040
rect 5092 34000 5132 34040
rect 5174 34000 5214 34040
rect 5256 34000 5296 34040
rect 4928 32488 4968 32528
rect 5010 32488 5050 32528
rect 5092 32488 5132 32528
rect 5174 32488 5214 32528
rect 5256 32488 5296 32528
rect 4928 30976 4968 31016
rect 5010 30976 5050 31016
rect 5092 30976 5132 31016
rect 5174 30976 5214 31016
rect 5256 30976 5296 31016
rect 5356 30136 5396 30176
rect 4928 29464 4968 29504
rect 5010 29464 5050 29504
rect 5092 29464 5132 29504
rect 5174 29464 5214 29504
rect 5256 29464 5296 29504
rect 4928 27952 4968 27992
rect 5010 27952 5050 27992
rect 5092 27952 5132 27992
rect 5174 27952 5214 27992
rect 5256 27952 5296 27992
rect 4492 21568 4532 21608
rect 4396 20560 4436 20600
rect 4928 26440 4968 26480
rect 5010 26440 5050 26480
rect 5092 26440 5132 26480
rect 5174 26440 5214 26480
rect 5256 26440 5296 26480
rect 5356 25684 5396 25724
rect 5548 33748 5588 33788
rect 5548 32740 5588 32780
rect 5548 30136 5588 30176
rect 6028 39208 6068 39248
rect 6124 39124 6164 39164
rect 5740 37108 5780 37148
rect 5932 36772 5972 36812
rect 4928 24928 4968 24968
rect 5010 24928 5050 24968
rect 5092 24928 5132 24968
rect 5174 24928 5214 24968
rect 5256 24928 5296 24968
rect 5356 23752 5396 23792
rect 4928 23416 4968 23456
rect 5010 23416 5050 23456
rect 5092 23416 5132 23456
rect 5174 23416 5214 23456
rect 5256 23416 5296 23456
rect 4928 21904 4968 21944
rect 5010 21904 5050 21944
rect 5092 21904 5132 21944
rect 5174 21904 5214 21944
rect 5256 21904 5296 21944
rect 4396 20392 4436 20432
rect 4204 19804 4244 19844
rect 3688 19636 3728 19676
rect 3770 19636 3810 19676
rect 3852 19636 3892 19676
rect 3934 19636 3974 19676
rect 4016 19636 4056 19676
rect 3688 18124 3728 18164
rect 3770 18124 3810 18164
rect 3852 18124 3892 18164
rect 3934 18124 3974 18164
rect 4016 18124 4056 18164
rect 3688 16612 3728 16652
rect 3770 16612 3810 16652
rect 3852 16612 3892 16652
rect 3934 16612 3974 16652
rect 4016 16612 4056 16652
rect 3052 14764 3092 14804
rect 2860 10984 2900 11024
rect 2668 6280 2708 6320
rect 2668 5524 2708 5564
rect 3148 12832 3188 12872
rect 3148 12580 3188 12620
rect 3148 4096 3188 4136
rect 3688 15100 3728 15140
rect 3770 15100 3810 15140
rect 3852 15100 3892 15140
rect 3934 15100 3974 15140
rect 4016 15100 4056 15140
rect 3820 14092 3860 14132
rect 3688 13588 3728 13628
rect 3770 13588 3810 13628
rect 3852 13588 3892 13628
rect 3934 13588 3974 13628
rect 4016 13588 4056 13628
rect 4300 12832 4340 12872
rect 4780 20560 4820 20600
rect 4928 20392 4968 20432
rect 5010 20392 5050 20432
rect 5092 20392 5132 20432
rect 5174 20392 5214 20432
rect 5256 20392 5296 20432
rect 4928 18880 4968 18920
rect 5010 18880 5050 18920
rect 5092 18880 5132 18920
rect 5174 18880 5214 18920
rect 5256 18880 5296 18920
rect 4928 17368 4968 17408
rect 5010 17368 5050 17408
rect 5092 17368 5132 17408
rect 5174 17368 5214 17408
rect 5256 17368 5296 17408
rect 4928 15856 4968 15896
rect 5010 15856 5050 15896
rect 5092 15856 5132 15896
rect 5174 15856 5214 15896
rect 5256 15856 5296 15896
rect 4928 14344 4968 14384
rect 5010 14344 5050 14384
rect 5092 14344 5132 14384
rect 5174 14344 5214 14384
rect 5256 14344 5296 14384
rect 3688 12076 3728 12116
rect 3770 12076 3810 12116
rect 3852 12076 3892 12116
rect 3934 12076 3974 12116
rect 4016 12076 4056 12116
rect 3724 11656 3764 11696
rect 3532 10984 3572 11024
rect 3436 3424 3476 3464
rect 3688 10564 3728 10604
rect 3770 10564 3810 10604
rect 3852 10564 3892 10604
rect 3934 10564 3974 10604
rect 4016 10564 4056 10604
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 4492 12076 4532 12116
rect 4108 2080 4148 2120
rect 3628 1828 3668 1868
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 3532 1324 3572 1364
rect 3724 1240 3764 1280
rect 4928 12832 4968 12872
rect 5010 12832 5050 12872
rect 5092 12832 5132 12872
rect 5174 12832 5214 12872
rect 5256 12832 5296 12872
rect 5644 26692 5684 26732
rect 5740 25852 5780 25892
rect 5644 25684 5684 25724
rect 5644 22408 5684 22448
rect 5740 21316 5780 21356
rect 6028 35260 6068 35300
rect 6124 35092 6164 35132
rect 6988 40468 7028 40508
rect 6220 31984 6260 32024
rect 5932 31312 5972 31352
rect 6796 38116 6836 38156
rect 6700 35092 6740 35132
rect 6508 34924 6548 34964
rect 6412 31144 6452 31184
rect 6316 26692 6356 26732
rect 6220 25348 6260 25388
rect 6220 22408 6260 22448
rect 6124 21652 6164 21692
rect 6124 21316 6164 21356
rect 5740 17788 5780 17828
rect 4928 11320 4968 11360
rect 5010 11320 5050 11360
rect 5092 11320 5132 11360
rect 5174 11320 5214 11360
rect 5256 11320 5296 11360
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 5452 9976 5492 10016
rect 4972 8632 5012 8672
rect 5356 8632 5396 8672
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 4780 5860 4820 5900
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 5452 7876 5492 7916
rect 5356 4600 5396 4640
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 4684 736 4724 776
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 5068 1324 5108 1364
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 5644 7456 5684 7496
rect 5548 3592 5588 3632
rect 5644 3508 5684 3548
rect 5452 3088 5492 3128
rect 5836 3592 5876 3632
rect 5644 1156 5684 1196
rect 6316 21400 6356 21440
rect 6124 14680 6164 14720
rect 6220 14092 6260 14132
rect 6220 7036 6260 7076
rect 6124 6952 6164 6992
rect 6124 6616 6164 6656
rect 5932 1912 5972 1952
rect 5932 820 5972 860
rect 6316 2248 6356 2288
rect 6316 1324 6356 1364
rect 6604 12076 6644 12116
rect 6508 6868 6548 6908
rect 6700 1240 6740 1280
rect 7084 36100 7124 36140
rect 7372 39712 7412 39752
rect 7276 36688 7316 36728
rect 7180 35260 7220 35300
rect 6892 27700 6932 27740
rect 6892 26860 6932 26900
rect 7372 36016 7412 36056
rect 7276 30052 7316 30092
rect 7180 26860 7220 26900
rect 7180 23752 7220 23792
rect 6988 22660 7028 22700
rect 7084 22324 7124 22364
rect 6988 21484 7028 21524
rect 6892 1828 6932 1868
rect 6604 316 6644 356
rect 7084 3340 7124 3380
rect 7564 33496 7604 33536
rect 7564 32908 7604 32948
rect 7468 22660 7508 22700
rect 7660 22240 7700 22280
rect 7660 21820 7700 21860
rect 7660 21652 7700 21692
rect 7276 6280 7316 6320
rect 7564 17620 7604 17660
rect 7660 15688 7700 15728
rect 7564 12580 7604 12620
rect 7468 11656 7508 11696
rect 7660 6700 7700 6740
rect 7564 3676 7604 3716
rect 7468 2668 7508 2708
rect 8236 40300 8276 40340
rect 8620 38872 8660 38912
rect 7948 37696 7988 37736
rect 8716 38032 8756 38072
rect 8428 37108 8468 37148
rect 8236 36604 8276 36644
rect 8332 36520 8372 36560
rect 7948 32572 7988 32612
rect 7948 28624 7988 28664
rect 7852 6616 7892 6656
rect 7852 2416 7892 2456
rect 8140 32572 8180 32612
rect 8524 36604 8564 36644
rect 8236 22072 8276 22112
rect 8236 21820 8276 21860
rect 8236 15688 8276 15728
rect 8716 36520 8756 36560
rect 8716 33748 8756 33788
rect 8620 26188 8660 26228
rect 8716 22912 8756 22952
rect 8716 21484 8756 21524
rect 8908 37696 8948 37736
rect 9388 36772 9428 36812
rect 9100 36688 9140 36728
rect 9196 34336 9236 34376
rect 9196 34000 9236 34040
rect 9196 32992 9236 33032
rect 9772 36520 9812 36560
rect 9388 36268 9428 36308
rect 9676 35176 9716 35216
rect 9580 32656 9620 32696
rect 9292 32068 9332 32108
rect 8428 3424 8468 3464
rect 8524 1240 8564 1280
rect 8908 16024 8948 16064
rect 8812 9724 8852 9764
rect 8812 8632 8852 8672
rect 8812 8464 8852 8504
rect 8716 8380 8756 8420
rect 8716 7876 8756 7916
rect 8716 7120 8756 7160
rect 8812 3760 8852 3800
rect 9580 25684 9620 25724
rect 9100 14428 9140 14468
rect 9100 8632 9140 8672
rect 9196 8380 9236 8420
rect 9004 3508 9044 3548
rect 9484 14428 9524 14468
rect 9484 9724 9524 9764
rect 9388 8548 9428 8588
rect 9580 8632 9620 8672
rect 9484 8464 9524 8504
rect 9484 8296 9524 8336
rect 9676 6952 9716 6992
rect 9292 2080 9332 2120
rect 10348 38872 10388 38912
rect 10060 34168 10100 34208
rect 10060 29632 10100 29672
rect 9964 29212 10004 29252
rect 9964 26776 10004 26816
rect 10252 24508 10292 24548
rect 9964 13168 10004 13208
rect 10732 39208 10772 39248
rect 10540 31984 10580 32024
rect 10444 26440 10484 26480
rect 10540 24508 10580 24548
rect 10636 22072 10676 22112
rect 9964 9892 10004 9932
rect 9868 3760 9908 3800
rect 10444 13420 10484 13460
rect 10444 13168 10484 13208
rect 10156 4600 10196 4640
rect 10252 4264 10292 4304
rect 10636 4264 10676 4304
rect 10636 3676 10676 3716
rect 10828 36520 10868 36560
rect 10924 32740 10964 32780
rect 10828 28960 10868 29000
rect 10828 12076 10868 12116
rect 11212 35092 11252 35132
rect 11116 29212 11156 29252
rect 11116 20812 11156 20852
rect 11308 28624 11348 28664
rect 11404 26440 11444 26480
rect 11308 12244 11348 12284
rect 11308 12076 11348 12116
rect 11116 3340 11156 3380
rect 10732 2332 10772 2372
rect 11404 11908 11444 11948
rect 11404 11740 11444 11780
rect 11596 25180 11636 25220
rect 12268 31480 12308 31520
rect 11788 13840 11828 13880
rect 11596 11740 11636 11780
rect 11404 5860 11444 5900
rect 268 148 308 188
rect 5260 148 5300 188
rect 10156 820 10196 860
rect 12076 21484 12116 21524
rect 11788 9388 11828 9428
rect 13708 40468 13748 40508
rect 12748 39460 12788 39500
rect 12748 37192 12788 37232
rect 13132 37612 13172 37652
rect 13132 37444 13172 37484
rect 13036 35428 13076 35468
rect 12652 27616 12692 27656
rect 13324 33580 13364 33620
rect 13516 35008 13556 35048
rect 13516 33580 13556 33620
rect 13420 32320 13460 32360
rect 13228 31228 13268 31268
rect 13324 31144 13364 31184
rect 12172 8128 12212 8168
rect 11980 3088 12020 3128
rect 11884 2668 11924 2708
rect 12652 11236 12692 11276
rect 12556 9892 12596 9932
rect 12460 3172 12500 3212
rect 12652 7036 12692 7076
rect 13132 10144 13172 10184
rect 13036 6280 13076 6320
rect 12844 5020 12884 5060
rect 13228 8128 13268 8168
rect 13132 5776 13172 5816
rect 12748 1240 12788 1280
rect 13612 28624 13652 28664
rect 13612 15352 13652 15392
rect 13612 15100 13652 15140
rect 13612 14680 13652 14720
rect 13324 4684 13364 4724
rect 13228 1996 13268 2036
rect 13612 10144 13652 10184
rect 13612 9976 13652 10016
rect 13612 8128 13652 8168
rect 12364 1072 12404 1112
rect 13996 37444 14036 37484
rect 13804 35092 13844 35132
rect 13804 32404 13844 32444
rect 14188 35176 14228 35216
rect 14380 39712 14420 39752
rect 13996 14848 14036 14888
rect 13900 8716 13940 8756
rect 14092 7456 14132 7496
rect 13900 5020 13940 5060
rect 13804 4936 13844 4976
rect 14668 39460 14708 39500
rect 14188 5692 14228 5732
rect 13996 2248 14036 2288
rect 14284 904 14324 944
rect 14572 11488 14612 11528
rect 14572 6112 14612 6152
rect 14572 3004 14612 3044
rect 14572 2332 14612 2372
rect 15148 40720 15188 40760
rect 15148 39376 15188 39416
rect 15148 36772 15188 36812
rect 15436 37612 15476 37652
rect 15340 35344 15380 35384
rect 14956 13420 14996 13460
rect 14380 652 14420 692
rect 16588 40468 16628 40508
rect 15628 35260 15668 35300
rect 15820 36436 15860 36476
rect 15724 35092 15764 35132
rect 15724 34000 15764 34040
rect 15244 28372 15284 28412
rect 15436 11404 15476 11444
rect 15436 10900 15476 10940
rect 15340 8296 15380 8336
rect 15244 6448 15284 6488
rect 15532 7288 15572 7328
rect 15436 5608 15476 5648
rect 15436 1660 15476 1700
rect 15916 32320 15956 32360
rect 15724 25936 15764 25976
rect 15724 7288 15764 7328
rect 15724 6700 15764 6740
rect 16012 12244 16052 12284
rect 16012 10900 16052 10940
rect 16396 36772 16436 36812
rect 16204 36436 16244 36476
rect 16300 35260 16340 35300
rect 16204 35008 16244 35048
rect 16300 34924 16340 34964
rect 16492 33916 16532 33956
rect 16684 32908 16724 32948
rect 16876 39712 16916 39752
rect 16300 22912 16340 22952
rect 16588 29212 16628 29252
rect 16876 31228 16916 31268
rect 16588 26692 16628 26732
rect 16684 25684 16724 25724
rect 16492 15940 16532 15980
rect 16492 15100 16532 15140
rect 16876 24592 16916 24632
rect 17548 40972 17588 41012
rect 17644 40636 17684 40676
rect 17260 35176 17300 35216
rect 17356 35092 17396 35132
rect 17452 31228 17492 31268
rect 17260 24592 17300 24632
rect 16780 20392 16820 20432
rect 16972 20392 17012 20432
rect 17164 22240 17204 22280
rect 17068 15940 17108 15980
rect 16972 15772 17012 15812
rect 16300 7372 16340 7412
rect 11500 148 11540 188
rect 6028 64 6068 104
rect 10060 64 10100 104
rect 17068 3172 17108 3212
rect 17452 26692 17492 26732
rect 17452 15772 17492 15812
rect 17644 33916 17684 33956
rect 17932 40720 17972 40760
rect 17932 40300 17972 40340
rect 17836 35596 17876 35636
rect 17644 25180 17684 25220
rect 18220 35596 18260 35636
rect 18124 28288 18164 28328
rect 18028 27616 18068 27656
rect 17932 24676 17972 24716
rect 18220 23920 18260 23960
rect 17836 4936 17876 4976
rect 20048 41560 20088 41600
rect 20130 41560 20170 41600
rect 20212 41560 20252 41600
rect 20294 41560 20334 41600
rect 20376 41560 20416 41600
rect 18412 39460 18452 39500
rect 18412 37696 18452 37736
rect 18508 32068 18548 32108
rect 18412 30808 18452 30848
rect 18808 40804 18848 40844
rect 18890 40804 18930 40844
rect 18972 40804 19012 40844
rect 19054 40804 19094 40844
rect 19136 40804 19176 40844
rect 18892 40636 18932 40676
rect 18808 39292 18848 39332
rect 18890 39292 18930 39332
rect 18972 39292 19012 39332
rect 19054 39292 19094 39332
rect 19136 39292 19176 39332
rect 18808 37780 18848 37820
rect 18890 37780 18930 37820
rect 18972 37780 19012 37820
rect 19054 37780 19094 37820
rect 19136 37780 19176 37820
rect 18808 36268 18848 36308
rect 18890 36268 18930 36308
rect 18972 36268 19012 36308
rect 19054 36268 19094 36308
rect 19136 36268 19176 36308
rect 18808 34756 18848 34796
rect 18890 34756 18930 34796
rect 18972 34756 19012 34796
rect 19054 34756 19094 34796
rect 19136 34756 19176 34796
rect 18808 33244 18848 33284
rect 18890 33244 18930 33284
rect 18972 33244 19012 33284
rect 19054 33244 19094 33284
rect 19136 33244 19176 33284
rect 18808 31732 18848 31772
rect 18890 31732 18930 31772
rect 18972 31732 19012 31772
rect 19054 31732 19094 31772
rect 19136 31732 19176 31772
rect 18796 30808 18836 30848
rect 18808 30220 18848 30260
rect 18890 30220 18930 30260
rect 18972 30220 19012 30260
rect 19054 30220 19094 30260
rect 19136 30220 19176 30260
rect 18808 28708 18848 28748
rect 18890 28708 18930 28748
rect 18972 28708 19012 28748
rect 19054 28708 19094 28748
rect 19136 28708 19176 28748
rect 18808 27196 18848 27236
rect 18890 27196 18930 27236
rect 18972 27196 19012 27236
rect 19054 27196 19094 27236
rect 19136 27196 19176 27236
rect 18808 25684 18848 25724
rect 18890 25684 18930 25724
rect 18972 25684 19012 25724
rect 19054 25684 19094 25724
rect 19136 25684 19176 25724
rect 18604 25180 18644 25220
rect 18604 24676 18644 24716
rect 18808 24172 18848 24212
rect 18890 24172 18930 24212
rect 18972 24172 19012 24212
rect 19054 24172 19094 24212
rect 19136 24172 19176 24212
rect 18808 22660 18848 22700
rect 18890 22660 18930 22700
rect 18972 22660 19012 22700
rect 19054 22660 19094 22700
rect 19136 22660 19176 22700
rect 18808 21148 18848 21188
rect 18890 21148 18930 21188
rect 18972 21148 19012 21188
rect 19054 21148 19094 21188
rect 19136 21148 19176 21188
rect 18808 19636 18848 19676
rect 18890 19636 18930 19676
rect 18972 19636 19012 19676
rect 19054 19636 19094 19676
rect 19136 19636 19176 19676
rect 18808 18124 18848 18164
rect 18890 18124 18930 18164
rect 18972 18124 19012 18164
rect 19054 18124 19094 18164
rect 19136 18124 19176 18164
rect 18808 16612 18848 16652
rect 18890 16612 18930 16652
rect 18972 16612 19012 16652
rect 19054 16612 19094 16652
rect 19136 16612 19176 16652
rect 18808 15100 18848 15140
rect 18890 15100 18930 15140
rect 18972 15100 19012 15140
rect 19054 15100 19094 15140
rect 19136 15100 19176 15140
rect 18316 9976 18356 10016
rect 18508 4096 18548 4136
rect 20048 40048 20088 40088
rect 20130 40048 20170 40088
rect 20212 40048 20252 40088
rect 20294 40048 20334 40088
rect 20376 40048 20416 40088
rect 20048 38536 20088 38576
rect 20130 38536 20170 38576
rect 20212 38536 20252 38576
rect 20294 38536 20334 38576
rect 20376 38536 20416 38576
rect 20048 37024 20088 37064
rect 20130 37024 20170 37064
rect 20212 37024 20252 37064
rect 20294 37024 20334 37064
rect 20376 37024 20416 37064
rect 20812 37192 20852 37232
rect 20716 36100 20756 36140
rect 20048 35512 20088 35552
rect 20130 35512 20170 35552
rect 20212 35512 20252 35552
rect 20294 35512 20334 35552
rect 20376 35512 20416 35552
rect 20048 34000 20088 34040
rect 20130 34000 20170 34040
rect 20212 34000 20252 34040
rect 20294 34000 20334 34040
rect 20376 34000 20416 34040
rect 19852 33580 19892 33620
rect 20048 32488 20088 32528
rect 20130 32488 20170 32528
rect 20212 32488 20252 32528
rect 20294 32488 20334 32528
rect 20376 32488 20416 32528
rect 20048 30976 20088 31016
rect 20130 30976 20170 31016
rect 20212 30976 20252 31016
rect 20294 30976 20334 31016
rect 20376 30976 20416 31016
rect 20048 29464 20088 29504
rect 20130 29464 20170 29504
rect 20212 29464 20252 29504
rect 20294 29464 20334 29504
rect 20376 29464 20416 29504
rect 20048 27952 20088 27992
rect 20130 27952 20170 27992
rect 20212 27952 20252 27992
rect 20294 27952 20334 27992
rect 20376 27952 20416 27992
rect 20048 26440 20088 26480
rect 20130 26440 20170 26480
rect 20212 26440 20252 26480
rect 20294 26440 20334 26480
rect 20376 26440 20416 26480
rect 20048 24928 20088 24968
rect 20130 24928 20170 24968
rect 20212 24928 20252 24968
rect 20294 24928 20334 24968
rect 20376 24928 20416 24968
rect 20812 36016 20852 36056
rect 21196 36520 21236 36560
rect 20048 23416 20088 23456
rect 20130 23416 20170 23456
rect 20212 23416 20252 23456
rect 20294 23416 20334 23456
rect 20376 23416 20416 23456
rect 20048 21904 20088 21944
rect 20130 21904 20170 21944
rect 20212 21904 20252 21944
rect 20294 21904 20334 21944
rect 20376 21904 20416 21944
rect 20048 20392 20088 20432
rect 20130 20392 20170 20432
rect 20212 20392 20252 20432
rect 20294 20392 20334 20432
rect 20376 20392 20416 20432
rect 20048 18880 20088 18920
rect 20130 18880 20170 18920
rect 20212 18880 20252 18920
rect 20294 18880 20334 18920
rect 20376 18880 20416 18920
rect 20048 17368 20088 17408
rect 20130 17368 20170 17408
rect 20212 17368 20252 17408
rect 20294 17368 20334 17408
rect 20376 17368 20416 17408
rect 18808 13588 18848 13628
rect 18890 13588 18930 13628
rect 18972 13588 19012 13628
rect 19054 13588 19094 13628
rect 19136 13588 19176 13628
rect 18808 12076 18848 12116
rect 18890 12076 18930 12116
rect 18972 12076 19012 12116
rect 19054 12076 19094 12116
rect 19136 12076 19176 12116
rect 18892 11404 18932 11444
rect 18988 11236 19028 11276
rect 18808 10564 18848 10604
rect 18890 10564 18930 10604
rect 18972 10564 19012 10604
rect 19054 10564 19094 10604
rect 19136 10564 19176 10604
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 18892 7372 18932 7412
rect 18892 6700 18932 6740
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 20048 15856 20088 15896
rect 20130 15856 20170 15896
rect 20212 15856 20252 15896
rect 20294 15856 20334 15896
rect 20376 15856 20416 15896
rect 20048 14344 20088 14384
rect 20130 14344 20170 14384
rect 20212 14344 20252 14384
rect 20294 14344 20334 14384
rect 20376 14344 20416 14384
rect 20048 12832 20088 12872
rect 20130 12832 20170 12872
rect 20212 12832 20252 12872
rect 20294 12832 20334 12872
rect 20376 12832 20416 12872
rect 20044 12244 20084 12284
rect 20044 11488 20084 11528
rect 20048 11320 20088 11360
rect 20130 11320 20170 11360
rect 20212 11320 20252 11360
rect 20294 11320 20334 11360
rect 20376 11320 20416 11360
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 18700 1408 18740 1448
rect 18700 820 18740 860
rect 21292 29044 21332 29084
rect 21196 20728 21236 20768
rect 20812 6448 20852 6488
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 19276 652 19316 692
<< metal5 >>
rect 4919 41623 5305 41642
rect 4919 41600 4985 41623
rect 5071 41600 5153 41623
rect 5239 41600 5305 41623
rect 4919 41560 4928 41600
rect 4968 41560 4985 41600
rect 5071 41560 5092 41600
rect 5132 41560 5153 41600
rect 5239 41560 5256 41600
rect 5296 41560 5305 41600
rect 4919 41537 4985 41560
rect 5071 41537 5153 41560
rect 5239 41537 5305 41560
rect 4919 41518 5305 41537
rect 20039 41623 20425 41642
rect 20039 41600 20105 41623
rect 20191 41600 20273 41623
rect 20359 41600 20425 41623
rect 20039 41560 20048 41600
rect 20088 41560 20105 41600
rect 20191 41560 20212 41600
rect 20252 41560 20273 41600
rect 20359 41560 20376 41600
rect 20416 41560 20425 41600
rect 20039 41537 20105 41560
rect 20191 41537 20273 41560
rect 20359 41537 20425 41560
rect 20039 41518 20425 41537
rect 1315 41140 1324 41180
rect 1364 41140 6700 41180
rect 6740 41140 6749 41180
rect 17138 41035 17262 41054
rect 17138 40949 17157 41035
rect 17243 41012 17262 41035
rect 17243 40972 17548 41012
rect 17588 40972 17597 41012
rect 17243 40949 17262 40972
rect 17138 40930 17262 40949
rect 3679 40867 4065 40886
rect 3679 40844 3745 40867
rect 3831 40844 3913 40867
rect 3999 40844 4065 40867
rect 3679 40804 3688 40844
rect 3728 40804 3745 40844
rect 3831 40804 3852 40844
rect 3892 40804 3913 40844
rect 3999 40804 4016 40844
rect 4056 40804 4065 40844
rect 3679 40781 3745 40804
rect 3831 40781 3913 40804
rect 3999 40781 4065 40804
rect 3679 40762 4065 40781
rect 18799 40867 19185 40886
rect 18799 40844 18865 40867
rect 18951 40844 19033 40867
rect 19119 40844 19185 40867
rect 18799 40804 18808 40844
rect 18848 40804 18865 40844
rect 18951 40804 18972 40844
rect 19012 40804 19033 40844
rect 19119 40804 19136 40844
rect 19176 40804 19185 40844
rect 18799 40781 18865 40804
rect 18951 40781 19033 40804
rect 19119 40781 19185 40804
rect 18799 40762 19185 40781
rect 15139 40720 15148 40760
rect 15188 40720 17932 40760
rect 17972 40720 17981 40760
rect 17635 40636 17644 40676
rect 17684 40636 18892 40676
rect 18932 40636 18941 40676
rect 5635 40468 5644 40508
rect 5684 40468 6988 40508
rect 7028 40468 7037 40508
rect 13699 40468 13708 40508
rect 13748 40468 16588 40508
rect 16628 40468 16637 40508
rect 14402 40363 14526 40382
rect 1411 40300 1420 40340
rect 1460 40300 8236 40340
rect 8276 40300 8285 40340
rect 14402 40277 14421 40363
rect 14507 40340 14526 40363
rect 14507 40300 17932 40340
rect 17972 40300 17981 40340
rect 14507 40277 14526 40300
rect 14402 40258 14526 40277
rect 4919 40111 5305 40130
rect 4919 40088 4985 40111
rect 5071 40088 5153 40111
rect 5239 40088 5305 40111
rect 4919 40048 4928 40088
rect 4968 40048 4985 40088
rect 5071 40048 5092 40088
rect 5132 40048 5153 40088
rect 5239 40048 5256 40088
rect 5296 40048 5305 40088
rect 4919 40025 4985 40048
rect 5071 40025 5153 40048
rect 5239 40025 5305 40048
rect 4919 40006 5305 40025
rect 20039 40111 20425 40130
rect 20039 40088 20105 40111
rect 20191 40088 20273 40111
rect 20359 40088 20425 40111
rect 20039 40048 20048 40088
rect 20088 40048 20105 40088
rect 20191 40048 20212 40088
rect 20252 40048 20273 40088
rect 20359 40048 20376 40088
rect 20416 40048 20425 40088
rect 20039 40025 20105 40048
rect 20191 40025 20273 40048
rect 20359 40025 20425 40048
rect 20039 40006 20425 40025
rect 3619 39796 3628 39836
rect 3668 39796 6028 39836
rect 6068 39796 6077 39836
rect 1699 39712 1708 39752
rect 1748 39712 4396 39752
rect 4436 39712 7372 39752
rect 7412 39712 7421 39752
rect 14371 39712 14380 39752
rect 14420 39712 16876 39752
rect 16916 39712 16925 39752
rect 4291 39460 4300 39500
rect 4340 39460 12748 39500
rect 12788 39460 12797 39500
rect 14659 39460 14668 39500
rect 14708 39460 18412 39500
rect 18452 39460 18461 39500
rect 13490 39439 13614 39458
rect 3679 39355 4065 39374
rect 3679 39332 3745 39355
rect 3831 39332 3913 39355
rect 3999 39332 4065 39355
rect 13490 39353 13509 39439
rect 13595 39416 13614 39439
rect 13595 39376 15148 39416
rect 15188 39376 15197 39416
rect 13595 39353 13614 39376
rect 13490 39334 13614 39353
rect 18799 39355 19185 39374
rect 3679 39292 3688 39332
rect 3728 39292 3745 39332
rect 3831 39292 3852 39332
rect 3892 39292 3913 39332
rect 3999 39292 4016 39332
rect 4056 39292 4065 39332
rect 3679 39269 3745 39292
rect 3831 39269 3913 39292
rect 3999 39269 4065 39292
rect 3679 39250 4065 39269
rect 18799 39332 18865 39355
rect 18951 39332 19033 39355
rect 19119 39332 19185 39355
rect 18799 39292 18808 39332
rect 18848 39292 18865 39332
rect 18951 39292 18972 39332
rect 19012 39292 19033 39332
rect 19119 39292 19136 39332
rect 19176 39292 19185 39332
rect 18799 39269 18865 39292
rect 18951 39269 19033 39292
rect 19119 39269 19185 39292
rect 18799 39250 19185 39269
rect 6019 39208 6028 39248
rect 6068 39208 10732 39248
rect 10772 39208 10781 39248
rect 355 39124 364 39164
rect 404 39124 6124 39164
rect 6164 39124 6173 39164
rect 8611 38872 8620 38912
rect 8660 38872 10348 38912
rect 10388 38872 10397 38912
rect 4919 38599 5305 38618
rect 4919 38576 4985 38599
rect 5071 38576 5153 38599
rect 5239 38576 5305 38599
rect 4919 38536 4928 38576
rect 4968 38536 4985 38576
rect 5071 38536 5092 38576
rect 5132 38536 5153 38576
rect 5239 38536 5256 38576
rect 5296 38536 5305 38576
rect 4919 38513 4985 38536
rect 5071 38513 5153 38536
rect 5239 38513 5305 38536
rect 4919 38494 5305 38513
rect 20039 38599 20425 38618
rect 20039 38576 20105 38599
rect 20191 38576 20273 38599
rect 20359 38576 20425 38599
rect 20039 38536 20048 38576
rect 20088 38536 20105 38576
rect 20191 38536 20212 38576
rect 20252 38536 20273 38576
rect 20359 38536 20376 38576
rect 20416 38536 20425 38576
rect 20039 38513 20105 38536
rect 20191 38513 20273 38536
rect 20359 38513 20425 38536
rect 20039 38494 20425 38513
rect 7106 38347 7230 38366
rect 7106 38324 7125 38347
rect 2371 38284 2380 38324
rect 2420 38284 7125 38324
rect 7106 38261 7125 38284
rect 7211 38261 7230 38347
rect 7106 38242 7230 38261
rect 3331 38116 3340 38156
rect 3380 38116 6796 38156
rect 6836 38116 6845 38156
rect 4867 38032 4876 38072
rect 4916 38032 8716 38072
rect 8756 38032 8765 38072
rect 3679 37843 4065 37862
rect 3679 37820 3745 37843
rect 3831 37820 3913 37843
rect 3999 37820 4065 37843
rect 3679 37780 3688 37820
rect 3728 37780 3745 37820
rect 3831 37780 3852 37820
rect 3892 37780 3913 37820
rect 3999 37780 4016 37820
rect 4056 37780 4065 37820
rect 3679 37757 3745 37780
rect 3831 37757 3913 37780
rect 3999 37757 4065 37780
rect 3679 37738 4065 37757
rect 18799 37843 19185 37862
rect 18799 37820 18865 37843
rect 18951 37820 19033 37843
rect 19119 37820 19185 37843
rect 18799 37780 18808 37820
rect 18848 37780 18865 37820
rect 18951 37780 18972 37820
rect 19012 37780 19033 37820
rect 19119 37780 19136 37820
rect 19176 37780 19185 37820
rect 18799 37757 18865 37780
rect 18951 37757 19033 37780
rect 19119 37757 19185 37780
rect 18799 37738 19185 37757
rect 4483 37696 4492 37736
rect 4532 37696 4684 37736
rect 4724 37696 7948 37736
rect 7988 37696 7997 37736
rect 8899 37696 8908 37736
rect 8948 37696 18412 37736
rect 18452 37696 18461 37736
rect 1603 37612 1612 37652
rect 1652 37612 13132 37652
rect 13172 37612 13181 37652
rect 13532 37612 15436 37652
rect 15476 37612 15485 37652
rect 13532 37568 13572 37612
rect 3715 37528 3724 37568
rect 3764 37528 13572 37568
rect 1315 37444 1324 37484
rect 1364 37444 4684 37484
rect 4724 37444 4733 37484
rect 13123 37444 13132 37484
rect 13172 37444 13996 37484
rect 14036 37444 14045 37484
rect 12739 37192 12748 37232
rect 12788 37192 20812 37232
rect 20852 37192 20861 37232
rect 5731 37108 5740 37148
rect 5780 37108 8428 37148
rect 8468 37108 8477 37148
rect 4919 37087 5305 37106
rect 4919 37064 4985 37087
rect 5071 37064 5153 37087
rect 5239 37064 5305 37087
rect 4919 37024 4928 37064
rect 4968 37024 4985 37064
rect 5071 37024 5092 37064
rect 5132 37024 5153 37064
rect 5239 37024 5256 37064
rect 5296 37024 5305 37064
rect 4919 37001 4985 37024
rect 5071 37001 5153 37024
rect 5239 37001 5305 37024
rect 4919 36982 5305 37001
rect 20039 37087 20425 37106
rect 20039 37064 20105 37087
rect 20191 37064 20273 37087
rect 20359 37064 20425 37087
rect 20039 37024 20048 37064
rect 20088 37024 20105 37064
rect 20191 37024 20212 37064
rect 20252 37024 20273 37064
rect 20359 37024 20376 37064
rect 20416 37024 20425 37064
rect 20039 37001 20105 37024
rect 20191 37001 20273 37024
rect 20359 37001 20425 37024
rect 20039 36982 20425 37001
rect 5923 36772 5932 36812
rect 5972 36772 9388 36812
rect 9428 36772 9437 36812
rect 15139 36772 15148 36812
rect 15188 36772 16396 36812
rect 16436 36772 16445 36812
rect 7267 36688 7276 36728
rect 7316 36688 9100 36728
rect 9140 36688 9149 36728
rect 8227 36604 8236 36644
rect 8276 36604 8524 36644
rect 8564 36604 8573 36644
rect 163 36520 172 36560
rect 212 36520 4108 36560
rect 4148 36520 4157 36560
rect 5251 36520 5260 36560
rect 5300 36520 8332 36560
rect 8372 36520 8381 36560
rect 8707 36520 8716 36560
rect 8756 36520 9772 36560
rect 9812 36520 9821 36560
rect 10819 36520 10828 36560
rect 10868 36520 21196 36560
rect 21236 36520 21245 36560
rect 15811 36436 15820 36476
rect 15860 36436 16204 36476
rect 16244 36436 16253 36476
rect 3679 36331 4065 36350
rect 3679 36308 3745 36331
rect 3831 36308 3913 36331
rect 3999 36308 4065 36331
rect 9386 36331 9510 36350
rect 9386 36308 9405 36331
rect 3679 36268 3688 36308
rect 3728 36268 3745 36308
rect 3831 36268 3852 36308
rect 3892 36268 3913 36308
rect 3999 36268 4016 36308
rect 4056 36268 4065 36308
rect 9379 36268 9388 36308
rect 3679 36245 3745 36268
rect 3831 36245 3913 36268
rect 3999 36245 4065 36268
rect 3679 36226 4065 36245
rect 9386 36245 9405 36268
rect 9491 36245 9510 36331
rect 9386 36226 9510 36245
rect 18799 36331 19185 36350
rect 18799 36308 18865 36331
rect 18951 36308 19033 36331
rect 19119 36308 19185 36331
rect 18799 36268 18808 36308
rect 18848 36268 18865 36308
rect 18951 36268 18972 36308
rect 19012 36268 19033 36308
rect 19119 36268 19136 36308
rect 19176 36268 19185 36308
rect 18799 36245 18865 36268
rect 18951 36245 19033 36268
rect 19119 36245 19185 36268
rect 18799 36226 19185 36245
rect 7075 36100 7084 36140
rect 7124 36100 20716 36140
rect 20756 36100 20765 36140
rect 7363 36016 7372 36056
rect 7412 36016 20812 36056
rect 20852 36016 20861 36056
rect 17827 35596 17836 35636
rect 17876 35596 18220 35636
rect 18260 35596 18269 35636
rect 4919 35575 5305 35594
rect 4919 35552 4985 35575
rect 5071 35552 5153 35575
rect 5239 35552 5305 35575
rect 4919 35512 4928 35552
rect 4968 35512 4985 35552
rect 5071 35512 5092 35552
rect 5132 35512 5153 35552
rect 5239 35512 5256 35552
rect 5296 35512 5305 35552
rect 4919 35489 4985 35512
rect 5071 35489 5153 35512
rect 5239 35489 5305 35512
rect 20039 35575 20425 35594
rect 20039 35552 20105 35575
rect 20191 35552 20273 35575
rect 20359 35552 20425 35575
rect 20039 35512 20048 35552
rect 20088 35512 20105 35552
rect 20191 35512 20212 35552
rect 20252 35512 20273 35552
rect 20359 35512 20376 35552
rect 20416 35512 20425 35552
rect 4919 35470 5305 35489
rect 15770 35491 15894 35510
rect 15770 35468 15789 35491
rect 13027 35428 13036 35468
rect 13076 35428 15789 35468
rect 15770 35405 15789 35428
rect 15875 35405 15894 35491
rect 20039 35489 20105 35512
rect 20191 35489 20273 35512
rect 20359 35489 20425 35512
rect 20039 35470 20425 35489
rect 15770 35386 15894 35405
rect 3331 35344 3340 35384
rect 3380 35344 4684 35384
rect 4724 35344 15340 35384
rect 15380 35344 15389 35384
rect 1178 35323 1302 35342
rect 1178 35237 1197 35323
rect 1283 35300 1302 35323
rect 1283 35260 6028 35300
rect 6068 35260 6077 35300
rect 7171 35260 7180 35300
rect 7220 35260 15628 35300
rect 15668 35260 16300 35300
rect 16340 35260 16349 35300
rect 1283 35237 1302 35260
rect 1178 35218 1302 35237
rect 2371 35176 2380 35216
rect 2420 35176 9676 35216
rect 9716 35176 9725 35216
rect 11320 35176 14188 35216
rect 14228 35176 17260 35216
rect 17300 35176 17309 35216
rect 11320 35132 11360 35176
rect 6115 35092 6124 35132
rect 6164 35092 6700 35132
rect 6740 35092 11212 35132
rect 11252 35092 11360 35132
rect 13795 35092 13804 35132
rect 13844 35092 15724 35132
rect 15764 35092 17356 35132
rect 17396 35092 17405 35132
rect 13507 35008 13516 35048
rect 13556 35008 16204 35048
rect 16244 35008 16253 35048
rect 6499 34924 6508 34964
rect 6548 34924 16300 34964
rect 16340 34924 16349 34964
rect 3679 34819 4065 34838
rect 3679 34796 3745 34819
rect 3831 34796 3913 34819
rect 3999 34796 4065 34819
rect 3679 34756 3688 34796
rect 3728 34756 3745 34796
rect 3831 34756 3852 34796
rect 3892 34756 3913 34796
rect 3999 34756 4016 34796
rect 4056 34756 4065 34796
rect 3679 34733 3745 34756
rect 3831 34733 3913 34756
rect 3999 34733 4065 34756
rect 3679 34714 4065 34733
rect 18799 34819 19185 34838
rect 18799 34796 18865 34819
rect 18951 34796 19033 34819
rect 19119 34796 19185 34819
rect 18799 34756 18808 34796
rect 18848 34756 18865 34796
rect 18951 34756 18972 34796
rect 19012 34756 19033 34796
rect 19119 34756 19136 34796
rect 19176 34756 19185 34796
rect 18799 34733 18865 34756
rect 18951 34733 19033 34756
rect 19119 34733 19185 34756
rect 18799 34714 19185 34733
rect 1507 34336 1516 34376
rect 1556 34336 2380 34376
rect 2420 34336 9196 34376
rect 9236 34336 9245 34376
rect 2500 34168 10060 34208
rect 10100 34168 10109 34208
rect 2500 34124 2540 34168
rect 1795 34084 1804 34124
rect 1844 34084 2092 34124
rect 2132 34084 2540 34124
rect 4919 34063 5305 34082
rect 4919 34040 4985 34063
rect 5071 34040 5153 34063
rect 5239 34040 5305 34063
rect 20039 34063 20425 34082
rect 20039 34040 20105 34063
rect 20191 34040 20273 34063
rect 20359 34040 20425 34063
rect 4919 34000 4928 34040
rect 4968 34000 4985 34040
rect 5071 34000 5092 34040
rect 5132 34000 5153 34040
rect 5239 34000 5256 34040
rect 5296 34000 5305 34040
rect 9187 34000 9196 34040
rect 9236 34000 15724 34040
rect 15764 34000 15773 34040
rect 20039 34000 20048 34040
rect 20088 34000 20105 34040
rect 20191 34000 20212 34040
rect 20252 34000 20273 34040
rect 20359 34000 20376 34040
rect 20416 34000 20425 34040
rect 4919 33977 4985 34000
rect 5071 33977 5153 34000
rect 5239 33977 5305 34000
rect 4919 33958 5305 33977
rect 20039 33977 20105 34000
rect 20191 33977 20273 34000
rect 20359 33977 20425 34000
rect 20039 33958 20425 33977
rect 16483 33916 16492 33956
rect 16532 33916 17644 33956
rect 17684 33916 17693 33956
rect 2500 33748 5548 33788
rect 5588 33748 8716 33788
rect 8756 33748 8765 33788
rect 2500 33704 2540 33748
rect 1219 33664 1228 33704
rect 1268 33664 2540 33704
rect 13315 33580 13324 33620
rect 13364 33580 13516 33620
rect 13556 33580 19852 33620
rect 19892 33580 19901 33620
rect 3619 33496 3628 33536
rect 3668 33496 7564 33536
rect 7604 33496 7613 33536
rect 3679 33307 4065 33326
rect 3679 33284 3745 33307
rect 3831 33284 3913 33307
rect 3999 33284 4065 33307
rect 3679 33244 3688 33284
rect 3728 33244 3745 33284
rect 3831 33244 3852 33284
rect 3892 33244 3913 33284
rect 3999 33244 4016 33284
rect 4056 33244 4065 33284
rect 3679 33221 3745 33244
rect 3831 33221 3913 33244
rect 3999 33221 4065 33244
rect 3679 33202 4065 33221
rect 18799 33307 19185 33326
rect 18799 33284 18865 33307
rect 18951 33284 19033 33307
rect 19119 33284 19185 33307
rect 18799 33244 18808 33284
rect 18848 33244 18865 33284
rect 18951 33244 18972 33284
rect 19012 33244 19033 33284
rect 19119 33244 19136 33284
rect 19176 33244 19185 33284
rect 18799 33221 18865 33244
rect 18951 33221 19033 33244
rect 19119 33221 19185 33244
rect 18799 33202 19185 33221
rect 931 32992 940 33032
rect 980 32992 1612 33032
rect 1652 32992 9196 33032
rect 9236 32992 9245 33032
rect 2083 32908 2092 32948
rect 2132 32908 4492 32948
rect 4532 32908 7564 32948
rect 7604 32908 7613 32948
rect 11320 32908 16684 32948
rect 16724 32908 16733 32948
rect 11320 32780 11360 32908
rect 5539 32740 5548 32780
rect 5588 32740 10924 32780
rect 10964 32740 11360 32780
rect 3523 32656 3532 32696
rect 3572 32656 9580 32696
rect 9620 32656 9629 32696
rect 7939 32572 7948 32612
rect 7988 32572 8140 32612
rect 8180 32572 8189 32612
rect 4919 32551 5305 32570
rect 4919 32528 4985 32551
rect 5071 32528 5153 32551
rect 5239 32528 5305 32551
rect 2755 32488 2764 32528
rect 2804 32488 3532 32528
rect 3572 32488 3581 32528
rect 4919 32488 4928 32528
rect 4968 32488 4985 32528
rect 5071 32488 5092 32528
rect 5132 32488 5153 32528
rect 5239 32488 5256 32528
rect 5296 32488 5305 32528
rect 4919 32465 4985 32488
rect 5071 32465 5153 32488
rect 5239 32465 5305 32488
rect 4919 32446 5305 32465
rect 20039 32551 20425 32570
rect 20039 32528 20105 32551
rect 20191 32528 20273 32551
rect 20359 32528 20425 32551
rect 20039 32488 20048 32528
rect 20088 32488 20105 32528
rect 20191 32488 20212 32528
rect 20252 32488 20273 32528
rect 20359 32488 20376 32528
rect 20416 32488 20425 32528
rect 20039 32465 20105 32488
rect 20191 32465 20273 32488
rect 20359 32465 20425 32488
rect 20039 32446 20425 32465
rect 2659 32404 2668 32444
rect 2708 32404 2956 32444
rect 2996 32404 3005 32444
rect 11320 32404 13804 32444
rect 13844 32404 13853 32444
rect 11320 32360 11360 32404
rect 3523 32320 3532 32360
rect 3572 32320 11360 32360
rect 13411 32320 13420 32360
rect 13460 32320 15916 32360
rect 15956 32320 15965 32360
rect 1507 32068 1516 32108
rect 1556 32068 2540 32108
rect 2659 32068 2668 32108
rect 2708 32068 9292 32108
rect 9332 32068 18508 32108
rect 18548 32068 18557 32108
rect 2500 32024 2540 32068
rect 2500 31984 6220 32024
rect 6260 31984 10540 32024
rect 10580 31984 10589 32024
rect 1507 31816 1516 31856
rect 1556 31816 2380 31856
rect 2420 31816 2429 31856
rect 3679 31795 4065 31814
rect 3679 31772 3745 31795
rect 3831 31772 3913 31795
rect 3999 31772 4065 31795
rect 3679 31732 3688 31772
rect 3728 31732 3745 31772
rect 3831 31732 3852 31772
rect 3892 31732 3913 31772
rect 3999 31732 4016 31772
rect 4056 31732 4065 31772
rect 3679 31709 3745 31732
rect 3831 31709 3913 31732
rect 3999 31709 4065 31732
rect 3679 31690 4065 31709
rect 18799 31795 19185 31814
rect 18799 31772 18865 31795
rect 18951 31772 19033 31795
rect 19119 31772 19185 31795
rect 18799 31732 18808 31772
rect 18848 31732 18865 31772
rect 18951 31732 18972 31772
rect 19012 31732 19033 31772
rect 19119 31732 19136 31772
rect 19176 31732 19185 31772
rect 18799 31709 18865 31732
rect 18951 31709 19033 31732
rect 19119 31709 19185 31732
rect 18799 31690 19185 31709
rect 2467 31648 2476 31688
rect 2516 31648 2668 31688
rect 2708 31648 2717 31688
rect 12164 31480 12268 31520
rect 12308 31480 12317 31520
rect 12164 31394 12204 31480
rect 12122 31375 12246 31394
rect 3331 31312 3340 31352
rect 3380 31312 5932 31352
rect 5972 31312 5981 31352
rect 12122 31289 12141 31375
rect 12227 31289 12246 31375
rect 12122 31270 12246 31289
rect 1219 31228 1228 31268
rect 1268 31228 11360 31268
rect 13219 31228 13228 31268
rect 13268 31228 16876 31268
rect 16916 31228 17452 31268
rect 17492 31228 17501 31268
rect 11320 31184 11360 31228
rect 1315 31144 1324 31184
rect 1364 31144 6412 31184
rect 6452 31144 6732 31184
rect 11320 31144 13324 31184
rect 13364 31144 13373 31184
rect 6692 31100 6732 31144
rect 10298 31123 10422 31142
rect 10298 31100 10317 31123
rect 1219 31060 1228 31100
rect 1268 31060 4108 31100
rect 4148 31060 4157 31100
rect 6692 31060 10317 31100
rect 4919 31039 5305 31058
rect 4919 31016 4985 31039
rect 5071 31016 5153 31039
rect 5239 31016 5305 31039
rect 10298 31037 10317 31060
rect 10403 31037 10422 31123
rect 10298 31018 10422 31037
rect 20039 31039 20425 31058
rect 4919 30976 4928 31016
rect 4968 30976 4985 31016
rect 5071 30976 5092 31016
rect 5132 30976 5153 31016
rect 5239 30976 5256 31016
rect 5296 30976 5305 31016
rect 4919 30953 4985 30976
rect 5071 30953 5153 30976
rect 5239 30953 5305 30976
rect 4919 30934 5305 30953
rect 20039 31016 20105 31039
rect 20191 31016 20273 31039
rect 20359 31016 20425 31039
rect 20039 30976 20048 31016
rect 20088 30976 20105 31016
rect 20191 30976 20212 31016
rect 20252 30976 20273 31016
rect 20359 30976 20376 31016
rect 20416 30976 20425 31016
rect 20039 30953 20105 30976
rect 20191 30953 20273 30976
rect 20359 30953 20425 30976
rect 20039 30934 20425 30953
rect 2467 30808 2476 30848
rect 2516 30808 18412 30848
rect 18452 30808 18796 30848
rect 18836 30808 18845 30848
rect 1411 30724 1420 30764
rect 1460 30724 1612 30764
rect 1652 30724 1661 30764
rect 1603 30556 1612 30596
rect 1652 30556 1804 30596
rect 1844 30556 1853 30596
rect 3679 30283 4065 30302
rect 3679 30260 3745 30283
rect 3831 30260 3913 30283
rect 3999 30260 4065 30283
rect 3679 30220 3688 30260
rect 3728 30220 3745 30260
rect 3831 30220 3852 30260
rect 3892 30220 3913 30260
rect 3999 30220 4016 30260
rect 4056 30220 4065 30260
rect 3679 30197 3745 30220
rect 3831 30197 3913 30220
rect 3999 30197 4065 30220
rect 3679 30178 4065 30197
rect 18799 30283 19185 30302
rect 18799 30260 18865 30283
rect 18951 30260 19033 30283
rect 19119 30260 19185 30283
rect 18799 30220 18808 30260
rect 18848 30220 18865 30260
rect 18951 30220 18972 30260
rect 19012 30220 19033 30260
rect 19119 30220 19136 30260
rect 19176 30220 19185 30260
rect 18799 30197 18865 30220
rect 18951 30197 19033 30220
rect 19119 30197 19185 30220
rect 18799 30178 19185 30197
rect 5347 30136 5356 30176
rect 5396 30136 5548 30176
rect 5588 30136 5597 30176
rect 1123 30052 1132 30092
rect 1172 30052 7276 30092
rect 7316 30052 7325 30092
rect 643 29632 652 29672
rect 692 29632 10060 29672
rect 10100 29632 10109 29672
rect 4919 29527 5305 29546
rect 4919 29504 4985 29527
rect 5071 29504 5153 29527
rect 5239 29504 5305 29527
rect 4919 29464 4928 29504
rect 4968 29464 4985 29504
rect 5071 29464 5092 29504
rect 5132 29464 5153 29504
rect 5239 29464 5256 29504
rect 5296 29464 5305 29504
rect 4919 29441 4985 29464
rect 5071 29441 5153 29464
rect 5239 29441 5305 29464
rect 4919 29422 5305 29441
rect 20039 29527 20425 29546
rect 20039 29504 20105 29527
rect 20191 29504 20273 29527
rect 20359 29504 20425 29527
rect 20039 29464 20048 29504
rect 20088 29464 20105 29504
rect 20191 29464 20212 29504
rect 20252 29464 20273 29504
rect 20359 29464 20376 29504
rect 20416 29464 20425 29504
rect 20039 29441 20105 29464
rect 20191 29441 20273 29464
rect 20359 29441 20425 29464
rect 20039 29422 20425 29441
rect 9955 29212 9964 29252
rect 10004 29212 11116 29252
rect 11156 29212 16588 29252
rect 16628 29212 16637 29252
rect 2659 29128 2668 29168
rect 2708 29128 11360 29168
rect 11320 29084 11360 29128
rect 739 29044 748 29084
rect 788 29044 3052 29084
rect 3092 29044 3101 29084
rect 11320 29044 21292 29084
rect 21332 29044 21341 29084
rect 1987 28960 1996 29000
rect 2036 28960 2668 29000
rect 2708 28960 2717 29000
rect 10796 28960 10828 29000
rect 10868 28960 10877 29000
rect 10796 28916 10836 28960
rect 3043 28876 3052 28916
rect 3092 28876 10836 28916
rect 3679 28771 4065 28790
rect 3679 28748 3745 28771
rect 3831 28748 3913 28771
rect 3999 28748 4065 28771
rect 3679 28708 3688 28748
rect 3728 28708 3745 28748
rect 3831 28708 3852 28748
rect 3892 28708 3913 28748
rect 3999 28708 4016 28748
rect 4056 28708 4065 28748
rect 3679 28685 3745 28708
rect 3831 28685 3913 28708
rect 3999 28685 4065 28708
rect 3679 28666 4065 28685
rect 18799 28771 19185 28790
rect 18799 28748 18865 28771
rect 18951 28748 19033 28771
rect 19119 28748 19185 28771
rect 18799 28708 18808 28748
rect 18848 28708 18865 28748
rect 18951 28708 18972 28748
rect 19012 28708 19033 28748
rect 19119 28708 19136 28748
rect 19176 28708 19185 28748
rect 18799 28685 18865 28708
rect 18951 28685 19033 28708
rect 19119 28685 19185 28708
rect 18799 28666 19185 28685
rect 7939 28624 7948 28664
rect 7988 28624 11308 28664
rect 11348 28624 13612 28664
rect 13652 28624 13661 28664
rect 3427 28372 3436 28412
rect 3476 28372 15244 28412
rect 15284 28372 15293 28412
rect 163 28288 172 28328
rect 212 28288 18124 28328
rect 18164 28288 18173 28328
rect 4919 28015 5305 28034
rect 4919 27992 4985 28015
rect 5071 27992 5153 28015
rect 5239 27992 5305 28015
rect 4919 27952 4928 27992
rect 4968 27952 4985 27992
rect 5071 27952 5092 27992
rect 5132 27952 5153 27992
rect 5239 27952 5256 27992
rect 5296 27952 5305 27992
rect 4919 27929 4985 27952
rect 5071 27929 5153 27952
rect 5239 27929 5305 27952
rect 4919 27910 5305 27929
rect 20039 28015 20425 28034
rect 20039 27992 20105 28015
rect 20191 27992 20273 28015
rect 20359 27992 20425 28015
rect 20039 27952 20048 27992
rect 20088 27952 20105 27992
rect 20191 27952 20212 27992
rect 20252 27952 20273 27992
rect 20359 27952 20376 27992
rect 20416 27952 20425 27992
rect 20039 27929 20105 27952
rect 20191 27929 20273 27952
rect 20359 27929 20425 27952
rect 20039 27910 20425 27929
rect 2090 27763 2214 27782
rect 2090 27677 2109 27763
rect 2195 27740 2214 27763
rect 2195 27700 6892 27740
rect 6932 27700 6941 27740
rect 2195 27677 2214 27700
rect 2090 27658 2214 27677
rect 12643 27616 12652 27656
rect 12692 27616 18028 27656
rect 18068 27616 18077 27656
rect 3679 27259 4065 27278
rect 3679 27236 3745 27259
rect 3831 27236 3913 27259
rect 3999 27236 4065 27259
rect 3679 27196 3688 27236
rect 3728 27196 3745 27236
rect 3831 27196 3852 27236
rect 3892 27196 3913 27236
rect 3999 27196 4016 27236
rect 4056 27196 4065 27236
rect 3679 27173 3745 27196
rect 3831 27173 3913 27196
rect 3999 27173 4065 27196
rect 3679 27154 4065 27173
rect 18799 27259 19185 27278
rect 18799 27236 18865 27259
rect 18951 27236 19033 27259
rect 19119 27236 19185 27259
rect 18799 27196 18808 27236
rect 18848 27196 18865 27236
rect 18951 27196 18972 27236
rect 19012 27196 19033 27236
rect 19119 27196 19136 27236
rect 19176 27196 19185 27236
rect 18799 27173 18865 27196
rect 18951 27173 19033 27196
rect 19119 27173 19185 27196
rect 18799 27154 19185 27173
rect 6883 26860 6892 26900
rect 6932 26860 7180 26900
rect 7220 26860 7229 26900
rect 4195 26776 4204 26816
rect 4244 26776 9964 26816
rect 10004 26776 11360 26816
rect 11320 26732 11360 26776
rect 5635 26692 5644 26732
rect 5684 26692 6316 26732
rect 6356 26692 6365 26732
rect 11320 26692 16588 26732
rect 16628 26692 17452 26732
rect 17492 26692 17501 26732
rect 2755 26524 2764 26564
rect 2804 26524 3340 26564
rect 3380 26524 3389 26564
rect 4919 26503 5305 26522
rect 4919 26480 4985 26503
rect 5071 26480 5153 26503
rect 5239 26480 5305 26503
rect 20039 26503 20425 26522
rect 20039 26480 20105 26503
rect 20191 26480 20273 26503
rect 20359 26480 20425 26503
rect 4919 26440 4928 26480
rect 4968 26440 4985 26480
rect 5071 26440 5092 26480
rect 5132 26440 5153 26480
rect 5239 26440 5256 26480
rect 5296 26440 5305 26480
rect 10435 26440 10444 26480
rect 10484 26440 11404 26480
rect 11444 26440 11453 26480
rect 20039 26440 20048 26480
rect 20088 26440 20105 26480
rect 20191 26440 20212 26480
rect 20252 26440 20273 26480
rect 20359 26440 20376 26480
rect 20416 26440 20425 26480
rect 4919 26417 4985 26440
rect 5071 26417 5153 26440
rect 5239 26417 5305 26440
rect 4919 26398 5305 26417
rect 20039 26417 20105 26440
rect 20191 26417 20273 26440
rect 20359 26417 20425 26440
rect 20039 26398 20425 26417
rect 2467 26356 2476 26396
rect 2516 26356 4492 26396
rect 4532 26356 4541 26396
rect 2179 26188 2188 26228
rect 2228 26188 8620 26228
rect 8660 26188 8669 26228
rect 3532 25936 3724 25976
rect 3764 25936 3773 25976
rect 4195 25936 4204 25976
rect 4244 25936 15724 25976
rect 15764 25936 15773 25976
rect 3532 25892 3572 25936
rect 3139 25852 3148 25892
rect 3188 25852 3572 25892
rect 3619 25852 3628 25892
rect 3668 25852 5740 25892
rect 5780 25852 5789 25892
rect 3679 25747 4065 25766
rect 3679 25724 3745 25747
rect 3831 25724 3913 25747
rect 3999 25724 4065 25747
rect 18799 25747 19185 25766
rect 18799 25724 18865 25747
rect 18951 25724 19033 25747
rect 19119 25724 19185 25747
rect 3679 25684 3688 25724
rect 3728 25684 3745 25724
rect 3831 25684 3852 25724
rect 3892 25684 3913 25724
rect 3999 25684 4016 25724
rect 4056 25684 4065 25724
rect 5347 25684 5356 25724
rect 5396 25684 5644 25724
rect 5684 25684 5693 25724
rect 9571 25684 9580 25724
rect 9620 25684 16684 25724
rect 16724 25684 16733 25724
rect 18799 25684 18808 25724
rect 18848 25684 18865 25724
rect 18951 25684 18972 25724
rect 19012 25684 19033 25724
rect 19119 25684 19136 25724
rect 19176 25684 19185 25724
rect 3679 25661 3745 25684
rect 3831 25661 3913 25684
rect 3999 25661 4065 25684
rect 3679 25642 4065 25661
rect 18799 25661 18865 25684
rect 18951 25661 19033 25684
rect 19119 25661 19185 25684
rect 18799 25642 19185 25661
rect 2275 25348 2284 25388
rect 2324 25348 6220 25388
rect 6260 25348 6269 25388
rect 11587 25180 11596 25220
rect 11636 25180 17644 25220
rect 17684 25180 18604 25220
rect 18644 25180 18653 25220
rect 4919 24991 5305 25010
rect 4919 24968 4985 24991
rect 5071 24968 5153 24991
rect 5239 24968 5305 24991
rect 4919 24928 4928 24968
rect 4968 24928 4985 24968
rect 5071 24928 5092 24968
rect 5132 24928 5153 24968
rect 5239 24928 5256 24968
rect 5296 24928 5305 24968
rect 4919 24905 4985 24928
rect 5071 24905 5153 24928
rect 5239 24905 5305 24928
rect 4919 24886 5305 24905
rect 20039 24991 20425 25010
rect 20039 24968 20105 24991
rect 20191 24968 20273 24991
rect 20359 24968 20425 24991
rect 20039 24928 20048 24968
rect 20088 24928 20105 24968
rect 20191 24928 20212 24968
rect 20252 24928 20273 24968
rect 20359 24928 20376 24968
rect 20416 24928 20425 24968
rect 20039 24905 20105 24928
rect 20191 24905 20273 24928
rect 20359 24905 20425 24928
rect 20039 24886 20425 24905
rect 2500 24676 17932 24716
rect 17972 24676 18604 24716
rect 18644 24676 18653 24716
rect 2500 24632 2540 24676
rect 1219 24592 1228 24632
rect 1268 24592 2540 24632
rect 16867 24592 16876 24632
rect 16916 24592 17260 24632
rect 17300 24592 17309 24632
rect 10243 24508 10252 24548
rect 10292 24508 10540 24548
rect 10580 24508 10589 24548
rect 3679 24235 4065 24254
rect 3679 24212 3745 24235
rect 3831 24212 3913 24235
rect 3999 24212 4065 24235
rect 3679 24172 3688 24212
rect 3728 24172 3745 24212
rect 3831 24172 3852 24212
rect 3892 24172 3913 24212
rect 3999 24172 4016 24212
rect 4056 24172 4065 24212
rect 3679 24149 3745 24172
rect 3831 24149 3913 24172
rect 3999 24149 4065 24172
rect 3679 24130 4065 24149
rect 18799 24235 19185 24254
rect 18799 24212 18865 24235
rect 18951 24212 19033 24235
rect 19119 24212 19185 24235
rect 18799 24172 18808 24212
rect 18848 24172 18865 24212
rect 18951 24172 18972 24212
rect 19012 24172 19033 24212
rect 19119 24172 19136 24212
rect 19176 24172 19185 24212
rect 18799 24149 18865 24172
rect 18951 24149 19033 24172
rect 19119 24149 19185 24172
rect 18799 24130 19185 24149
rect 2659 23920 2668 23960
rect 2708 23920 3724 23960
rect 3764 23920 18220 23960
rect 18260 23920 18269 23960
rect 1891 23752 1900 23792
rect 1940 23752 5356 23792
rect 5396 23752 7180 23792
rect 7220 23752 7229 23792
rect 4919 23479 5305 23498
rect 4919 23456 4985 23479
rect 5071 23456 5153 23479
rect 5239 23456 5305 23479
rect 4919 23416 4928 23456
rect 4968 23416 4985 23456
rect 5071 23416 5092 23456
rect 5132 23416 5153 23456
rect 5239 23416 5256 23456
rect 5296 23416 5305 23456
rect 4919 23393 4985 23416
rect 5071 23393 5153 23416
rect 5239 23393 5305 23416
rect 4919 23374 5305 23393
rect 20039 23479 20425 23498
rect 20039 23456 20105 23479
rect 20191 23456 20273 23479
rect 20359 23456 20425 23479
rect 20039 23416 20048 23456
rect 20088 23416 20105 23456
rect 20191 23416 20212 23456
rect 20252 23416 20273 23456
rect 20359 23416 20376 23456
rect 20416 23416 20425 23456
rect 20039 23393 20105 23416
rect 20191 23393 20273 23416
rect 20359 23393 20425 23416
rect 20039 23374 20425 23393
rect 8707 22912 8716 22952
rect 8756 22912 16300 22952
rect 16340 22912 16349 22952
rect 3679 22723 4065 22742
rect 3679 22700 3745 22723
rect 3831 22700 3913 22723
rect 3999 22700 4065 22723
rect 18799 22723 19185 22742
rect 18799 22700 18865 22723
rect 18951 22700 19033 22723
rect 19119 22700 19185 22723
rect 3679 22660 3688 22700
rect 3728 22660 3745 22700
rect 3831 22660 3852 22700
rect 3892 22660 3913 22700
rect 3999 22660 4016 22700
rect 4056 22660 4065 22700
rect 6979 22660 6988 22700
rect 7028 22660 7468 22700
rect 7508 22660 7517 22700
rect 18799 22660 18808 22700
rect 18848 22660 18865 22700
rect 18951 22660 18972 22700
rect 19012 22660 19033 22700
rect 19119 22660 19136 22700
rect 19176 22660 19185 22700
rect 3679 22637 3745 22660
rect 3831 22637 3913 22660
rect 3999 22637 4065 22660
rect 3679 22618 4065 22637
rect 18799 22637 18865 22660
rect 18951 22637 19033 22660
rect 19119 22637 19185 22660
rect 18799 22618 19185 22637
rect 1219 22408 1228 22448
rect 1268 22408 5644 22448
rect 5684 22408 6220 22448
rect 6260 22408 6269 22448
rect 4195 22324 4204 22364
rect 4244 22324 7084 22364
rect 7124 22324 7133 22364
rect 7651 22240 7660 22280
rect 7700 22240 17164 22280
rect 17204 22240 17213 22280
rect 259 22156 268 22196
rect 308 22156 4204 22196
rect 4244 22156 4253 22196
rect 8227 22072 8236 22112
rect 8276 22072 10636 22112
rect 10676 22072 10685 22112
rect 4919 21967 5305 21986
rect 4919 21944 4985 21967
rect 5071 21944 5153 21967
rect 5239 21944 5305 21967
rect 4919 21904 4928 21944
rect 4968 21904 4985 21944
rect 5071 21904 5092 21944
rect 5132 21904 5153 21944
rect 5239 21904 5256 21944
rect 5296 21904 5305 21944
rect 4919 21881 4985 21904
rect 5071 21881 5153 21904
rect 5239 21881 5305 21904
rect 4919 21862 5305 21881
rect 20039 21967 20425 21986
rect 20039 21944 20105 21967
rect 20191 21944 20273 21967
rect 20359 21944 20425 21967
rect 20039 21904 20048 21944
rect 20088 21904 20105 21944
rect 20191 21904 20212 21944
rect 20252 21904 20273 21944
rect 20359 21904 20376 21944
rect 20416 21904 20425 21944
rect 20039 21881 20105 21904
rect 20191 21881 20273 21904
rect 20359 21881 20425 21904
rect 20039 21862 20425 21881
rect 7651 21820 7660 21860
rect 7700 21820 8236 21860
rect 8276 21820 8285 21860
rect 67 21736 76 21776
rect 116 21736 3916 21776
rect 3956 21736 3965 21776
rect 6115 21652 6124 21692
rect 6164 21652 7660 21692
rect 7700 21652 7709 21692
rect 3619 21568 3628 21608
rect 3668 21568 4492 21608
rect 4532 21568 4541 21608
rect 3427 21484 3436 21524
rect 3476 21484 6988 21524
rect 7028 21484 7037 21524
rect 8707 21484 8716 21524
rect 8756 21484 12076 21524
rect 12116 21484 12125 21524
rect 8474 21463 8598 21482
rect 8474 21440 8493 21463
rect 547 21400 556 21440
rect 596 21400 6316 21440
rect 6356 21400 8493 21440
rect 8474 21377 8493 21400
rect 8579 21377 8598 21463
rect 8474 21358 8598 21377
rect 3500 21316 3628 21356
rect 3668 21316 3677 21356
rect 5731 21316 5740 21356
rect 5780 21316 6124 21356
rect 6164 21316 6173 21356
rect 3500 21272 3540 21316
rect 3331 21232 3340 21272
rect 3380 21232 3540 21272
rect 3679 21211 4065 21230
rect 3679 21188 3745 21211
rect 3831 21188 3913 21211
rect 3999 21188 4065 21211
rect 3679 21148 3688 21188
rect 3728 21148 3745 21188
rect 3831 21148 3852 21188
rect 3892 21148 3913 21188
rect 3999 21148 4016 21188
rect 4056 21148 4065 21188
rect 3679 21125 3745 21148
rect 3831 21125 3913 21148
rect 3999 21125 4065 21148
rect 3679 21106 4065 21125
rect 18799 21211 19185 21230
rect 18799 21188 18865 21211
rect 18951 21188 19033 21211
rect 19119 21188 19185 21211
rect 18799 21148 18808 21188
rect 18848 21148 18865 21188
rect 18951 21148 18972 21188
rect 19012 21148 19033 21188
rect 19119 21148 19136 21188
rect 19176 21148 19185 21188
rect 18799 21125 18865 21148
rect 18951 21125 19033 21148
rect 19119 21125 19185 21148
rect 18799 21106 19185 21125
rect 1603 20812 1612 20852
rect 1652 20812 11116 20852
rect 11156 20812 11165 20852
rect 3523 20728 3532 20768
rect 3572 20728 21196 20768
rect 21236 20728 21245 20768
rect 4387 20560 4396 20600
rect 4436 20560 4780 20600
rect 4820 20560 4829 20600
rect 4919 20455 5305 20474
rect 4919 20432 4985 20455
rect 5071 20432 5153 20455
rect 5239 20432 5305 20455
rect 20039 20455 20425 20474
rect 20039 20432 20105 20455
rect 20191 20432 20273 20455
rect 20359 20432 20425 20455
rect 4195 20392 4204 20432
rect 4244 20392 4396 20432
rect 4436 20392 4445 20432
rect 4919 20392 4928 20432
rect 4968 20392 4985 20432
rect 5071 20392 5092 20432
rect 5132 20392 5153 20432
rect 5239 20392 5256 20432
rect 5296 20392 5305 20432
rect 16771 20392 16780 20432
rect 16820 20392 16972 20432
rect 17012 20392 17021 20432
rect 20039 20392 20048 20432
rect 20088 20392 20105 20432
rect 20191 20392 20212 20432
rect 20252 20392 20273 20432
rect 20359 20392 20376 20432
rect 20416 20392 20425 20432
rect 4919 20369 4985 20392
rect 5071 20369 5153 20392
rect 5239 20369 5305 20392
rect 4919 20350 5305 20369
rect 20039 20369 20105 20392
rect 20191 20369 20273 20392
rect 20359 20369 20425 20392
rect 20039 20350 20425 20369
rect 1411 19804 1420 19844
rect 1460 19804 4204 19844
rect 4244 19804 4253 19844
rect 3679 19699 4065 19718
rect 3679 19676 3745 19699
rect 3831 19676 3913 19699
rect 3999 19676 4065 19699
rect 3679 19636 3688 19676
rect 3728 19636 3745 19676
rect 3831 19636 3852 19676
rect 3892 19636 3913 19676
rect 3999 19636 4016 19676
rect 4056 19636 4065 19676
rect 3679 19613 3745 19636
rect 3831 19613 3913 19636
rect 3999 19613 4065 19636
rect 3679 19594 4065 19613
rect 18799 19699 19185 19718
rect 18799 19676 18865 19699
rect 18951 19676 19033 19699
rect 19119 19676 19185 19699
rect 18799 19636 18808 19676
rect 18848 19636 18865 19676
rect 18951 19636 18972 19676
rect 19012 19636 19033 19676
rect 19119 19636 19136 19676
rect 19176 19636 19185 19676
rect 18799 19613 18865 19636
rect 18951 19613 19033 19636
rect 19119 19613 19185 19636
rect 18799 19594 19185 19613
rect 4919 18943 5305 18962
rect 4919 18920 4985 18943
rect 5071 18920 5153 18943
rect 5239 18920 5305 18943
rect 4919 18880 4928 18920
rect 4968 18880 4985 18920
rect 5071 18880 5092 18920
rect 5132 18880 5153 18920
rect 5239 18880 5256 18920
rect 5296 18880 5305 18920
rect 4919 18857 4985 18880
rect 5071 18857 5153 18880
rect 5239 18857 5305 18880
rect 4919 18838 5305 18857
rect 20039 18943 20425 18962
rect 20039 18920 20105 18943
rect 20191 18920 20273 18943
rect 20359 18920 20425 18943
rect 20039 18880 20048 18920
rect 20088 18880 20105 18920
rect 20191 18880 20212 18920
rect 20252 18880 20273 18920
rect 20359 18880 20376 18920
rect 20416 18880 20425 18920
rect 20039 18857 20105 18880
rect 20191 18857 20273 18880
rect 20359 18857 20425 18880
rect 20039 18838 20425 18857
rect 3679 18187 4065 18206
rect 3679 18164 3745 18187
rect 3831 18164 3913 18187
rect 3999 18164 4065 18187
rect 3679 18124 3688 18164
rect 3728 18124 3745 18164
rect 3831 18124 3852 18164
rect 3892 18124 3913 18164
rect 3999 18124 4016 18164
rect 4056 18124 4065 18164
rect 3679 18101 3745 18124
rect 3831 18101 3913 18124
rect 3999 18101 4065 18124
rect 3679 18082 4065 18101
rect 18799 18187 19185 18206
rect 18799 18164 18865 18187
rect 18951 18164 19033 18187
rect 19119 18164 19185 18187
rect 18799 18124 18808 18164
rect 18848 18124 18865 18164
rect 18951 18124 18972 18164
rect 19012 18124 19033 18164
rect 19119 18124 19136 18164
rect 19176 18124 19185 18164
rect 18799 18101 18865 18124
rect 18951 18101 19033 18124
rect 19119 18101 19185 18124
rect 18799 18082 19185 18101
rect 1219 17788 1228 17828
rect 1268 17788 5740 17828
rect 5780 17788 5789 17828
rect 1315 17704 1324 17744
rect 1364 17704 2540 17744
rect 2500 17660 2540 17704
rect 2500 17620 7564 17660
rect 7604 17620 7613 17660
rect 4919 17431 5305 17450
rect 4919 17408 4985 17431
rect 5071 17408 5153 17431
rect 5239 17408 5305 17431
rect 4919 17368 4928 17408
rect 4968 17368 4985 17408
rect 5071 17368 5092 17408
rect 5132 17368 5153 17408
rect 5239 17368 5256 17408
rect 5296 17368 5305 17408
rect 4919 17345 4985 17368
rect 5071 17345 5153 17368
rect 5239 17345 5305 17368
rect 4919 17326 5305 17345
rect 20039 17431 20425 17450
rect 20039 17408 20105 17431
rect 20191 17408 20273 17431
rect 20359 17408 20425 17431
rect 20039 17368 20048 17408
rect 20088 17368 20105 17408
rect 20191 17368 20212 17408
rect 20252 17368 20273 17408
rect 20359 17368 20376 17408
rect 20416 17368 20425 17408
rect 20039 17345 20105 17368
rect 20191 17345 20273 17368
rect 20359 17345 20425 17368
rect 20039 17326 20425 17345
rect 3679 16675 4065 16694
rect 3679 16652 3745 16675
rect 3831 16652 3913 16675
rect 3999 16652 4065 16675
rect 3679 16612 3688 16652
rect 3728 16612 3745 16652
rect 3831 16612 3852 16652
rect 3892 16612 3913 16652
rect 3999 16612 4016 16652
rect 4056 16612 4065 16652
rect 3679 16589 3745 16612
rect 3831 16589 3913 16612
rect 3999 16589 4065 16612
rect 3679 16570 4065 16589
rect 18799 16675 19185 16694
rect 18799 16652 18865 16675
rect 18951 16652 19033 16675
rect 19119 16652 19185 16675
rect 18799 16612 18808 16652
rect 18848 16612 18865 16652
rect 18951 16612 18972 16652
rect 19012 16612 19033 16652
rect 19119 16612 19136 16652
rect 19176 16612 19185 16652
rect 18799 16589 18865 16612
rect 18951 16589 19033 16612
rect 19119 16589 19185 16612
rect 18799 16570 19185 16589
rect 1315 16192 1324 16232
rect 1364 16192 1516 16232
rect 1556 16192 1565 16232
rect 1507 16024 1516 16064
rect 1556 16024 8908 16064
rect 8948 16024 8957 16064
rect 16483 15940 16492 15980
rect 16532 15940 17068 15980
rect 17108 15940 17117 15980
rect 4919 15919 5305 15938
rect 4919 15896 4985 15919
rect 5071 15896 5153 15919
rect 5239 15896 5305 15919
rect 4919 15856 4928 15896
rect 4968 15856 4985 15896
rect 5071 15856 5092 15896
rect 5132 15856 5153 15896
rect 5239 15856 5256 15896
rect 5296 15856 5305 15896
rect 4919 15833 4985 15856
rect 5071 15833 5153 15856
rect 5239 15833 5305 15856
rect 4919 15814 5305 15833
rect 20039 15919 20425 15938
rect 20039 15896 20105 15919
rect 20191 15896 20273 15919
rect 20359 15896 20425 15919
rect 20039 15856 20048 15896
rect 20088 15856 20105 15896
rect 20191 15856 20212 15896
rect 20252 15856 20273 15896
rect 20359 15856 20376 15896
rect 20416 15856 20425 15896
rect 20039 15833 20105 15856
rect 20191 15833 20273 15856
rect 20359 15833 20425 15856
rect 20039 15814 20425 15833
rect 16963 15772 16972 15812
rect 17012 15772 17452 15812
rect 17492 15772 17501 15812
rect 7651 15688 7660 15728
rect 7700 15688 8236 15728
rect 8276 15688 8285 15728
rect 13490 15415 13614 15434
rect 13490 15329 13509 15415
rect 13595 15392 13614 15415
rect 13595 15352 13612 15392
rect 13652 15352 13661 15392
rect 13595 15329 13614 15352
rect 13490 15310 13614 15329
rect 3679 15163 4065 15182
rect 3679 15140 3745 15163
rect 3831 15140 3913 15163
rect 3999 15140 4065 15163
rect 18799 15163 19185 15182
rect 18799 15140 18865 15163
rect 18951 15140 19033 15163
rect 19119 15140 19185 15163
rect 3679 15100 3688 15140
rect 3728 15100 3745 15140
rect 3831 15100 3852 15140
rect 3892 15100 3913 15140
rect 3999 15100 4016 15140
rect 4056 15100 4065 15140
rect 13603 15100 13612 15140
rect 13652 15100 16492 15140
rect 16532 15100 16541 15140
rect 18799 15100 18808 15140
rect 18848 15100 18865 15140
rect 18951 15100 18972 15140
rect 19012 15100 19033 15140
rect 19119 15100 19136 15140
rect 19176 15100 19185 15140
rect 3679 15077 3745 15100
rect 3831 15077 3913 15100
rect 3999 15077 4065 15100
rect 3679 15058 4065 15077
rect 18799 15077 18865 15100
rect 18951 15077 19033 15100
rect 19119 15077 19185 15100
rect 18799 15058 19185 15077
rect 11320 14848 13996 14888
rect 14036 14848 14045 14888
rect 11320 14804 11360 14848
rect 3043 14764 3052 14804
rect 3092 14764 11360 14804
rect 13490 14743 13614 14762
rect 1411 14680 1420 14720
rect 1460 14680 6124 14720
rect 6164 14680 6173 14720
rect 13490 14657 13509 14743
rect 13595 14720 13614 14743
rect 13595 14680 13612 14720
rect 13652 14680 13661 14720
rect 13595 14657 13614 14680
rect 13490 14638 13614 14657
rect 9091 14428 9100 14468
rect 9140 14428 9484 14468
rect 9524 14428 9533 14468
rect 4919 14407 5305 14426
rect 4919 14384 4985 14407
rect 5071 14384 5153 14407
rect 5239 14384 5305 14407
rect 4919 14344 4928 14384
rect 4968 14344 4985 14384
rect 5071 14344 5092 14384
rect 5132 14344 5153 14384
rect 5239 14344 5256 14384
rect 5296 14344 5305 14384
rect 4919 14321 4985 14344
rect 5071 14321 5153 14344
rect 5239 14321 5305 14344
rect 4919 14302 5305 14321
rect 20039 14407 20425 14426
rect 20039 14384 20105 14407
rect 20191 14384 20273 14407
rect 20359 14384 20425 14407
rect 20039 14344 20048 14384
rect 20088 14344 20105 14384
rect 20191 14344 20212 14384
rect 20252 14344 20273 14384
rect 20359 14344 20376 14384
rect 20416 14344 20425 14384
rect 20039 14321 20105 14344
rect 20191 14321 20273 14344
rect 20359 14321 20425 14344
rect 20039 14302 20425 14321
rect 3811 14092 3820 14132
rect 3860 14092 6220 14132
rect 6260 14092 6269 14132
rect 2371 13840 2380 13880
rect 2420 13840 11788 13880
rect 11828 13840 11837 13880
rect 3679 13651 4065 13670
rect 3679 13628 3745 13651
rect 3831 13628 3913 13651
rect 3999 13628 4065 13651
rect 3679 13588 3688 13628
rect 3728 13588 3745 13628
rect 3831 13588 3852 13628
rect 3892 13588 3913 13628
rect 3999 13588 4016 13628
rect 4056 13588 4065 13628
rect 3679 13565 3745 13588
rect 3831 13565 3913 13588
rect 3999 13565 4065 13588
rect 3679 13546 4065 13565
rect 18799 13651 19185 13670
rect 18799 13628 18865 13651
rect 18951 13628 19033 13651
rect 19119 13628 19185 13651
rect 18799 13588 18808 13628
rect 18848 13588 18865 13628
rect 18951 13588 18972 13628
rect 19012 13588 19033 13628
rect 19119 13588 19136 13628
rect 19176 13588 19185 13628
rect 18799 13565 18865 13588
rect 18951 13565 19033 13588
rect 19119 13565 19185 13588
rect 18799 13546 19185 13565
rect 10435 13420 10444 13460
rect 10484 13420 14956 13460
rect 14996 13420 15005 13460
rect 9955 13168 9964 13208
rect 10004 13168 10444 13208
rect 10484 13168 10493 13208
rect 4919 12895 5305 12914
rect 4919 12872 4985 12895
rect 5071 12872 5153 12895
rect 5239 12872 5305 12895
rect 3139 12832 3148 12872
rect 3188 12832 4300 12872
rect 4340 12832 4349 12872
rect 4919 12832 4928 12872
rect 4968 12832 4985 12872
rect 5071 12832 5092 12872
rect 5132 12832 5153 12872
rect 5239 12832 5256 12872
rect 5296 12832 5305 12872
rect 4919 12809 4985 12832
rect 5071 12809 5153 12832
rect 5239 12809 5305 12832
rect 4919 12790 5305 12809
rect 20039 12895 20425 12914
rect 20039 12872 20105 12895
rect 20191 12872 20273 12895
rect 20359 12872 20425 12895
rect 20039 12832 20048 12872
rect 20088 12832 20105 12872
rect 20191 12832 20212 12872
rect 20252 12832 20273 12872
rect 20359 12832 20376 12872
rect 20416 12832 20425 12872
rect 20039 12809 20105 12832
rect 20191 12809 20273 12832
rect 20359 12809 20425 12832
rect 20039 12790 20425 12809
rect 3139 12580 3148 12620
rect 3188 12580 7564 12620
rect 7604 12580 7613 12620
rect 259 12244 268 12284
rect 308 12244 11308 12284
rect 11348 12244 11357 12284
rect 16003 12244 16012 12284
rect 16052 12244 20044 12284
rect 20084 12244 20093 12284
rect 3679 12139 4065 12158
rect 3679 12116 3745 12139
rect 3831 12116 3913 12139
rect 3999 12116 4065 12139
rect 18799 12139 19185 12158
rect 18799 12116 18865 12139
rect 18951 12116 19033 12139
rect 19119 12116 19185 12139
rect 3679 12076 3688 12116
rect 3728 12076 3745 12116
rect 3831 12076 3852 12116
rect 3892 12076 3913 12116
rect 3999 12076 4016 12116
rect 4056 12076 4065 12116
rect 4483 12076 4492 12116
rect 4532 12076 6604 12116
rect 6644 12076 6653 12116
rect 10819 12076 10828 12116
rect 10868 12076 11308 12116
rect 11348 12076 11357 12116
rect 18799 12076 18808 12116
rect 18848 12076 18865 12116
rect 18951 12076 18972 12116
rect 19012 12076 19033 12116
rect 19119 12076 19136 12116
rect 19176 12076 19185 12116
rect 3679 12053 3745 12076
rect 3831 12053 3913 12076
rect 3999 12053 4065 12076
rect 3679 12034 4065 12053
rect 18799 12053 18865 12076
rect 18951 12053 19033 12076
rect 19119 12053 19185 12076
rect 18799 12034 19185 12053
rect 451 11908 460 11948
rect 500 11908 11404 11948
rect 11444 11908 11453 11948
rect 11395 11740 11404 11780
rect 11444 11740 11596 11780
rect 11636 11740 11645 11780
rect 3715 11656 3724 11696
rect 3764 11656 7468 11696
rect 7508 11656 7517 11696
rect 14563 11488 14572 11528
rect 14612 11488 20044 11528
rect 20084 11488 20093 11528
rect 15427 11404 15436 11444
rect 15476 11404 18892 11444
rect 18932 11404 18941 11444
rect 4919 11383 5305 11402
rect 4919 11360 4985 11383
rect 5071 11360 5153 11383
rect 5239 11360 5305 11383
rect 4919 11320 4928 11360
rect 4968 11320 4985 11360
rect 5071 11320 5092 11360
rect 5132 11320 5153 11360
rect 5239 11320 5256 11360
rect 5296 11320 5305 11360
rect 4919 11297 4985 11320
rect 5071 11297 5153 11320
rect 5239 11297 5305 11320
rect 4919 11278 5305 11297
rect 20039 11383 20425 11402
rect 20039 11360 20105 11383
rect 20191 11360 20273 11383
rect 20359 11360 20425 11383
rect 20039 11320 20048 11360
rect 20088 11320 20105 11360
rect 20191 11320 20212 11360
rect 20252 11320 20273 11360
rect 20359 11320 20376 11360
rect 20416 11320 20425 11360
rect 20039 11297 20105 11320
rect 20191 11297 20273 11320
rect 20359 11297 20425 11320
rect 20039 11278 20425 11297
rect 12643 11236 12652 11276
rect 12692 11236 18988 11276
rect 19028 11236 19037 11276
rect 2851 10984 2860 11024
rect 2900 10984 3532 11024
rect 3572 10984 3581 11024
rect 15427 10900 15436 10940
rect 15476 10900 16012 10940
rect 16052 10900 16061 10940
rect 3679 10627 4065 10646
rect 3679 10604 3745 10627
rect 3831 10604 3913 10627
rect 3999 10604 4065 10627
rect 3679 10564 3688 10604
rect 3728 10564 3745 10604
rect 3831 10564 3852 10604
rect 3892 10564 3913 10604
rect 3999 10564 4016 10604
rect 4056 10564 4065 10604
rect 3679 10541 3745 10564
rect 3831 10541 3913 10564
rect 3999 10541 4065 10564
rect 3679 10522 4065 10541
rect 18799 10627 19185 10646
rect 18799 10604 18865 10627
rect 18951 10604 19033 10627
rect 19119 10604 19185 10627
rect 18799 10564 18808 10604
rect 18848 10564 18865 10604
rect 18951 10564 18972 10604
rect 19012 10564 19033 10604
rect 19119 10564 19136 10604
rect 19176 10564 19185 10604
rect 18799 10541 18865 10564
rect 18951 10541 19033 10564
rect 19119 10541 19185 10564
rect 18799 10522 19185 10541
rect 13123 10144 13132 10184
rect 13172 10144 13612 10184
rect 13652 10144 13661 10184
rect 5443 9976 5452 10016
rect 5492 9976 13612 10016
rect 13652 9976 18316 10016
rect 18356 9976 18365 10016
rect 9955 9892 9964 9932
rect 10004 9892 12556 9932
rect 12596 9892 12605 9932
rect 4919 9871 5305 9890
rect 4919 9848 4985 9871
rect 5071 9848 5153 9871
rect 5239 9848 5305 9871
rect 4919 9808 4928 9848
rect 4968 9808 4985 9848
rect 5071 9808 5092 9848
rect 5132 9808 5153 9848
rect 5239 9808 5256 9848
rect 5296 9808 5305 9848
rect 4919 9785 4985 9808
rect 5071 9785 5153 9808
rect 5239 9785 5305 9808
rect 4919 9766 5305 9785
rect 20039 9871 20425 9890
rect 20039 9848 20105 9871
rect 20191 9848 20273 9871
rect 20359 9848 20425 9871
rect 20039 9808 20048 9848
rect 20088 9808 20105 9848
rect 20191 9808 20212 9848
rect 20252 9808 20273 9848
rect 20359 9808 20376 9848
rect 20416 9808 20425 9848
rect 20039 9785 20105 9808
rect 20191 9785 20273 9808
rect 20359 9785 20425 9808
rect 20039 9766 20425 9785
rect 8803 9724 8812 9764
rect 8852 9724 9484 9764
rect 9524 9724 9533 9764
rect 2083 9388 2092 9428
rect 2132 9388 11788 9428
rect 11828 9388 11837 9428
rect 3679 9115 4065 9134
rect 3679 9092 3745 9115
rect 3831 9092 3913 9115
rect 3999 9092 4065 9115
rect 3679 9052 3688 9092
rect 3728 9052 3745 9092
rect 3831 9052 3852 9092
rect 3892 9052 3913 9092
rect 3999 9052 4016 9092
rect 4056 9052 4065 9092
rect 3679 9029 3745 9052
rect 3831 9029 3913 9052
rect 3999 9029 4065 9052
rect 3679 9010 4065 9029
rect 18799 9115 19185 9134
rect 18799 9092 18865 9115
rect 18951 9092 19033 9115
rect 19119 9092 19185 9115
rect 18799 9052 18808 9092
rect 18848 9052 18865 9092
rect 18951 9052 18972 9092
rect 19012 9052 19033 9092
rect 19119 9052 19136 9092
rect 19176 9052 19185 9092
rect 18799 9029 18865 9052
rect 18951 9029 19033 9052
rect 19119 9029 19185 9052
rect 18799 9010 19185 9029
rect 1795 8716 1804 8756
rect 1844 8716 13900 8756
rect 13940 8716 13949 8756
rect 4963 8632 4972 8672
rect 5012 8632 5356 8672
rect 5396 8632 5405 8672
rect 8803 8632 8812 8672
rect 8852 8632 8861 8672
rect 9091 8632 9100 8672
rect 9140 8632 9580 8672
rect 9620 8632 9629 8672
rect 8812 8588 8852 8632
rect 8812 8548 9388 8588
rect 9428 8548 9437 8588
rect 8803 8464 8812 8504
rect 8852 8464 9484 8504
rect 9524 8464 9533 8504
rect 8707 8380 8716 8420
rect 8756 8380 9196 8420
rect 9236 8380 9245 8420
rect 4919 8359 5305 8378
rect 4919 8336 4985 8359
rect 5071 8336 5153 8359
rect 5239 8336 5305 8359
rect 20039 8359 20425 8378
rect 20039 8336 20105 8359
rect 20191 8336 20273 8359
rect 20359 8336 20425 8359
rect 4919 8296 4928 8336
rect 4968 8296 4985 8336
rect 5071 8296 5092 8336
rect 5132 8296 5153 8336
rect 5239 8296 5256 8336
rect 5296 8296 5305 8336
rect 9475 8296 9484 8336
rect 9524 8296 15340 8336
rect 15380 8296 15389 8336
rect 20039 8296 20048 8336
rect 20088 8296 20105 8336
rect 20191 8296 20212 8336
rect 20252 8296 20273 8336
rect 20359 8296 20376 8336
rect 20416 8296 20425 8336
rect 4919 8273 4985 8296
rect 5071 8273 5153 8296
rect 5239 8273 5305 8296
rect 4919 8254 5305 8273
rect 20039 8273 20105 8296
rect 20191 8273 20273 8296
rect 20359 8273 20425 8296
rect 20039 8254 20425 8273
rect 1219 8128 1228 8168
rect 1268 8128 12172 8168
rect 12212 8128 12221 8168
rect 13219 8128 13228 8168
rect 13268 8128 13612 8168
rect 13652 8128 13661 8168
rect 5443 7876 5452 7916
rect 5492 7876 8716 7916
rect 8756 7876 8765 7916
rect 3679 7603 4065 7622
rect 3679 7580 3745 7603
rect 3831 7580 3913 7603
rect 3999 7580 4065 7603
rect 3679 7540 3688 7580
rect 3728 7540 3745 7580
rect 3831 7540 3852 7580
rect 3892 7540 3913 7580
rect 3999 7540 4016 7580
rect 4056 7540 4065 7580
rect 3679 7517 3745 7540
rect 3831 7517 3913 7540
rect 3999 7517 4065 7540
rect 3679 7498 4065 7517
rect 18799 7603 19185 7622
rect 18799 7580 18865 7603
rect 18951 7580 19033 7603
rect 19119 7580 19185 7603
rect 18799 7540 18808 7580
rect 18848 7540 18865 7580
rect 18951 7540 18972 7580
rect 19012 7540 19033 7580
rect 19119 7540 19136 7580
rect 19176 7540 19185 7580
rect 18799 7517 18865 7540
rect 18951 7517 19033 7540
rect 19119 7517 19185 7540
rect 18799 7498 19185 7517
rect 5635 7456 5644 7496
rect 5684 7456 14092 7496
rect 14132 7456 14141 7496
rect 16291 7372 16300 7412
rect 16340 7372 18892 7412
rect 18932 7372 18941 7412
rect 15523 7288 15532 7328
rect 15572 7288 15724 7328
rect 15764 7288 15773 7328
rect 2500 7120 8716 7160
rect 8756 7120 8765 7160
rect 2500 7076 2540 7120
rect 1603 7036 1612 7076
rect 1652 7036 2540 7076
rect 6211 7036 6220 7076
rect 6260 7036 12652 7076
rect 12692 7036 12701 7076
rect 6115 6952 6124 6992
rect 6164 6952 9676 6992
rect 9716 6952 9725 6992
rect 6499 6868 6508 6908
rect 6548 6868 7644 6908
rect 4919 6847 5305 6866
rect 4919 6824 4985 6847
rect 5071 6824 5153 6847
rect 5239 6824 5305 6847
rect 4919 6784 4928 6824
rect 4968 6784 4985 6824
rect 5071 6784 5092 6824
rect 5132 6784 5153 6824
rect 5239 6784 5256 6824
rect 5296 6784 5305 6824
rect 4919 6761 4985 6784
rect 5071 6761 5153 6784
rect 5239 6761 5305 6784
rect 4919 6742 5305 6761
rect 7604 6740 7644 6868
rect 20039 6847 20425 6866
rect 20039 6824 20105 6847
rect 20191 6824 20273 6847
rect 20359 6824 20425 6847
rect 20039 6784 20048 6824
rect 20088 6784 20105 6824
rect 20191 6784 20212 6824
rect 20252 6784 20273 6824
rect 20359 6784 20376 6824
rect 20416 6784 20425 6824
rect 20039 6761 20105 6784
rect 20191 6761 20273 6784
rect 20359 6761 20425 6784
rect 20039 6742 20425 6761
rect 7604 6700 7660 6740
rect 7700 6700 7709 6740
rect 15715 6700 15724 6740
rect 15764 6700 18892 6740
rect 18932 6700 18941 6740
rect 6115 6616 6124 6656
rect 6164 6616 7852 6656
rect 7892 6616 7901 6656
rect 15235 6448 15244 6488
rect 15284 6448 20812 6488
rect 20852 6448 20861 6488
rect 17138 6343 17262 6362
rect 17138 6320 17157 6343
rect 2659 6280 2668 6320
rect 2708 6280 7276 6320
rect 7316 6280 7325 6320
rect 13027 6280 13036 6320
rect 13076 6280 17157 6320
rect 17138 6257 17157 6280
rect 17243 6257 17262 6343
rect 17138 6238 17262 6257
rect 643 6196 652 6236
rect 692 6196 11360 6236
rect 11320 6152 11360 6196
rect 11320 6112 14572 6152
rect 14612 6112 14621 6152
rect 3679 6091 4065 6110
rect 3679 6068 3745 6091
rect 3831 6068 3913 6091
rect 3999 6068 4065 6091
rect 3679 6028 3688 6068
rect 3728 6028 3745 6068
rect 3831 6028 3852 6068
rect 3892 6028 3913 6068
rect 3999 6028 4016 6068
rect 4056 6028 4065 6068
rect 3679 6005 3745 6028
rect 3831 6005 3913 6028
rect 3999 6005 4065 6028
rect 3679 5986 4065 6005
rect 18799 6091 19185 6110
rect 18799 6068 18865 6091
rect 18951 6068 19033 6091
rect 19119 6068 19185 6091
rect 18799 6028 18808 6068
rect 18848 6028 18865 6068
rect 18951 6028 18972 6068
rect 19012 6028 19033 6068
rect 19119 6028 19136 6068
rect 19176 6028 19185 6068
rect 18799 6005 18865 6028
rect 18951 6005 19033 6028
rect 19119 6005 19185 6028
rect 18799 5986 19185 6005
rect 4771 5860 4780 5900
rect 4820 5860 11404 5900
rect 11444 5860 11453 5900
rect 1507 5776 1516 5816
rect 1556 5776 13132 5816
rect 13172 5776 13181 5816
rect 2371 5692 2380 5732
rect 2420 5692 14188 5732
rect 14228 5692 14237 5732
rect 266 5671 390 5690
rect 266 5585 285 5671
rect 371 5648 390 5671
rect 371 5608 15436 5648
rect 15476 5608 15485 5648
rect 371 5585 390 5608
rect 266 5566 390 5585
rect 931 5524 940 5564
rect 980 5524 2668 5564
rect 2708 5524 2717 5564
rect 1178 5419 1302 5438
rect 1178 5396 1197 5419
rect 1027 5356 1036 5396
rect 1076 5356 1197 5396
rect 1178 5333 1197 5356
rect 1283 5333 1302 5419
rect 1178 5314 1302 5333
rect 4919 5335 5305 5354
rect 4919 5312 4985 5335
rect 5071 5312 5153 5335
rect 5239 5312 5305 5335
rect 4919 5272 4928 5312
rect 4968 5272 4985 5312
rect 5071 5272 5092 5312
rect 5132 5272 5153 5312
rect 5239 5272 5256 5312
rect 5296 5272 5305 5312
rect 4919 5249 4985 5272
rect 5071 5249 5153 5272
rect 5239 5249 5305 5272
rect 4919 5230 5305 5249
rect 20039 5335 20425 5354
rect 20039 5312 20105 5335
rect 20191 5312 20273 5335
rect 20359 5312 20425 5335
rect 20039 5272 20048 5312
rect 20088 5272 20105 5312
rect 20191 5272 20212 5312
rect 20252 5272 20273 5312
rect 20359 5272 20376 5312
rect 20416 5272 20425 5312
rect 20039 5249 20105 5272
rect 20191 5249 20273 5272
rect 20359 5249 20425 5272
rect 20039 5230 20425 5249
rect 1219 5188 1228 5228
rect 1268 5188 1277 5228
rect 1228 5144 1268 5188
rect 1027 5104 1036 5144
rect 1076 5104 1268 5144
rect 12835 5020 12844 5060
rect 12884 5020 13900 5060
rect 13940 5020 13949 5060
rect 13795 4936 13804 4976
rect 13844 4936 17836 4976
rect 17876 4936 17885 4976
rect 1219 4684 1228 4724
rect 1268 4684 13324 4724
rect 13364 4684 13373 4724
rect 5347 4600 5356 4640
rect 5396 4600 10156 4640
rect 10196 4600 10205 4640
rect 3679 4579 4065 4598
rect 3679 4556 3745 4579
rect 3831 4556 3913 4579
rect 3999 4556 4065 4579
rect 3679 4516 3688 4556
rect 3728 4516 3745 4556
rect 3831 4516 3852 4556
rect 3892 4516 3913 4556
rect 3999 4516 4016 4556
rect 4056 4516 4065 4556
rect 3679 4493 3745 4516
rect 3831 4493 3913 4516
rect 3999 4493 4065 4516
rect 3679 4474 4065 4493
rect 18799 4579 19185 4598
rect 18799 4556 18865 4579
rect 18951 4556 19033 4579
rect 19119 4556 19185 4579
rect 18799 4516 18808 4556
rect 18848 4516 18865 4556
rect 18951 4516 18972 4556
rect 19012 4516 19033 4556
rect 19119 4516 19136 4556
rect 19176 4516 19185 4556
rect 18799 4493 18865 4516
rect 18951 4493 19033 4516
rect 19119 4493 19185 4516
rect 18799 4474 19185 4493
rect 10243 4264 10252 4304
rect 10292 4264 10636 4304
rect 10676 4264 10685 4304
rect 3139 4096 3148 4136
rect 3188 4096 18508 4136
rect 18548 4096 18557 4136
rect 4919 3823 5305 3842
rect 4919 3800 4985 3823
rect 5071 3800 5153 3823
rect 5239 3800 5305 3823
rect 20039 3823 20425 3842
rect 20039 3800 20105 3823
rect 20191 3800 20273 3823
rect 20359 3800 20425 3823
rect 4919 3760 4928 3800
rect 4968 3760 4985 3800
rect 5071 3760 5092 3800
rect 5132 3760 5153 3800
rect 5239 3760 5256 3800
rect 5296 3760 5305 3800
rect 8803 3760 8812 3800
rect 8852 3760 9868 3800
rect 9908 3760 9917 3800
rect 20039 3760 20048 3800
rect 20088 3760 20105 3800
rect 20191 3760 20212 3800
rect 20252 3760 20273 3800
rect 20359 3760 20376 3800
rect 20416 3760 20425 3800
rect 4919 3737 4985 3760
rect 5071 3737 5153 3760
rect 5239 3737 5305 3760
rect 4919 3718 5305 3737
rect 20039 3737 20105 3760
rect 20191 3737 20273 3760
rect 20359 3737 20425 3760
rect 20039 3718 20425 3737
rect 7555 3676 7564 3716
rect 7604 3676 10636 3716
rect 10676 3676 10685 3716
rect 5539 3592 5548 3632
rect 5588 3592 5836 3632
rect 5876 3592 5885 3632
rect 5635 3508 5644 3548
rect 5684 3508 9004 3548
rect 9044 3508 9053 3548
rect 3427 3424 3436 3464
rect 3476 3424 8428 3464
rect 8468 3424 8477 3464
rect 7075 3340 7084 3380
rect 7124 3340 11116 3380
rect 11156 3340 11165 3380
rect 12451 3172 12460 3212
rect 12500 3172 17068 3212
rect 17108 3172 17117 3212
rect 5443 3088 5452 3128
rect 5492 3088 11980 3128
rect 12020 3088 12029 3128
rect 3679 3067 4065 3086
rect 3679 3044 3745 3067
rect 3831 3044 3913 3067
rect 3999 3044 4065 3067
rect 3679 3004 3688 3044
rect 3728 3004 3745 3044
rect 3831 3004 3852 3044
rect 3892 3004 3913 3044
rect 3999 3004 4016 3044
rect 4056 3004 4065 3044
rect 3679 2981 3745 3004
rect 3831 2981 3913 3004
rect 3999 2981 4065 3004
rect 3679 2962 4065 2981
rect 12122 3067 12246 3086
rect 12122 2981 12141 3067
rect 12227 3044 12246 3067
rect 18799 3067 19185 3086
rect 18799 3044 18865 3067
rect 18951 3044 19033 3067
rect 19119 3044 19185 3067
rect 12227 3004 14572 3044
rect 14612 3004 14621 3044
rect 18799 3004 18808 3044
rect 18848 3004 18865 3044
rect 18951 3004 18972 3044
rect 19012 3004 19033 3044
rect 19119 3004 19136 3044
rect 19176 3004 19185 3044
rect 12227 2981 12246 3004
rect 12122 2962 12246 2981
rect 18799 2981 18865 3004
rect 18951 2981 19033 3004
rect 19119 2981 19185 3004
rect 18799 2962 19185 2981
rect 7459 2668 7468 2708
rect 7508 2668 11884 2708
rect 11924 2668 11933 2708
rect 10298 2479 10422 2498
rect 10298 2456 10317 2479
rect 1219 2416 1228 2456
rect 1268 2416 7852 2456
rect 7892 2416 7901 2456
rect 8524 2416 10317 2456
rect 8524 2372 8564 2416
rect 10298 2393 10317 2416
rect 10403 2393 10422 2479
rect 10298 2374 10422 2393
rect 5780 2332 8564 2372
rect 10723 2332 10732 2372
rect 10772 2332 14572 2372
rect 14612 2332 14621 2372
rect 4919 2311 5305 2330
rect 4919 2288 4985 2311
rect 5071 2288 5153 2311
rect 5239 2288 5305 2311
rect 4919 2248 4928 2288
rect 4968 2248 4985 2288
rect 5071 2248 5092 2288
rect 5132 2248 5153 2288
rect 5239 2248 5256 2288
rect 5296 2248 5305 2288
rect 4919 2225 4985 2248
rect 5071 2225 5153 2248
rect 5239 2225 5305 2248
rect 4919 2206 5305 2225
rect 5780 2120 5820 2332
rect 20039 2311 20425 2330
rect 20039 2288 20105 2311
rect 20191 2288 20273 2311
rect 20359 2288 20425 2311
rect 6307 2248 6316 2288
rect 6356 2248 13996 2288
rect 14036 2248 14045 2288
rect 20039 2248 20048 2288
rect 20088 2248 20105 2288
rect 20191 2248 20212 2288
rect 20252 2248 20273 2288
rect 20359 2248 20376 2288
rect 20416 2248 20425 2288
rect 20039 2225 20105 2248
rect 20191 2225 20273 2248
rect 20359 2225 20425 2248
rect 20039 2206 20425 2225
rect 9386 2143 9510 2162
rect 9386 2120 9405 2143
rect 4099 2080 4108 2120
rect 4148 2080 5820 2120
rect 9283 2080 9292 2120
rect 9332 2080 9405 2120
rect 9386 2057 9405 2080
rect 9491 2057 9510 2143
rect 9386 2038 9510 2057
rect 11320 1996 13228 2036
rect 13268 1996 13277 2036
rect 11320 1952 11360 1996
rect 5923 1912 5932 1952
rect 5972 1912 11360 1952
rect 3619 1828 3628 1868
rect 3668 1828 6892 1868
rect 6932 1828 6941 1868
rect 1411 1660 1420 1700
rect 1460 1660 15436 1700
rect 15476 1660 15485 1700
rect 3679 1555 4065 1574
rect 3679 1532 3745 1555
rect 3831 1532 3913 1555
rect 3999 1532 4065 1555
rect 3679 1492 3688 1532
rect 3728 1492 3745 1532
rect 3831 1492 3852 1532
rect 3892 1492 3913 1532
rect 3999 1492 4016 1532
rect 4056 1492 4065 1532
rect 3679 1469 3745 1492
rect 3831 1469 3913 1492
rect 3999 1469 4065 1492
rect 3679 1450 4065 1469
rect 18799 1555 19185 1574
rect 18799 1532 18865 1555
rect 18951 1532 19033 1555
rect 19119 1532 19185 1555
rect 18799 1492 18808 1532
rect 18848 1492 18865 1532
rect 18951 1492 18972 1532
rect 19012 1492 19033 1532
rect 19119 1492 19136 1532
rect 19176 1492 19185 1532
rect 18799 1469 18865 1492
rect 18951 1469 19033 1492
rect 19119 1469 19185 1492
rect 18799 1450 19185 1469
rect 4412 1408 18700 1448
rect 18740 1408 18749 1448
rect 4412 1364 4452 1408
rect 3523 1324 3532 1364
rect 3572 1324 4452 1364
rect 5059 1324 5068 1364
rect 5108 1324 6316 1364
rect 6356 1324 6365 1364
rect 8474 1303 8598 1322
rect 3715 1240 3724 1280
rect 3764 1240 6700 1280
rect 6740 1240 6749 1280
rect 8474 1217 8493 1303
rect 8579 1217 8598 1303
rect 13490 1303 13614 1322
rect 13490 1280 13509 1303
rect 12739 1240 12748 1280
rect 12788 1240 13509 1280
rect 8474 1198 8598 1217
rect 13490 1217 13509 1240
rect 13595 1217 13614 1303
rect 13490 1198 13614 1217
rect 5635 1156 5644 1196
rect 5684 1156 8100 1196
rect 8060 1112 8100 1156
rect 8060 1072 12364 1112
rect 12404 1072 12413 1112
rect 14402 967 14526 986
rect 14402 944 14421 967
rect 14275 904 14284 944
rect 14324 904 14421 944
rect 14402 881 14421 904
rect 14507 881 14526 967
rect 14402 862 14526 881
rect 15770 883 15894 902
rect 5923 820 5932 860
rect 5972 820 10156 860
rect 10196 820 10205 860
rect 2090 799 2214 818
rect 2090 713 2109 799
rect 2195 776 2214 799
rect 4919 799 5305 818
rect 4919 776 4985 799
rect 5071 776 5153 799
rect 5239 776 5305 799
rect 15770 797 15789 883
rect 15875 860 15894 883
rect 15875 820 18700 860
rect 18740 820 18749 860
rect 15875 797 15894 820
rect 15770 778 15894 797
rect 20039 799 20425 818
rect 2195 736 4684 776
rect 4724 736 4733 776
rect 4919 736 4928 776
rect 4968 736 4985 776
rect 5071 736 5092 776
rect 5132 736 5153 776
rect 5239 736 5256 776
rect 5296 736 5305 776
rect 2195 713 2214 736
rect 2090 694 2214 713
rect 4919 713 4985 736
rect 5071 713 5153 736
rect 5239 713 5305 736
rect 4919 694 5305 713
rect 20039 776 20105 799
rect 20191 776 20273 799
rect 20359 776 20425 799
rect 20039 736 20048 776
rect 20088 736 20105 776
rect 20191 736 20212 776
rect 20252 736 20273 776
rect 20359 736 20376 776
rect 20416 736 20425 776
rect 20039 713 20105 736
rect 20191 713 20273 736
rect 20359 713 20425 736
rect 20039 694 20425 713
rect 14371 652 14380 692
rect 14420 652 19276 692
rect 19316 652 19325 692
rect 7106 379 7230 398
rect 7106 356 7125 379
rect 6595 316 6604 356
rect 6644 316 7125 356
rect 7106 293 7125 316
rect 7211 293 7230 379
rect 7106 274 7230 293
rect 266 211 390 230
rect 266 188 285 211
rect 259 148 268 188
rect 266 125 285 148
rect 371 125 390 211
rect 5251 148 5260 188
rect 5300 148 11500 188
rect 11540 148 11549 188
rect 266 106 390 125
rect 6019 64 6028 104
rect 6068 64 10060 104
rect 10100 64 10109 104
<< via5 >>
rect 4985 41600 5071 41623
rect 5153 41600 5239 41623
rect 4985 41560 5010 41600
rect 5010 41560 5050 41600
rect 5050 41560 5071 41600
rect 5153 41560 5174 41600
rect 5174 41560 5214 41600
rect 5214 41560 5239 41600
rect 4985 41537 5071 41560
rect 5153 41537 5239 41560
rect 20105 41600 20191 41623
rect 20273 41600 20359 41623
rect 20105 41560 20130 41600
rect 20130 41560 20170 41600
rect 20170 41560 20191 41600
rect 20273 41560 20294 41600
rect 20294 41560 20334 41600
rect 20334 41560 20359 41600
rect 20105 41537 20191 41560
rect 20273 41537 20359 41560
rect 17157 40949 17243 41035
rect 3745 40844 3831 40867
rect 3913 40844 3999 40867
rect 3745 40804 3770 40844
rect 3770 40804 3810 40844
rect 3810 40804 3831 40844
rect 3913 40804 3934 40844
rect 3934 40804 3974 40844
rect 3974 40804 3999 40844
rect 3745 40781 3831 40804
rect 3913 40781 3999 40804
rect 18865 40844 18951 40867
rect 19033 40844 19119 40867
rect 18865 40804 18890 40844
rect 18890 40804 18930 40844
rect 18930 40804 18951 40844
rect 19033 40804 19054 40844
rect 19054 40804 19094 40844
rect 19094 40804 19119 40844
rect 18865 40781 18951 40804
rect 19033 40781 19119 40804
rect 14421 40277 14507 40363
rect 4985 40088 5071 40111
rect 5153 40088 5239 40111
rect 4985 40048 5010 40088
rect 5010 40048 5050 40088
rect 5050 40048 5071 40088
rect 5153 40048 5174 40088
rect 5174 40048 5214 40088
rect 5214 40048 5239 40088
rect 4985 40025 5071 40048
rect 5153 40025 5239 40048
rect 20105 40088 20191 40111
rect 20273 40088 20359 40111
rect 20105 40048 20130 40088
rect 20130 40048 20170 40088
rect 20170 40048 20191 40088
rect 20273 40048 20294 40088
rect 20294 40048 20334 40088
rect 20334 40048 20359 40088
rect 20105 40025 20191 40048
rect 20273 40025 20359 40048
rect 3745 39332 3831 39355
rect 3913 39332 3999 39355
rect 13509 39353 13595 39439
rect 3745 39292 3770 39332
rect 3770 39292 3810 39332
rect 3810 39292 3831 39332
rect 3913 39292 3934 39332
rect 3934 39292 3974 39332
rect 3974 39292 3999 39332
rect 3745 39269 3831 39292
rect 3913 39269 3999 39292
rect 18865 39332 18951 39355
rect 19033 39332 19119 39355
rect 18865 39292 18890 39332
rect 18890 39292 18930 39332
rect 18930 39292 18951 39332
rect 19033 39292 19054 39332
rect 19054 39292 19094 39332
rect 19094 39292 19119 39332
rect 18865 39269 18951 39292
rect 19033 39269 19119 39292
rect 4985 38576 5071 38599
rect 5153 38576 5239 38599
rect 4985 38536 5010 38576
rect 5010 38536 5050 38576
rect 5050 38536 5071 38576
rect 5153 38536 5174 38576
rect 5174 38536 5214 38576
rect 5214 38536 5239 38576
rect 4985 38513 5071 38536
rect 5153 38513 5239 38536
rect 20105 38576 20191 38599
rect 20273 38576 20359 38599
rect 20105 38536 20130 38576
rect 20130 38536 20170 38576
rect 20170 38536 20191 38576
rect 20273 38536 20294 38576
rect 20294 38536 20334 38576
rect 20334 38536 20359 38576
rect 20105 38513 20191 38536
rect 20273 38513 20359 38536
rect 7125 38261 7211 38347
rect 3745 37820 3831 37843
rect 3913 37820 3999 37843
rect 3745 37780 3770 37820
rect 3770 37780 3810 37820
rect 3810 37780 3831 37820
rect 3913 37780 3934 37820
rect 3934 37780 3974 37820
rect 3974 37780 3999 37820
rect 3745 37757 3831 37780
rect 3913 37757 3999 37780
rect 18865 37820 18951 37843
rect 19033 37820 19119 37843
rect 18865 37780 18890 37820
rect 18890 37780 18930 37820
rect 18930 37780 18951 37820
rect 19033 37780 19054 37820
rect 19054 37780 19094 37820
rect 19094 37780 19119 37820
rect 18865 37757 18951 37780
rect 19033 37757 19119 37780
rect 4985 37064 5071 37087
rect 5153 37064 5239 37087
rect 4985 37024 5010 37064
rect 5010 37024 5050 37064
rect 5050 37024 5071 37064
rect 5153 37024 5174 37064
rect 5174 37024 5214 37064
rect 5214 37024 5239 37064
rect 4985 37001 5071 37024
rect 5153 37001 5239 37024
rect 20105 37064 20191 37087
rect 20273 37064 20359 37087
rect 20105 37024 20130 37064
rect 20130 37024 20170 37064
rect 20170 37024 20191 37064
rect 20273 37024 20294 37064
rect 20294 37024 20334 37064
rect 20334 37024 20359 37064
rect 20105 37001 20191 37024
rect 20273 37001 20359 37024
rect 3745 36308 3831 36331
rect 3913 36308 3999 36331
rect 9405 36308 9491 36331
rect 3745 36268 3770 36308
rect 3770 36268 3810 36308
rect 3810 36268 3831 36308
rect 3913 36268 3934 36308
rect 3934 36268 3974 36308
rect 3974 36268 3999 36308
rect 9405 36268 9428 36308
rect 9428 36268 9491 36308
rect 3745 36245 3831 36268
rect 3913 36245 3999 36268
rect 9405 36245 9491 36268
rect 18865 36308 18951 36331
rect 19033 36308 19119 36331
rect 18865 36268 18890 36308
rect 18890 36268 18930 36308
rect 18930 36268 18951 36308
rect 19033 36268 19054 36308
rect 19054 36268 19094 36308
rect 19094 36268 19119 36308
rect 18865 36245 18951 36268
rect 19033 36245 19119 36268
rect 4985 35552 5071 35575
rect 5153 35552 5239 35575
rect 4985 35512 5010 35552
rect 5010 35512 5050 35552
rect 5050 35512 5071 35552
rect 5153 35512 5174 35552
rect 5174 35512 5214 35552
rect 5214 35512 5239 35552
rect 4985 35489 5071 35512
rect 5153 35489 5239 35512
rect 20105 35552 20191 35575
rect 20273 35552 20359 35575
rect 20105 35512 20130 35552
rect 20130 35512 20170 35552
rect 20170 35512 20191 35552
rect 20273 35512 20294 35552
rect 20294 35512 20334 35552
rect 20334 35512 20359 35552
rect 15789 35405 15875 35491
rect 20105 35489 20191 35512
rect 20273 35489 20359 35512
rect 1197 35237 1283 35323
rect 3745 34796 3831 34819
rect 3913 34796 3999 34819
rect 3745 34756 3770 34796
rect 3770 34756 3810 34796
rect 3810 34756 3831 34796
rect 3913 34756 3934 34796
rect 3934 34756 3974 34796
rect 3974 34756 3999 34796
rect 3745 34733 3831 34756
rect 3913 34733 3999 34756
rect 18865 34796 18951 34819
rect 19033 34796 19119 34819
rect 18865 34756 18890 34796
rect 18890 34756 18930 34796
rect 18930 34756 18951 34796
rect 19033 34756 19054 34796
rect 19054 34756 19094 34796
rect 19094 34756 19119 34796
rect 18865 34733 18951 34756
rect 19033 34733 19119 34756
rect 4985 34040 5071 34063
rect 5153 34040 5239 34063
rect 20105 34040 20191 34063
rect 20273 34040 20359 34063
rect 4985 34000 5010 34040
rect 5010 34000 5050 34040
rect 5050 34000 5071 34040
rect 5153 34000 5174 34040
rect 5174 34000 5214 34040
rect 5214 34000 5239 34040
rect 20105 34000 20130 34040
rect 20130 34000 20170 34040
rect 20170 34000 20191 34040
rect 20273 34000 20294 34040
rect 20294 34000 20334 34040
rect 20334 34000 20359 34040
rect 4985 33977 5071 34000
rect 5153 33977 5239 34000
rect 20105 33977 20191 34000
rect 20273 33977 20359 34000
rect 3745 33284 3831 33307
rect 3913 33284 3999 33307
rect 3745 33244 3770 33284
rect 3770 33244 3810 33284
rect 3810 33244 3831 33284
rect 3913 33244 3934 33284
rect 3934 33244 3974 33284
rect 3974 33244 3999 33284
rect 3745 33221 3831 33244
rect 3913 33221 3999 33244
rect 18865 33284 18951 33307
rect 19033 33284 19119 33307
rect 18865 33244 18890 33284
rect 18890 33244 18930 33284
rect 18930 33244 18951 33284
rect 19033 33244 19054 33284
rect 19054 33244 19094 33284
rect 19094 33244 19119 33284
rect 18865 33221 18951 33244
rect 19033 33221 19119 33244
rect 4985 32528 5071 32551
rect 5153 32528 5239 32551
rect 4985 32488 5010 32528
rect 5010 32488 5050 32528
rect 5050 32488 5071 32528
rect 5153 32488 5174 32528
rect 5174 32488 5214 32528
rect 5214 32488 5239 32528
rect 4985 32465 5071 32488
rect 5153 32465 5239 32488
rect 20105 32528 20191 32551
rect 20273 32528 20359 32551
rect 20105 32488 20130 32528
rect 20130 32488 20170 32528
rect 20170 32488 20191 32528
rect 20273 32488 20294 32528
rect 20294 32488 20334 32528
rect 20334 32488 20359 32528
rect 20105 32465 20191 32488
rect 20273 32465 20359 32488
rect 3745 31772 3831 31795
rect 3913 31772 3999 31795
rect 3745 31732 3770 31772
rect 3770 31732 3810 31772
rect 3810 31732 3831 31772
rect 3913 31732 3934 31772
rect 3934 31732 3974 31772
rect 3974 31732 3999 31772
rect 3745 31709 3831 31732
rect 3913 31709 3999 31732
rect 18865 31772 18951 31795
rect 19033 31772 19119 31795
rect 18865 31732 18890 31772
rect 18890 31732 18930 31772
rect 18930 31732 18951 31772
rect 19033 31732 19054 31772
rect 19054 31732 19094 31772
rect 19094 31732 19119 31772
rect 18865 31709 18951 31732
rect 19033 31709 19119 31732
rect 12141 31289 12227 31375
rect 4985 31016 5071 31039
rect 5153 31016 5239 31039
rect 10317 31037 10403 31123
rect 4985 30976 5010 31016
rect 5010 30976 5050 31016
rect 5050 30976 5071 31016
rect 5153 30976 5174 31016
rect 5174 30976 5214 31016
rect 5214 30976 5239 31016
rect 4985 30953 5071 30976
rect 5153 30953 5239 30976
rect 20105 31016 20191 31039
rect 20273 31016 20359 31039
rect 20105 30976 20130 31016
rect 20130 30976 20170 31016
rect 20170 30976 20191 31016
rect 20273 30976 20294 31016
rect 20294 30976 20334 31016
rect 20334 30976 20359 31016
rect 20105 30953 20191 30976
rect 20273 30953 20359 30976
rect 3745 30260 3831 30283
rect 3913 30260 3999 30283
rect 3745 30220 3770 30260
rect 3770 30220 3810 30260
rect 3810 30220 3831 30260
rect 3913 30220 3934 30260
rect 3934 30220 3974 30260
rect 3974 30220 3999 30260
rect 3745 30197 3831 30220
rect 3913 30197 3999 30220
rect 18865 30260 18951 30283
rect 19033 30260 19119 30283
rect 18865 30220 18890 30260
rect 18890 30220 18930 30260
rect 18930 30220 18951 30260
rect 19033 30220 19054 30260
rect 19054 30220 19094 30260
rect 19094 30220 19119 30260
rect 18865 30197 18951 30220
rect 19033 30197 19119 30220
rect 4985 29504 5071 29527
rect 5153 29504 5239 29527
rect 4985 29464 5010 29504
rect 5010 29464 5050 29504
rect 5050 29464 5071 29504
rect 5153 29464 5174 29504
rect 5174 29464 5214 29504
rect 5214 29464 5239 29504
rect 4985 29441 5071 29464
rect 5153 29441 5239 29464
rect 20105 29504 20191 29527
rect 20273 29504 20359 29527
rect 20105 29464 20130 29504
rect 20130 29464 20170 29504
rect 20170 29464 20191 29504
rect 20273 29464 20294 29504
rect 20294 29464 20334 29504
rect 20334 29464 20359 29504
rect 20105 29441 20191 29464
rect 20273 29441 20359 29464
rect 3745 28748 3831 28771
rect 3913 28748 3999 28771
rect 3745 28708 3770 28748
rect 3770 28708 3810 28748
rect 3810 28708 3831 28748
rect 3913 28708 3934 28748
rect 3934 28708 3974 28748
rect 3974 28708 3999 28748
rect 3745 28685 3831 28708
rect 3913 28685 3999 28708
rect 18865 28748 18951 28771
rect 19033 28748 19119 28771
rect 18865 28708 18890 28748
rect 18890 28708 18930 28748
rect 18930 28708 18951 28748
rect 19033 28708 19054 28748
rect 19054 28708 19094 28748
rect 19094 28708 19119 28748
rect 18865 28685 18951 28708
rect 19033 28685 19119 28708
rect 4985 27992 5071 28015
rect 5153 27992 5239 28015
rect 4985 27952 5010 27992
rect 5010 27952 5050 27992
rect 5050 27952 5071 27992
rect 5153 27952 5174 27992
rect 5174 27952 5214 27992
rect 5214 27952 5239 27992
rect 4985 27929 5071 27952
rect 5153 27929 5239 27952
rect 20105 27992 20191 28015
rect 20273 27992 20359 28015
rect 20105 27952 20130 27992
rect 20130 27952 20170 27992
rect 20170 27952 20191 27992
rect 20273 27952 20294 27992
rect 20294 27952 20334 27992
rect 20334 27952 20359 27992
rect 20105 27929 20191 27952
rect 20273 27929 20359 27952
rect 2109 27677 2195 27763
rect 3745 27236 3831 27259
rect 3913 27236 3999 27259
rect 3745 27196 3770 27236
rect 3770 27196 3810 27236
rect 3810 27196 3831 27236
rect 3913 27196 3934 27236
rect 3934 27196 3974 27236
rect 3974 27196 3999 27236
rect 3745 27173 3831 27196
rect 3913 27173 3999 27196
rect 18865 27236 18951 27259
rect 19033 27236 19119 27259
rect 18865 27196 18890 27236
rect 18890 27196 18930 27236
rect 18930 27196 18951 27236
rect 19033 27196 19054 27236
rect 19054 27196 19094 27236
rect 19094 27196 19119 27236
rect 18865 27173 18951 27196
rect 19033 27173 19119 27196
rect 4985 26480 5071 26503
rect 5153 26480 5239 26503
rect 20105 26480 20191 26503
rect 20273 26480 20359 26503
rect 4985 26440 5010 26480
rect 5010 26440 5050 26480
rect 5050 26440 5071 26480
rect 5153 26440 5174 26480
rect 5174 26440 5214 26480
rect 5214 26440 5239 26480
rect 20105 26440 20130 26480
rect 20130 26440 20170 26480
rect 20170 26440 20191 26480
rect 20273 26440 20294 26480
rect 20294 26440 20334 26480
rect 20334 26440 20359 26480
rect 4985 26417 5071 26440
rect 5153 26417 5239 26440
rect 20105 26417 20191 26440
rect 20273 26417 20359 26440
rect 3745 25724 3831 25747
rect 3913 25724 3999 25747
rect 18865 25724 18951 25747
rect 19033 25724 19119 25747
rect 3745 25684 3770 25724
rect 3770 25684 3810 25724
rect 3810 25684 3831 25724
rect 3913 25684 3934 25724
rect 3934 25684 3974 25724
rect 3974 25684 3999 25724
rect 18865 25684 18890 25724
rect 18890 25684 18930 25724
rect 18930 25684 18951 25724
rect 19033 25684 19054 25724
rect 19054 25684 19094 25724
rect 19094 25684 19119 25724
rect 3745 25661 3831 25684
rect 3913 25661 3999 25684
rect 18865 25661 18951 25684
rect 19033 25661 19119 25684
rect 4985 24968 5071 24991
rect 5153 24968 5239 24991
rect 4985 24928 5010 24968
rect 5010 24928 5050 24968
rect 5050 24928 5071 24968
rect 5153 24928 5174 24968
rect 5174 24928 5214 24968
rect 5214 24928 5239 24968
rect 4985 24905 5071 24928
rect 5153 24905 5239 24928
rect 20105 24968 20191 24991
rect 20273 24968 20359 24991
rect 20105 24928 20130 24968
rect 20130 24928 20170 24968
rect 20170 24928 20191 24968
rect 20273 24928 20294 24968
rect 20294 24928 20334 24968
rect 20334 24928 20359 24968
rect 20105 24905 20191 24928
rect 20273 24905 20359 24928
rect 3745 24212 3831 24235
rect 3913 24212 3999 24235
rect 3745 24172 3770 24212
rect 3770 24172 3810 24212
rect 3810 24172 3831 24212
rect 3913 24172 3934 24212
rect 3934 24172 3974 24212
rect 3974 24172 3999 24212
rect 3745 24149 3831 24172
rect 3913 24149 3999 24172
rect 18865 24212 18951 24235
rect 19033 24212 19119 24235
rect 18865 24172 18890 24212
rect 18890 24172 18930 24212
rect 18930 24172 18951 24212
rect 19033 24172 19054 24212
rect 19054 24172 19094 24212
rect 19094 24172 19119 24212
rect 18865 24149 18951 24172
rect 19033 24149 19119 24172
rect 4985 23456 5071 23479
rect 5153 23456 5239 23479
rect 4985 23416 5010 23456
rect 5010 23416 5050 23456
rect 5050 23416 5071 23456
rect 5153 23416 5174 23456
rect 5174 23416 5214 23456
rect 5214 23416 5239 23456
rect 4985 23393 5071 23416
rect 5153 23393 5239 23416
rect 20105 23456 20191 23479
rect 20273 23456 20359 23479
rect 20105 23416 20130 23456
rect 20130 23416 20170 23456
rect 20170 23416 20191 23456
rect 20273 23416 20294 23456
rect 20294 23416 20334 23456
rect 20334 23416 20359 23456
rect 20105 23393 20191 23416
rect 20273 23393 20359 23416
rect 3745 22700 3831 22723
rect 3913 22700 3999 22723
rect 18865 22700 18951 22723
rect 19033 22700 19119 22723
rect 3745 22660 3770 22700
rect 3770 22660 3810 22700
rect 3810 22660 3831 22700
rect 3913 22660 3934 22700
rect 3934 22660 3974 22700
rect 3974 22660 3999 22700
rect 18865 22660 18890 22700
rect 18890 22660 18930 22700
rect 18930 22660 18951 22700
rect 19033 22660 19054 22700
rect 19054 22660 19094 22700
rect 19094 22660 19119 22700
rect 3745 22637 3831 22660
rect 3913 22637 3999 22660
rect 18865 22637 18951 22660
rect 19033 22637 19119 22660
rect 4985 21944 5071 21967
rect 5153 21944 5239 21967
rect 4985 21904 5010 21944
rect 5010 21904 5050 21944
rect 5050 21904 5071 21944
rect 5153 21904 5174 21944
rect 5174 21904 5214 21944
rect 5214 21904 5239 21944
rect 4985 21881 5071 21904
rect 5153 21881 5239 21904
rect 20105 21944 20191 21967
rect 20273 21944 20359 21967
rect 20105 21904 20130 21944
rect 20130 21904 20170 21944
rect 20170 21904 20191 21944
rect 20273 21904 20294 21944
rect 20294 21904 20334 21944
rect 20334 21904 20359 21944
rect 20105 21881 20191 21904
rect 20273 21881 20359 21904
rect 8493 21377 8579 21463
rect 3745 21188 3831 21211
rect 3913 21188 3999 21211
rect 3745 21148 3770 21188
rect 3770 21148 3810 21188
rect 3810 21148 3831 21188
rect 3913 21148 3934 21188
rect 3934 21148 3974 21188
rect 3974 21148 3999 21188
rect 3745 21125 3831 21148
rect 3913 21125 3999 21148
rect 18865 21188 18951 21211
rect 19033 21188 19119 21211
rect 18865 21148 18890 21188
rect 18890 21148 18930 21188
rect 18930 21148 18951 21188
rect 19033 21148 19054 21188
rect 19054 21148 19094 21188
rect 19094 21148 19119 21188
rect 18865 21125 18951 21148
rect 19033 21125 19119 21148
rect 4985 20432 5071 20455
rect 5153 20432 5239 20455
rect 20105 20432 20191 20455
rect 20273 20432 20359 20455
rect 4985 20392 5010 20432
rect 5010 20392 5050 20432
rect 5050 20392 5071 20432
rect 5153 20392 5174 20432
rect 5174 20392 5214 20432
rect 5214 20392 5239 20432
rect 20105 20392 20130 20432
rect 20130 20392 20170 20432
rect 20170 20392 20191 20432
rect 20273 20392 20294 20432
rect 20294 20392 20334 20432
rect 20334 20392 20359 20432
rect 4985 20369 5071 20392
rect 5153 20369 5239 20392
rect 20105 20369 20191 20392
rect 20273 20369 20359 20392
rect 3745 19676 3831 19699
rect 3913 19676 3999 19699
rect 3745 19636 3770 19676
rect 3770 19636 3810 19676
rect 3810 19636 3831 19676
rect 3913 19636 3934 19676
rect 3934 19636 3974 19676
rect 3974 19636 3999 19676
rect 3745 19613 3831 19636
rect 3913 19613 3999 19636
rect 18865 19676 18951 19699
rect 19033 19676 19119 19699
rect 18865 19636 18890 19676
rect 18890 19636 18930 19676
rect 18930 19636 18951 19676
rect 19033 19636 19054 19676
rect 19054 19636 19094 19676
rect 19094 19636 19119 19676
rect 18865 19613 18951 19636
rect 19033 19613 19119 19636
rect 4985 18920 5071 18943
rect 5153 18920 5239 18943
rect 4985 18880 5010 18920
rect 5010 18880 5050 18920
rect 5050 18880 5071 18920
rect 5153 18880 5174 18920
rect 5174 18880 5214 18920
rect 5214 18880 5239 18920
rect 4985 18857 5071 18880
rect 5153 18857 5239 18880
rect 20105 18920 20191 18943
rect 20273 18920 20359 18943
rect 20105 18880 20130 18920
rect 20130 18880 20170 18920
rect 20170 18880 20191 18920
rect 20273 18880 20294 18920
rect 20294 18880 20334 18920
rect 20334 18880 20359 18920
rect 20105 18857 20191 18880
rect 20273 18857 20359 18880
rect 3745 18164 3831 18187
rect 3913 18164 3999 18187
rect 3745 18124 3770 18164
rect 3770 18124 3810 18164
rect 3810 18124 3831 18164
rect 3913 18124 3934 18164
rect 3934 18124 3974 18164
rect 3974 18124 3999 18164
rect 3745 18101 3831 18124
rect 3913 18101 3999 18124
rect 18865 18164 18951 18187
rect 19033 18164 19119 18187
rect 18865 18124 18890 18164
rect 18890 18124 18930 18164
rect 18930 18124 18951 18164
rect 19033 18124 19054 18164
rect 19054 18124 19094 18164
rect 19094 18124 19119 18164
rect 18865 18101 18951 18124
rect 19033 18101 19119 18124
rect 4985 17408 5071 17431
rect 5153 17408 5239 17431
rect 4985 17368 5010 17408
rect 5010 17368 5050 17408
rect 5050 17368 5071 17408
rect 5153 17368 5174 17408
rect 5174 17368 5214 17408
rect 5214 17368 5239 17408
rect 4985 17345 5071 17368
rect 5153 17345 5239 17368
rect 20105 17408 20191 17431
rect 20273 17408 20359 17431
rect 20105 17368 20130 17408
rect 20130 17368 20170 17408
rect 20170 17368 20191 17408
rect 20273 17368 20294 17408
rect 20294 17368 20334 17408
rect 20334 17368 20359 17408
rect 20105 17345 20191 17368
rect 20273 17345 20359 17368
rect 3745 16652 3831 16675
rect 3913 16652 3999 16675
rect 3745 16612 3770 16652
rect 3770 16612 3810 16652
rect 3810 16612 3831 16652
rect 3913 16612 3934 16652
rect 3934 16612 3974 16652
rect 3974 16612 3999 16652
rect 3745 16589 3831 16612
rect 3913 16589 3999 16612
rect 18865 16652 18951 16675
rect 19033 16652 19119 16675
rect 18865 16612 18890 16652
rect 18890 16612 18930 16652
rect 18930 16612 18951 16652
rect 19033 16612 19054 16652
rect 19054 16612 19094 16652
rect 19094 16612 19119 16652
rect 18865 16589 18951 16612
rect 19033 16589 19119 16612
rect 4985 15896 5071 15919
rect 5153 15896 5239 15919
rect 4985 15856 5010 15896
rect 5010 15856 5050 15896
rect 5050 15856 5071 15896
rect 5153 15856 5174 15896
rect 5174 15856 5214 15896
rect 5214 15856 5239 15896
rect 4985 15833 5071 15856
rect 5153 15833 5239 15856
rect 20105 15896 20191 15919
rect 20273 15896 20359 15919
rect 20105 15856 20130 15896
rect 20130 15856 20170 15896
rect 20170 15856 20191 15896
rect 20273 15856 20294 15896
rect 20294 15856 20334 15896
rect 20334 15856 20359 15896
rect 20105 15833 20191 15856
rect 20273 15833 20359 15856
rect 13509 15329 13595 15415
rect 3745 15140 3831 15163
rect 3913 15140 3999 15163
rect 18865 15140 18951 15163
rect 19033 15140 19119 15163
rect 3745 15100 3770 15140
rect 3770 15100 3810 15140
rect 3810 15100 3831 15140
rect 3913 15100 3934 15140
rect 3934 15100 3974 15140
rect 3974 15100 3999 15140
rect 18865 15100 18890 15140
rect 18890 15100 18930 15140
rect 18930 15100 18951 15140
rect 19033 15100 19054 15140
rect 19054 15100 19094 15140
rect 19094 15100 19119 15140
rect 3745 15077 3831 15100
rect 3913 15077 3999 15100
rect 18865 15077 18951 15100
rect 19033 15077 19119 15100
rect 13509 14657 13595 14743
rect 4985 14384 5071 14407
rect 5153 14384 5239 14407
rect 4985 14344 5010 14384
rect 5010 14344 5050 14384
rect 5050 14344 5071 14384
rect 5153 14344 5174 14384
rect 5174 14344 5214 14384
rect 5214 14344 5239 14384
rect 4985 14321 5071 14344
rect 5153 14321 5239 14344
rect 20105 14384 20191 14407
rect 20273 14384 20359 14407
rect 20105 14344 20130 14384
rect 20130 14344 20170 14384
rect 20170 14344 20191 14384
rect 20273 14344 20294 14384
rect 20294 14344 20334 14384
rect 20334 14344 20359 14384
rect 20105 14321 20191 14344
rect 20273 14321 20359 14344
rect 3745 13628 3831 13651
rect 3913 13628 3999 13651
rect 3745 13588 3770 13628
rect 3770 13588 3810 13628
rect 3810 13588 3831 13628
rect 3913 13588 3934 13628
rect 3934 13588 3974 13628
rect 3974 13588 3999 13628
rect 3745 13565 3831 13588
rect 3913 13565 3999 13588
rect 18865 13628 18951 13651
rect 19033 13628 19119 13651
rect 18865 13588 18890 13628
rect 18890 13588 18930 13628
rect 18930 13588 18951 13628
rect 19033 13588 19054 13628
rect 19054 13588 19094 13628
rect 19094 13588 19119 13628
rect 18865 13565 18951 13588
rect 19033 13565 19119 13588
rect 4985 12872 5071 12895
rect 5153 12872 5239 12895
rect 4985 12832 5010 12872
rect 5010 12832 5050 12872
rect 5050 12832 5071 12872
rect 5153 12832 5174 12872
rect 5174 12832 5214 12872
rect 5214 12832 5239 12872
rect 4985 12809 5071 12832
rect 5153 12809 5239 12832
rect 20105 12872 20191 12895
rect 20273 12872 20359 12895
rect 20105 12832 20130 12872
rect 20130 12832 20170 12872
rect 20170 12832 20191 12872
rect 20273 12832 20294 12872
rect 20294 12832 20334 12872
rect 20334 12832 20359 12872
rect 20105 12809 20191 12832
rect 20273 12809 20359 12832
rect 3745 12116 3831 12139
rect 3913 12116 3999 12139
rect 18865 12116 18951 12139
rect 19033 12116 19119 12139
rect 3745 12076 3770 12116
rect 3770 12076 3810 12116
rect 3810 12076 3831 12116
rect 3913 12076 3934 12116
rect 3934 12076 3974 12116
rect 3974 12076 3999 12116
rect 18865 12076 18890 12116
rect 18890 12076 18930 12116
rect 18930 12076 18951 12116
rect 19033 12076 19054 12116
rect 19054 12076 19094 12116
rect 19094 12076 19119 12116
rect 3745 12053 3831 12076
rect 3913 12053 3999 12076
rect 18865 12053 18951 12076
rect 19033 12053 19119 12076
rect 4985 11360 5071 11383
rect 5153 11360 5239 11383
rect 4985 11320 5010 11360
rect 5010 11320 5050 11360
rect 5050 11320 5071 11360
rect 5153 11320 5174 11360
rect 5174 11320 5214 11360
rect 5214 11320 5239 11360
rect 4985 11297 5071 11320
rect 5153 11297 5239 11320
rect 20105 11360 20191 11383
rect 20273 11360 20359 11383
rect 20105 11320 20130 11360
rect 20130 11320 20170 11360
rect 20170 11320 20191 11360
rect 20273 11320 20294 11360
rect 20294 11320 20334 11360
rect 20334 11320 20359 11360
rect 20105 11297 20191 11320
rect 20273 11297 20359 11320
rect 3745 10604 3831 10627
rect 3913 10604 3999 10627
rect 3745 10564 3770 10604
rect 3770 10564 3810 10604
rect 3810 10564 3831 10604
rect 3913 10564 3934 10604
rect 3934 10564 3974 10604
rect 3974 10564 3999 10604
rect 3745 10541 3831 10564
rect 3913 10541 3999 10564
rect 18865 10604 18951 10627
rect 19033 10604 19119 10627
rect 18865 10564 18890 10604
rect 18890 10564 18930 10604
rect 18930 10564 18951 10604
rect 19033 10564 19054 10604
rect 19054 10564 19094 10604
rect 19094 10564 19119 10604
rect 18865 10541 18951 10564
rect 19033 10541 19119 10564
rect 4985 9848 5071 9871
rect 5153 9848 5239 9871
rect 4985 9808 5010 9848
rect 5010 9808 5050 9848
rect 5050 9808 5071 9848
rect 5153 9808 5174 9848
rect 5174 9808 5214 9848
rect 5214 9808 5239 9848
rect 4985 9785 5071 9808
rect 5153 9785 5239 9808
rect 20105 9848 20191 9871
rect 20273 9848 20359 9871
rect 20105 9808 20130 9848
rect 20130 9808 20170 9848
rect 20170 9808 20191 9848
rect 20273 9808 20294 9848
rect 20294 9808 20334 9848
rect 20334 9808 20359 9848
rect 20105 9785 20191 9808
rect 20273 9785 20359 9808
rect 3745 9092 3831 9115
rect 3913 9092 3999 9115
rect 3745 9052 3770 9092
rect 3770 9052 3810 9092
rect 3810 9052 3831 9092
rect 3913 9052 3934 9092
rect 3934 9052 3974 9092
rect 3974 9052 3999 9092
rect 3745 9029 3831 9052
rect 3913 9029 3999 9052
rect 18865 9092 18951 9115
rect 19033 9092 19119 9115
rect 18865 9052 18890 9092
rect 18890 9052 18930 9092
rect 18930 9052 18951 9092
rect 19033 9052 19054 9092
rect 19054 9052 19094 9092
rect 19094 9052 19119 9092
rect 18865 9029 18951 9052
rect 19033 9029 19119 9052
rect 4985 8336 5071 8359
rect 5153 8336 5239 8359
rect 20105 8336 20191 8359
rect 20273 8336 20359 8359
rect 4985 8296 5010 8336
rect 5010 8296 5050 8336
rect 5050 8296 5071 8336
rect 5153 8296 5174 8336
rect 5174 8296 5214 8336
rect 5214 8296 5239 8336
rect 20105 8296 20130 8336
rect 20130 8296 20170 8336
rect 20170 8296 20191 8336
rect 20273 8296 20294 8336
rect 20294 8296 20334 8336
rect 20334 8296 20359 8336
rect 4985 8273 5071 8296
rect 5153 8273 5239 8296
rect 20105 8273 20191 8296
rect 20273 8273 20359 8296
rect 3745 7580 3831 7603
rect 3913 7580 3999 7603
rect 3745 7540 3770 7580
rect 3770 7540 3810 7580
rect 3810 7540 3831 7580
rect 3913 7540 3934 7580
rect 3934 7540 3974 7580
rect 3974 7540 3999 7580
rect 3745 7517 3831 7540
rect 3913 7517 3999 7540
rect 18865 7580 18951 7603
rect 19033 7580 19119 7603
rect 18865 7540 18890 7580
rect 18890 7540 18930 7580
rect 18930 7540 18951 7580
rect 19033 7540 19054 7580
rect 19054 7540 19094 7580
rect 19094 7540 19119 7580
rect 18865 7517 18951 7540
rect 19033 7517 19119 7540
rect 4985 6824 5071 6847
rect 5153 6824 5239 6847
rect 4985 6784 5010 6824
rect 5010 6784 5050 6824
rect 5050 6784 5071 6824
rect 5153 6784 5174 6824
rect 5174 6784 5214 6824
rect 5214 6784 5239 6824
rect 4985 6761 5071 6784
rect 5153 6761 5239 6784
rect 20105 6824 20191 6847
rect 20273 6824 20359 6847
rect 20105 6784 20130 6824
rect 20130 6784 20170 6824
rect 20170 6784 20191 6824
rect 20273 6784 20294 6824
rect 20294 6784 20334 6824
rect 20334 6784 20359 6824
rect 20105 6761 20191 6784
rect 20273 6761 20359 6784
rect 17157 6257 17243 6343
rect 3745 6068 3831 6091
rect 3913 6068 3999 6091
rect 3745 6028 3770 6068
rect 3770 6028 3810 6068
rect 3810 6028 3831 6068
rect 3913 6028 3934 6068
rect 3934 6028 3974 6068
rect 3974 6028 3999 6068
rect 3745 6005 3831 6028
rect 3913 6005 3999 6028
rect 18865 6068 18951 6091
rect 19033 6068 19119 6091
rect 18865 6028 18890 6068
rect 18890 6028 18930 6068
rect 18930 6028 18951 6068
rect 19033 6028 19054 6068
rect 19054 6028 19094 6068
rect 19094 6028 19119 6068
rect 18865 6005 18951 6028
rect 19033 6005 19119 6028
rect 285 5585 371 5671
rect 1197 5333 1283 5419
rect 4985 5312 5071 5335
rect 5153 5312 5239 5335
rect 4985 5272 5010 5312
rect 5010 5272 5050 5312
rect 5050 5272 5071 5312
rect 5153 5272 5174 5312
rect 5174 5272 5214 5312
rect 5214 5272 5239 5312
rect 4985 5249 5071 5272
rect 5153 5249 5239 5272
rect 20105 5312 20191 5335
rect 20273 5312 20359 5335
rect 20105 5272 20130 5312
rect 20130 5272 20170 5312
rect 20170 5272 20191 5312
rect 20273 5272 20294 5312
rect 20294 5272 20334 5312
rect 20334 5272 20359 5312
rect 20105 5249 20191 5272
rect 20273 5249 20359 5272
rect 3745 4556 3831 4579
rect 3913 4556 3999 4579
rect 3745 4516 3770 4556
rect 3770 4516 3810 4556
rect 3810 4516 3831 4556
rect 3913 4516 3934 4556
rect 3934 4516 3974 4556
rect 3974 4516 3999 4556
rect 3745 4493 3831 4516
rect 3913 4493 3999 4516
rect 18865 4556 18951 4579
rect 19033 4556 19119 4579
rect 18865 4516 18890 4556
rect 18890 4516 18930 4556
rect 18930 4516 18951 4556
rect 19033 4516 19054 4556
rect 19054 4516 19094 4556
rect 19094 4516 19119 4556
rect 18865 4493 18951 4516
rect 19033 4493 19119 4516
rect 4985 3800 5071 3823
rect 5153 3800 5239 3823
rect 20105 3800 20191 3823
rect 20273 3800 20359 3823
rect 4985 3760 5010 3800
rect 5010 3760 5050 3800
rect 5050 3760 5071 3800
rect 5153 3760 5174 3800
rect 5174 3760 5214 3800
rect 5214 3760 5239 3800
rect 20105 3760 20130 3800
rect 20130 3760 20170 3800
rect 20170 3760 20191 3800
rect 20273 3760 20294 3800
rect 20294 3760 20334 3800
rect 20334 3760 20359 3800
rect 4985 3737 5071 3760
rect 5153 3737 5239 3760
rect 20105 3737 20191 3760
rect 20273 3737 20359 3760
rect 3745 3044 3831 3067
rect 3913 3044 3999 3067
rect 3745 3004 3770 3044
rect 3770 3004 3810 3044
rect 3810 3004 3831 3044
rect 3913 3004 3934 3044
rect 3934 3004 3974 3044
rect 3974 3004 3999 3044
rect 3745 2981 3831 3004
rect 3913 2981 3999 3004
rect 12141 2981 12227 3067
rect 18865 3044 18951 3067
rect 19033 3044 19119 3067
rect 18865 3004 18890 3044
rect 18890 3004 18930 3044
rect 18930 3004 18951 3044
rect 19033 3004 19054 3044
rect 19054 3004 19094 3044
rect 19094 3004 19119 3044
rect 18865 2981 18951 3004
rect 19033 2981 19119 3004
rect 10317 2393 10403 2479
rect 4985 2288 5071 2311
rect 5153 2288 5239 2311
rect 4985 2248 5010 2288
rect 5010 2248 5050 2288
rect 5050 2248 5071 2288
rect 5153 2248 5174 2288
rect 5174 2248 5214 2288
rect 5214 2248 5239 2288
rect 4985 2225 5071 2248
rect 5153 2225 5239 2248
rect 20105 2288 20191 2311
rect 20273 2288 20359 2311
rect 20105 2248 20130 2288
rect 20130 2248 20170 2288
rect 20170 2248 20191 2288
rect 20273 2248 20294 2288
rect 20294 2248 20334 2288
rect 20334 2248 20359 2288
rect 20105 2225 20191 2248
rect 20273 2225 20359 2248
rect 9405 2057 9491 2143
rect 3745 1532 3831 1555
rect 3913 1532 3999 1555
rect 3745 1492 3770 1532
rect 3770 1492 3810 1532
rect 3810 1492 3831 1532
rect 3913 1492 3934 1532
rect 3934 1492 3974 1532
rect 3974 1492 3999 1532
rect 3745 1469 3831 1492
rect 3913 1469 3999 1492
rect 18865 1532 18951 1555
rect 19033 1532 19119 1555
rect 18865 1492 18890 1532
rect 18890 1492 18930 1532
rect 18930 1492 18951 1532
rect 19033 1492 19054 1532
rect 19054 1492 19094 1532
rect 19094 1492 19119 1532
rect 18865 1469 18951 1492
rect 19033 1469 19119 1492
rect 8493 1280 8579 1303
rect 8493 1240 8524 1280
rect 8524 1240 8564 1280
rect 8564 1240 8579 1280
rect 8493 1217 8579 1240
rect 13509 1217 13595 1303
rect 14421 881 14507 967
rect 2109 713 2195 799
rect 4985 776 5071 799
rect 5153 776 5239 799
rect 15789 797 15875 883
rect 4985 736 5010 776
rect 5010 736 5050 776
rect 5050 736 5071 776
rect 5153 736 5174 776
rect 5174 736 5214 776
rect 5214 736 5239 776
rect 4985 713 5071 736
rect 5153 713 5239 736
rect 20105 776 20191 799
rect 20273 776 20359 799
rect 20105 736 20130 776
rect 20130 736 20170 776
rect 20170 736 20191 776
rect 20273 736 20294 776
rect 20294 736 20334 776
rect 20334 736 20359 776
rect 20105 713 20191 736
rect 20273 713 20359 736
rect 7125 293 7211 379
rect 285 188 371 211
rect 285 148 308 188
rect 308 148 371 188
rect 285 125 371 148
<< metal6 >>
rect 3652 40867 4092 43008
rect 3652 40781 3745 40867
rect 3831 40781 3913 40867
rect 3999 40781 4092 40867
rect 3652 39355 4092 40781
rect 3652 39269 3745 39355
rect 3831 39269 3913 39355
rect 3999 39269 4092 39355
rect 3652 37843 4092 39269
rect 3652 37757 3745 37843
rect 3831 37757 3913 37843
rect 3999 37757 4092 37843
rect 3652 36331 4092 37757
rect 3652 36245 3745 36331
rect 3831 36245 3913 36331
rect 3999 36245 4092 36331
rect 1076 35323 1404 35444
rect 1076 35237 1197 35323
rect 1283 35237 1404 35323
rect 164 5671 492 5792
rect 164 5585 285 5671
rect 371 5585 492 5671
rect 164 211 492 5585
rect 1076 5419 1404 35237
rect 3652 34819 4092 36245
rect 3652 34733 3745 34819
rect 3831 34733 3913 34819
rect 3999 34733 4092 34819
rect 3652 33307 4092 34733
rect 3652 33221 3745 33307
rect 3831 33221 3913 33307
rect 3999 33221 4092 33307
rect 3652 31795 4092 33221
rect 3652 31709 3745 31795
rect 3831 31709 3913 31795
rect 3999 31709 4092 31795
rect 3652 30283 4092 31709
rect 3652 30197 3745 30283
rect 3831 30197 3913 30283
rect 3999 30197 4092 30283
rect 3652 28771 4092 30197
rect 3652 28685 3745 28771
rect 3831 28685 3913 28771
rect 3999 28685 4092 28771
rect 1076 5333 1197 5419
rect 1283 5333 1404 5419
rect 1076 5212 1404 5333
rect 1988 27763 2316 27884
rect 1988 27677 2109 27763
rect 2195 27677 2316 27763
rect 1988 799 2316 27677
rect 1988 713 2109 799
rect 2195 713 2316 799
rect 1988 592 2316 713
rect 3652 27259 4092 28685
rect 3652 27173 3745 27259
rect 3831 27173 3913 27259
rect 3999 27173 4092 27259
rect 3652 25747 4092 27173
rect 3652 25661 3745 25747
rect 3831 25661 3913 25747
rect 3999 25661 4092 25747
rect 3652 24235 4092 25661
rect 3652 24149 3745 24235
rect 3831 24149 3913 24235
rect 3999 24149 4092 24235
rect 3652 22723 4092 24149
rect 3652 22637 3745 22723
rect 3831 22637 3913 22723
rect 3999 22637 4092 22723
rect 3652 21211 4092 22637
rect 3652 21125 3745 21211
rect 3831 21125 3913 21211
rect 3999 21125 4092 21211
rect 3652 19699 4092 21125
rect 3652 19613 3745 19699
rect 3831 19613 3913 19699
rect 3999 19613 4092 19699
rect 3652 18187 4092 19613
rect 3652 18101 3745 18187
rect 3831 18101 3913 18187
rect 3999 18101 4092 18187
rect 3652 16675 4092 18101
rect 3652 16589 3745 16675
rect 3831 16589 3913 16675
rect 3999 16589 4092 16675
rect 3652 15163 4092 16589
rect 3652 15077 3745 15163
rect 3831 15077 3913 15163
rect 3999 15077 4092 15163
rect 3652 13651 4092 15077
rect 3652 13565 3745 13651
rect 3831 13565 3913 13651
rect 3999 13565 4092 13651
rect 3652 12139 4092 13565
rect 3652 12053 3745 12139
rect 3831 12053 3913 12139
rect 3999 12053 4092 12139
rect 3652 10627 4092 12053
rect 3652 10541 3745 10627
rect 3831 10541 3913 10627
rect 3999 10541 4092 10627
rect 3652 9115 4092 10541
rect 3652 9029 3745 9115
rect 3831 9029 3913 9115
rect 3999 9029 4092 9115
rect 3652 7603 4092 9029
rect 3652 7517 3745 7603
rect 3831 7517 3913 7603
rect 3999 7517 4092 7603
rect 3652 6091 4092 7517
rect 3652 6005 3745 6091
rect 3831 6005 3913 6091
rect 3999 6005 4092 6091
rect 3652 4579 4092 6005
rect 3652 4493 3745 4579
rect 3831 4493 3913 4579
rect 3999 4493 4092 4579
rect 3652 3067 4092 4493
rect 3652 2981 3745 3067
rect 3831 2981 3913 3067
rect 3999 2981 4092 3067
rect 3652 1555 4092 2981
rect 3652 1469 3745 1555
rect 3831 1469 3913 1555
rect 3999 1469 4092 1555
rect 164 125 285 211
rect 371 125 492 211
rect 164 4 492 125
rect 3652 0 4092 1469
rect 4892 41623 5332 43008
rect 4892 41537 4985 41623
rect 5071 41537 5153 41623
rect 5239 41537 5332 41623
rect 4892 40111 5332 41537
rect 17036 41035 17364 41156
rect 17036 40949 17157 41035
rect 17243 40949 17364 41035
rect 4892 40025 4985 40111
rect 5071 40025 5153 40111
rect 5239 40025 5332 40111
rect 4892 38599 5332 40025
rect 14300 40363 14628 40484
rect 14300 40277 14421 40363
rect 14507 40277 14628 40363
rect 4892 38513 4985 38599
rect 5071 38513 5153 38599
rect 5239 38513 5332 38599
rect 4892 37087 5332 38513
rect 13388 39439 13716 39560
rect 13388 39353 13509 39439
rect 13595 39353 13716 39439
rect 4892 37001 4985 37087
rect 5071 37001 5153 37087
rect 5239 37001 5332 37087
rect 4892 35575 5332 37001
rect 4892 35489 4985 35575
rect 5071 35489 5153 35575
rect 5239 35489 5332 35575
rect 4892 34063 5332 35489
rect 4892 33977 4985 34063
rect 5071 33977 5153 34063
rect 5239 33977 5332 34063
rect 4892 32551 5332 33977
rect 4892 32465 4985 32551
rect 5071 32465 5153 32551
rect 5239 32465 5332 32551
rect 4892 31039 5332 32465
rect 4892 30953 4985 31039
rect 5071 30953 5153 31039
rect 5239 30953 5332 31039
rect 4892 29527 5332 30953
rect 4892 29441 4985 29527
rect 5071 29441 5153 29527
rect 5239 29441 5332 29527
rect 4892 28015 5332 29441
rect 4892 27929 4985 28015
rect 5071 27929 5153 28015
rect 5239 27929 5332 28015
rect 4892 26503 5332 27929
rect 4892 26417 4985 26503
rect 5071 26417 5153 26503
rect 5239 26417 5332 26503
rect 4892 24991 5332 26417
rect 4892 24905 4985 24991
rect 5071 24905 5153 24991
rect 5239 24905 5332 24991
rect 4892 23479 5332 24905
rect 4892 23393 4985 23479
rect 5071 23393 5153 23479
rect 5239 23393 5332 23479
rect 4892 21967 5332 23393
rect 4892 21881 4985 21967
rect 5071 21881 5153 21967
rect 5239 21881 5332 21967
rect 4892 20455 5332 21881
rect 4892 20369 4985 20455
rect 5071 20369 5153 20455
rect 5239 20369 5332 20455
rect 4892 18943 5332 20369
rect 4892 18857 4985 18943
rect 5071 18857 5153 18943
rect 5239 18857 5332 18943
rect 4892 17431 5332 18857
rect 4892 17345 4985 17431
rect 5071 17345 5153 17431
rect 5239 17345 5332 17431
rect 4892 15919 5332 17345
rect 4892 15833 4985 15919
rect 5071 15833 5153 15919
rect 5239 15833 5332 15919
rect 4892 14407 5332 15833
rect 4892 14321 4985 14407
rect 5071 14321 5153 14407
rect 5239 14321 5332 14407
rect 4892 12895 5332 14321
rect 4892 12809 4985 12895
rect 5071 12809 5153 12895
rect 5239 12809 5332 12895
rect 4892 11383 5332 12809
rect 4892 11297 4985 11383
rect 5071 11297 5153 11383
rect 5239 11297 5332 11383
rect 4892 9871 5332 11297
rect 4892 9785 4985 9871
rect 5071 9785 5153 9871
rect 5239 9785 5332 9871
rect 4892 8359 5332 9785
rect 4892 8273 4985 8359
rect 5071 8273 5153 8359
rect 5239 8273 5332 8359
rect 4892 6847 5332 8273
rect 4892 6761 4985 6847
rect 5071 6761 5153 6847
rect 5239 6761 5332 6847
rect 4892 5335 5332 6761
rect 4892 5249 4985 5335
rect 5071 5249 5153 5335
rect 5239 5249 5332 5335
rect 4892 3823 5332 5249
rect 4892 3737 4985 3823
rect 5071 3737 5153 3823
rect 5239 3737 5332 3823
rect 4892 2311 5332 3737
rect 4892 2225 4985 2311
rect 5071 2225 5153 2311
rect 5239 2225 5332 2311
rect 4892 799 5332 2225
rect 4892 713 4985 799
rect 5071 713 5153 799
rect 5239 713 5332 799
rect 4892 0 5332 713
rect 7004 38347 7332 38468
rect 7004 38261 7125 38347
rect 7211 38261 7332 38347
rect 7004 379 7332 38261
rect 9284 36331 9612 36452
rect 9284 36245 9405 36331
rect 9491 36245 9612 36331
rect 8372 21463 8700 21584
rect 8372 21377 8493 21463
rect 8579 21377 8700 21463
rect 8372 1303 8700 21377
rect 9284 2143 9612 36245
rect 12020 31375 12348 31496
rect 12020 31289 12141 31375
rect 12227 31289 12348 31375
rect 10196 31123 10524 31244
rect 10196 31037 10317 31123
rect 10403 31037 10524 31123
rect 10196 2479 10524 31037
rect 12020 3067 12348 31289
rect 13388 15415 13716 39353
rect 13388 15329 13509 15415
rect 13595 15329 13716 15415
rect 13388 15208 13716 15329
rect 12020 2981 12141 3067
rect 12227 2981 12348 3067
rect 12020 2860 12348 2981
rect 13388 14743 13716 14864
rect 13388 14657 13509 14743
rect 13595 14657 13716 14743
rect 10196 2393 10317 2479
rect 10403 2393 10524 2479
rect 10196 2272 10524 2393
rect 9284 2057 9405 2143
rect 9491 2057 9612 2143
rect 9284 1936 9612 2057
rect 8372 1217 8493 1303
rect 8579 1217 8700 1303
rect 8372 1096 8700 1217
rect 13388 1303 13716 14657
rect 13388 1217 13509 1303
rect 13595 1217 13716 1303
rect 13388 1096 13716 1217
rect 14300 967 14628 40277
rect 14300 881 14421 967
rect 14507 881 14628 967
rect 14300 760 14628 881
rect 15668 35491 15996 35612
rect 15668 35405 15789 35491
rect 15875 35405 15996 35491
rect 15668 883 15996 35405
rect 17036 6343 17364 40949
rect 17036 6257 17157 6343
rect 17243 6257 17364 6343
rect 17036 6136 17364 6257
rect 18772 40867 19212 43008
rect 18772 40781 18865 40867
rect 18951 40781 19033 40867
rect 19119 40781 19212 40867
rect 18772 39355 19212 40781
rect 18772 39269 18865 39355
rect 18951 39269 19033 39355
rect 19119 39269 19212 39355
rect 18772 37843 19212 39269
rect 18772 37757 18865 37843
rect 18951 37757 19033 37843
rect 19119 37757 19212 37843
rect 18772 36331 19212 37757
rect 18772 36245 18865 36331
rect 18951 36245 19033 36331
rect 19119 36245 19212 36331
rect 18772 34819 19212 36245
rect 18772 34733 18865 34819
rect 18951 34733 19033 34819
rect 19119 34733 19212 34819
rect 18772 33307 19212 34733
rect 18772 33221 18865 33307
rect 18951 33221 19033 33307
rect 19119 33221 19212 33307
rect 18772 31795 19212 33221
rect 18772 31709 18865 31795
rect 18951 31709 19033 31795
rect 19119 31709 19212 31795
rect 18772 30283 19212 31709
rect 18772 30197 18865 30283
rect 18951 30197 19033 30283
rect 19119 30197 19212 30283
rect 18772 28771 19212 30197
rect 18772 28685 18865 28771
rect 18951 28685 19033 28771
rect 19119 28685 19212 28771
rect 18772 27259 19212 28685
rect 18772 27173 18865 27259
rect 18951 27173 19033 27259
rect 19119 27173 19212 27259
rect 18772 25747 19212 27173
rect 18772 25661 18865 25747
rect 18951 25661 19033 25747
rect 19119 25661 19212 25747
rect 18772 24235 19212 25661
rect 18772 24149 18865 24235
rect 18951 24149 19033 24235
rect 19119 24149 19212 24235
rect 18772 22723 19212 24149
rect 18772 22637 18865 22723
rect 18951 22637 19033 22723
rect 19119 22637 19212 22723
rect 18772 21211 19212 22637
rect 18772 21125 18865 21211
rect 18951 21125 19033 21211
rect 19119 21125 19212 21211
rect 18772 19699 19212 21125
rect 18772 19613 18865 19699
rect 18951 19613 19033 19699
rect 19119 19613 19212 19699
rect 18772 18187 19212 19613
rect 18772 18101 18865 18187
rect 18951 18101 19033 18187
rect 19119 18101 19212 18187
rect 18772 16675 19212 18101
rect 18772 16589 18865 16675
rect 18951 16589 19033 16675
rect 19119 16589 19212 16675
rect 18772 15163 19212 16589
rect 18772 15077 18865 15163
rect 18951 15077 19033 15163
rect 19119 15077 19212 15163
rect 18772 13651 19212 15077
rect 18772 13565 18865 13651
rect 18951 13565 19033 13651
rect 19119 13565 19212 13651
rect 18772 12139 19212 13565
rect 18772 12053 18865 12139
rect 18951 12053 19033 12139
rect 19119 12053 19212 12139
rect 18772 10627 19212 12053
rect 18772 10541 18865 10627
rect 18951 10541 19033 10627
rect 19119 10541 19212 10627
rect 18772 9115 19212 10541
rect 18772 9029 18865 9115
rect 18951 9029 19033 9115
rect 19119 9029 19212 9115
rect 18772 7603 19212 9029
rect 18772 7517 18865 7603
rect 18951 7517 19033 7603
rect 19119 7517 19212 7603
rect 15668 797 15789 883
rect 15875 797 15996 883
rect 15668 676 15996 797
rect 18772 6091 19212 7517
rect 18772 6005 18865 6091
rect 18951 6005 19033 6091
rect 19119 6005 19212 6091
rect 18772 4579 19212 6005
rect 18772 4493 18865 4579
rect 18951 4493 19033 4579
rect 19119 4493 19212 4579
rect 18772 3067 19212 4493
rect 18772 2981 18865 3067
rect 18951 2981 19033 3067
rect 19119 2981 19212 3067
rect 18772 1555 19212 2981
rect 18772 1469 18865 1555
rect 18951 1469 19033 1555
rect 19119 1469 19212 1555
rect 7004 293 7125 379
rect 7211 293 7332 379
rect 7004 172 7332 293
rect 18772 0 19212 1469
rect 20012 41623 20452 43008
rect 20012 41537 20105 41623
rect 20191 41537 20273 41623
rect 20359 41537 20452 41623
rect 20012 40111 20452 41537
rect 20012 40025 20105 40111
rect 20191 40025 20273 40111
rect 20359 40025 20452 40111
rect 20012 38599 20452 40025
rect 20012 38513 20105 38599
rect 20191 38513 20273 38599
rect 20359 38513 20452 38599
rect 20012 37087 20452 38513
rect 20012 37001 20105 37087
rect 20191 37001 20273 37087
rect 20359 37001 20452 37087
rect 20012 35575 20452 37001
rect 20012 35489 20105 35575
rect 20191 35489 20273 35575
rect 20359 35489 20452 35575
rect 20012 34063 20452 35489
rect 20012 33977 20105 34063
rect 20191 33977 20273 34063
rect 20359 33977 20452 34063
rect 20012 32551 20452 33977
rect 20012 32465 20105 32551
rect 20191 32465 20273 32551
rect 20359 32465 20452 32551
rect 20012 31039 20452 32465
rect 20012 30953 20105 31039
rect 20191 30953 20273 31039
rect 20359 30953 20452 31039
rect 20012 29527 20452 30953
rect 20012 29441 20105 29527
rect 20191 29441 20273 29527
rect 20359 29441 20452 29527
rect 20012 28015 20452 29441
rect 20012 27929 20105 28015
rect 20191 27929 20273 28015
rect 20359 27929 20452 28015
rect 20012 26503 20452 27929
rect 20012 26417 20105 26503
rect 20191 26417 20273 26503
rect 20359 26417 20452 26503
rect 20012 24991 20452 26417
rect 20012 24905 20105 24991
rect 20191 24905 20273 24991
rect 20359 24905 20452 24991
rect 20012 23479 20452 24905
rect 20012 23393 20105 23479
rect 20191 23393 20273 23479
rect 20359 23393 20452 23479
rect 20012 21967 20452 23393
rect 20012 21881 20105 21967
rect 20191 21881 20273 21967
rect 20359 21881 20452 21967
rect 20012 20455 20452 21881
rect 20012 20369 20105 20455
rect 20191 20369 20273 20455
rect 20359 20369 20452 20455
rect 20012 18943 20452 20369
rect 20012 18857 20105 18943
rect 20191 18857 20273 18943
rect 20359 18857 20452 18943
rect 20012 17431 20452 18857
rect 20012 17345 20105 17431
rect 20191 17345 20273 17431
rect 20359 17345 20452 17431
rect 20012 15919 20452 17345
rect 20012 15833 20105 15919
rect 20191 15833 20273 15919
rect 20359 15833 20452 15919
rect 20012 14407 20452 15833
rect 20012 14321 20105 14407
rect 20191 14321 20273 14407
rect 20359 14321 20452 14407
rect 20012 12895 20452 14321
rect 20012 12809 20105 12895
rect 20191 12809 20273 12895
rect 20359 12809 20452 12895
rect 20012 11383 20452 12809
rect 20012 11297 20105 11383
rect 20191 11297 20273 11383
rect 20359 11297 20452 11383
rect 20012 9871 20452 11297
rect 20012 9785 20105 9871
rect 20191 9785 20273 9871
rect 20359 9785 20452 9871
rect 20012 8359 20452 9785
rect 20012 8273 20105 8359
rect 20191 8273 20273 8359
rect 20359 8273 20452 8359
rect 20012 6847 20452 8273
rect 20012 6761 20105 6847
rect 20191 6761 20273 6847
rect 20359 6761 20452 6847
rect 20012 5335 20452 6761
rect 20012 5249 20105 5335
rect 20191 5249 20273 5335
rect 20359 5249 20452 5335
rect 20012 3823 20452 5249
rect 20012 3737 20105 3823
rect 20191 3737 20273 3823
rect 20359 3737 20452 3823
rect 20012 2311 20452 3737
rect 20012 2225 20105 2311
rect 20191 2225 20273 2311
rect 20359 2225 20452 2311
rect 20012 799 20452 2225
rect 20012 713 20105 799
rect 20191 713 20273 799
rect 20359 713 20452 799
rect 20012 0 20452 713
use sg13g2_inv_1  _0381_
timestamp 1676382929
transform 1 0 1152 0 -1 32508
box -48 -56 336 834
use sg13g2_inv_1  _0382_
timestamp 1676382929
transform 1 0 6144 0 -1 29484
box -48 -56 336 834
use sg13g2_inv_1  _0383_
timestamp 1676382929
transform 1 0 8640 0 1 26460
box -48 -56 336 834
use sg13g2_inv_1  _0384_
timestamp 1676382929
transform -1 0 5856 0 1 24948
box -48 -56 336 834
use sg13g2_inv_1  _0385_
timestamp 1676382929
transform 1 0 5760 0 -1 37044
box -48 -56 336 834
use sg13g2_inv_1  _0386_
timestamp 1676382929
transform 1 0 11712 0 -1 26460
box -48 -56 336 834
use sg13g2_inv_1  _0387_
timestamp 1676382929
transform 1 0 20064 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _0388_
timestamp 1676382929
transform 1 0 13248 0 -1 29484
box -48 -56 336 834
use sg13g2_inv_1  _0389_
timestamp 1676382929
transform 1 0 20064 0 1 21924
box -48 -56 336 834
use sg13g2_inv_1  _0390_
timestamp 1676382929
transform -1 0 3072 0 1 11340
box -48 -56 336 834
use sg13g2_inv_1  _0391_
timestamp 1676382929
transform 1 0 11424 0 -1 23436
box -48 -56 336 834
use sg13g2_inv_1  _0392_
timestamp 1676382929
transform -1 0 1440 0 -1 26460
box -48 -56 336 834
use sg13g2_inv_1  _0393_
timestamp 1676382929
transform -1 0 13920 0 1 26460
box -48 -56 336 834
use sg13g2_inv_1  _0394_
timestamp 1676382929
transform 1 0 17184 0 1 26460
box -48 -56 336 834
use sg13g2_inv_1  _0395_
timestamp 1676382929
transform 1 0 2784 0 -1 20412
box -48 -56 336 834
use sg13g2_inv_1  _0396_
timestamp 1676382929
transform -1 0 10368 0 -1 41580
box -48 -56 336 834
use sg13g2_inv_1  _0397_
timestamp 1676382929
transform -1 0 14496 0 1 26460
box -48 -56 336 834
use sg13g2_inv_1  _0398_
timestamp 1676382929
transform -1 0 6624 0 1 23436
box -48 -56 336 834
use sg13g2_inv_1  _0399_
timestamp 1676382929
transform -1 0 2016 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  _0400_
timestamp 1676382929
transform -1 0 5472 0 -1 40068
box -48 -56 336 834
use sg13g2_inv_1  _0401_
timestamp 1676382929
transform -1 0 14208 0 1 26460
box -48 -56 336 834
use sg13g2_inv_1  _0402_
timestamp 1676382929
transform 1 0 4320 0 1 20412
box -48 -56 336 834
use sg13g2_inv_1  _0403_
timestamp 1676382929
transform -1 0 15264 0 1 9828
box -48 -56 336 834
use sg13g2_inv_1  _0404_
timestamp 1676382929
transform -1 0 20352 0 1 6804
box -48 -56 336 834
use sg13g2_inv_1  _0405_
timestamp 1676382929
transform -1 0 20352 0 1 5292
box -48 -56 336 834
use sg13g2_inv_1  _0406_
timestamp 1676382929
transform 1 0 12960 0 -1 8316
box -48 -56 336 834
use sg13g2_inv_1  _0407_
timestamp 1676382929
transform -1 0 11712 0 -1 5292
box -48 -56 336 834
use sg13g2_inv_1  _0408_
timestamp 1676382929
transform -1 0 5664 0 -1 11340
box -48 -56 336 834
use sg13g2_inv_1  _0409_
timestamp 1676382929
transform -1 0 20352 0 -1 11340
box -48 -56 336 834
use sg13g2_inv_1  _0410_
timestamp 1676382929
transform 1 0 20064 0 1 8316
box -48 -56 336 834
use sg13g2_inv_1  _0411_
timestamp 1676382929
transform -1 0 4512 0 -1 3780
box -48 -56 336 834
use sg13g2_inv_1  _0412_
timestamp 1676382929
transform -1 0 10080 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  _0413_
timestamp 1676382929
transform -1 0 14304 0 -1 30996
box -48 -56 336 834
use sg13g2_inv_1  _0414_
timestamp 1676382929
transform -1 0 3168 0 1 32508
box -48 -56 336 834
use sg13g2_inv_1  _0415_
timestamp 1676382929
transform -1 0 10176 0 -1 38556
box -48 -56 336 834
use sg13g2_inv_1  _0416_
timestamp 1676382929
transform 1 0 18144 0 -1 35532
box -48 -56 336 834
use sg13g2_inv_1  _0417_
timestamp 1676382929
transform 1 0 2976 0 -1 24948
box -48 -56 336 834
use sg13g2_mux4_1  _0418_
timestamp 1677257233
transform 1 0 6048 0 -1 34020
box -48 -56 2064 834
use sg13g2_inv_1  _0419_
timestamp 1676382929
transform 1 0 14400 0 1 40068
box -48 -56 336 834
use sg13g2_nor2_1  _0420_
timestamp 1676627187
transform 1 0 3552 0 1 32508
box -48 -56 432 834
use sg13g2_mux4_1  _0421_
timestamp 1677257233
transform -1 0 7968 0 1 34020
box -48 -56 2064 834
use sg13g2_a21oi_1  _0422_
timestamp 1683973020
transform -1 0 4800 0 -1 35532
box -48 -56 528 834
use sg13g2_o21ai_1  _0423_
timestamp 1685175443
transform 1 0 6624 0 1 35532
box -48 -56 538 834
use sg13g2_o21ai_1  _0424_
timestamp 1685175443
transform 1 0 3936 0 1 32508
box -48 -56 538 834
use sg13g2_a22oi_1  _0425_
timestamp 1685173987
transform 1 0 9120 0 1 35532
box -48 -56 624 834
use sg13g2_nand3_1  _0426_
timestamp 1683988354
transform -1 0 10464 0 -1 34020
box -48 -56 528 834
use sg13g2_nand2b_1  _0427_
timestamp 1676567195
transform 1 0 7488 0 -1 40068
box -48 -56 528 834
use sg13g2_a22oi_1  _0428_
timestamp 1685173987
transform 1 0 8544 0 1 34020
box -48 -56 624 834
use sg13g2_nand2b_1  _0429_
timestamp 1676567195
transform -1 0 9312 0 1 37044
box -48 -56 528 834
use sg13g2_a21oi_1  _0430_
timestamp 1683973020
transform 1 0 6144 0 1 35532
box -48 -56 528 834
use sg13g2_nand2_1  _0431_
timestamp 1676557249
transform -1 0 8352 0 1 30996
box -48 -56 432 834
use sg13g2_o21ai_1  _0432_
timestamp 1685175443
transform 1 0 9984 0 1 32508
box -48 -56 538 834
use sg13g2_mux4_1  _0433_
timestamp 1677257233
transform 1 0 9120 0 -1 20412
box -48 -56 2064 834
use sg13g2_mux4_1  _0434_
timestamp 1677257233
transform 1 0 5472 0 -1 40068
box -48 -56 2064 834
use sg13g2_inv_1  _0435_
timestamp 1676382929
transform 1 0 5856 0 1 14364
box -48 -56 336 834
use sg13g2_nand3_1  _0436_
timestamp 1683988354
transform 1 0 5856 0 1 24948
box -48 -56 528 834
use sg13g2_mux2_1  _0437_
timestamp 1677247768
transform 1 0 5856 0 -1 26460
box -48 -56 1008 834
use sg13g2_nor2_1  _0438_
timestamp 1676627187
transform 1 0 3936 0 1 26460
box -48 -56 432 834
use sg13g2_a221oi_1  _0439_
timestamp 1685197497
transform -1 0 7584 0 -1 26460
box -48 -56 816 834
use sg13g2_mux2_1  _0440_
timestamp 1677247768
transform 1 0 4896 0 -1 26460
box -48 -56 1008 834
use sg13g2_a22oi_1  _0441_
timestamp 1685173987
transform 1 0 6048 0 1 26460
box -48 -56 624 834
use sg13g2_a22oi_1  _0442_
timestamp 1685173987
transform 1 0 6144 0 1 27972
box -48 -56 624 834
use sg13g2_mux4_1  _0443_
timestamp 1677257233
transform 1 0 11328 0 -1 35532
box -48 -56 2064 834
use sg13g2_mux4_1  _0444_
timestamp 1677257233
transform 1 0 9792 0 1 40068
box -48 -56 2064 834
use sg13g2_inv_1  _0445_
timestamp 1676382929
transform 1 0 14592 0 1 30996
box -48 -56 336 834
use sg13g2_nand3_1  _0446_
timestamp 1683988354
transform 1 0 19680 0 -1 30996
box -48 -56 528 834
use sg13g2_mux2_1  _0447_
timestamp 1677247768
transform 1 0 17472 0 1 32508
box -48 -56 1008 834
use sg13g2_nor2_1  _0448_
timestamp 1676627187
transform 1 0 19872 0 -1 40068
box -48 -56 432 834
use sg13g2_a221oi_1  _0449_
timestamp 1685197497
transform -1 0 19392 0 1 30996
box -48 -56 816 834
use sg13g2_mux2_1  _0450_
timestamp 1677247768
transform 1 0 17568 0 1 30996
box -48 -56 1008 834
use sg13g2_a22oi_1  _0451_
timestamp 1685173987
transform 1 0 19680 0 1 32508
box -48 -56 624 834
use sg13g2_a22oi_1  _0452_
timestamp 1685173987
transform -1 0 19968 0 1 30996
box -48 -56 624 834
use sg13g2_mux4_1  _0453_
timestamp 1677257233
transform 1 0 12000 0 1 24948
box -48 -56 2064 834
use sg13g2_mux4_1  _0454_
timestamp 1677257233
transform 1 0 7968 0 1 38556
box -48 -56 2064 834
use sg13g2_inv_1  _0455_
timestamp 1676382929
transform 1 0 17856 0 -1 8316
box -48 -56 336 834
use sg13g2_nand3_1  _0456_
timestamp 1683988354
transform 1 0 19776 0 -1 21924
box -48 -56 528 834
use sg13g2_mux2_1  _0457_
timestamp 1677247768
transform 1 0 17952 0 1 23436
box -48 -56 1008 834
use sg13g2_nor2_1  _0458_
timestamp 1676627187
transform 1 0 19968 0 -1 23436
box -48 -56 432 834
use sg13g2_a221oi_1  _0459_
timestamp 1685197497
transform -1 0 19680 0 1 23436
box -48 -56 816 834
use sg13g2_mux2_1  _0460_
timestamp 1677247768
transform 1 0 17472 0 1 21924
box -48 -56 1008 834
use sg13g2_a22oi_1  _0461_
timestamp 1685173987
transform 1 0 18624 0 -1 21924
box -48 -56 624 834
use sg13g2_a22oi_1  _0462_
timestamp 1685173987
transform -1 0 19776 0 -1 21924
box -48 -56 624 834
use sg13g2_mux4_1  _0463_
timestamp 1677257233
transform 1 0 9792 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _0464_
timestamp 1677257233
transform -1 0 6720 0 1 37044
box -48 -56 2064 834
use sg13g2_inv_1  _0465_
timestamp 1676382929
transform -1 0 5184 0 1 15876
box -48 -56 336 834
use sg13g2_nand3_1  _0466_
timestamp 1683988354
transform 1 0 9792 0 1 23436
box -48 -56 528 834
use sg13g2_mux2_1  _0467_
timestamp 1677247768
transform 1 0 10848 0 1 21924
box -48 -56 1008 834
use sg13g2_nor2_1  _0468_
timestamp 1676627187
transform -1 0 12192 0 1 21924
box -48 -56 432 834
use sg13g2_a221oi_1  _0469_
timestamp 1685197497
transform 1 0 10656 0 -1 23436
box -48 -56 816 834
use sg13g2_mux2_1  _0470_
timestamp 1677247768
transform -1 0 9792 0 1 23436
box -48 -56 1008 834
use sg13g2_a22oi_1  _0471_
timestamp 1685173987
transform 1 0 8640 0 1 21924
box -48 -56 624 834
use sg13g2_a22oi_1  _0472_
timestamp 1685173987
transform 1 0 9888 0 -1 21924
box -48 -56 624 834
use sg13g2_mux4_1  _0473_
timestamp 1677257233
transform 1 0 8928 0 1 18900
box -48 -56 2064 834
use sg13g2_mux4_1  _0474_
timestamp 1677257233
transform 1 0 7104 0 1 35532
box -48 -56 2064 834
use sg13g2_nand3_1  _0475_
timestamp 1683988354
transform 1 0 3744 0 -1 27972
box -48 -56 528 834
use sg13g2_mux2_1  _0476_
timestamp 1677247768
transform 1 0 2976 0 1 26460
box -48 -56 1008 834
use sg13g2_nor2_1  _0477_
timestamp 1676627187
transform -1 0 4896 0 -1 26460
box -48 -56 432 834
use sg13g2_a221oi_1  _0478_
timestamp 1685197497
transform 1 0 3168 0 -1 26460
box -48 -56 816 834
use sg13g2_mux2_1  _0479_
timestamp 1677247768
transform -1 0 3744 0 -1 27972
box -48 -56 1008 834
use sg13g2_a22oi_1  _0480_
timestamp 1685173987
transform 1 0 2976 0 1 24948
box -48 -56 624 834
use sg13g2_a22oi_1  _0481_
timestamp 1685173987
transform -1 0 4512 0 -1 26460
box -48 -56 624 834
use sg13g2_mux4_1  _0482_
timestamp 1677257233
transform 1 0 10944 0 -1 38556
box -48 -56 2064 834
use sg13g2_mux4_1  _0483_
timestamp 1677257233
transform 1 0 8352 0 -1 37044
box -48 -56 2064 834
use sg13g2_nand3_1  _0484_
timestamp 1683988354
transform 1 0 15744 0 -1 37044
box -48 -56 528 834
use sg13g2_mux2_1  _0485_
timestamp 1677247768
transform 1 0 14880 0 -1 35532
box -48 -56 1008 834
use sg13g2_nor2_1  _0486_
timestamp 1676627187
transform 1 0 10176 0 -1 38556
box -48 -56 432 834
use sg13g2_a221oi_1  _0487_
timestamp 1685197497
transform -1 0 17568 0 -1 35532
box -48 -56 816 834
use sg13g2_mux2_1  _0488_
timestamp 1677247768
transform -1 0 16800 0 -1 35532
box -48 -56 1008 834
use sg13g2_a22oi_1  _0489_
timestamp 1685173987
transform -1 0 15552 0 -1 37044
box -48 -56 624 834
use sg13g2_a22oi_1  _0490_
timestamp 1685173987
transform -1 0 18144 0 -1 35532
box -48 -56 624 834
use sg13g2_mux4_1  _0491_
timestamp 1677257233
transform 1 0 14496 0 -1 21924
box -48 -56 2064 834
use sg13g2_mux4_1  _0492_
timestamp 1677257233
transform 1 0 4128 0 1 35532
box -48 -56 2064 834
use sg13g2_nand3_1  _0493_
timestamp 1683988354
transform -1 0 17184 0 1 26460
box -48 -56 528 834
use sg13g2_mux2_1  _0494_
timestamp 1677247768
transform 1 0 15648 0 1 24948
box -48 -56 1008 834
use sg13g2_nor2_1  _0495_
timestamp 1676627187
transform -1 0 17664 0 -1 26460
box -48 -56 432 834
use sg13g2_a221oi_1  _0496_
timestamp 1685197497
transform -1 0 17280 0 -1 26460
box -48 -56 816 834
use sg13g2_mux2_1  _0497_
timestamp 1677247768
transform 1 0 15552 0 -1 26460
box -48 -56 1008 834
use sg13g2_a22oi_1  _0498_
timestamp 1685173987
transform 1 0 16128 0 1 26460
box -48 -56 624 834
use sg13g2_a22oi_1  _0499_
timestamp 1685173987
transform 1 0 16608 0 1 24948
box -48 -56 624 834
use sg13g2_mux4_1  _0500_
timestamp 1677257233
transform 1 0 10656 0 1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _0501_
timestamp 1677257233
transform 1 0 3840 0 1 38556
box -48 -56 2064 834
use sg13g2_nand3_1  _0502_
timestamp 1683988354
transform 1 0 3264 0 1 18900
box -48 -56 528 834
use sg13g2_mux2_1  _0503_
timestamp 1677247768
transform 1 0 3072 0 1 17388
box -48 -56 1008 834
use sg13g2_nor2_1  _0504_
timestamp 1676627187
transform 1 0 3744 0 -1 18900
box -48 -56 432 834
use sg13g2_a221oi_1  _0505_
timestamp 1685197497
transform -1 0 6144 0 -1 17388
box -48 -56 816 834
use sg13g2_mux2_1  _0506_
timestamp 1677247768
transform 1 0 1536 0 1 15876
box -48 -56 1008 834
use sg13g2_a22oi_1  _0507_
timestamp 1685173987
transform 1 0 4224 0 1 21924
box -48 -56 624 834
use sg13g2_a22oi_1  _0508_
timestamp 1685173987
transform -1 0 7968 0 1 18900
box -48 -56 624 834
use sg13g2_nor2_1  _0509_
timestamp 1676627187
transform -1 0 11232 0 1 27972
box -48 -56 432 834
use sg13g2_mux4_1  _0510_
timestamp 1677257233
transform 1 0 8160 0 1 17388
box -48 -56 2064 834
use sg13g2_nand3b_1  _0511_
timestamp 1676573470
transform 1 0 8640 0 -1 27972
box -48 -56 720 834
use sg13g2_and2_1  _0512_
timestamp 1676901763
transform 1 0 8928 0 1 26460
box -48 -56 528 834
use sg13g2_a21oi_1  _0513_
timestamp 1683973020
transform -1 0 8640 0 -1 27972
box -48 -56 528 834
use sg13g2_nand2b_1  _0514_
timestamp 1676567195
transform 1 0 9312 0 -1 27972
box -48 -56 528 834
use sg13g2_mux4_1  _0515_
timestamp 1677257233
transform 1 0 6624 0 1 26460
box -48 -56 2064 834
use sg13g2_nor2_1  _0516_
timestamp 1676627187
transform 1 0 6240 0 -1 24948
box -48 -56 432 834
use sg13g2_a21oi_1  _0517_
timestamp 1683973020
transform 1 0 9408 0 1 26460
box -48 -56 528 834
use sg13g2_mux4_1  _0518_
timestamp 1677257233
transform 1 0 10656 0 1 38556
box -48 -56 2064 834
use sg13g2_nand3_1  _0519_
timestamp 1683988354
transform -1 0 19872 0 1 35532
box -48 -56 528 834
use sg13g2_mux2_1  _0520_
timestamp 1677247768
transform 1 0 18240 0 -1 34020
box -48 -56 1008 834
use sg13g2_nor2_1  _0521_
timestamp 1676627187
transform 1 0 19488 0 1 40068
box -48 -56 432 834
use sg13g2_a221oi_1  _0522_
timestamp 1685197497
transform -1 0 19584 0 1 34020
box -48 -56 816 834
use sg13g2_mux2_1  _0523_
timestamp 1677247768
transform 1 0 17856 0 1 34020
box -48 -56 1008 834
use sg13g2_a22oi_1  _0524_
timestamp 1685173987
transform -1 0 20160 0 1 34020
box -48 -56 624 834
use sg13g2_a22oi_1  _0525_
timestamp 1685173987
transform -1 0 19776 0 -1 34020
box -48 -56 624 834
use sg13g2_mux4_1  _0526_
timestamp 1677257233
transform 1 0 14304 0 1 23436
box -48 -56 2064 834
use sg13g2_nand3_1  _0527_
timestamp 1683988354
transform 1 0 18624 0 1 26460
box -48 -56 528 834
use sg13g2_mux2_1  _0528_
timestamp 1677247768
transform 1 0 18048 0 -1 24948
box -48 -56 1008 834
use sg13g2_nor2_1  _0529_
timestamp 1676627187
transform 1 0 19104 0 1 26460
box -48 -56 432 834
use sg13g2_a221oi_1  _0530_
timestamp 1685197497
transform -1 0 19776 0 -1 24948
box -48 -56 816 834
use sg13g2_mux2_1  _0531_
timestamp 1677247768
transform 1 0 18816 0 1 24948
box -48 -56 1008 834
use sg13g2_a22oi_1  _0532_
timestamp 1685173987
transform -1 0 20352 0 1 24948
box -48 -56 624 834
use sg13g2_a22oi_1  _0533_
timestamp 1685173987
transform -1 0 19872 0 -1 26460
box -48 -56 624 834
use sg13g2_mux4_1  _0534_
timestamp 1677257233
transform 1 0 9120 0 1 8316
box -48 -56 2064 834
use sg13g2_nand3_1  _0535_
timestamp 1683988354
transform 1 0 7680 0 -1 26460
box -48 -56 528 834
use sg13g2_mux2_1  _0536_
timestamp 1677247768
transform 1 0 8352 0 -1 24948
box -48 -56 1008 834
use sg13g2_nor2_1  _0537_
timestamp 1676627187
transform 1 0 8448 0 1 23436
box -48 -56 432 834
use sg13g2_a221oi_1  _0538_
timestamp 1685197497
transform -1 0 10080 0 -1 24948
box -48 -56 816 834
use sg13g2_mux2_1  _0539_
timestamp 1677247768
transform 1 0 8160 0 1 24948
box -48 -56 1008 834
use sg13g2_a22oi_1  _0540_
timestamp 1685173987
transform 1 0 9120 0 1 24948
box -48 -56 624 834
use sg13g2_a22oi_1  _0541_
timestamp 1685173987
transform 1 0 8448 0 -1 23436
box -48 -56 624 834
use sg13g2_mux4_1  _0542_
timestamp 1677257233
transform 1 0 7776 0 1 14364
box -48 -56 2064 834
use sg13g2_nand3_1  _0543_
timestamp 1683988354
transform 1 0 2016 0 1 30996
box -48 -56 528 834
use sg13g2_mux2_1  _0544_
timestamp 1677247768
transform 1 0 3168 0 -1 30996
box -48 -56 1008 834
use sg13g2_nor2_1  _0545_
timestamp 1676627187
transform 1 0 2784 0 -1 30996
box -48 -56 432 834
use sg13g2_a221oi_1  _0546_
timestamp 1685197497
transform 1 0 3840 0 -1 32508
box -48 -56 816 834
use sg13g2_mux2_1  _0547_
timestamp 1677247768
transform -1 0 6144 0 -1 29484
box -48 -56 1008 834
use sg13g2_a22oi_1  _0548_
timestamp 1685173987
transform -1 0 4416 0 1 27972
box -48 -56 624 834
use sg13g2_a22oi_1  _0549_
timestamp 1685173987
transform 1 0 1344 0 -1 29484
box -48 -56 624 834
use sg13g2_mux4_1  _0550_
timestamp 1677257233
transform 1 0 11328 0 1 37044
box -48 -56 2064 834
use sg13g2_nand3_1  _0551_
timestamp 1683988354
transform -1 0 16608 0 -1 34020
box -48 -56 528 834
use sg13g2_mux2_1  _0552_
timestamp 1677247768
transform -1 0 15264 0 -1 32508
box -48 -56 1008 834
use sg13g2_nor2_1  _0553_
timestamp 1676627187
transform 1 0 15168 0 1 32508
box -48 -56 432 834
use sg13g2_a221oi_1  _0554_
timestamp 1685197497
transform 1 0 14112 0 -1 34020
box -48 -56 816 834
use sg13g2_mux2_1  _0555_
timestamp 1677247768
transform -1 0 16128 0 -1 34020
box -48 -56 1008 834
use sg13g2_a22oi_1  _0556_
timestamp 1685173987
transform -1 0 15840 0 -1 32508
box -48 -56 624 834
use sg13g2_a22oi_1  _0557_
timestamp 1685173987
transform -1 0 15552 0 -1 30996
box -48 -56 624 834
use sg13g2_mux4_1  _0558_
timestamp 1677257233
transform 1 0 14400 0 -1 23436
box -48 -56 2064 834
use sg13g2_nand3_1  _0559_
timestamp 1683988354
transform 1 0 14496 0 -1 27972
box -48 -56 528 834
use sg13g2_mux2_1  _0560_
timestamp 1677247768
transform 1 0 15360 0 -1 29484
box -48 -56 1008 834
use sg13g2_nor2_1  _0561_
timestamp 1676627187
transform -1 0 16896 0 -1 27972
box -48 -56 432 834
use sg13g2_a221oi_1  _0562_
timestamp 1685197497
transform 1 0 15360 0 1 27972
box -48 -56 816 834
use sg13g2_mux2_1  _0563_
timestamp 1677247768
transform 1 0 14976 0 -1 27972
box -48 -56 1008 834
use sg13g2_a22oi_1  _0564_
timestamp 1685173987
transform 1 0 15936 0 -1 27972
box -48 -56 624 834
use sg13g2_a22oi_1  _0565_
timestamp 1685173987
transform -1 0 16896 0 -1 29484
box -48 -56 624 834
use sg13g2_mux4_1  _0566_
timestamp 1677257233
transform 1 0 9408 0 -1 5292
box -48 -56 2064 834
use sg13g2_nand3_1  _0567_
timestamp 1683988354
transform -1 0 4224 0 -1 23436
box -48 -56 528 834
use sg13g2_mux2_1  _0568_
timestamp 1677247768
transform 1 0 3168 0 -1 20412
box -48 -56 1008 834
use sg13g2_nor2_1  _0569_
timestamp 1676627187
transform 1 0 4128 0 -1 21924
box -48 -56 432 834
use sg13g2_a221oi_1  _0570_
timestamp 1685197497
transform 1 0 3456 0 1 21924
box -48 -56 816 834
use sg13g2_mux2_1  _0571_
timestamp 1677247768
transform 1 0 2784 0 -1 18900
box -48 -56 1008 834
use sg13g2_a22oi_1  _0572_
timestamp 1685173987
transform 1 0 3744 0 1 20412
box -48 -56 624 834
use sg13g2_a22oi_1  _0573_
timestamp 1685173987
transform 1 0 2880 0 1 21924
box -48 -56 624 834
use sg13g2_o21ai_1  _0574_
timestamp 1685175443
transform 1 0 6336 0 1 5292
box -48 -56 538 834
use sg13g2_a21oi_1  _0575_
timestamp 1683973020
transform 1 0 5280 0 -1 9828
box -48 -56 528 834
use sg13g2_nor2b_1  _0576_
timestamp 1685181386
transform 1 0 5856 0 1 5292
box -54 -56 528 834
use sg13g2_a21oi_1  _0577_
timestamp 1683973020
transform 1 0 6336 0 -1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _0578_
timestamp 1685175443
transform -1 0 7296 0 -1 6804
box -48 -56 538 834
use sg13g2_nor2_1  _0579_
timestamp 1676627187
transform -1 0 5280 0 1 8316
box -48 -56 432 834
use sg13g2_mux4_1  _0580_
timestamp 1677257233
transform 1 0 5760 0 -1 9828
box -48 -56 2064 834
use sg13g2_nor2_1  _0581_
timestamp 1676627187
transform -1 0 8160 0 -1 9828
box -48 -56 432 834
use sg13g2_nor2_1  _0582_
timestamp 1676627187
transform 1 0 4896 0 1 6804
box -48 -56 432 834
use sg13g2_o21ai_1  _0583_
timestamp 1685175443
transform -1 0 17952 0 -1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  _0584_
timestamp 1683973020
transform -1 0 17664 0 1 17388
box -48 -56 528 834
use sg13g2_nor2b_1  _0585_
timestamp 1685181386
transform 1 0 16704 0 -1 17388
box -54 -56 528 834
use sg13g2_a21oi_1  _0586_
timestamp 1683973020
transform 1 0 17376 0 1 18900
box -48 -56 528 834
use sg13g2_o21ai_1  _0587_
timestamp 1685175443
transform -1 0 17376 0 1 18900
box -48 -56 538 834
use sg13g2_nor2_1  _0588_
timestamp 1676627187
transform -1 0 17568 0 -1 17388
box -48 -56 432 834
use sg13g2_mux4_1  _0589_
timestamp 1677257233
transform -1 0 17472 0 -1 18900
box -48 -56 2064 834
use sg13g2_nor2_1  _0590_
timestamp 1676627187
transform 1 0 15072 0 -1 18900
box -48 -56 432 834
use sg13g2_nor2_1  _0591_
timestamp 1676627187
transform -1 0 17952 0 -1 17388
box -48 -56 432 834
use sg13g2_o21ai_1  _0592_
timestamp 1685175443
transform 1 0 16800 0 1 8316
box -48 -56 538 834
use sg13g2_a21oi_1  _0593_
timestamp 1683973020
transform 1 0 17376 0 -1 8316
box -48 -56 528 834
use sg13g2_nor2b_1  _0594_
timestamp 1685181386
transform -1 0 17760 0 1 8316
box -54 -56 528 834
use sg13g2_a21oi_1  _0595_
timestamp 1683973020
transform -1 0 17376 0 -1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _0596_
timestamp 1685175443
transform 1 0 16896 0 -1 9828
box -48 -56 538 834
use sg13g2_nor2_1  _0597_
timestamp 1676627187
transform -1 0 18144 0 1 8316
box -48 -56 432 834
use sg13g2_mux4_1  _0598_
timestamp 1677257233
transform 1 0 14880 0 -1 9828
box -48 -56 2064 834
use sg13g2_nor2_1  _0599_
timestamp 1676627187
transform -1 0 17760 0 -1 9828
box -48 -56 432 834
use sg13g2_nor2_1  _0600_
timestamp 1676627187
transform -1 0 16032 0 -1 6804
box -48 -56 432 834
use sg13g2_o21ai_1  _0601_
timestamp 1685175443
transform -1 0 5856 0 1 14364
box -48 -56 538 834
use sg13g2_a21oi_1  _0602_
timestamp 1683973020
transform -1 0 5088 0 -1 14364
box -48 -56 528 834
use sg13g2_nor2b_1  _0603_
timestamp 1685181386
transform -1 0 8064 0 -1 15876
box -54 -56 528 834
use sg13g2_a21oi_1  _0604_
timestamp 1683973020
transform -1 0 5664 0 -1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _0605_
timestamp 1685175443
transform -1 0 5568 0 -1 14364
box -48 -56 538 834
use sg13g2_nor2_1  _0606_
timestamp 1676627187
transform 1 0 4800 0 -1 12852
box -48 -56 432 834
use sg13g2_mux4_1  _0607_
timestamp 1677257233
transform 1 0 5568 0 -1 14364
box -48 -56 2064 834
use sg13g2_nor2_1  _0608_
timestamp 1676627187
transform 1 0 7200 0 1 11340
box -48 -56 432 834
use sg13g2_nor2_1  _0609_
timestamp 1676627187
transform 1 0 6144 0 -1 17388
box -48 -56 432 834
use sg13g2_o21ai_1  _0610_
timestamp 1685175443
transform 1 0 2016 0 -1 14364
box -48 -56 538 834
use sg13g2_a21oi_1  _0611_
timestamp 1683973020
transform 1 0 4704 0 1 11340
box -48 -56 528 834
use sg13g2_nor2b_1  _0612_
timestamp 1685181386
transform 1 0 1248 0 -1 11340
box -54 -56 528 834
use sg13g2_a21oi_1  _0613_
timestamp 1683973020
transform 1 0 1536 0 -1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _0614_
timestamp 1685175443
transform 1 0 2208 0 -1 15876
box -48 -56 538 834
use sg13g2_nor2_1  _0615_
timestamp 1676627187
transform -1 0 4992 0 1 9828
box -48 -56 432 834
use sg13g2_mux4_1  _0616_
timestamp 1677257233
transform -1 0 4800 0 -1 12852
box -48 -56 2064 834
use sg13g2_nor2_1  _0617_
timestamp 1676627187
transform 1 0 1152 0 -1 9828
box -48 -56 432 834
use sg13g2_nor2_1  _0618_
timestamp 1676627187
transform -1 0 3744 0 -1 8316
box -48 -56 432 834
use sg13g2_o21ai_1  _0619_
timestamp 1685175443
transform 1 0 17952 0 1 5292
box -48 -56 538 834
use sg13g2_a21oi_1  _0620_
timestamp 1683973020
transform -1 0 18720 0 -1 6804
box -48 -56 528 834
use sg13g2_nor2b_1  _0621_
timestamp 1685181386
transform 1 0 17088 0 -1 3780
box -54 -56 528 834
use sg13g2_a21oi_1  _0622_
timestamp 1683973020
transform 1 0 17760 0 -1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _0623_
timestamp 1685175443
transform 1 0 19584 0 -1 3780
box -48 -56 538 834
use sg13g2_nor2_1  _0624_
timestamp 1676627187
transform -1 0 20352 0 -1 6804
box -48 -56 432 834
use sg13g2_mux4_1  _0625_
timestamp 1677257233
transform 1 0 16320 0 1 6804
box -48 -56 2064 834
use sg13g2_nor2_1  _0626_
timestamp 1676627187
transform -1 0 19872 0 -1 2268
box -48 -56 432 834
use sg13g2_nor2_1  _0627_
timestamp 1676627187
transform -1 0 15168 0 -1 12852
box -48 -56 432 834
use sg13g2_o21ai_1  _0628_
timestamp 1685175443
transform 1 0 19200 0 -1 20412
box -48 -56 538 834
use sg13g2_a21oi_1  _0629_
timestamp 1683973020
transform -1 0 20256 0 1 18900
box -48 -56 528 834
use sg13g2_nor2b_1  _0630_
timestamp 1685181386
transform 1 0 17856 0 1 17388
box -54 -56 528 834
use sg13g2_a21oi_1  _0631_
timestamp 1683973020
transform -1 0 20160 0 -1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  _0632_
timestamp 1685175443
transform 1 0 19872 0 1 20412
box -48 -56 538 834
use sg13g2_nor2_1  _0633_
timestamp 1676627187
transform 1 0 19968 0 1 17388
box -48 -56 432 834
use sg13g2_mux4_1  _0634_
timestamp 1677257233
transform 1 0 18144 0 -1 18900
box -48 -56 2064 834
use sg13g2_nor2_1  _0635_
timestamp 1676627187
transform 1 0 16608 0 1 21924
box -48 -56 432 834
use sg13g2_nor2_1  _0636_
timestamp 1676627187
transform -1 0 18240 0 1 20412
box -48 -56 432 834
use sg13g2_o21ai_1  _0637_
timestamp 1685175443
transform -1 0 5856 0 -1 2268
box -48 -56 538 834
use sg13g2_a21oi_1  _0638_
timestamp 1683973020
transform 1 0 5376 0 1 5292
box -48 -56 528 834
use sg13g2_nor2b_1  _0639_
timestamp 1685181386
transform 1 0 2784 0 1 5292
box -54 -56 528 834
use sg13g2_a21oi_1  _0640_
timestamp 1683973020
transform 1 0 6240 0 -1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  _0641_
timestamp 1685175443
transform -1 0 3744 0 1 5292
box -48 -56 538 834
use sg13g2_nor2_1  _0642_
timestamp 1676627187
transform -1 0 3360 0 1 2268
box -48 -56 432 834
use sg13g2_mux4_1  _0643_
timestamp 1677257233
transform -1 0 6336 0 -1 6804
box -48 -56 2064 834
use sg13g2_nor2_1  _0644_
timestamp 1676627187
transform -1 0 2688 0 -1 6804
box -48 -56 432 834
use sg13g2_nor2_1  _0645_
timestamp 1676627187
transform 1 0 1920 0 -1 6804
box -48 -56 432 834
use sg13g2_nor3_1  _0646_
timestamp 1676639442
transform 1 0 9312 0 1 2268
box -48 -56 528 834
use sg13g2_nand2b_1  _0647_
timestamp 1676567195
transform 1 0 3936 0 -1 2268
box -48 -56 528 834
use sg13g2_a221oi_1  _0648_
timestamp 1685197497
transform 1 0 10944 0 -1 3780
box -48 -56 816 834
use sg13g2_mux4_1  _0649_
timestamp 1677257233
transform 1 0 6624 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _0650_
timestamp 1677257233
transform 1 0 6720 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux2_1  _0651_
timestamp 1677247768
transform 1 0 8448 0 1 5292
box -48 -56 1008 834
use sg13g2_nand2b_1  _0652_
timestamp 1676567195
transform 1 0 19104 0 1 15876
box -48 -56 528 834
use sg13g2_nand2_1  _0653_
timestamp 1676557249
transform -1 0 20352 0 -1 14364
box -48 -56 432 834
use sg13g2_a21oi_1  _0654_
timestamp 1683973020
transform 1 0 19872 0 -1 15876
box -48 -56 528 834
use sg13g2_nor3_1  _0655_
timestamp 1676639442
transform 1 0 12768 0 -1 29484
box -48 -56 528 834
use sg13g2_nand2b_1  _0656_
timestamp 1676567195
transform 1 0 13440 0 -1 27972
box -48 -56 528 834
use sg13g2_a221oi_1  _0657_
timestamp 1685197497
transform 1 0 12960 0 1 27972
box -48 -56 816 834
use sg13g2_inv_1  _0658_
timestamp 1676382929
transform 1 0 20064 0 -1 27972
box -48 -56 336 834
use sg13g2_o21ai_1  _0659_
timestamp 1685175443
transform -1 0 19680 0 1 14364
box -48 -56 538 834
use sg13g2_a21o_1  _0660_
timestamp 1677175127
transform 1 0 18240 0 -1 15876
box -48 -56 720 834
use sg13g2_nor2b_1  _0661_
timestamp 1685181386
transform 1 0 17760 0 -1 15876
box -54 -56 528 834
use sg13g2_a21oi_1  _0662_
timestamp 1683973020
transform 1 0 19680 0 1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _0663_
timestamp 1685175443
transform 1 0 18144 0 1 14364
box -48 -56 538 834
use sg13g2_mux2_1  _0664_
timestamp 1677247768
transform 1 0 18912 0 -1 15876
box -48 -56 1008 834
use sg13g2_a21oi_1  _0665_
timestamp 1683973020
transform 1 0 19584 0 1 15876
box -48 -56 528 834
use sg13g2_a22oi_1  _0666_
timestamp 1685173987
transform 1 0 18624 0 1 14364
box -48 -56 624 834
use sg13g2_mux2_1  _0667_
timestamp 1677247768
transform -1 0 19104 0 1 8316
box -48 -56 1008 834
use sg13g2_nand2b_1  _0668_
timestamp 1676567195
transform 1 0 15840 0 1 3780
box -48 -56 528 834
use sg13g2_nand2b_1  _0669_
timestamp 1676567195
transform 1 0 14976 0 -1 40068
box -48 -56 528 834
use sg13g2_nor3_1  _0670_
timestamp 1676639442
transform 1 0 14496 0 -1 40068
box -48 -56 528 834
use sg13g2_a221oi_1  _0671_
timestamp 1685197497
transform -1 0 14400 0 1 40068
box -48 -56 816 834
use sg13g2_mux2_1  _0672_
timestamp 1677247768
transform -1 0 19488 0 1 6804
box -48 -56 1008 834
use sg13g2_a21oi_1  _0673_
timestamp 1683973020
transform -1 0 14688 0 1 6804
box -48 -56 528 834
use sg13g2_a21oi_1  _0674_
timestamp 1683973020
transform 1 0 16032 0 -1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _0675_
timestamp 1685175443
transform -1 0 20352 0 1 2268
box -48 -56 538 834
use sg13g2_mux2_1  _0676_
timestamp 1677247768
transform 1 0 19008 0 -1 6804
box -48 -56 1008 834
use sg13g2_a21oi_1  _0677_
timestamp 1683973020
transform -1 0 20352 0 -1 2268
box -48 -56 528 834
use sg13g2_a22oi_1  _0678_
timestamp 1685173987
transform -1 0 20064 0 1 6804
box -48 -56 624 834
use sg13g2_mux2_1  _0679_
timestamp 1677247768
transform 1 0 11904 0 1 9828
box -48 -56 1008 834
use sg13g2_nand2b_1  _0680_
timestamp 1676567195
transform -1 0 12960 0 -1 8316
box -48 -56 528 834
use sg13g2_nand2b_1  _0681_
timestamp 1676567195
transform 1 0 9504 0 1 32508
box -48 -56 528 834
use sg13g2_nor3_1  _0682_
timestamp 1676639442
transform 1 0 8256 0 -1 32508
box -48 -56 528 834
use sg13g2_a221oi_1  _0683_
timestamp 1685197497
transform 1 0 9504 0 -1 30996
box -48 -56 816 834
use sg13g2_mux2_1  _0684_
timestamp 1677247768
transform 1 0 9408 0 1 11340
box -48 -56 1008 834
use sg13g2_a21oi_1  _0685_
timestamp 1683973020
transform -1 0 11712 0 1 8316
box -48 -56 528 834
use sg13g2_a21oi_1  _0686_
timestamp 1683973020
transform 1 0 12864 0 1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _0687_
timestamp 1685175443
transform 1 0 8640 0 1 8316
box -48 -56 538 834
use sg13g2_mux2_1  _0688_
timestamp 1677247768
transform 1 0 11712 0 1 8316
box -48 -56 1008 834
use sg13g2_a21oi_1  _0689_
timestamp 1683973020
transform -1 0 13152 0 1 8316
box -48 -56 528 834
use sg13g2_a22oi_1  _0690_
timestamp 1685173987
transform 1 0 10848 0 -1 9828
box -48 -56 624 834
use sg13g2_mux2_1  _0691_
timestamp 1677247768
transform 1 0 8928 0 -1 11340
box -48 -56 1008 834
use sg13g2_mux2_1  _0692_
timestamp 1677247768
transform -1 0 9120 0 -1 9828
box -48 -56 1008 834
use sg13g2_nand2b_1  _0693_
timestamp 1676567195
transform 1 0 7584 0 1 9828
box -48 -56 528 834
use sg13g2_a21oi_1  _0694_
timestamp 1683973020
transform 1 0 10368 0 -1 12852
box -48 -56 528 834
use sg13g2_a21oi_1  _0695_
timestamp 1683973020
transform -1 0 7488 0 -1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _0696_
timestamp 1685175443
transform 1 0 7104 0 1 9828
box -48 -56 538 834
use sg13g2_mux2_1  _0697_
timestamp 1677247768
transform -1 0 10368 0 -1 12852
box -48 -56 1008 834
use sg13g2_a21oi_1  _0698_
timestamp 1683973020
transform 1 0 7488 0 1 12852
box -48 -56 528 834
use sg13g2_a22oi_1  _0699_
timestamp 1685173987
transform 1 0 9696 0 1 9828
box -48 -56 624 834
use sg13g2_mux2_1  _0700_
timestamp 1677247768
transform -1 0 19968 0 1 9828
box -48 -56 1008 834
use sg13g2_mux2_1  _0701_
timestamp 1677247768
transform 1 0 18528 0 -1 11340
box -48 -56 1008 834
use sg13g2_nand2b_1  _0702_
timestamp 1676567195
transform 1 0 19776 0 -1 8316
box -48 -56 528 834
use sg13g2_a21oi_1  _0703_
timestamp 1683973020
transform -1 0 18432 0 1 3780
box -48 -56 528 834
use sg13g2_a21oi_1  _0704_
timestamp 1683973020
transform -1 0 17376 0 1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _0705_
timestamp 1685175443
transform 1 0 19584 0 1 8316
box -48 -56 538 834
use sg13g2_mux2_1  _0706_
timestamp 1677247768
transform -1 0 19968 0 1 11340
box -48 -56 1008 834
use sg13g2_a21oi_1  _0707_
timestamp 1683973020
transform -1 0 18432 0 -1 5292
box -48 -56 528 834
use sg13g2_a22oi_1  _0708_
timestamp 1685173987
transform -1 0 20064 0 -1 11340
box -48 -56 624 834
use sg13g2_o21ai_1  _0709_
timestamp 1685175443
transform 1 0 17664 0 1 14364
box -48 -56 538 834
use sg13g2_a21o_1  _0710_
timestamp 1677175127
transform -1 0 19488 0 -1 12852
box -48 -56 720 834
use sg13g2_nand2b_1  _0711_
timestamp 1676567195
transform -1 0 19968 0 -1 12852
box -48 -56 528 834
use sg13g2_nand2_1  _0712_
timestamp 1676557249
transform -1 0 20352 0 1 12852
box -48 -56 432 834
use sg13g2_a21oi_1  _0713_
timestamp 1683973020
transform 1 0 19104 0 1 8316
box -48 -56 528 834
use sg13g2_nor2b_1  _0714_
timestamp 1685181386
transform -1 0 20160 0 -1 17388
box -54 -56 528 834
use sg13g2_a21oi_1  _0715_
timestamp 1683973020
transform 1 0 17760 0 -1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _0716_
timestamp 1685175443
transform 1 0 17280 0 -1 15876
box -48 -56 538 834
use sg13g2_mux2_1  _0717_
timestamp 1677247768
transform 1 0 19008 0 1 12852
box -48 -56 1008 834
use sg13g2_a21oi_1  _0718_
timestamp 1683973020
transform -1 0 20352 0 -1 9828
box -48 -56 528 834
use sg13g2_a22oi_1  _0719_
timestamp 1685173987
transform 1 0 19392 0 -1 14364
box -48 -56 624 834
use sg13g2_nor2_1  _0720_
timestamp 1676627187
transform 1 0 10848 0 1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _0721_
timestamp 1676627187
transform -1 0 10368 0 -1 6804
box -48 -56 432 834
use sg13g2_nor3_1  _0722_
timestamp 1676639442
transform 1 0 9408 0 1 5292
box -48 -56 528 834
use sg13g2_o21ai_1  _0723_
timestamp 1685175443
transform 1 0 6144 0 1 3780
box -48 -56 538 834
use sg13g2_a21o_1  _0724_
timestamp 1677175127
transform 1 0 7872 0 -1 6804
box -48 -56 720 834
use sg13g2_nor2b_1  _0725_
timestamp 1685181386
transform -1 0 9984 0 -1 6804
box -54 -56 528 834
use sg13g2_a21oi_1  _0726_
timestamp 1683973020
transform -1 0 9408 0 1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _0727_
timestamp 1685175443
transform -1 0 10848 0 1 3780
box -48 -56 538 834
use sg13g2_mux2_1  _0728_
timestamp 1677247768
transform 1 0 8544 0 -1 6804
box -48 -56 1008 834
use sg13g2_a21oi_1  _0729_
timestamp 1683973020
transform -1 0 9888 0 1 6804
box -48 -56 528 834
use sg13g2_a22oi_1  _0730_
timestamp 1685173987
transform 1 0 7296 0 -1 6804
box -48 -56 624 834
use sg13g2_mux4_1  _0731_
timestamp 1677257233
transform 1 0 11712 0 -1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _0732_
timestamp 1677257233
transform 1 0 11232 0 1 3780
box -48 -56 2064 834
use sg13g2_mux2_1  _0733_
timestamp 1677247768
transform 1 0 13344 0 -1 3780
box -48 -56 1008 834
use sg13g2_mux4_1  _0734_
timestamp 1677257233
transform 1 0 13728 0 -1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _0735_
timestamp 1677257233
transform 1 0 13344 0 1 5292
box -48 -56 2064 834
use sg13g2_mux2_1  _0736_
timestamp 1677247768
transform -1 0 16320 0 1 5292
box -48 -56 1008 834
use sg13g2_mux4_1  _0737_
timestamp 1677257233
transform 1 0 17856 0 1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _0738_
timestamp 1677257233
transform 1 0 17568 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux2_1  _0739_
timestamp 1677247768
transform 1 0 19200 0 1 756
box -48 -56 1008 834
use sg13g2_mux4_1  _0740_
timestamp 1677257233
transform 1 0 15072 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _0741_
timestamp 1677257233
transform 1 0 14784 0 1 2268
box -48 -56 2064 834
use sg13g2_mux2_1  _0742_
timestamp 1677247768
transform 1 0 16800 0 -1 6804
box -48 -56 1008 834
use sg13g2_o21ai_1  _0743_
timestamp 1685175443
transform 1 0 10272 0 1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  _0744_
timestamp 1683973020
transform -1 0 9024 0 -1 29484
box -48 -56 528 834
use sg13g2_or2_1  _0745_
timestamp 1684236171
transform 1 0 6432 0 -1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  _0746_
timestamp 1685175443
transform -1 0 8928 0 1 27972
box -48 -56 538 834
use sg13g2_o21ai_1  _0747_
timestamp 1685175443
transform 1 0 9888 0 1 27972
box -48 -56 538 834
use sg13g2_nor2_1  _0748_
timestamp 1676627187
transform -1 0 14976 0 -1 30996
box -48 -56 432 834
use sg13g2_a21oi_1  _0749_
timestamp 1683973020
transform -1 0 10848 0 1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  _0750_
timestamp 1685175443
transform 1 0 9312 0 1 29484
box -48 -56 538 834
use sg13g2_mux2_1  _0751_
timestamp 1677247768
transform 1 0 8928 0 1 27972
box -48 -56 1008 834
use sg13g2_a21oi_1  _0752_
timestamp 1683973020
transform -1 0 9504 0 -1 29484
box -48 -56 528 834
use sg13g2_a21oi_1  _0753_
timestamp 1683973020
transform -1 0 10272 0 1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  _0754_
timestamp 1685175443
transform 1 0 17280 0 -1 37044
box -48 -56 538 834
use sg13g2_a21oi_1  _0755_
timestamp 1683973020
transform 1 0 19392 0 1 37044
box -48 -56 528 834
use sg13g2_or2_1  _0756_
timestamp 1684236171
transform -1 0 20352 0 1 35532
box -48 -56 528 834
use sg13g2_o21ai_1  _0757_
timestamp 1685175443
transform 1 0 19200 0 -1 37044
box -48 -56 538 834
use sg13g2_o21ai_1  _0758_
timestamp 1685175443
transform 1 0 19872 0 -1 38556
box -48 -56 538 834
use sg13g2_nor2_1  _0759_
timestamp 1676627187
transform 1 0 18720 0 1 38556
box -48 -56 432 834
use sg13g2_a21oi_1  _0760_
timestamp 1683973020
transform -1 0 19872 0 -1 38556
box -48 -56 528 834
use sg13g2_o21ai_1  _0761_
timestamp 1685175443
transform 1 0 18912 0 1 37044
box -48 -56 538 834
use sg13g2_mux2_1  _0762_
timestamp 1677247768
transform 1 0 17760 0 -1 37044
box -48 -56 1008 834
use sg13g2_a21oi_1  _0763_
timestamp 1683973020
transform -1 0 20352 0 -1 37044
box -48 -56 528 834
use sg13g2_a21oi_1  _0764_
timestamp 1683973020
transform 1 0 19872 0 1 37044
box -48 -56 528 834
use sg13g2_mux4_1  _0765_
timestamp 1677257233
transform 1 0 17760 0 1 27972
box -48 -56 2064 834
use sg13g2_mux4_1  _0766_
timestamp 1677257233
transform 1 0 17664 0 -1 27972
box -48 -56 2064 834
use sg13g2_mux2_1  _0767_
timestamp 1677247768
transform 1 0 19392 0 1 29484
box -48 -56 1008 834
use sg13g2_mux4_1  _0768_
timestamp 1677257233
transform 1 0 10176 0 -1 24948
box -48 -56 2064 834
use sg13g2_mux4_1  _0769_
timestamp 1677257233
transform 1 0 10272 0 1 23436
box -48 -56 2064 834
use sg13g2_mux2_1  _0770_
timestamp 1677247768
transform 1 0 11808 0 -1 23436
box -48 -56 1008 834
use sg13g2_mux2_1  _0771_
timestamp 1677247768
transform 1 0 6528 0 1 29484
box -48 -56 1008 834
use sg13g2_or2_1  _0772_
timestamp 1684236171
transform -1 0 11232 0 1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  _0773_
timestamp 1685175443
transform 1 0 8064 0 1 34020
box -48 -56 538 834
use sg13g2_o21ai_1  _0774_
timestamp 1685175443
transform -1 0 7872 0 -1 30996
box -48 -56 538 834
use sg13g2_a21oi_1  _0775_
timestamp 1683973020
transform 1 0 7680 0 -1 27972
box -48 -56 528 834
use sg13g2_mux4_1  _0776_
timestamp 1677257233
transform -1 0 6528 0 1 29484
box -48 -56 2064 834
use sg13g2_nor2_1  _0777_
timestamp 1676627187
transform 1 0 3168 0 1 32508
box -48 -56 432 834
use sg13g2_nor2_1  _0778_
timestamp 1676627187
transform -1 0 4320 0 -1 35532
box -48 -56 432 834
use sg13g2_mux2_1  _0779_
timestamp 1677247768
transform 1 0 15936 0 1 37044
box -48 -56 1008 834
use sg13g2_or2_1  _0780_
timestamp 1684236171
transform 1 0 15360 0 -1 38556
box -48 -56 528 834
use sg13g2_o21ai_1  _0781_
timestamp 1685175443
transform -1 0 16704 0 -1 37044
box -48 -56 538 834
use sg13g2_o21ai_1  _0782_
timestamp 1685175443
transform 1 0 15840 0 -1 38556
box -48 -56 538 834
use sg13g2_a21oi_1  _0783_
timestamp 1683973020
transform 1 0 16320 0 -1 38556
box -48 -56 528 834
use sg13g2_a21oi_1  _0784_
timestamp 1683973020
transform 1 0 16992 0 -1 38556
box -48 -56 528 834
use sg13g2_o21ai_1  _0785_
timestamp 1685175443
transform 1 0 18720 0 -1 37044
box -48 -56 538 834
use sg13g2_mux2_1  _0786_
timestamp 1677247768
transform 1 0 14976 0 1 37044
box -48 -56 1008 834
use sg13g2_a21oi_1  _0787_
timestamp 1683973020
transform -1 0 17184 0 -1 37044
box -48 -56 528 834
use sg13g2_a21oi_1  _0788_
timestamp 1683973020
transform -1 0 18336 0 1 38556
box -48 -56 528 834
use sg13g2_mux2_1  _0789_
timestamp 1677247768
transform -1 0 17568 0 1 30996
box -48 -56 1008 834
use sg13g2_or2_1  _0790_
timestamp 1684236171
transform -1 0 18048 0 -1 30996
box -48 -56 528 834
use sg13g2_o21ai_1  _0791_
timestamp 1685175443
transform -1 0 13824 0 1 30996
box -48 -56 538 834
use sg13g2_o21ai_1  _0792_
timestamp 1685175443
transform -1 0 14112 0 1 29484
box -48 -56 538 834
use sg13g2_a21oi_1  _0793_
timestamp 1683973020
transform 1 0 13824 0 1 30996
box -48 -56 528 834
use sg13g2_mux4_1  _0794_
timestamp 1677257233
transform 1 0 15552 0 -1 30996
box -48 -56 2064 834
use sg13g2_nor2_1  _0795_
timestamp 1676627187
transform 1 0 17376 0 1 29484
box -48 -56 432 834
use sg13g2_nor2_1  _0796_
timestamp 1676627187
transform -1 0 18144 0 -1 32508
box -48 -56 432 834
use sg13g2_mux2_1  _0797_
timestamp 1677247768
transform 1 0 4224 0 -1 24948
box -48 -56 1008 834
use sg13g2_or2_1  _0798_
timestamp 1684236171
transform 1 0 3264 0 -1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  _0799_
timestamp 1685175443
transform -1 0 4704 0 -1 23436
box -48 -56 538 834
use sg13g2_o21ai_1  _0800_
timestamp 1685175443
transform 1 0 3744 0 -1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  _0801_
timestamp 1683973020
transform -1 0 5664 0 -1 24948
box -48 -56 528 834
use sg13g2_mux4_1  _0802_
timestamp 1677257233
transform 1 0 2304 0 1 23436
box -48 -56 2064 834
use sg13g2_nor2_1  _0803_
timestamp 1676627187
transform 1 0 5184 0 1 24948
box -48 -56 432 834
use sg13g2_nor2_1  _0804_
timestamp 1676627187
transform -1 0 6048 0 -1 24948
box -48 -56 432 834
use sg13g2_o21ai_1  _0805_
timestamp 1685175443
transform -1 0 17856 0 1 20412
box -48 -56 538 834
use sg13g2_nand2b_1  _0806_
timestamp 1676567195
transform 1 0 16992 0 1 21924
box -48 -56 528 834
use sg13g2_o21ai_1  _0807_
timestamp 1685175443
transform 1 0 18144 0 -1 21924
box -48 -56 538 834
use sg13g2_mux4_1  _0808_
timestamp 1677257233
transform -1 0 4512 0 1 15876
box -48 -56 2064 834
use sg13g2_mux4_1  _0809_
timestamp 1677257233
transform -1 0 17472 0 1 15876
box -48 -56 2064 834
use sg13g2_mux4_1  _0810_
timestamp 1677257233
transform 1 0 12864 0 1 17388
box -48 -56 2064 834
use sg13g2_mux4_1  _0811_
timestamp 1677257233
transform -1 0 5376 0 -1 17388
box -48 -56 2064 834
use sg13g2_mux4_1  _0812_
timestamp 1677257233
transform -1 0 4512 0 -1 14364
box -48 -56 2064 834
use sg13g2_mux4_1  _0813_
timestamp 1677257233
transform -1 0 17376 0 1 14364
box -48 -56 2064 834
use sg13g2_mux4_1  _0814_
timestamp 1677257233
transform 1 0 11904 0 1 14364
box -48 -56 2064 834
use sg13g2_mux4_1  _0815_
timestamp 1677257233
transform 1 0 3264 0 1 14364
box -48 -56 2064 834
use sg13g2_mux4_1  _0816_
timestamp 1677257233
transform 1 0 9312 0 -1 14364
box -48 -56 2064 834
use sg13g2_mux4_1  _0817_
timestamp 1677257233
transform 1 0 12000 0 -1 30996
box -48 -56 2064 834
use sg13g2_mux4_1  _0818_
timestamp 1677257233
transform 1 0 12096 0 -1 21924
box -48 -56 2064 834
use sg13g2_mux4_1  _0819_
timestamp 1677257233
transform 1 0 9984 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _0820_
timestamp 1677257233
transform -1 0 3936 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _0821_
timestamp 1677257233
transform -1 0 17184 0 -1 12852
box -48 -56 2064 834
use sg13g2_mux4_1  _0822_
timestamp 1677257233
transform 1 0 12000 0 1 11340
box -48 -56 2064 834
use sg13g2_mux4_1  _0823_
timestamp 1677257233
transform 1 0 5184 0 1 11340
box -48 -56 2064 834
use sg13g2_mux4_1  _0824_
timestamp 1677257233
transform 1 0 2304 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _0825_
timestamp 1677257233
transform 1 0 14880 0 1 11340
box -48 -56 2064 834
use sg13g2_mux4_1  _0826_
timestamp 1677257233
transform 1 0 12480 0 -1 14364
box -48 -56 2064 834
use sg13g2_mux4_1  _0827_
timestamp 1677257233
transform -1 0 5184 0 -1 9828
box -48 -56 2064 834
use sg13g2_mux4_1  _0828_
timestamp 1677257233
transform 1 0 2400 0 -1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _0829_
timestamp 1677257233
transform -1 0 15264 0 -1 11340
box -48 -56 2064 834
use sg13g2_mux4_1  _0830_
timestamp 1677257233
transform 1 0 12096 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _0831_
timestamp 1677257233
transform 1 0 2880 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _0832_
timestamp 1677257233
transform 1 0 4896 0 1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _0833_
timestamp 1677257233
transform -1 0 16896 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _0834_
timestamp 1677257233
transform 1 0 13344 0 1 15876
box -48 -56 2064 834
use sg13g2_mux4_1  _0835_
timestamp 1677257233
transform 1 0 5280 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _0836_
timestamp 1677257233
transform 1 0 5664 0 1 17388
box -48 -56 2064 834
use sg13g2_mux4_1  _0837_
timestamp 1677257233
transform 1 0 10656 0 1 17388
box -48 -56 2064 834
use sg13g2_mux4_1  _0838_
timestamp 1677257233
transform 1 0 9792 0 1 15876
box -48 -56 2064 834
use sg13g2_mux4_1  _0839_
timestamp 1677257233
transform -1 0 8832 0 1 15876
box -48 -56 2064 834
use sg13g2_mux4_1  _0840_
timestamp 1677257233
transform 1 0 6336 0 1 21924
box -48 -56 2064 834
use sg13g2_mux4_1  _0841_
timestamp 1677257233
transform 1 0 12096 0 -1 20412
box -48 -56 2064 834
use sg13g2_mux4_1  _0842_
timestamp 1677257233
transform 1 0 10368 0 -1 32508
box -48 -56 2064 834
use sg13g2_mux4_1  _0843_
timestamp 1677257233
transform 1 0 6144 0 -1 20412
box -48 -56 2064 834
use sg13g2_mux4_1  _0844_
timestamp 1677257233
transform 1 0 6144 0 -1 21924
box -48 -56 2064 834
use sg13g2_mux4_1  _0845_
timestamp 1677257233
transform 1 0 13152 0 1 18900
box -48 -56 2064 834
use sg13g2_mux4_1  _0846_
timestamp 1677257233
transform 1 0 11520 0 1 26460
box -48 -56 2064 834
use sg13g2_mux4_1  _0847_
timestamp 1677257233
transform 1 0 5376 0 1 18900
box -48 -56 2064 834
use sg13g2_mux4_1  _0848_
timestamp 1677257233
transform -1 0 3840 0 1 37044
box -48 -56 2064 834
use sg13g2_mux4_1  _0849_
timestamp 1677257233
transform 1 0 10464 0 -1 34020
box -48 -56 2064 834
use sg13g2_mux4_1  _0850_
timestamp 1677257233
transform -1 0 3360 0 -1 40068
box -48 -56 2064 834
use sg13g2_mux4_1  _0851_
timestamp 1677257233
transform -1 0 4128 0 1 34020
box -48 -56 2064 834
use sg13g2_mux4_1  _0852_
timestamp 1677257233
transform 1 0 1152 0 -1 35532
box -48 -56 2064 834
use sg13g2_mux4_1  _0853_
timestamp 1677257233
transform 1 0 1824 0 -1 32508
box -48 -56 2064 834
use sg13g2_mux4_1  _0854_
timestamp 1677257233
transform -1 0 6048 0 -1 34020
box -48 -56 2064 834
use sg13g2_mux4_1  _0855_
timestamp 1677257233
transform 1 0 1824 0 1 27972
box -48 -56 2064 834
use sg13g2_mux4_1  _0856_
timestamp 1677257233
transform 1 0 5952 0 1 30996
box -48 -56 2064 834
use sg13g2_mux4_1  _0857_
timestamp 1677257233
transform 1 0 15936 0 -1 40068
box -48 -56 2064 834
use sg13g2_mux4_1  _0858_
timestamp 1677257233
transform 1 0 11424 0 1 29484
box -48 -56 2064 834
use sg13g2_mux4_1  _0859_
timestamp 1677257233
transform 1 0 4320 0 1 23436
box -48 -56 2064 834
use sg13g2_dlhq_1  _0860_
timestamp 1678805552
transform 1 0 1824 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _0861_
timestamp 1678805552
transform 1 0 4800 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _0862_
timestamp 1678805552
transform 1 0 9984 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _0863_
timestamp 1678805552
transform 1 0 11616 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _0864_
timestamp 1678805552
transform 1 0 14688 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _0865_
timestamp 1678805552
transform 1 0 16224 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _0866_
timestamp 1678805552
transform 1 0 4128 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _0867_
timestamp 1678805552
transform 1 0 6336 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _0868_
timestamp 1678805552
transform 1 0 1152 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _0869_
timestamp 1678805552
transform 1 0 1920 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _0870_
timestamp 1678805552
transform -1 0 7680 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _0871_
timestamp 1678805552
transform 1 0 4416 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _0872_
timestamp 1678805552
transform -1 0 4416 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _0873_
timestamp 1678805552
transform -1 0 3744 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _0874_
timestamp 1678805552
transform -1 0 9984 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _0875_
timestamp 1678805552
transform -1 0 7392 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _0876_
timestamp 1678805552
transform 1 0 1632 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _0877_
timestamp 1678805552
transform 1 0 2112 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _0878_
timestamp 1678805552
transform -1 0 11328 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _0879_
timestamp 1678805552
transform -1 0 13824 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _0880_
timestamp 1678805552
transform 1 0 10752 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _0881_
timestamp 1678805552
transform 1 0 9120 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _0882_
timestamp 1678805552
transform -1 0 5184 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _0883_
timestamp 1678805552
transform -1 0 17088 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _0884_
timestamp 1678805552
transform 1 0 1152 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _0885_
timestamp 1678805552
transform 1 0 3552 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _0886_
timestamp 1678805552
transform 1 0 1344 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _0887_
timestamp 1678805552
transform -1 0 16512 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _0888_
timestamp 1678805552
transform -1 0 17184 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _0889_
timestamp 1678805552
transform 1 0 15744 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _0890_
timestamp 1678805552
transform 1 0 14304 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _0891_
timestamp 1678805552
transform 1 0 13728 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _0892_
timestamp 1678805552
transform 1 0 13344 0 1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _0893_
timestamp 1678805552
transform 1 0 2496 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _0894_
timestamp 1678805552
transform 1 0 4704 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _0895_
timestamp 1678805552
transform 1 0 4128 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _0896_
timestamp 1678805552
transform 1 0 4128 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _0897_
timestamp 1678805552
transform 1 0 4512 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _0898_
timestamp 1678805552
transform 1 0 10080 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _0899_
timestamp 1678805552
transform 1 0 11808 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _0900_
timestamp 1678805552
transform 1 0 11520 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _0901_
timestamp 1678805552
transform -1 0 15744 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _0902_
timestamp 1678805552
transform 1 0 4608 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _0903_
timestamp 1678805552
transform 1 0 6240 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _0904_
timestamp 1678805552
transform 1 0 3744 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _0905_
timestamp 1678805552
transform 1 0 6048 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _0906_
timestamp 1678805552
transform 1 0 8736 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _0907_
timestamp 1678805552
transform 1 0 10560 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _0908_
timestamp 1678805552
transform 1 0 12576 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _0909_
timestamp 1678805552
transform 1 0 10944 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _0910_
timestamp 1678805552
transform 1 0 6624 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _0911_
timestamp 1678805552
transform 1 0 4512 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _0912_
timestamp 1678805552
transform 1 0 5184 0 1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _0913_
timestamp 1678805552
transform 1 0 4320 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _0914_
timestamp 1678805552
transform 1 0 6144 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _0915_
timestamp 1678805552
transform 1 0 10176 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _0916_
timestamp 1678805552
transform 1 0 8160 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _0917_
timestamp 1678805552
transform 1 0 10944 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _0918_
timestamp 1678805552
transform 1 0 5856 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _0919_
timestamp 1678805552
transform 1 0 4032 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _0920_
timestamp 1678805552
transform 1 0 9792 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _0921_
timestamp 1678805552
transform -1 0 13920 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _0922_
timestamp 1678805552
transform 1 0 9792 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _0923_
timestamp 1678805552
transform 1 0 16992 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _0924_
timestamp 1678805552
transform 1 0 17760 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _0925_
timestamp 1678805552
transform 1 0 16128 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _0926_
timestamp 1678805552
transform 1 0 17280 0 1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _0927_
timestamp 1678805552
transform 1 0 17568 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _0928_
timestamp 1678805552
transform 1 0 16512 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _0929_
timestamp 1678805552
transform 1 0 7488 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _0930_
timestamp 1678805552
transform -1 0 11136 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _0931_
timestamp 1678805552
transform 1 0 6912 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _0932_
timestamp 1678805552
transform 1 0 13728 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _0933_
timestamp 1678805552
transform 1 0 15648 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _0934_
timestamp 1678805552
transform 1 0 15168 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _0935_
timestamp 1678805552
transform -1 0 19200 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _0936_
timestamp 1678805552
transform 1 0 18432 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _0937_
timestamp 1678805552
transform 1 0 17856 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _0938_
timestamp 1678805552
transform 1 0 11712 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _0939_
timestamp 1678805552
transform 1 0 14016 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _0940_
timestamp 1678805552
transform 1 0 14016 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _0941_
timestamp 1678805552
transform 1 0 10080 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _0942_
timestamp 1678805552
transform 1 0 11712 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _0943_
timestamp 1678805552
transform 1 0 12672 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _0944_
timestamp 1678805552
transform 1 0 6816 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _0945_
timestamp 1678805552
transform -1 0 8928 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _0946_
timestamp 1678805552
transform 1 0 7488 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _0947_
timestamp 1678805552
transform 1 0 17088 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _0948_
timestamp 1678805552
transform 1 0 17760 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _0949_
timestamp 1678805552
transform 1 0 17280 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _0950_
timestamp 1678805552
transform 1 0 16896 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _0951_
timestamp 1678805552
transform 1 0 17376 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _0952_
timestamp 1678805552
transform 1 0 18240 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _0953_
timestamp 1678805552
transform 1 0 7296 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _0954_
timestamp 1678805552
transform -1 0 9216 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _0955_
timestamp 1678805552
transform -1 0 9408 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _0956_
timestamp 1678805552
transform -1 0 11616 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _0957_
timestamp 1678805552
transform 1 0 10272 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _0958_
timestamp 1678805552
transform 1 0 11424 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _0959_
timestamp 1678805552
transform 1 0 18432 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _0960_
timestamp 1678805552
transform 1 0 18144 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _0961_
timestamp 1678805552
transform 1 0 18432 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _0962_
timestamp 1678805552
transform 1 0 18336 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _0963_
timestamp 1678805552
transform 1 0 18048 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _0964_
timestamp 1678805552
transform 1 0 17472 0 1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _0965_
timestamp 1678805552
transform 1 0 5856 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _0966_
timestamp 1678805552
transform 1 0 6048 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _0967_
timestamp 1678805552
transform 1 0 2976 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _0968_
timestamp 1678805552
transform 1 0 2880 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _0969_
timestamp 1678805552
transform 1 0 4512 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _0970_
timestamp 1678805552
transform -1 0 6048 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _0971_
timestamp 1678805552
transform 1 0 17568 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _0972_
timestamp 1678805552
transform 1 0 18240 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _0973_
timestamp 1678805552
transform 1 0 18144 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _0974_
timestamp 1678805552
transform 1 0 16032 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _0975_
timestamp 1678805552
transform 1 0 16320 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _0976_
timestamp 1678805552
transform 1 0 16320 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _0977_
timestamp 1678805552
transform 1 0 1536 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _0978_
timestamp 1678805552
transform -1 0 4608 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _0979_
timestamp 1678805552
transform 1 0 1536 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _0980_
timestamp 1678805552
transform -1 0 7296 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _0981_
timestamp 1678805552
transform 1 0 4224 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _0982_
timestamp 1678805552
transform 1 0 3072 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _0983_
timestamp 1678805552
transform 1 0 15168 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _0984_
timestamp 1678805552
transform 1 0 13536 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _0985_
timestamp 1678805552
transform 1 0 15264 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _0986_
timestamp 1678805552
transform 1 0 15168 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _0987_
timestamp 1678805552
transform 1 0 15744 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _0988_
timestamp 1678805552
transform -1 0 17184 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _0989_
timestamp 1678805552
transform 1 0 3744 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _0990_
timestamp 1678805552
transform 1 0 5280 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _0991_
timestamp 1678805552
transform -1 0 8544 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _0992_
timestamp 1678805552
transform 1 0 5376 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _0993_
timestamp 1678805552
transform 1 0 3744 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _0994_
timestamp 1678805552
transform 1 0 13632 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _0995_
timestamp 1678805552
transform 1 0 11904 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _0996_
timestamp 1678805552
transform -1 0 16320 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _0997_
timestamp 1678805552
transform 1 0 13248 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _0998_
timestamp 1678805552
transform -1 0 12576 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _0999_
timestamp 1678805552
transform -1 0 10944 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _1000_
timestamp 1678805552
transform 1 0 2688 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1001_
timestamp 1678805552
transform 1 0 1344 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1002_
timestamp 1678805552
transform 1 0 12384 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1003_
timestamp 1678805552
transform 1 0 10848 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1004_
timestamp 1678805552
transform -1 0 14880 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1005_
timestamp 1678805552
transform 1 0 11616 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1006_
timestamp 1678805552
transform -1 0 10368 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _1007_
timestamp 1678805552
transform -1 0 7680 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1008_
timestamp 1678805552
transform 1 0 2112 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1009_
timestamp 1678805552
transform 1 0 1248 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _1010_
timestamp 1678805552
transform -1 0 15168 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1011_
timestamp 1678805552
transform 1 0 11040 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1012_
timestamp 1678805552
transform 1 0 15168 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1013_
timestamp 1678805552
transform 1 0 13344 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1014_
timestamp 1678805552
transform 1 0 1248 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1015_
timestamp 1678805552
transform 1 0 1152 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1016_
timestamp 1678805552
transform 1 0 5376 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1017_
timestamp 1678805552
transform 1 0 3744 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1018_
timestamp 1678805552
transform 1 0 12672 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1019_
timestamp 1678805552
transform 1 0 10368 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1020_
timestamp 1678805552
transform -1 0 18816 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1021_
timestamp 1678805552
transform 1 0 15264 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1022_
timestamp 1678805552
transform -1 0 9312 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1023_
timestamp 1678805552
transform -1 0 6144 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _1024_
timestamp 1678805552
transform 1 0 9120 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1025_
timestamp 1678805552
transform 1 0 10368 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1026_
timestamp 1678805552
transform 1 0 10464 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1027_
timestamp 1678805552
transform 1 0 12192 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1028_
timestamp 1678805552
transform 1 0 10368 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1029_
timestamp 1678805552
transform 1 0 12672 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1030_
timestamp 1678805552
transform 1 0 8064 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1031_
timestamp 1678805552
transform 1 0 9792 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1032_
timestamp 1678805552
transform 1 0 1632 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1033_
timestamp 1678805552
transform 1 0 1344 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1034_
timestamp 1678805552
transform 1 0 11904 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1035_
timestamp 1678805552
transform 1 0 10272 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1036_
timestamp 1678805552
transform -1 0 17760 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1037_
timestamp 1678805552
transform 1 0 14496 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1038_
timestamp 1678805552
transform 1 0 1152 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1039_
timestamp 1678805552
transform 1 0 1152 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1040_
timestamp 1678805552
transform 1 0 2688 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1041_
timestamp 1678805552
transform 1 0 1440 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1042_
timestamp 1678805552
transform 1 0 13248 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1043_
timestamp 1678805552
transform 1 0 11616 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1044_
timestamp 1678805552
transform -1 0 17184 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1045_
timestamp 1678805552
transform 1 0 14880 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1046_
timestamp 1678805552
transform 1 0 1728 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1047_
timestamp 1678805552
transform 1 0 1152 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1048_
timestamp 1678805552
transform 1 0 1536 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1049_
timestamp 1678805552
transform 1 0 1152 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1050_
timestamp 1678805552
transform 1 0 1152 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1051_
timestamp 1678805552
transform 1 0 14112 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1052_
timestamp 1678805552
transform 1 0 13536 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1053_
timestamp 1678805552
transform -1 0 15360 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1054_
timestamp 1678805552
transform -1 0 16032 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1055_
timestamp 1678805552
transform 1 0 12480 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1056_
timestamp 1678805552
transform -1 0 14208 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1057_
timestamp 1678805552
transform 1 0 1536 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1058_
timestamp 1678805552
transform 1 0 1152 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1059_
timestamp 1678805552
transform 1 0 1248 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1060_
timestamp 1678805552
transform 1 0 6816 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1061_
timestamp 1678805552
transform 1 0 6528 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1062_
timestamp 1678805552
transform -1 0 8256 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1063_
timestamp 1678805552
transform 1 0 17664 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1064_
timestamp 1678805552
transform 1 0 16416 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1065_
timestamp 1678805552
transform -1 0 18816 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1066_
timestamp 1678805552
transform 1 0 18432 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1067_
timestamp 1678805552
transform 1 0 16128 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1068_
timestamp 1678805552
transform -1 0 18240 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1069_
timestamp 1678805552
transform 1 0 6048 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1070_
timestamp 1678805552
transform 1 0 6816 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1071_
timestamp 1678805552
transform -1 0 9792 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1072_
timestamp 1678805552
transform 1 0 1632 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1073_
timestamp 1678805552
transform 1 0 1152 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1074_
timestamp 1678805552
transform 1 0 1152 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1075_
timestamp 1678805552
transform 1 0 14496 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1076_
timestamp 1678805552
transform 1 0 13920 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1077_
timestamp 1678805552
transform 1 0 14016 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1078_
timestamp 1678805552
transform 1 0 14880 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1079_
timestamp 1678805552
transform 1 0 13344 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1080_
timestamp 1678805552
transform 1 0 13248 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1081_
timestamp 1678805552
transform 1 0 1440 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1082_
timestamp 1678805552
transform 1 0 1152 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1083_
timestamp 1678805552
transform 1 0 1152 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1084_
timestamp 1678805552
transform 1 0 9216 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1085_
timestamp 1678805552
transform 1 0 8160 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1086_
timestamp 1678805552
transform 1 0 9024 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1087_
timestamp 1678805552
transform 1 0 18336 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1088_
timestamp 1678805552
transform 1 0 16512 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1089_
timestamp 1678805552
transform 1 0 18432 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1090_
timestamp 1678805552
transform 1 0 18144 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1091_
timestamp 1678805552
transform 1 0 16128 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1092_
timestamp 1678805552
transform 1 0 18048 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1093_
timestamp 1678805552
transform 1 0 4416 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1094_
timestamp 1678805552
transform 1 0 4224 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1095_
timestamp 1678805552
transform 1 0 4320 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1096_
timestamp 1678805552
transform 1 0 15744 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1097_
timestamp 1678805552
transform 1 0 16512 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1098_
timestamp 1678805552
transform 1 0 4992 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1099_
timestamp 1678805552
transform 1 0 4800 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1100_
timestamp 1678805552
transform 1 0 6432 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1101_
timestamp 1678805552
transform -1 0 9696 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1102_
timestamp 1678805552
transform 1 0 7680 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1103_
timestamp 1678805552
transform 1 0 8736 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _1104_
timestamp 1678805552
transform 1 0 12768 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1105_
timestamp 1678805552
transform -1 0 17952 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1106_
timestamp 1678805552
transform 1 0 9696 0 1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1107_
timestamp 1678805552
transform 1 0 11712 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1108_
timestamp 1678805552
transform 1 0 6144 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1109_
timestamp 1678805552
transform 1 0 7680 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1110_
timestamp 1678805552
transform 1 0 8064 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1111_
timestamp 1678805552
transform 1 0 9120 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1112_
timestamp 1678805552
transform 1 0 12960 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1113_
timestamp 1678805552
transform 1 0 14784 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1114_
timestamp 1678805552
transform 1 0 7968 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1115_
timestamp 1678805552
transform 1 0 10560 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1116_
timestamp 1678805552
transform 1 0 5952 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1117_
timestamp 1678805552
transform 1 0 8160 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1118_
timestamp 1678805552
transform 1 0 7488 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1119_
timestamp 1678805552
transform -1 0 13536 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1120_
timestamp 1678805552
transform 1 0 13344 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1121_
timestamp 1678805552
transform 1 0 14784 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1122_
timestamp 1678805552
transform 1 0 8160 0 -1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1123_
timestamp 1678805552
transform 1 0 11232 0 -1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1124_
timestamp 1678805552
transform 1 0 6528 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1125_
timestamp 1678805552
transform 1 0 9312 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1126_
timestamp 1678805552
transform 1 0 7680 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _1127_
timestamp 1678805552
transform -1 0 14400 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _1128_
timestamp 1678805552
transform 1 0 9888 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1129_
timestamp 1678805552
transform 1 0 12288 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1130_
timestamp 1678805552
transform 1 0 9888 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1131_
timestamp 1678805552
transform 1 0 11520 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1132_
timestamp 1678805552
transform 1 0 7680 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1133_
timestamp 1678805552
transform 1 0 9312 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1134_
timestamp 1678805552
transform -1 0 14304 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1135_
timestamp 1678805552
transform -1 0 15456 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1136_
timestamp 1678805552
transform 1 0 2208 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1137_
timestamp 1678805552
transform 1 0 3072 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1138_
timestamp 1678805552
transform 1 0 8256 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1139_
timestamp 1678805552
transform 1 0 7104 0 1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1140_
timestamp 1678805552
transform 1 0 6432 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1141_
timestamp 1678805552
transform 1 0 5856 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1142_
timestamp 1678805552
transform -1 0 9312 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1143_
timestamp 1678805552
transform 1 0 3264 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1144_
timestamp 1678805552
transform 1 0 5952 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1145_
timestamp 1678805552
transform 1 0 6528 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1146_
timestamp 1678805552
transform 1 0 4896 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1147_
timestamp 1678805552
transform 1 0 8160 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1148_
timestamp 1678805552
transform 1 0 4128 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1149_
timestamp 1678805552
transform 1 0 3840 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1150_
timestamp 1678805552
transform 1 0 1344 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _1151_
timestamp 1678805552
transform 1 0 2304 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1152_
timestamp 1678805552
transform 1 0 11136 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1153_
timestamp 1678805552
transform 1 0 11328 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1154_
timestamp 1678805552
transform 1 0 12000 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1155_
timestamp 1678805552
transform 1 0 12864 0 -1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1156_
timestamp 1678805552
transform 1 0 7872 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1157_
timestamp 1678805552
transform 1 0 8352 0 1 30996
box -50 -56 1692 834
use sg13g2_buf_1  _1158_
timestamp 1676381911
transform 1 0 19680 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  _1159_
timestamp 1676381911
transform 1 0 19776 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  _1160_
timestamp 1676381911
transform 1 0 19872 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  _1161_
timestamp 1676381911
transform 1 0 19488 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  _1162_
timestamp 1676381911
transform 1 0 19872 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  _1163_
timestamp 1676381911
transform 1 0 18240 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  _1164_
timestamp 1676381911
transform 1 0 19680 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_1  _1165_
timestamp 1676381911
transform 1 0 19776 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  _1166_
timestamp 1676381911
transform 1 0 18624 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_1  _1167_
timestamp 1676381911
transform 1 0 19968 0 1 30996
box -48 -56 432 834
use sg13g2_buf_1  _1168_
timestamp 1676381911
transform 1 0 19776 0 -1 32508
box -48 -56 432 834
use sg13g2_buf_1  _1169_
timestamp 1676381911
transform 1 0 19776 0 -1 34020
box -48 -56 432 834
use sg13g2_buf_1  _1170_
timestamp 1676381911
transform 1 0 17280 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_1  _1171_
timestamp 1676381911
transform 1 0 19776 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1172_
timestamp 1676381911
transform 1 0 19296 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1173_
timestamp 1676381911
transform 1 0 19488 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1174_
timestamp 1676381911
transform 1 0 18336 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1175_
timestamp 1676381911
transform 1 0 19104 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1176_
timestamp 1676381911
transform 1 0 3072 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1177_
timestamp 1676381911
transform 1 0 2304 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1178_
timestamp 1676381911
transform 1 0 3456 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1179_
timestamp 1676381911
transform 1 0 4992 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1180_
timestamp 1676381911
transform 1 0 13344 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  _1181_
timestamp 1676381911
transform 1 0 10080 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1182_
timestamp 1676381911
transform 1 0 11328 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1183_
timestamp 1676381911
transform 1 0 19104 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1184_
timestamp 1676381911
transform 1 0 4032 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1185_
timestamp 1676381911
transform 1 0 10560 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1186_
timestamp 1676381911
transform 1 0 18720 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1187_
timestamp 1676381911
transform 1 0 12768 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  _1188_
timestamp 1676381911
transform 1 0 17856 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  _1189_
timestamp 1676381911
transform 1 0 16896 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_1  _1190_
timestamp 1676381911
transform 1 0 16896 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1191_
timestamp 1676381911
transform -1 0 19104 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1192_
timestamp 1676381911
transform -1 0 19872 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1193_
timestamp 1676381911
transform -1 0 18336 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1194_
timestamp 1676381911
transform 1 0 14400 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  _1195_
timestamp 1676381911
transform -1 0 20256 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1196_
timestamp 1676381911
transform 1 0 15360 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  _1197_
timestamp 1676381911
transform 1 0 14688 0 -1 18900
box -48 -56 432 834
use sg13g2_buf_1  _1198_
timestamp 1676381911
transform 1 0 10560 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1199_
timestamp 1676381911
transform 1 0 10944 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1200_
timestamp 1676381911
transform 1 0 13344 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  _1201_
timestamp 1676381911
transform -1 0 18720 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1202_
timestamp 1676381911
transform 1 0 12384 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  _1203_
timestamp 1676381911
transform 1 0 9312 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1204_
timestamp 1676381911
transform 1 0 3648 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1205_
timestamp 1676381911
transform 1 0 17472 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  _1206_
timestamp 1676381911
transform 1 0 12960 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1207_
timestamp 1676381911
transform 1 0 14496 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  _1208_
timestamp 1676381911
transform 1 0 13344 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1209_
timestamp 1676381911
transform 1 0 14112 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  _1210_
timestamp 1676381911
transform 1 0 13728 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  _1211_
timestamp 1676381911
transform -1 0 3936 0 -1 34020
box -48 -56 432 834
use sg13g2_buf_1  _1212_
timestamp 1676381911
transform 1 0 1152 0 -1 34020
box -48 -56 432 834
use sg13g2_buf_1  _1213_
timestamp 1676381911
transform -1 0 19488 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1214_
timestamp 1676381911
transform 1 0 1440 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1215_
timestamp 1676381911
transform 1 0 1344 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  _1216_
timestamp 1676381911
transform 1 0 1728 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  _1217_
timestamp 1676381911
transform -1 0 4896 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1218_
timestamp 1676381911
transform -1 0 3840 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  _1219_
timestamp 1676381911
transform 1 0 1440 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  _1220_
timestamp 1676381911
transform 1 0 1440 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1221_
timestamp 1676381911
transform -1 0 10656 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1222_
timestamp 1676381911
transform 1 0 1152 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1223_
timestamp 1676381911
transform 1 0 1152 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1224_
timestamp 1676381911
transform 1 0 4128 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1225_
timestamp 1676381911
transform 1 0 1248 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1226_
timestamp 1676381911
transform 1 0 3744 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  _1227_
timestamp 1676381911
transform 1 0 3744 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1228_
timestamp 1676381911
transform 1 0 1344 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1229_
timestamp 1676381911
transform 1 0 1536 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1230_
timestamp 1676381911
transform 1 0 1440 0 -1 32508
box -48 -56 432 834
use sg13g2_buf_1  _1231_
timestamp 1676381911
transform 1 0 4032 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1232_
timestamp 1676381911
transform 1 0 2304 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1233_
timestamp 1676381911
transform 1 0 2688 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1234_
timestamp 1676381911
transform -1 0 6432 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1235_
timestamp 1676381911
transform 1 0 5376 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1236_
timestamp 1676381911
transform -1 0 7968 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1237_
timestamp 1676381911
transform 1 0 4800 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1238_
timestamp 1676381911
transform -1 0 7872 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1239_
timestamp 1676381911
transform 1 0 6816 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1240_
timestamp 1676381911
transform 1 0 4416 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1241_
timestamp 1676381911
transform 1 0 1824 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1242_
timestamp 1676381911
transform 1 0 1920 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1243_
timestamp 1676381911
transform 1 0 3168 0 -1 34020
box -48 -56 432 834
use sg13g2_buf_1  _1244_
timestamp 1676381911
transform 1 0 5568 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1245_
timestamp 1676381911
transform -1 0 20256 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1246_
timestamp 1676381911
transform 1 0 2688 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1247_
timestamp 1676381911
transform -1 0 10272 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1248_
timestamp 1676381911
transform -1 0 17184 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1249_
timestamp 1676381911
transform -1 0 17568 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1250_
timestamp 1676381911
transform -1 0 15072 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1251_
timestamp 1676381911
transform 1 0 4992 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1252_
timestamp 1676381911
transform -1 0 14688 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1253_
timestamp 1676381911
transform -1 0 14784 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  _1254_
timestamp 1676381911
transform -1 0 10656 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1255_
timestamp 1676381911
transform 1 0 6912 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1256_
timestamp 1676381911
transform 1 0 1920 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1257_
timestamp 1676381911
transform -1 0 14880 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  _1258_
timestamp 1676381911
transform 1 0 2016 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _1259_
timestamp 1676381911
transform 1 0 1536 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1260_
timestamp 1676381911
transform 1 0 7296 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1261_
timestamp 1676381911
transform 1 0 4992 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1262_
timestamp 1676381911
transform -1 0 17184 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1263_
timestamp 1676381911
transform 1 0 9408 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1264_
timestamp 1676381911
transform -1 0 17664 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1265_
timestamp 1676381911
transform 1 0 4608 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1266_
timestamp 1676381911
transform -1 0 15072 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1267_
timestamp 1676381911
transform -1 0 16704 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1268_
timestamp 1676381911
transform -1 0 17472 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1269_
timestamp 1676381911
transform -1 0 17856 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1270_
timestamp 1676381911
transform -1 0 15840 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1271_
timestamp 1676381911
transform -1 0 17472 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1272_
timestamp 1676381911
transform -1 0 18240 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1273_
timestamp 1676381911
transform -1 0 17088 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1274_
timestamp 1676381911
transform -1 0 17856 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1275_
timestamp 1676381911
transform -1 0 18624 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1276_
timestamp 1676381911
transform -1 0 18240 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1277_
timestamp 1676381911
transform -1 0 19008 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1278_
timestamp 1676381911
transform -1 0 18720 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1279_
timestamp 1676381911
transform 1 0 14304 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1280_
timestamp 1676381911
transform -1 0 20352 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  _1281_
timestamp 1676381911
transform 1 0 3552 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1282_
timestamp 1676381911
transform 1 0 1152 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1283_
timestamp 1676381911
transform 1 0 14784 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  _1284_
timestamp 1676381911
transform -1 0 20352 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  _1285_
timestamp 1676381911
transform -1 0 20352 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  _1286_
timestamp 1676381911
transform -1 0 14016 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1287_
timestamp 1676381911
transform -1 0 17280 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  _1288_
timestamp 1676381911
transform -1 0 12480 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  _1289_
timestamp 1676381911
transform -1 0 14400 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  _1290_
timestamp 1676381911
transform -1 0 12096 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  _1291_
timestamp 1676381911
transform -1 0 9600 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  _1292_
timestamp 1676381911
transform -1 0 1728 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  _1293_
timestamp 1676381911
transform -1 0 11712 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  _1294_
timestamp 1676381911
transform -1 0 11808 0 1 12852
box -48 -56 432 834
use sg13g2_buf_1  _1295_
timestamp 1676381911
transform -1 0 9216 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  _1296_
timestamp 1676381911
transform -1 0 4512 0 -1 20412
box -48 -56 432 834
use sg13g2_buf_1  _1297_
timestamp 1676381911
transform -1 0 1632 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  _1298_
timestamp 1676381911
transform -1 0 13632 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1299_
timestamp 1676381911
transform -1 0 10752 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1300_
timestamp 1676381911
transform -1 0 6048 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  _1301_
timestamp 1676381911
transform -1 0 3168 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  _1302_
timestamp 1676381911
transform -1 0 2208 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  _1303_
timestamp 1676381911
transform -1 0 4032 0 1 12852
box -48 -56 432 834
use sg13g2_buf_1  _1304_
timestamp 1676381911
transform -1 0 2304 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _1305_
timestamp 1676381911
transform -1 0 1536 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  _1306_
timestamp 1676381911
transform -1 0 14304 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_1  _1307_
timestamp 1676381911
transform -1 0 1536 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _1308_
timestamp 1676381911
transform -1 0 4896 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  _1309_
timestamp 1676381911
transform -1 0 1536 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _1310_
timestamp 1676381911
transform -1 0 1536 0 1 12852
box -48 -56 432 834
use sg13g2_buf_1  _1311_
timestamp 1676381911
transform -1 0 1536 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  _1312_
timestamp 1676381911
transform -1 0 1536 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  _1313_
timestamp 1676381911
transform -1 0 15264 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  _1314_
timestamp 1676381911
transform -1 0 1824 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  _1315_
timestamp 1676381911
transform -1 0 1728 0 -1 17388
box -48 -56 432 834
use sg13g2_buf_1  _1316_
timestamp 1676381911
transform -1 0 5376 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  _1317_
timestamp 1676381911
transform -1 0 13536 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _1318_
timestamp 1676381911
transform -1 0 3648 0 1 12852
box -48 -56 432 834
use sg13g2_buf_1  _1319_
timestamp 1676381911
transform -1 0 8064 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  _1320_
timestamp 1676381911
transform -1 0 2016 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _1321_
timestamp 1676381911
transform -1 0 1920 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _1322_
timestamp 1676381911
transform -1 0 2112 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  _1323_
timestamp 1676381911
transform -1 0 12384 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _1324_
timestamp 1676381911
transform -1 0 1536 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _1325_
timestamp 1676381911
transform -1 0 1632 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1326_
timestamp 1676381911
transform -1 0 5760 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1327_
timestamp 1676381911
transform -1 0 4704 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _1328_
timestamp 1676381911
transform -1 0 4320 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1329_
timestamp 1676381911
transform -1 0 1536 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _1330_
timestamp 1676381911
transform -1 0 1920 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _1331_
timestamp 1676381911
transform -1 0 1824 0 -1 23436
box -48 -56 432 834
use sg13g2_antennanp  ANTENNA_1
timestamp 1679999689
transform -1 0 11712 0 1 24948
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_2
timestamp 1679999689
transform -1 0 12576 0 1 32508
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_3
timestamp 1679999689
transform -1 0 2304 0 1 23436
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_4
timestamp 1679999689
transform 1 0 15840 0 -1 32508
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_5
timestamp 1679999689
transform 1 0 20064 0 -1 3780
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_6
timestamp 1679999689
transform -1 0 1440 0 1 30996
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_7
timestamp 1679999689
transform 1 0 12384 0 -1 32508
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_8
timestamp 1679999689
transform -1 0 4032 0 -1 21924
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_9
timestamp 1679999689
transform -1 0 3456 0 -1 21924
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_10
timestamp 1679999689
transform -1 0 2016 0 1 23436
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_11
timestamp 1679999689
transform 1 0 10464 0 -1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_12
timestamp 1679999689
transform 1 0 8064 0 -1 34020
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_13
timestamp 1679999689
transform 1 0 1536 0 1 27972
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_14
timestamp 1679999689
transform 1 0 15744 0 -1 5292
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_15
timestamp 1679999689
transform 1 0 3168 0 -1 35532
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_16
timestamp 1679999689
transform 1 0 5376 0 1 21924
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_17
timestamp 1679999689
transform 1 0 17280 0 1 756
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_18
timestamp 1679999689
transform 1 0 7968 0 -1 32508
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_19
timestamp 1679999689
transform 1 0 1248 0 1 27972
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_20
timestamp 1679999689
transform -1 0 1440 0 -1 15876
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_21
timestamp 1679999689
transform 1 0 2784 0 1 20412
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_22
timestamp 1679999689
transform 1 0 15360 0 -1 2268
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_23
timestamp 1679999689
transform -1 0 1728 0 1 30996
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_24
timestamp 1679999689
transform 1 0 4320 0 1 2268
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_25
timestamp 1679999689
transform 1 0 15936 0 1 38556
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_26
timestamp 1679999689
transform 1 0 14304 0 1 30996
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_27
timestamp 1679999689
transform 1 0 9792 0 -1 15876
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_28
timestamp 1679999689
transform 1 0 5664 0 1 21924
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_29
timestamp 1679999689
transform 1 0 20064 0 -1 35532
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_30
timestamp 1679999689
transform 1 0 14880 0 -1 34020
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_31
timestamp 1679999689
transform 1 0 9792 0 -1 17388
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_32
timestamp 1679999689
transform 1 0 1152 0 1 17388
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_33
timestamp 1679999689
transform 1 0 17184 0 1 32508
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_34
timestamp 1679999689
transform 1 0 14304 0 -1 30996
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_35
timestamp 1679999689
transform -1 0 10080 0 1 14364
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_36
timestamp 1679999689
transform 1 0 3072 0 1 20412
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_37
timestamp 1679999689
transform -1 0 4992 0 -1 38556
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_38
timestamp 1679999689
transform 1 0 11424 0 -1 26460
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_39
timestamp 1679999689
transform 1 0 7968 0 -1 38556
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_40
timestamp 1679999689
transform 1 0 5952 0 1 21924
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_41
timestamp 1679999689
transform 1 0 1536 0 -1 37044
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_42
timestamp 1679999689
transform -1 0 1440 0 1 35532
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_43
timestamp 1679999689
transform 1 0 4800 0 1 21924
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_44
timestamp 1679999689
transform -1 0 1440 0 -1 23436
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_45
timestamp 1679999689
transform -1 0 1440 0 1 37044
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_46
timestamp 1679999689
transform 1 0 5088 0 1 21924
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_47
timestamp 1679999689
transform 1 0 3456 0 -1 21924
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_48
timestamp 1679999689
transform -1 0 6048 0 1 756
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_49
timestamp 1679999689
transform 1 0 1824 0 -1 37044
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_50
timestamp 1679999689
transform 1 0 3456 0 -1 23436
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_51
timestamp 1679999689
transform 1 0 16512 0 -1 6804
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_52
timestamp 1679999689
transform -1 0 1440 0 -1 38556
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_53
timestamp 1679999689
transform 1 0 3456 0 1 20412
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_54
timestamp 1679999689
transform 1 0 3936 0 -1 3780
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_55
timestamp 1679999689
transform 1 0 1824 0 1 35532
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_56
timestamp 1679999689
transform 1 0 14112 0 1 34020
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_57
timestamp 1679999689
transform 1 0 13728 0 1 34020
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_58
timestamp 1679999689
transform 1 0 12000 0 -1 26460
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_59
timestamp 1679999689
transform 1 0 9984 0 1 38556
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_60
timestamp 1679999689
transform 1 0 8352 0 1 21924
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_61
timestamp 1679999689
transform -1 0 7680 0 -1 38556
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_62
timestamp 1679999689
transform 1 0 6816 0 1 37044
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_63
timestamp 1679999689
transform -1 0 2304 0 -1 38556
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_64
timestamp 1679999689
transform -1 0 7968 0 -1 38556
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_65
timestamp 1679999689
transform 1 0 17664 0 -1 5292
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_66
timestamp 1679999689
transform 1 0 10752 0 -1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_67
timestamp 1679999689
transform 1 0 17568 0 1 2268
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_68
timestamp 1679999689
transform -1 0 4704 0 1 37044
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_69
timestamp 1679999689
transform 1 0 9120 0 -1 2268
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_70
timestamp 1679999689
transform 1 0 9792 0 -1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_71
timestamp 1679999689
transform -1 0 1920 0 -1 3780
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_72
timestamp 1679999689
transform 1 0 9792 0 -1 41580
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_73
timestamp 1679999689
transform 1 0 4608 0 1 2268
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_74
timestamp 1679999689
transform -1 0 3648 0 -1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_75
timestamp 1679999689
transform -1 0 14688 0 1 756
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_76
timestamp 1679999689
transform 1 0 8064 0 -1 37044
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_77
timestamp 1679999689
transform -1 0 4992 0 1 756
box -48 -56 336 834
use sg13g2_buf_8  clkbuf_0_UserCLK
timestamp 1676451365
transform 1 0 18432 0 1 32508
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_1_0__f_UserCLK
timestamp 1676451365
transform 1 0 19008 0 -1 29484
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_1_1__f_UserCLK
timestamp 1676451365
transform -1 0 19392 0 1 35532
box -48 -56 1296 834
use sg13g2_fill_2  FILLER_0_0
timestamp 1677580104
transform 1 0 1152 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_36
timestamp 1677579658
transform 1 0 4608 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_119
timestamp 1677580104
transform 1 0 12576 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_145
timestamp 1677579658
transform 1 0 15072 0 1 756
box -48 -56 144 834
use sg13g2_fill_1  FILLER_0_167
timestamp 1677579658
transform 1 0 17184 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_198
timestamp 1677580104
transform 1 0 20160 0 1 756
box -48 -56 240 834
use sg13g2_fill_2  FILLER_1_34
timestamp 1677580104
transform 1 0 4416 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_111
timestamp 1677579658
transform 1 0 11808 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_129
timestamp 1677580104
transform 1 0 13536 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_1_172
timestamp 1677580104
transform 1 0 17664 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_0
timestamp 1677580104
transform 1 0 1152 0 1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_23
timestamp 1677580104
transform 1 0 3360 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_90
timestamp 1677579658
transform 1 0 9792 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_141
timestamp 1677579658
transform 1 0 14688 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_0
timestamp 1677579658
transform 1 0 1152 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_52
timestamp 1677579658
transform 1 0 6144 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_100
timestamp 1677580104
transform 1 0 10752 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_0
timestamp 1677579658
transform 1 0 1152 0 1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_78
timestamp 1677579658
transform 1 0 8640 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_151
timestamp 1677580104
transform 1 0 15648 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_197
timestamp 1677580104
transform 1 0 20064 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_199
timestamp 1677579658
transform 1 0 20256 0 1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_4
timestamp 1677579658
transform 1 0 1536 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_85
timestamp 1677579658
transform 1 0 9312 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_197
timestamp 1677580104
transform 1 0 20064 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_199
timestamp 1677579658
transform 1 0 20256 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_91
timestamp 1677580104
transform 1 0 9888 0 1 5292
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_183
timestamp 1677580104
transform 1 0 18720 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_185
timestamp 1677579658
transform 1 0 18912 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_0
timestamp 1677579658
transform 1 0 1152 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_91
timestamp 1677579658
transform 1 0 9888 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_113
timestamp 1677579658
transform 1 0 12000 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_135
timestamp 1677579658
transform 1 0 14112 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_179
timestamp 1677580104
transform 1 0 18336 0 1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_21
timestamp 1677580104
transform 1 0 3168 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_100
timestamp 1677579658
transform 1 0 10752 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_199
timestamp 1677579658
transform 1 0 20256 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_37
timestamp 1677580104
transform 1 0 4704 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_77
timestamp 1677579658
transform 1 0 8544 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_104
timestamp 1677579658
transform 1 0 11136 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_42
timestamp 1677579658
transform 1 0 5184 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_100
timestamp 1677579658
transform 1 0 10752 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_124
timestamp 1677580104
transform 1 0 13056 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_12_0
timestamp 1677580104
transform 1 0 1152 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_61
timestamp 1677579658
transform 1 0 7008 0 1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_13_0
timestamp 1677579658
transform 1 0 1152 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_13_91
timestamp 1677579658
transform 1 0 9888 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_84
timestamp 1677580104
transform 1 0 9216 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_14_138
timestamp 1677579658
transform 1 0 14400 0 1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_185
timestamp 1677579658
transform 1 0 18912 0 1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_15_51
timestamp 1677579658
transform 1 0 6048 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_101
timestamp 1677580104
transform 1 0 10848 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_137
timestamp 1677579658
transform 1 0 14304 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_16_4
timestamp 1677579658
transform 1 0 1536 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_30
timestamp 1677580104
transform 1 0 4032 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_71
timestamp 1677579658
transform 1 0 7968 0 1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_16_89
timestamp 1677579658
transform 1 0 9696 0 1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_16_111
timestamp 1677579658
transform 1 0 11808 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_163
timestamp 1677580104
transform 1 0 16800 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_165
timestamp 1677579658
transform 1 0 16992 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_183
timestamp 1677580104
transform 1 0 18720 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_185
timestamp 1677579658
transform 1 0 18912 0 1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_17_35
timestamp 1677579658
transform 1 0 4512 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_17_67
timestamp 1677579658
transform 1 0 7584 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_21
timestamp 1677579658
transform 1 0 3168 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_43
timestamp 1677579658
transform 1 0 5280 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_93
timestamp 1677580104
transform 1 0 10080 0 1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_133
timestamp 1679581782
transform 1 0 13920 0 1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_18_140
timestamp 1679581782
transform 1 0 14592 0 1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_18_147
timestamp 1677579658
transform 1 0 15264 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_169
timestamp 1677580104
transform 1 0 17376 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_171
timestamp 1677579658
transform 1 0 17568 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_198
timestamp 1677580104
transform 1 0 20160 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_72
timestamp 1677579658
transform 1 0 8064 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_19_93
timestamp 1677579658
transform 1 0 10080 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_19_111
timestamp 1677579658
transform 1 0 11808 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_19_129
timestamp 1677579658
transform 1 0 13536 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_147
timestamp 1677580104
transform 1 0 15264 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_149
timestamp 1677579658
transform 1 0 15456 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_19_167
timestamp 1677579658
transform 1 0 17184 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_88
timestamp 1677580104
transform 1 0 9600 0 1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_20_111
timestamp 1679581782
transform 1 0 11808 0 1 15876
box -48 -56 720 834
use sg13g2_decap_8  FILLER_20_118
timestamp 1679581782
transform 1 0 12480 0 1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_20_125
timestamp 1677580104
transform 1 0 13152 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_148
timestamp 1677579658
transform 1 0 15360 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_197
timestamp 1677580104
transform 1 0 20064 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_199
timestamp 1677579658
transform 1 0 20256 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_0
timestamp 1677580104
transform 1 0 1152 0 -1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_21_93
timestamp 1679581782
transform 1 0 10080 0 -1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_21_100
timestamp 1679581782
transform 1 0 10752 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_21_107
timestamp 1677580104
transform 1 0 11424 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_21_160
timestamp 1677580104
transform 1 0 16512 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_175
timestamp 1677579658
transform 1 0 17952 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_198
timestamp 1677580104
transform 1 0 20160 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_72
timestamp 1677579658
transform 1 0 8064 0 1 17388
box -48 -56 144 834
use sg13g2_decap_4  FILLER_22_94
timestamp 1679577901
transform 1 0 10176 0 1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_22_98
timestamp 1677579658
transform 1 0 10560 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_120
timestamp 1677580104
transform 1 0 12672 0 1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_22_147
timestamp 1677580104
transform 1 0 15264 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_149
timestamp 1677579658
transform 1 0 15456 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_172
timestamp 1677580104
transform 1 0 17664 0 1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_23_48
timestamp 1677580104
transform 1 0 5760 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_50
timestamp 1677579658
transform 1 0 5952 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_4  FILLER_23_136
timestamp 1679577901
transform 1 0 14208 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_23_140
timestamp 1677579658
transform 1 0 14592 0 -1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_175
timestamp 1677580104
transform 1 0 17952 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_23_198
timestamp 1677580104
transform 1 0 20160 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_0
timestamp 1677579658
transform 1 0 1152 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_71
timestamp 1679581782
transform 1 0 7968 0 1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_24_78
timestamp 1677580104
transform 1 0 8640 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_80
timestamp 1677579658
transform 1 0 8832 0 1 18900
box -48 -56 144 834
use sg13g2_decap_4  FILLER_24_102
timestamp 1679577901
transform 1 0 10944 0 1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_24_106
timestamp 1677580104
transform 1 0 11328 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_163
timestamp 1677579658
transform 1 0 16800 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_174
timestamp 1677580104
transform 1 0 17856 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_176
timestamp 1677579658
transform 1 0 18048 0 1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_24_199
timestamp 1677579658
transform 1 0 20256 0 1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_25_20
timestamp 1677579658
transform 1 0 3072 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_73
timestamp 1679581782
transform 1 0 8160 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_80
timestamp 1677580104
transform 1 0 8832 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_82
timestamp 1677579658
transform 1 0 9024 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_104
timestamp 1679581782
transform 1 0 11136 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_111
timestamp 1677580104
transform 1 0 11808 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_113
timestamp 1677579658
transform 1 0 12000 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_25_169
timestamp 1677580104
transform 1 0 17376 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_2  FILLER_25_198
timestamp 1677580104
transform 1 0 20160 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_23
timestamp 1677579658
transform 1 0 3360 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_70
timestamp 1679581782
transform 1 0 7872 0 1 20412
box -48 -56 720 834
use sg13g2_decap_8  FILLER_26_77
timestamp 1679581782
transform 1 0 8544 0 1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_26_84
timestamp 1677579658
transform 1 0 9216 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_119
timestamp 1679581782
transform 1 0 12576 0 1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_26_126
timestamp 1677579658
transform 1 0 13248 0 1 20412
box -48 -56 144 834
use sg13g2_decap_4  FILLER_26_144
timestamp 1679577901
transform 1 0 14976 0 1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_30
timestamp 1677579658
transform 1 0 4032 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_27_90
timestamp 1677579658
transform 1 0 9792 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_4  FILLER_27_135
timestamp 1679577901
transform 1 0 14112 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_199
timestamp 1677579658
transform 1 0 20256 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_28_17
timestamp 1677579658
transform 1 0 2784 0 1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_28_53
timestamp 1677579658
transform 1 0 6240 0 1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_132
timestamp 1679581782
transform 1 0 13824 0 1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_28_139
timestamp 1677580104
transform 1 0 14496 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_141
timestamp 1677579658
transform 1 0 14688 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_159
timestamp 1677580104
transform 1 0 16416 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_37
timestamp 1677579658
transform 1 0 4704 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_55
timestamp 1677580104
transform 1 0 6432 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_29_74
timestamp 1677580104
transform 1 0 8256 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_110
timestamp 1677579658
transform 1 0 11712 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_159
timestamp 1677579658
transform 1 0 16416 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_177
timestamp 1677580104
transform 1 0 18144 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_30_0
timestamp 1677580104
transform 1 0 1152 0 1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_30_57
timestamp 1677580104
transform 1 0 6624 0 1 23436
box -48 -56 240 834
use sg13g2_decap_4  FILLER_30_133
timestamp 1679577901
transform 1 0 13920 0 1 23436
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_0
timestamp 1677580104
transform 1 0 1152 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_51
timestamp 1677580104
transform 1 0 6048 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_74
timestamp 1677579658
transform 1 0 8256 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_31_93
timestamp 1677579658
transform 1 0 10080 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_31_115
timestamp 1679581782
transform 1 0 12192 0 -1 24948
box -48 -56 720 834
use sg13g2_fill_1  FILLER_31_122
timestamp 1677579658
transform 1 0 12864 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_31_140
timestamp 1677580104
transform 1 0 14592 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_198
timestamp 1677580104
transform 1 0 20160 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_32_17
timestamp 1677580104
transform 1 0 2784 0 1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_32_54
timestamp 1677580104
transform 1 0 6336 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_89
timestamp 1677579658
transform 1 0 9696 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_110
timestamp 1677580104
transform 1 0 11712 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_112
timestamp 1677579658
transform 1 0 11904 0 1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_33_20
timestamp 1677579658
transform 1 0 3072 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_33_67
timestamp 1677579658
transform 1 0 7584 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_33_199
timestamp 1677579658
transform 1 0 20256 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_34_17
timestamp 1677580104
transform 1 0 2784 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_50
timestamp 1677579658
transform 1 0 5952 0 1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_34_129
timestamp 1677579658
transform 1 0 13536 0 1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_34_199
timestamp 1677579658
transform 1 0 20256 0 1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_35_49
timestamp 1677580104
transform 1 0 5856 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_110
timestamp 1677579658
transform 1 0 11712 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_35_137
timestamp 1677580104
transform 1 0 14304 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_0
timestamp 1677579658
transform 1 0 1152 0 1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_36_51
timestamp 1677579658
transform 1 0 6048 0 1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_36_58
timestamp 1677579658
transform 1 0 6720 0 1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_36_105
timestamp 1677579658
transform 1 0 11232 0 1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_36_198
timestamp 1677580104
transform 1 0 20160 0 1 27972
box -48 -56 240 834
use sg13g2_fill_2  FILLER_37_0
timestamp 1677580104
transform 1 0 1152 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_37_146
timestamp 1677580104
transform 1 0 15168 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_164
timestamp 1677579658
transform 1 0 16896 0 -1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_37_199
timestamp 1677579658
transform 1 0 20256 0 -1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_38_34
timestamp 1677579658
transform 1 0 4416 0 1 29484
box -48 -56 144 834
use sg13g2_fill_2  FILLER_38_83
timestamp 1677580104
transform 1 0 9120 0 1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_38_105
timestamp 1677580104
transform 1 0 11232 0 1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_38_128
timestamp 1677580104
transform 1 0 13440 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_95
timestamp 1677579658
transform 1 0 10272 0 -1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_39_198
timestamp 1677580104
transform 1 0 20160 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_2  FILLER_40_48
timestamp 1677580104
transform 1 0 5760 0 1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_126
timestamp 1677579658
transform 1 0 13248 0 1 30996
box -48 -56 144 834
use sg13g2_fill_1  FILLER_40_160
timestamp 1677579658
transform 1 0 16512 0 1 30996
box -48 -56 144 834
use sg13g2_fill_1  FILLER_40_181
timestamp 1677579658
transform 1 0 18528 0 1 30996
box -48 -56 144 834
use sg13g2_fill_1  FILLER_41_36
timestamp 1677579658
transform 1 0 4608 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_41_198
timestamp 1677580104
transform 1 0 20160 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_0
timestamp 1677579658
transform 1 0 1152 0 1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_42_85
timestamp 1677580104
transform 1 0 9312 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_97
timestamp 1677579658
transform 1 0 10464 0 1 32508
box -48 -56 144 834
use sg13g2_fill_1  FILLER_42_115
timestamp 1677579658
transform 1 0 12192 0 1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_42_136
timestamp 1677580104
transform 1 0 14208 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_199
timestamp 1677579658
transform 1 0 20256 0 1 32508
box -48 -56 144 834
use sg13g2_fill_1  FILLER_43_29
timestamp 1677579658
transform 1 0 3936 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_43_198
timestamp 1677580104
transform 1 0 20160 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_44_0
timestamp 1677580104
transform 1 0 1152 0 1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_44_48
timestamp 1677580104
transform 1 0 5760 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_71
timestamp 1677579658
transform 1 0 7968 0 1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_44_125
timestamp 1677580104
transform 1 0 13152 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_134
timestamp 1677579658
transform 1 0 14016 0 1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_44_155
timestamp 1677579658
transform 1 0 16032 0 1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_44_173
timestamp 1677579658
transform 1 0 17760 0 1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_44_198
timestamp 1677580104
transform 1 0 20160 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_45_28
timestamp 1677579658
transform 1 0 3840 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_46_89
timestamp 1677580104
transform 1 0 9696 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_125
timestamp 1677579658
transform 1 0 13152 0 1 35532
box -48 -56 144 834
use sg13g2_fill_1  FILLER_47_39
timestamp 1677579658
transform 1 0 4896 0 -1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_47_96
timestamp 1677580104
transform 1 0 10368 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_2  FILLER_47_150
timestamp 1677580104
transform 1 0 15552 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_47_167
timestamp 1677579658
transform 1 0 17184 0 -1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_47_193
timestamp 1677580104
transform 1 0 19680 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_2  FILLER_48_28
timestamp 1677580104
transform 1 0 3840 0 1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_48_58
timestamp 1677579658
transform 1 0 6720 0 1 37044
box -48 -56 144 834
use sg13g2_fill_1  FILLER_48_79
timestamp 1677579658
transform 1 0 8736 0 1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_49_7
timestamp 1677580104
transform 1 0 1824 0 -1 38556
box -48 -56 240 834
use sg13g2_fill_2  FILLER_49_57
timestamp 1677580104
transform 1 0 6624 0 -1 38556
box -48 -56 240 834
use sg13g2_fill_2  FILLER_49_63
timestamp 1677580104
transform 1 0 7200 0 -1 38556
box -48 -56 240 834
use sg13g2_fill_2  FILLER_49_163
timestamp 1677580104
transform 1 0 16800 0 -1 38556
box -48 -56 240 834
use sg13g2_fill_1  FILLER_49_170
timestamp 1677579658
transform 1 0 17472 0 -1 38556
box -48 -56 144 834
use sg13g2_fill_2  FILLER_49_188
timestamp 1677580104
transform 1 0 19200 0 -1 38556
box -48 -56 240 834
use sg13g2_fill_1  FILLER_50_70
timestamp 1677579658
transform 1 0 7872 0 1 38556
box -48 -56 144 834
use sg13g2_fill_2  FILLER_50_187
timestamp 1677580104
transform 1 0 19104 0 1 38556
box -48 -56 240 834
use sg13g2_fill_1  FILLER_50_193
timestamp 1677579658
transform 1 0 19680 0 1 38556
box -48 -56 144 834
use sg13g2_fill_2  FILLER_50_198
timestamp 1677580104
transform 1 0 20160 0 1 38556
box -48 -56 240 834
use sg13g2_fill_2  FILLER_51_0
timestamp 1677580104
transform 1 0 1152 0 -1 40068
box -48 -56 240 834
use sg13g2_fill_2  FILLER_51_71
timestamp 1677580104
transform 1 0 7968 0 -1 40068
box -48 -56 240 834
use sg13g2_fill_2  FILLER_51_103
timestamp 1677580104
transform 1 0 11040 0 -1 40068
box -48 -56 240 834
use sg13g2_fill_1  FILLER_51_153
timestamp 1677579658
transform 1 0 15840 0 -1 40068
box -48 -56 144 834
use sg13g2_fill_1  FILLER_51_199
timestamp 1677579658
transform 1 0 20256 0 -1 40068
box -48 -56 144 834
use sg13g2_fill_2  FILLER_52_0
timestamp 1677580104
transform 1 0 1152 0 1 40068
box -48 -56 240 834
use sg13g2_fill_1  FILLER_52_6
timestamp 1677579658
transform 1 0 1728 0 1 40068
box -48 -56 144 834
use sg13g2_fill_1  FILLER_52_45
timestamp 1677579658
transform 1 0 5472 0 1 40068
box -48 -56 144 834
use sg13g2_fill_2  FILLER_52_88
timestamp 1677580104
transform 1 0 9600 0 1 40068
box -48 -56 240 834
use sg13g2_fill_2  FILLER_52_111
timestamp 1677580104
transform 1 0 11808 0 1 40068
box -48 -56 240 834
use sg13g2_fill_1  FILLER_52_178
timestamp 1677579658
transform 1 0 18240 0 1 40068
box -48 -56 144 834
use sg13g2_fill_1  FILLER_52_199
timestamp 1677579658
transform 1 0 20256 0 1 40068
box -48 -56 144 834
use sg13g2_fill_1  FILLER_53_0
timestamp 1677579658
transform 1 0 1152 0 -1 41580
box -48 -56 144 834
use sg13g2_fill_2  FILLER_53_96
timestamp 1677580104
transform 1 0 10368 0 -1 41580
box -48 -56 240 834
use sg13g2_fill_1  FILLER_53_186
timestamp 1677579658
transform 1 0 19008 0 -1 41580
box -48 -56 144 834
use sg13g2_fill_1  FILLER_53_199
timestamp 1677579658
transform 1 0 20256 0 -1 41580
box -48 -56 144 834
<< labels >>
flabel metal3 s 21424 23396 21504 23476 0 FreeSans 320 0 0 0 CLK_TT_PROJECT
port 0 nsew signal output
flabel metal3 s 0 16172 80 16252 0 FreeSans 320 0 0 0 E1END[0]
port 1 nsew signal input
flabel metal3 s 0 16508 80 16588 0 FreeSans 320 0 0 0 E1END[1]
port 2 nsew signal input
flabel metal3 s 0 16844 80 16924 0 FreeSans 320 0 0 0 E1END[2]
port 3 nsew signal input
flabel metal3 s 0 17180 80 17260 0 FreeSans 320 0 0 0 E1END[3]
port 4 nsew signal input
flabel metal3 s 0 20204 80 20284 0 FreeSans 320 0 0 0 E2END[0]
port 5 nsew signal input
flabel metal3 s 0 20540 80 20620 0 FreeSans 320 0 0 0 E2END[1]
port 6 nsew signal input
flabel metal3 s 0 20876 80 20956 0 FreeSans 320 0 0 0 E2END[2]
port 7 nsew signal input
flabel metal3 s 0 21212 80 21292 0 FreeSans 320 0 0 0 E2END[3]
port 8 nsew signal input
flabel metal3 s 0 21548 80 21628 0 FreeSans 320 0 0 0 E2END[4]
port 9 nsew signal input
flabel metal3 s 0 21884 80 21964 0 FreeSans 320 0 0 0 E2END[5]
port 10 nsew signal input
flabel metal3 s 0 22220 80 22300 0 FreeSans 320 0 0 0 E2END[6]
port 11 nsew signal input
flabel metal3 s 0 22556 80 22636 0 FreeSans 320 0 0 0 E2END[7]
port 12 nsew signal input
flabel metal3 s 0 17516 80 17596 0 FreeSans 320 0 0 0 E2MID[0]
port 13 nsew signal input
flabel metal3 s 0 17852 80 17932 0 FreeSans 320 0 0 0 E2MID[1]
port 14 nsew signal input
flabel metal3 s 0 18188 80 18268 0 FreeSans 320 0 0 0 E2MID[2]
port 15 nsew signal input
flabel metal3 s 0 18524 80 18604 0 FreeSans 320 0 0 0 E2MID[3]
port 16 nsew signal input
flabel metal3 s 0 18860 80 18940 0 FreeSans 320 0 0 0 E2MID[4]
port 17 nsew signal input
flabel metal3 s 0 19196 80 19276 0 FreeSans 320 0 0 0 E2MID[5]
port 18 nsew signal input
flabel metal3 s 0 19532 80 19612 0 FreeSans 320 0 0 0 E2MID[6]
port 19 nsew signal input
flabel metal3 s 0 19868 80 19948 0 FreeSans 320 0 0 0 E2MID[7]
port 20 nsew signal input
flabel metal3 s 0 28268 80 28348 0 FreeSans 320 0 0 0 E6END[0]
port 21 nsew signal input
flabel metal3 s 0 31628 80 31708 0 FreeSans 320 0 0 0 E6END[10]
port 22 nsew signal input
flabel metal3 s 0 31964 80 32044 0 FreeSans 320 0 0 0 E6END[11]
port 23 nsew signal input
flabel metal3 s 0 28604 80 28684 0 FreeSans 320 0 0 0 E6END[1]
port 24 nsew signal input
flabel metal3 s 0 28940 80 29020 0 FreeSans 320 0 0 0 E6END[2]
port 25 nsew signal input
flabel metal3 s 0 29276 80 29356 0 FreeSans 320 0 0 0 E6END[3]
port 26 nsew signal input
flabel metal3 s 0 29612 80 29692 0 FreeSans 320 0 0 0 E6END[4]
port 27 nsew signal input
flabel metal3 s 0 29948 80 30028 0 FreeSans 320 0 0 0 E6END[5]
port 28 nsew signal input
flabel metal3 s 0 30284 80 30364 0 FreeSans 320 0 0 0 E6END[6]
port 29 nsew signal input
flabel metal3 s 0 30620 80 30700 0 FreeSans 320 0 0 0 E6END[7]
port 30 nsew signal input
flabel metal3 s 0 30956 80 31036 0 FreeSans 320 0 0 0 E6END[8]
port 31 nsew signal input
flabel metal3 s 0 31292 80 31372 0 FreeSans 320 0 0 0 E6END[9]
port 32 nsew signal input
flabel metal3 s 0 22892 80 22972 0 FreeSans 320 0 0 0 EE4END[0]
port 33 nsew signal input
flabel metal3 s 0 26252 80 26332 0 FreeSans 320 0 0 0 EE4END[10]
port 34 nsew signal input
flabel metal3 s 0 26588 80 26668 0 FreeSans 320 0 0 0 EE4END[11]
port 35 nsew signal input
flabel metal3 s 0 26924 80 27004 0 FreeSans 320 0 0 0 EE4END[12]
port 36 nsew signal input
flabel metal3 s 0 27260 80 27340 0 FreeSans 320 0 0 0 EE4END[13]
port 37 nsew signal input
flabel metal3 s 0 27596 80 27676 0 FreeSans 320 0 0 0 EE4END[14]
port 38 nsew signal input
flabel metal3 s 0 27932 80 28012 0 FreeSans 320 0 0 0 EE4END[15]
port 39 nsew signal input
flabel metal3 s 0 23228 80 23308 0 FreeSans 320 0 0 0 EE4END[1]
port 40 nsew signal input
flabel metal3 s 0 23564 80 23644 0 FreeSans 320 0 0 0 EE4END[2]
port 41 nsew signal input
flabel metal3 s 0 23900 80 23980 0 FreeSans 320 0 0 0 EE4END[3]
port 42 nsew signal input
flabel metal3 s 0 24236 80 24316 0 FreeSans 320 0 0 0 EE4END[4]
port 43 nsew signal input
flabel metal3 s 0 24572 80 24652 0 FreeSans 320 0 0 0 EE4END[5]
port 44 nsew signal input
flabel metal3 s 0 24908 80 24988 0 FreeSans 320 0 0 0 EE4END[6]
port 45 nsew signal input
flabel metal3 s 0 25244 80 25324 0 FreeSans 320 0 0 0 EE4END[7]
port 46 nsew signal input
flabel metal3 s 0 25580 80 25660 0 FreeSans 320 0 0 0 EE4END[8]
port 47 nsew signal input
flabel metal3 s 0 25916 80 25996 0 FreeSans 320 0 0 0 EE4END[9]
port 48 nsew signal input
flabel metal3 s 21424 22892 21504 22972 0 FreeSans 320 0 0 0 ENA_TT_PROJECT
port 49 nsew signal output
flabel metal3 s 0 32300 80 32380 0 FreeSans 320 0 0 0 FrameData[0]
port 50 nsew signal input
flabel metal3 s 0 35660 80 35740 0 FreeSans 320 0 0 0 FrameData[10]
port 51 nsew signal input
flabel metal3 s 0 35996 80 36076 0 FreeSans 320 0 0 0 FrameData[11]
port 52 nsew signal input
flabel metal3 s 0 36332 80 36412 0 FreeSans 320 0 0 0 FrameData[12]
port 53 nsew signal input
flabel metal3 s 0 36668 80 36748 0 FreeSans 320 0 0 0 FrameData[13]
port 54 nsew signal input
flabel metal3 s 0 37004 80 37084 0 FreeSans 320 0 0 0 FrameData[14]
port 55 nsew signal input
flabel metal3 s 0 37340 80 37420 0 FreeSans 320 0 0 0 FrameData[15]
port 56 nsew signal input
flabel metal3 s 0 37676 80 37756 0 FreeSans 320 0 0 0 FrameData[16]
port 57 nsew signal input
flabel metal3 s 0 38012 80 38092 0 FreeSans 320 0 0 0 FrameData[17]
port 58 nsew signal input
flabel metal3 s 0 38348 80 38428 0 FreeSans 320 0 0 0 FrameData[18]
port 59 nsew signal input
flabel metal3 s 0 38684 80 38764 0 FreeSans 320 0 0 0 FrameData[19]
port 60 nsew signal input
flabel metal3 s 0 32636 80 32716 0 FreeSans 320 0 0 0 FrameData[1]
port 61 nsew signal input
flabel metal3 s 0 39020 80 39100 0 FreeSans 320 0 0 0 FrameData[20]
port 62 nsew signal input
flabel metal3 s 0 39356 80 39436 0 FreeSans 320 0 0 0 FrameData[21]
port 63 nsew signal input
flabel metal3 s 0 39692 80 39772 0 FreeSans 320 0 0 0 FrameData[22]
port 64 nsew signal input
flabel metal3 s 0 40028 80 40108 0 FreeSans 320 0 0 0 FrameData[23]
port 65 nsew signal input
flabel metal3 s 0 40364 80 40444 0 FreeSans 320 0 0 0 FrameData[24]
port 66 nsew signal input
flabel metal3 s 0 40700 80 40780 0 FreeSans 320 0 0 0 FrameData[25]
port 67 nsew signal input
flabel metal3 s 0 41036 80 41116 0 FreeSans 320 0 0 0 FrameData[26]
port 68 nsew signal input
flabel metal3 s 0 41372 80 41452 0 FreeSans 320 0 0 0 FrameData[27]
port 69 nsew signal input
flabel metal3 s 0 41708 80 41788 0 FreeSans 320 0 0 0 FrameData[28]
port 70 nsew signal input
flabel metal3 s 0 42044 80 42124 0 FreeSans 320 0 0 0 FrameData[29]
port 71 nsew signal input
flabel metal3 s 0 32972 80 33052 0 FreeSans 320 0 0 0 FrameData[2]
port 72 nsew signal input
flabel metal3 s 0 42380 80 42460 0 FreeSans 320 0 0 0 FrameData[30]
port 73 nsew signal input
flabel metal3 s 0 42716 80 42796 0 FreeSans 320 0 0 0 FrameData[31]
port 74 nsew signal input
flabel metal3 s 0 33308 80 33388 0 FreeSans 320 0 0 0 FrameData[3]
port 75 nsew signal input
flabel metal3 s 0 33644 80 33724 0 FreeSans 320 0 0 0 FrameData[4]
port 76 nsew signal input
flabel metal3 s 0 33980 80 34060 0 FreeSans 320 0 0 0 FrameData[5]
port 77 nsew signal input
flabel metal3 s 0 34316 80 34396 0 FreeSans 320 0 0 0 FrameData[6]
port 78 nsew signal input
flabel metal3 s 0 34652 80 34732 0 FreeSans 320 0 0 0 FrameData[7]
port 79 nsew signal input
flabel metal3 s 0 34988 80 35068 0 FreeSans 320 0 0 0 FrameData[8]
port 80 nsew signal input
flabel metal3 s 0 35324 80 35404 0 FreeSans 320 0 0 0 FrameData[9]
port 81 nsew signal input
flabel metal3 s 21424 24404 21504 24484 0 FreeSans 320 0 0 0 FrameData_O[0]
port 82 nsew signal output
flabel metal3 s 21424 29444 21504 29524 0 FreeSans 320 0 0 0 FrameData_O[10]
port 83 nsew signal output
flabel metal3 s 21424 29948 21504 30028 0 FreeSans 320 0 0 0 FrameData_O[11]
port 84 nsew signal output
flabel metal3 s 21424 30452 21504 30532 0 FreeSans 320 0 0 0 FrameData_O[12]
port 85 nsew signal output
flabel metal3 s 21424 30956 21504 31036 0 FreeSans 320 0 0 0 FrameData_O[13]
port 86 nsew signal output
flabel metal3 s 21424 31460 21504 31540 0 FreeSans 320 0 0 0 FrameData_O[14]
port 87 nsew signal output
flabel metal3 s 21424 31964 21504 32044 0 FreeSans 320 0 0 0 FrameData_O[15]
port 88 nsew signal output
flabel metal3 s 21424 32468 21504 32548 0 FreeSans 320 0 0 0 FrameData_O[16]
port 89 nsew signal output
flabel metal3 s 21424 32972 21504 33052 0 FreeSans 320 0 0 0 FrameData_O[17]
port 90 nsew signal output
flabel metal3 s 21424 33476 21504 33556 0 FreeSans 320 0 0 0 FrameData_O[18]
port 91 nsew signal output
flabel metal3 s 21424 33980 21504 34060 0 FreeSans 320 0 0 0 FrameData_O[19]
port 92 nsew signal output
flabel metal3 s 21424 24908 21504 24988 0 FreeSans 320 0 0 0 FrameData_O[1]
port 93 nsew signal output
flabel metal3 s 21424 34484 21504 34564 0 FreeSans 320 0 0 0 FrameData_O[20]
port 94 nsew signal output
flabel metal3 s 21424 34988 21504 35068 0 FreeSans 320 0 0 0 FrameData_O[21]
port 95 nsew signal output
flabel metal3 s 21424 35492 21504 35572 0 FreeSans 320 0 0 0 FrameData_O[22]
port 96 nsew signal output
flabel metal3 s 21424 35996 21504 36076 0 FreeSans 320 0 0 0 FrameData_O[23]
port 97 nsew signal output
flabel metal3 s 21424 36500 21504 36580 0 FreeSans 320 0 0 0 FrameData_O[24]
port 98 nsew signal output
flabel metal3 s 21424 37004 21504 37084 0 FreeSans 320 0 0 0 FrameData_O[25]
port 99 nsew signal output
flabel metal3 s 21424 37508 21504 37588 0 FreeSans 320 0 0 0 FrameData_O[26]
port 100 nsew signal output
flabel metal3 s 21424 38012 21504 38092 0 FreeSans 320 0 0 0 FrameData_O[27]
port 101 nsew signal output
flabel metal3 s 21424 38516 21504 38596 0 FreeSans 320 0 0 0 FrameData_O[28]
port 102 nsew signal output
flabel metal3 s 21424 39020 21504 39100 0 FreeSans 320 0 0 0 FrameData_O[29]
port 103 nsew signal output
flabel metal3 s 21424 25412 21504 25492 0 FreeSans 320 0 0 0 FrameData_O[2]
port 104 nsew signal output
flabel metal3 s 21424 39524 21504 39604 0 FreeSans 320 0 0 0 FrameData_O[30]
port 105 nsew signal output
flabel metal3 s 21424 40028 21504 40108 0 FreeSans 320 0 0 0 FrameData_O[31]
port 106 nsew signal output
flabel metal3 s 21424 25916 21504 25996 0 FreeSans 320 0 0 0 FrameData_O[3]
port 107 nsew signal output
flabel metal3 s 21424 26420 21504 26500 0 FreeSans 320 0 0 0 FrameData_O[4]
port 108 nsew signal output
flabel metal3 s 21424 26924 21504 27004 0 FreeSans 320 0 0 0 FrameData_O[5]
port 109 nsew signal output
flabel metal3 s 21424 27428 21504 27508 0 FreeSans 320 0 0 0 FrameData_O[6]
port 110 nsew signal output
flabel metal3 s 21424 27932 21504 28012 0 FreeSans 320 0 0 0 FrameData_O[7]
port 111 nsew signal output
flabel metal3 s 21424 28436 21504 28516 0 FreeSans 320 0 0 0 FrameData_O[8]
port 112 nsew signal output
flabel metal3 s 21424 28940 21504 29020 0 FreeSans 320 0 0 0 FrameData_O[9]
port 113 nsew signal output
flabel metal2 s 15800 0 15880 80 0 FreeSans 320 0 0 0 FrameStrobe[0]
port 114 nsew signal input
flabel metal2 s 17720 0 17800 80 0 FreeSans 320 0 0 0 FrameStrobe[10]
port 115 nsew signal input
flabel metal2 s 17912 0 17992 80 0 FreeSans 320 0 0 0 FrameStrobe[11]
port 116 nsew signal input
flabel metal2 s 18104 0 18184 80 0 FreeSans 320 0 0 0 FrameStrobe[12]
port 117 nsew signal input
flabel metal2 s 18296 0 18376 80 0 FreeSans 320 0 0 0 FrameStrobe[13]
port 118 nsew signal input
flabel metal2 s 18488 0 18568 80 0 FreeSans 320 0 0 0 FrameStrobe[14]
port 119 nsew signal input
flabel metal2 s 18680 0 18760 80 0 FreeSans 320 0 0 0 FrameStrobe[15]
port 120 nsew signal input
flabel metal2 s 18872 0 18952 80 0 FreeSans 320 0 0 0 FrameStrobe[16]
port 121 nsew signal input
flabel metal2 s 19064 0 19144 80 0 FreeSans 320 0 0 0 FrameStrobe[17]
port 122 nsew signal input
flabel metal2 s 19256 0 19336 80 0 FreeSans 320 0 0 0 FrameStrobe[18]
port 123 nsew signal input
flabel metal2 s 19448 0 19528 80 0 FreeSans 320 0 0 0 FrameStrobe[19]
port 124 nsew signal input
flabel metal2 s 15992 0 16072 80 0 FreeSans 320 0 0 0 FrameStrobe[1]
port 125 nsew signal input
flabel metal2 s 16184 0 16264 80 0 FreeSans 320 0 0 0 FrameStrobe[2]
port 126 nsew signal input
flabel metal2 s 16376 0 16456 80 0 FreeSans 320 0 0 0 FrameStrobe[3]
port 127 nsew signal input
flabel metal2 s 16568 0 16648 80 0 FreeSans 320 0 0 0 FrameStrobe[4]
port 128 nsew signal input
flabel metal2 s 16760 0 16840 80 0 FreeSans 320 0 0 0 FrameStrobe[5]
port 129 nsew signal input
flabel metal2 s 16952 0 17032 80 0 FreeSans 320 0 0 0 FrameStrobe[6]
port 130 nsew signal input
flabel metal2 s 17144 0 17224 80 0 FreeSans 320 0 0 0 FrameStrobe[7]
port 131 nsew signal input
flabel metal2 s 17336 0 17416 80 0 FreeSans 320 0 0 0 FrameStrobe[8]
port 132 nsew signal input
flabel metal2 s 17528 0 17608 80 0 FreeSans 320 0 0 0 FrameStrobe[9]
port 133 nsew signal input
flabel metal2 s 15800 42928 15880 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[0]
port 134 nsew signal output
flabel metal2 s 17720 42928 17800 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[10]
port 135 nsew signal output
flabel metal2 s 17912 42928 17992 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[11]
port 136 nsew signal output
flabel metal2 s 18104 42928 18184 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[12]
port 137 nsew signal output
flabel metal2 s 18296 42928 18376 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[13]
port 138 nsew signal output
flabel metal2 s 18488 42928 18568 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[14]
port 139 nsew signal output
flabel metal2 s 18680 42928 18760 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[15]
port 140 nsew signal output
flabel metal2 s 18872 42928 18952 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[16]
port 141 nsew signal output
flabel metal2 s 19064 42928 19144 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[17]
port 142 nsew signal output
flabel metal2 s 19256 42928 19336 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[18]
port 143 nsew signal output
flabel metal2 s 19448 42928 19528 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[19]
port 144 nsew signal output
flabel metal2 s 15992 42928 16072 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[1]
port 145 nsew signal output
flabel metal2 s 16184 42928 16264 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[2]
port 146 nsew signal output
flabel metal2 s 16376 42928 16456 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[3]
port 147 nsew signal output
flabel metal2 s 16568 42928 16648 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[4]
port 148 nsew signal output
flabel metal2 s 16760 42928 16840 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[5]
port 149 nsew signal output
flabel metal2 s 16952 42928 17032 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[6]
port 150 nsew signal output
flabel metal2 s 17144 42928 17224 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[7]
port 151 nsew signal output
flabel metal2 s 17336 42928 17416 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[8]
port 152 nsew signal output
flabel metal2 s 17528 42928 17608 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[9]
port 153 nsew signal output
flabel metal2 s 1784 42928 1864 43008 0 FreeSans 320 0 0 0 N1BEG[0]
port 154 nsew signal output
flabel metal2 s 1976 42928 2056 43008 0 FreeSans 320 0 0 0 N1BEG[1]
port 155 nsew signal output
flabel metal2 s 2168 42928 2248 43008 0 FreeSans 320 0 0 0 N1BEG[2]
port 156 nsew signal output
flabel metal2 s 2360 42928 2440 43008 0 FreeSans 320 0 0 0 N1BEG[3]
port 157 nsew signal output
flabel metal2 s 1784 0 1864 80 0 FreeSans 320 0 0 0 N1END[0]
port 158 nsew signal input
flabel metal2 s 1976 0 2056 80 0 FreeSans 320 0 0 0 N1END[1]
port 159 nsew signal input
flabel metal2 s 2168 0 2248 80 0 FreeSans 320 0 0 0 N1END[2]
port 160 nsew signal input
flabel metal2 s 2360 0 2440 80 0 FreeSans 320 0 0 0 N1END[3]
port 161 nsew signal input
flabel metal2 s 2552 42928 2632 43008 0 FreeSans 320 0 0 0 N2BEG[0]
port 162 nsew signal output
flabel metal2 s 2744 42928 2824 43008 0 FreeSans 320 0 0 0 N2BEG[1]
port 163 nsew signal output
flabel metal2 s 2936 42928 3016 43008 0 FreeSans 320 0 0 0 N2BEG[2]
port 164 nsew signal output
flabel metal2 s 3128 42928 3208 43008 0 FreeSans 320 0 0 0 N2BEG[3]
port 165 nsew signal output
flabel metal2 s 3320 42928 3400 43008 0 FreeSans 320 0 0 0 N2BEG[4]
port 166 nsew signal output
flabel metal2 s 3512 42928 3592 43008 0 FreeSans 320 0 0 0 N2BEG[5]
port 167 nsew signal output
flabel metal2 s 3704 42928 3784 43008 0 FreeSans 320 0 0 0 N2BEG[6]
port 168 nsew signal output
flabel metal2 s 3896 42928 3976 43008 0 FreeSans 320 0 0 0 N2BEG[7]
port 169 nsew signal output
flabel metal2 s 4088 42928 4168 43008 0 FreeSans 320 0 0 0 N2BEGb[0]
port 170 nsew signal output
flabel metal2 s 4280 42928 4360 43008 0 FreeSans 320 0 0 0 N2BEGb[1]
port 171 nsew signal output
flabel metal2 s 4472 42928 4552 43008 0 FreeSans 320 0 0 0 N2BEGb[2]
port 172 nsew signal output
flabel metal2 s 4664 42928 4744 43008 0 FreeSans 320 0 0 0 N2BEGb[3]
port 173 nsew signal output
flabel metal2 s 4856 42928 4936 43008 0 FreeSans 320 0 0 0 N2BEGb[4]
port 174 nsew signal output
flabel metal2 s 5048 42928 5128 43008 0 FreeSans 320 0 0 0 N2BEGb[5]
port 175 nsew signal output
flabel metal2 s 5240 42928 5320 43008 0 FreeSans 320 0 0 0 N2BEGb[6]
port 176 nsew signal output
flabel metal2 s 5432 42928 5512 43008 0 FreeSans 320 0 0 0 N2BEGb[7]
port 177 nsew signal output
flabel metal2 s 4088 0 4168 80 0 FreeSans 320 0 0 0 N2END[0]
port 178 nsew signal input
flabel metal2 s 4280 0 4360 80 0 FreeSans 320 0 0 0 N2END[1]
port 179 nsew signal input
flabel metal2 s 4472 0 4552 80 0 FreeSans 320 0 0 0 N2END[2]
port 180 nsew signal input
flabel metal2 s 4664 0 4744 80 0 FreeSans 320 0 0 0 N2END[3]
port 181 nsew signal input
flabel metal2 s 4856 0 4936 80 0 FreeSans 320 0 0 0 N2END[4]
port 182 nsew signal input
flabel metal2 s 5048 0 5128 80 0 FreeSans 320 0 0 0 N2END[5]
port 183 nsew signal input
flabel metal2 s 5240 0 5320 80 0 FreeSans 320 0 0 0 N2END[6]
port 184 nsew signal input
flabel metal2 s 5432 0 5512 80 0 FreeSans 320 0 0 0 N2END[7]
port 185 nsew signal input
flabel metal2 s 2552 0 2632 80 0 FreeSans 320 0 0 0 N2MID[0]
port 186 nsew signal input
flabel metal2 s 2744 0 2824 80 0 FreeSans 320 0 0 0 N2MID[1]
port 187 nsew signal input
flabel metal2 s 2936 0 3016 80 0 FreeSans 320 0 0 0 N2MID[2]
port 188 nsew signal input
flabel metal2 s 3128 0 3208 80 0 FreeSans 320 0 0 0 N2MID[3]
port 189 nsew signal input
flabel metal2 s 3320 0 3400 80 0 FreeSans 320 0 0 0 N2MID[4]
port 190 nsew signal input
flabel metal2 s 3512 0 3592 80 0 FreeSans 320 0 0 0 N2MID[5]
port 191 nsew signal input
flabel metal2 s 3704 0 3784 80 0 FreeSans 320 0 0 0 N2MID[6]
port 192 nsew signal input
flabel metal2 s 3896 0 3976 80 0 FreeSans 320 0 0 0 N2MID[7]
port 193 nsew signal input
flabel metal2 s 5624 42928 5704 43008 0 FreeSans 320 0 0 0 N4BEG[0]
port 194 nsew signal output
flabel metal2 s 7544 42928 7624 43008 0 FreeSans 320 0 0 0 N4BEG[10]
port 195 nsew signal output
flabel metal2 s 7736 42928 7816 43008 0 FreeSans 320 0 0 0 N4BEG[11]
port 196 nsew signal output
flabel metal2 s 7928 42928 8008 43008 0 FreeSans 320 0 0 0 N4BEG[12]
port 197 nsew signal output
flabel metal2 s 8120 42928 8200 43008 0 FreeSans 320 0 0 0 N4BEG[13]
port 198 nsew signal output
flabel metal2 s 8312 42928 8392 43008 0 FreeSans 320 0 0 0 N4BEG[14]
port 199 nsew signal output
flabel metal2 s 8504 42928 8584 43008 0 FreeSans 320 0 0 0 N4BEG[15]
port 200 nsew signal output
flabel metal2 s 5816 42928 5896 43008 0 FreeSans 320 0 0 0 N4BEG[1]
port 201 nsew signal output
flabel metal2 s 6008 42928 6088 43008 0 FreeSans 320 0 0 0 N4BEG[2]
port 202 nsew signal output
flabel metal2 s 6200 42928 6280 43008 0 FreeSans 320 0 0 0 N4BEG[3]
port 203 nsew signal output
flabel metal2 s 6392 42928 6472 43008 0 FreeSans 320 0 0 0 N4BEG[4]
port 204 nsew signal output
flabel metal2 s 6584 42928 6664 43008 0 FreeSans 320 0 0 0 N4BEG[5]
port 205 nsew signal output
flabel metal2 s 6776 42928 6856 43008 0 FreeSans 320 0 0 0 N4BEG[6]
port 206 nsew signal output
flabel metal2 s 6968 42928 7048 43008 0 FreeSans 320 0 0 0 N4BEG[7]
port 207 nsew signal output
flabel metal2 s 7160 42928 7240 43008 0 FreeSans 320 0 0 0 N4BEG[8]
port 208 nsew signal output
flabel metal2 s 7352 42928 7432 43008 0 FreeSans 320 0 0 0 N4BEG[9]
port 209 nsew signal output
flabel metal2 s 5624 0 5704 80 0 FreeSans 320 0 0 0 N4END[0]
port 210 nsew signal input
flabel metal2 s 7544 0 7624 80 0 FreeSans 320 0 0 0 N4END[10]
port 211 nsew signal input
flabel metal2 s 7736 0 7816 80 0 FreeSans 320 0 0 0 N4END[11]
port 212 nsew signal input
flabel metal2 s 7928 0 8008 80 0 FreeSans 320 0 0 0 N4END[12]
port 213 nsew signal input
flabel metal2 s 8120 0 8200 80 0 FreeSans 320 0 0 0 N4END[13]
port 214 nsew signal input
flabel metal2 s 8312 0 8392 80 0 FreeSans 320 0 0 0 N4END[14]
port 215 nsew signal input
flabel metal2 s 8504 0 8584 80 0 FreeSans 320 0 0 0 N4END[15]
port 216 nsew signal input
flabel metal2 s 5816 0 5896 80 0 FreeSans 320 0 0 0 N4END[1]
port 217 nsew signal input
flabel metal2 s 6008 0 6088 80 0 FreeSans 320 0 0 0 N4END[2]
port 218 nsew signal input
flabel metal2 s 6200 0 6280 80 0 FreeSans 320 0 0 0 N4END[3]
port 219 nsew signal input
flabel metal2 s 6392 0 6472 80 0 FreeSans 320 0 0 0 N4END[4]
port 220 nsew signal input
flabel metal2 s 6584 0 6664 80 0 FreeSans 320 0 0 0 N4END[5]
port 221 nsew signal input
flabel metal2 s 6776 0 6856 80 0 FreeSans 320 0 0 0 N4END[6]
port 222 nsew signal input
flabel metal2 s 6968 0 7048 80 0 FreeSans 320 0 0 0 N4END[7]
port 223 nsew signal input
flabel metal2 s 7160 0 7240 80 0 FreeSans 320 0 0 0 N4END[8]
port 224 nsew signal input
flabel metal2 s 7352 0 7432 80 0 FreeSans 320 0 0 0 N4END[9]
port 225 nsew signal input
flabel metal3 s 21424 23900 21504 23980 0 FreeSans 320 0 0 0 RST_N_TT_PROJECT
port 226 nsew signal output
flabel metal2 s 8696 0 8776 80 0 FreeSans 320 0 0 0 S1BEG[0]
port 227 nsew signal output
flabel metal2 s 8888 0 8968 80 0 FreeSans 320 0 0 0 S1BEG[1]
port 228 nsew signal output
flabel metal2 s 9080 0 9160 80 0 FreeSans 320 0 0 0 S1BEG[2]
port 229 nsew signal output
flabel metal2 s 9272 0 9352 80 0 FreeSans 320 0 0 0 S1BEG[3]
port 230 nsew signal output
flabel metal2 s 8696 42928 8776 43008 0 FreeSans 320 0 0 0 S1END[0]
port 231 nsew signal input
flabel metal2 s 8888 42928 8968 43008 0 FreeSans 320 0 0 0 S1END[1]
port 232 nsew signal input
flabel metal2 s 9080 42928 9160 43008 0 FreeSans 320 0 0 0 S1END[2]
port 233 nsew signal input
flabel metal2 s 9272 42928 9352 43008 0 FreeSans 320 0 0 0 S1END[3]
port 234 nsew signal input
flabel metal2 s 9464 0 9544 80 0 FreeSans 320 0 0 0 S2BEG[0]
port 235 nsew signal output
flabel metal2 s 9656 0 9736 80 0 FreeSans 320 0 0 0 S2BEG[1]
port 236 nsew signal output
flabel metal2 s 9848 0 9928 80 0 FreeSans 320 0 0 0 S2BEG[2]
port 237 nsew signal output
flabel metal2 s 10040 0 10120 80 0 FreeSans 320 0 0 0 S2BEG[3]
port 238 nsew signal output
flabel metal2 s 10232 0 10312 80 0 FreeSans 320 0 0 0 S2BEG[4]
port 239 nsew signal output
flabel metal2 s 10424 0 10504 80 0 FreeSans 320 0 0 0 S2BEG[5]
port 240 nsew signal output
flabel metal2 s 10616 0 10696 80 0 FreeSans 320 0 0 0 S2BEG[6]
port 241 nsew signal output
flabel metal2 s 10808 0 10888 80 0 FreeSans 320 0 0 0 S2BEG[7]
port 242 nsew signal output
flabel metal2 s 11000 0 11080 80 0 FreeSans 320 0 0 0 S2BEGb[0]
port 243 nsew signal output
flabel metal2 s 11192 0 11272 80 0 FreeSans 320 0 0 0 S2BEGb[1]
port 244 nsew signal output
flabel metal2 s 11384 0 11464 80 0 FreeSans 320 0 0 0 S2BEGb[2]
port 245 nsew signal output
flabel metal2 s 11576 0 11656 80 0 FreeSans 320 0 0 0 S2BEGb[3]
port 246 nsew signal output
flabel metal2 s 11768 0 11848 80 0 FreeSans 320 0 0 0 S2BEGb[4]
port 247 nsew signal output
flabel metal2 s 11960 0 12040 80 0 FreeSans 320 0 0 0 S2BEGb[5]
port 248 nsew signal output
flabel metal2 s 12152 0 12232 80 0 FreeSans 320 0 0 0 S2BEGb[6]
port 249 nsew signal output
flabel metal2 s 12344 0 12424 80 0 FreeSans 320 0 0 0 S2BEGb[7]
port 250 nsew signal output
flabel metal2 s 11000 42928 11080 43008 0 FreeSans 320 0 0 0 S2END[0]
port 251 nsew signal input
flabel metal2 s 11192 42928 11272 43008 0 FreeSans 320 0 0 0 S2END[1]
port 252 nsew signal input
flabel metal2 s 11384 42928 11464 43008 0 FreeSans 320 0 0 0 S2END[2]
port 253 nsew signal input
flabel metal2 s 11576 42928 11656 43008 0 FreeSans 320 0 0 0 S2END[3]
port 254 nsew signal input
flabel metal2 s 11768 42928 11848 43008 0 FreeSans 320 0 0 0 S2END[4]
port 255 nsew signal input
flabel metal2 s 11960 42928 12040 43008 0 FreeSans 320 0 0 0 S2END[5]
port 256 nsew signal input
flabel metal2 s 12152 42928 12232 43008 0 FreeSans 320 0 0 0 S2END[6]
port 257 nsew signal input
flabel metal2 s 12344 42928 12424 43008 0 FreeSans 320 0 0 0 S2END[7]
port 258 nsew signal input
flabel metal2 s 9464 42928 9544 43008 0 FreeSans 320 0 0 0 S2MID[0]
port 259 nsew signal input
flabel metal2 s 9656 42928 9736 43008 0 FreeSans 320 0 0 0 S2MID[1]
port 260 nsew signal input
flabel metal2 s 9848 42928 9928 43008 0 FreeSans 320 0 0 0 S2MID[2]
port 261 nsew signal input
flabel metal2 s 10040 42928 10120 43008 0 FreeSans 320 0 0 0 S2MID[3]
port 262 nsew signal input
flabel metal2 s 10232 42928 10312 43008 0 FreeSans 320 0 0 0 S2MID[4]
port 263 nsew signal input
flabel metal2 s 10424 42928 10504 43008 0 FreeSans 320 0 0 0 S2MID[5]
port 264 nsew signal input
flabel metal2 s 10616 42928 10696 43008 0 FreeSans 320 0 0 0 S2MID[6]
port 265 nsew signal input
flabel metal2 s 10808 42928 10888 43008 0 FreeSans 320 0 0 0 S2MID[7]
port 266 nsew signal input
flabel metal2 s 12536 0 12616 80 0 FreeSans 320 0 0 0 S4BEG[0]
port 267 nsew signal output
flabel metal2 s 14456 0 14536 80 0 FreeSans 320 0 0 0 S4BEG[10]
port 268 nsew signal output
flabel metal2 s 14648 0 14728 80 0 FreeSans 320 0 0 0 S4BEG[11]
port 269 nsew signal output
flabel metal2 s 14840 0 14920 80 0 FreeSans 320 0 0 0 S4BEG[12]
port 270 nsew signal output
flabel metal2 s 15032 0 15112 80 0 FreeSans 320 0 0 0 S4BEG[13]
port 271 nsew signal output
flabel metal2 s 15224 0 15304 80 0 FreeSans 320 0 0 0 S4BEG[14]
port 272 nsew signal output
flabel metal2 s 15416 0 15496 80 0 FreeSans 320 0 0 0 S4BEG[15]
port 273 nsew signal output
flabel metal2 s 12728 0 12808 80 0 FreeSans 320 0 0 0 S4BEG[1]
port 274 nsew signal output
flabel metal2 s 12920 0 13000 80 0 FreeSans 320 0 0 0 S4BEG[2]
port 275 nsew signal output
flabel metal2 s 13112 0 13192 80 0 FreeSans 320 0 0 0 S4BEG[3]
port 276 nsew signal output
flabel metal2 s 13304 0 13384 80 0 FreeSans 320 0 0 0 S4BEG[4]
port 277 nsew signal output
flabel metal2 s 13496 0 13576 80 0 FreeSans 320 0 0 0 S4BEG[5]
port 278 nsew signal output
flabel metal2 s 13688 0 13768 80 0 FreeSans 320 0 0 0 S4BEG[6]
port 279 nsew signal output
flabel metal2 s 13880 0 13960 80 0 FreeSans 320 0 0 0 S4BEG[7]
port 280 nsew signal output
flabel metal2 s 14072 0 14152 80 0 FreeSans 320 0 0 0 S4BEG[8]
port 281 nsew signal output
flabel metal2 s 14264 0 14344 80 0 FreeSans 320 0 0 0 S4BEG[9]
port 282 nsew signal output
flabel metal2 s 12536 42928 12616 43008 0 FreeSans 320 0 0 0 S4END[0]
port 283 nsew signal input
flabel metal2 s 14456 42928 14536 43008 0 FreeSans 320 0 0 0 S4END[10]
port 284 nsew signal input
flabel metal2 s 14648 42928 14728 43008 0 FreeSans 320 0 0 0 S4END[11]
port 285 nsew signal input
flabel metal2 s 14840 42928 14920 43008 0 FreeSans 320 0 0 0 S4END[12]
port 286 nsew signal input
flabel metal2 s 15032 42928 15112 43008 0 FreeSans 320 0 0 0 S4END[13]
port 287 nsew signal input
flabel metal2 s 15224 42928 15304 43008 0 FreeSans 320 0 0 0 S4END[14]
port 288 nsew signal input
flabel metal2 s 15416 42928 15496 43008 0 FreeSans 320 0 0 0 S4END[15]
port 289 nsew signal input
flabel metal2 s 12728 42928 12808 43008 0 FreeSans 320 0 0 0 S4END[1]
port 290 nsew signal input
flabel metal2 s 12920 42928 13000 43008 0 FreeSans 320 0 0 0 S4END[2]
port 291 nsew signal input
flabel metal2 s 13112 42928 13192 43008 0 FreeSans 320 0 0 0 S4END[3]
port 292 nsew signal input
flabel metal2 s 13304 42928 13384 43008 0 FreeSans 320 0 0 0 S4END[4]
port 293 nsew signal input
flabel metal2 s 13496 42928 13576 43008 0 FreeSans 320 0 0 0 S4END[5]
port 294 nsew signal input
flabel metal2 s 13688 42928 13768 43008 0 FreeSans 320 0 0 0 S4END[6]
port 295 nsew signal input
flabel metal2 s 13880 42928 13960 43008 0 FreeSans 320 0 0 0 S4END[7]
port 296 nsew signal input
flabel metal2 s 14072 42928 14152 43008 0 FreeSans 320 0 0 0 S4END[8]
port 297 nsew signal input
flabel metal2 s 14264 42928 14344 43008 0 FreeSans 320 0 0 0 S4END[9]
port 298 nsew signal input
flabel metal3 s 21424 18860 21504 18940 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT0
port 299 nsew signal output
flabel metal3 s 21424 19364 21504 19444 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT1
port 300 nsew signal output
flabel metal3 s 21424 19868 21504 19948 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT2
port 301 nsew signal output
flabel metal3 s 21424 20372 21504 20452 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT3
port 302 nsew signal output
flabel metal3 s 21424 20876 21504 20956 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT4
port 303 nsew signal output
flabel metal3 s 21424 21380 21504 21460 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT5
port 304 nsew signal output
flabel metal3 s 21424 21884 21504 21964 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT6
port 305 nsew signal output
flabel metal3 s 21424 22388 21504 22468 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT7
port 306 nsew signal output
flabel metal3 s 21424 10796 21504 10876 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT0
port 307 nsew signal input
flabel metal3 s 21424 11300 21504 11380 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT1
port 308 nsew signal input
flabel metal3 s 21424 11804 21504 11884 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT2
port 309 nsew signal input
flabel metal3 s 21424 12308 21504 12388 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT3
port 310 nsew signal input
flabel metal3 s 21424 12812 21504 12892 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT4
port 311 nsew signal input
flabel metal3 s 21424 13316 21504 13396 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT5
port 312 nsew signal input
flabel metal3 s 21424 13820 21504 13900 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT6
port 313 nsew signal input
flabel metal3 s 21424 14324 21504 14404 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT7
port 314 nsew signal input
flabel metal3 s 21424 6764 21504 6844 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT0
port 315 nsew signal input
flabel metal3 s 21424 7268 21504 7348 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT1
port 316 nsew signal input
flabel metal3 s 21424 7772 21504 7852 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT2
port 317 nsew signal input
flabel metal3 s 21424 8276 21504 8356 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT3
port 318 nsew signal input
flabel metal3 s 21424 8780 21504 8860 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT4
port 319 nsew signal input
flabel metal3 s 21424 9284 21504 9364 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT5
port 320 nsew signal input
flabel metal3 s 21424 9788 21504 9868 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT6
port 321 nsew signal input
flabel metal3 s 21424 10292 21504 10372 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT7
port 322 nsew signal input
flabel metal3 s 21424 14828 21504 14908 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT0
port 323 nsew signal output
flabel metal3 s 21424 15332 21504 15412 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT1
port 324 nsew signal output
flabel metal3 s 21424 15836 21504 15916 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT2
port 325 nsew signal output
flabel metal3 s 21424 16340 21504 16420 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT3
port 326 nsew signal output
flabel metal3 s 21424 16844 21504 16924 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT4
port 327 nsew signal output
flabel metal3 s 21424 17348 21504 17428 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT5
port 328 nsew signal output
flabel metal3 s 21424 17852 21504 17932 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT6
port 329 nsew signal output
flabel metal3 s 21424 18356 21504 18436 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT7
port 330 nsew signal output
flabel metal3 s 21424 2732 21504 2812 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT0
port 331 nsew signal input
flabel metal3 s 21424 3236 21504 3316 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT1
port 332 nsew signal input
flabel metal3 s 21424 3740 21504 3820 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT2
port 333 nsew signal input
flabel metal3 s 21424 4244 21504 4324 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT3
port 334 nsew signal input
flabel metal3 s 21424 4748 21504 4828 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT4
port 335 nsew signal input
flabel metal3 s 21424 5252 21504 5332 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT5
port 336 nsew signal input
flabel metal3 s 21424 5756 21504 5836 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT6
port 337 nsew signal input
flabel metal3 s 21424 6260 21504 6340 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT7
port 338 nsew signal input
flabel metal2 s 15608 0 15688 80 0 FreeSans 320 0 0 0 UserCLK
port 339 nsew signal input
flabel metal2 s 15608 42928 15688 43008 0 FreeSans 320 0 0 0 UserCLKo
port 340 nsew signal output
flabel metal6 s 4892 0 5332 43008 0 FreeSans 2624 90 0 0 VGND
port 341 nsew ground bidirectional
flabel metal6 s 4892 0 5332 328 0 FreeSans 2624 0 0 0 VGND
port 341 nsew ground bidirectional
flabel metal6 s 4892 42680 5332 43008 0 FreeSans 2624 0 0 0 VGND
port 341 nsew ground bidirectional
flabel metal6 s 20012 0 20452 43008 0 FreeSans 2624 90 0 0 VGND
port 341 nsew ground bidirectional
flabel metal6 s 20012 0 20452 328 0 FreeSans 2624 0 0 0 VGND
port 341 nsew ground bidirectional
flabel metal6 s 20012 42680 20452 43008 0 FreeSans 2624 0 0 0 VGND
port 341 nsew ground bidirectional
flabel metal6 s 3652 0 4092 43008 0 FreeSans 2624 90 0 0 VPWR
port 342 nsew power bidirectional
flabel metal6 s 3652 0 4092 328 0 FreeSans 2624 0 0 0 VPWR
port 342 nsew power bidirectional
flabel metal6 s 3652 42680 4092 43008 0 FreeSans 2624 0 0 0 VPWR
port 342 nsew power bidirectional
flabel metal6 s 18772 0 19212 43008 0 FreeSans 2624 90 0 0 VPWR
port 342 nsew power bidirectional
flabel metal6 s 18772 0 19212 328 0 FreeSans 2624 0 0 0 VPWR
port 342 nsew power bidirectional
flabel metal6 s 18772 42680 19212 43008 0 FreeSans 2624 0 0 0 VPWR
port 342 nsew power bidirectional
flabel metal3 s 0 44 80 124 0 FreeSans 320 0 0 0 W1BEG[0]
port 343 nsew signal output
flabel metal3 s 0 380 80 460 0 FreeSans 320 0 0 0 W1BEG[1]
port 344 nsew signal output
flabel metal3 s 0 716 80 796 0 FreeSans 320 0 0 0 W1BEG[2]
port 345 nsew signal output
flabel metal3 s 0 1052 80 1132 0 FreeSans 320 0 0 0 W1BEG[3]
port 346 nsew signal output
flabel metal3 s 0 1388 80 1468 0 FreeSans 320 0 0 0 W2BEG[0]
port 347 nsew signal output
flabel metal3 s 0 1724 80 1804 0 FreeSans 320 0 0 0 W2BEG[1]
port 348 nsew signal output
flabel metal3 s 0 2060 80 2140 0 FreeSans 320 0 0 0 W2BEG[2]
port 349 nsew signal output
flabel metal3 s 0 2396 80 2476 0 FreeSans 320 0 0 0 W2BEG[3]
port 350 nsew signal output
flabel metal3 s 0 2732 80 2812 0 FreeSans 320 0 0 0 W2BEG[4]
port 351 nsew signal output
flabel metal3 s 0 3068 80 3148 0 FreeSans 320 0 0 0 W2BEG[5]
port 352 nsew signal output
flabel metal3 s 0 3404 80 3484 0 FreeSans 320 0 0 0 W2BEG[6]
port 353 nsew signal output
flabel metal3 s 0 3740 80 3820 0 FreeSans 320 0 0 0 W2BEG[7]
port 354 nsew signal output
flabel metal3 s 0 4076 80 4156 0 FreeSans 320 0 0 0 W2BEGb[0]
port 355 nsew signal output
flabel metal3 s 0 4412 80 4492 0 FreeSans 320 0 0 0 W2BEGb[1]
port 356 nsew signal output
flabel metal3 s 0 4748 80 4828 0 FreeSans 320 0 0 0 W2BEGb[2]
port 357 nsew signal output
flabel metal3 s 0 5084 80 5164 0 FreeSans 320 0 0 0 W2BEGb[3]
port 358 nsew signal output
flabel metal3 s 0 5420 80 5500 0 FreeSans 320 0 0 0 W2BEGb[4]
port 359 nsew signal output
flabel metal3 s 0 5756 80 5836 0 FreeSans 320 0 0 0 W2BEGb[5]
port 360 nsew signal output
flabel metal3 s 0 6092 80 6172 0 FreeSans 320 0 0 0 W2BEGb[6]
port 361 nsew signal output
flabel metal3 s 0 6428 80 6508 0 FreeSans 320 0 0 0 W2BEGb[7]
port 362 nsew signal output
flabel metal3 s 0 12140 80 12220 0 FreeSans 320 0 0 0 W6BEG[0]
port 363 nsew signal output
flabel metal3 s 0 15500 80 15580 0 FreeSans 320 0 0 0 W6BEG[10]
port 364 nsew signal output
flabel metal3 s 0 15836 80 15916 0 FreeSans 320 0 0 0 W6BEG[11]
port 365 nsew signal output
flabel metal3 s 0 12476 80 12556 0 FreeSans 320 0 0 0 W6BEG[1]
port 366 nsew signal output
flabel metal3 s 0 12812 80 12892 0 FreeSans 320 0 0 0 W6BEG[2]
port 367 nsew signal output
flabel metal3 s 0 13148 80 13228 0 FreeSans 320 0 0 0 W6BEG[3]
port 368 nsew signal output
flabel metal3 s 0 13484 80 13564 0 FreeSans 320 0 0 0 W6BEG[4]
port 369 nsew signal output
flabel metal3 s 0 13820 80 13900 0 FreeSans 320 0 0 0 W6BEG[5]
port 370 nsew signal output
flabel metal3 s 0 14156 80 14236 0 FreeSans 320 0 0 0 W6BEG[6]
port 371 nsew signal output
flabel metal3 s 0 14492 80 14572 0 FreeSans 320 0 0 0 W6BEG[7]
port 372 nsew signal output
flabel metal3 s 0 14828 80 14908 0 FreeSans 320 0 0 0 W6BEG[8]
port 373 nsew signal output
flabel metal3 s 0 15164 80 15244 0 FreeSans 320 0 0 0 W6BEG[9]
port 374 nsew signal output
flabel metal3 s 0 6764 80 6844 0 FreeSans 320 0 0 0 WW4BEG[0]
port 375 nsew signal output
flabel metal3 s 0 10124 80 10204 0 FreeSans 320 0 0 0 WW4BEG[10]
port 376 nsew signal output
flabel metal3 s 0 10460 80 10540 0 FreeSans 320 0 0 0 WW4BEG[11]
port 377 nsew signal output
flabel metal3 s 0 10796 80 10876 0 FreeSans 320 0 0 0 WW4BEG[12]
port 378 nsew signal output
flabel metal3 s 0 11132 80 11212 0 FreeSans 320 0 0 0 WW4BEG[13]
port 379 nsew signal output
flabel metal3 s 0 11468 80 11548 0 FreeSans 320 0 0 0 WW4BEG[14]
port 380 nsew signal output
flabel metal3 s 0 11804 80 11884 0 FreeSans 320 0 0 0 WW4BEG[15]
port 381 nsew signal output
flabel metal3 s 0 7100 80 7180 0 FreeSans 320 0 0 0 WW4BEG[1]
port 382 nsew signal output
flabel metal3 s 0 7436 80 7516 0 FreeSans 320 0 0 0 WW4BEG[2]
port 383 nsew signal output
flabel metal3 s 0 7772 80 7852 0 FreeSans 320 0 0 0 WW4BEG[3]
port 384 nsew signal output
flabel metal3 s 0 8108 80 8188 0 FreeSans 320 0 0 0 WW4BEG[4]
port 385 nsew signal output
flabel metal3 s 0 8444 80 8524 0 FreeSans 320 0 0 0 WW4BEG[5]
port 386 nsew signal output
flabel metal3 s 0 8780 80 8860 0 FreeSans 320 0 0 0 WW4BEG[6]
port 387 nsew signal output
flabel metal3 s 0 9116 80 9196 0 FreeSans 320 0 0 0 WW4BEG[7]
port 388 nsew signal output
flabel metal3 s 0 9452 80 9532 0 FreeSans 320 0 0 0 WW4BEG[8]
port 389 nsew signal output
flabel metal3 s 0 9788 80 9868 0 FreeSans 320 0 0 0 WW4BEG[9]
port 390 nsew signal output
rlabel metal1 10802 41580 10802 41580 0 VGND
rlabel metal1 10752 40824 10752 40824 0 VPWR
rlabel metal3 21426 23436 21426 23436 0 CLK_TT_PROJECT
rlabel metal2 8544 16086 8544 16086 0 E1END[0]
rlabel metal2 11424 16338 11424 16338 0 E1END[1]
rlabel metal3 654 16884 654 16884 0 E1END[2]
rlabel metal3 2430 17220 2430 17220 0 E1END[3]
rlabel metal2 2016 16086 2016 16086 0 E2END[0]
rlabel metal3 15504 18816 15504 18816 0 E2END[1]
rlabel metal2 16320 35280 16320 35280 0 E2END[2]
rlabel metal2 1248 31962 1248 31962 0 E2END[3]
rlabel metal2 1920 35364 1920 35364 0 E2END[4]
rlabel metal4 16560 14952 16560 14952 0 E2END[5]
rlabel metal2 18480 18564 18480 18564 0 E2END[6]
rlabel metal3 942 22596 942 22596 0 E2END[7]
rlabel metal3 1806 17556 1806 17556 0 E2MID[0]
rlabel metal2 15264 18396 15264 18396 0 E2MID[1]
rlabel metal2 2304 18480 2304 18480 0 E2MID[2]
rlabel metal2 8112 17052 8112 17052 0 E2MID[3]
rlabel metal3 1086 18900 1086 18900 0 E2MID[4]
rlabel metal3 1086 19236 1086 19236 0 E2MID[5]
rlabel metal2 17760 20664 17760 20664 0 E2MID[6]
rlabel metal2 6432 19908 6432 19908 0 E2MID[7]
rlabel metal2 1872 35700 1872 35700 0 E6END[0]
rlabel metal2 13824 19194 13824 19194 0 E6END[10]
rlabel metal3 414 32004 414 32004 0 E6END[11]
rlabel metal2 13632 27678 13632 27678 0 E6END[1]
rlabel metal3 126 28980 126 28980 0 E6END[2]
rlabel metal3 510 29316 510 29316 0 E6END[3]
rlabel metal2 4944 23772 4944 23772 0 E6END[4]
rlabel metal2 2112 30408 2112 30408 0 E6END[5]
rlabel metal3 606 30324 606 30324 0 E6END[6]
rlabel metal3 1632 30534 1632 30534 0 E6END[7]
rlabel metal3 462 30996 462 30996 0 E6END[8]
rlabel metal3 17568 30660 17568 30660 0 E6END[9]
rlabel metal2 3648 17850 3648 17850 0 EE4END[0]
rlabel metal3 15408 33684 15408 33684 0 EE4END[10]
rlabel metal3 4272 27720 4272 27720 0 EE4END[11]
rlabel metal3 126 26964 126 26964 0 EE4END[12]
rlabel metal2 18336 27426 18336 27426 0 EE4END[13]
rlabel metal2 19200 31080 19200 31080 0 EE4END[14]
rlabel metal3 1290 27972 1290 27972 0 EE4END[15]
rlabel metal2 16080 29232 16080 29232 0 EE4END[1]
rlabel metal2 14688 31920 14688 31920 0 EE4END[2]
rlabel metal3 366 23940 366 23940 0 EE4END[3]
rlabel metal2 8928 24444 8928 24444 0 EE4END[4]
rlabel metal3 654 24612 654 24612 0 EE4END[5]
rlabel metal3 126 24948 126 24948 0 EE4END[6]
rlabel metal2 5472 26040 5472 26040 0 EE4END[7]
rlabel metal2 2112 17430 2112 17430 0 EE4END[8]
rlabel metal3 126 25956 126 25956 0 EE4END[9]
rlabel metal2 18480 21756 18480 21756 0 ENA_TT_PROJECT
rlabel metal3 13872 1092 13872 1092 0 FrameData[0]
rlabel metal2 1728 19194 1728 19194 0 FrameData[10]
rlabel metal3 1584 17724 1584 17724 0 FrameData[11]
rlabel metal2 1344 19908 1344 19908 0 FrameData[12]
rlabel metal2 14400 17094 14400 17094 0 FrameData[13]
rlabel metal3 126 37044 126 37044 0 FrameData[14]
rlabel metal3 13776 12012 13776 12012 0 FrameData[15]
rlabel metal2 1920 17892 1920 17892 0 FrameData[16]
rlabel metal3 1296 14700 1296 14700 0 FrameData[17]
rlabel metal3 13248 35868 13248 35868 0 FrameData[18]
rlabel metal3 1248 37212 1248 37212 0 FrameData[19]
rlabel metal3 654 32676 654 32676 0 FrameData[1]
rlabel metal2 1248 27678 1248 27678 0 FrameData[20]
rlabel metal3 2112 31080 2112 31080 0 FrameData[21]
rlabel metal2 11904 15036 11904 15036 0 FrameData[22]
rlabel metal2 11424 36246 11424 36246 0 FrameData[23]
rlabel metal2 1536 1554 1536 1554 0 FrameData[24]
rlabel metal2 12576 33621 12576 33621 0 FrameData[25]
rlabel metal2 14112 32760 14112 32760 0 FrameData[26]
rlabel metal2 1632 34020 1632 34020 0 FrameData[27]
rlabel metal2 2448 36456 2448 36456 0 FrameData[28]
rlabel metal2 1248 32844 1248 32844 0 FrameData[29]
rlabel metal3 654 33012 654 33012 0 FrameData[2]
rlabel metal2 1248 29862 1248 29862 0 FrameData[30]
rlabel metal2 2064 29148 2064 29148 0 FrameData[31]
rlabel metal3 18048 1932 18048 1932 0 FrameData[3]
rlabel metal3 654 33684 654 33684 0 FrameData[4]
rlabel metal3 17184 18816 17184 18816 0 FrameData[5]
rlabel metal3 510 34356 510 34356 0 FrameData[6]
rlabel metal2 2256 36708 2256 36708 0 FrameData[7]
rlabel metal2 1344 12264 1344 12264 0 FrameData[8]
rlabel metal2 1296 11676 1296 11676 0 FrameData[9]
rlabel metal3 20754 24444 20754 24444 0 FrameData_O[0]
rlabel metal3 21042 29484 21042 29484 0 FrameData_O[10]
rlabel metal2 17568 28602 17568 28602 0 FrameData_O[11]
rlabel via3 21426 30492 21426 30492 0 FrameData_O[12]
rlabel metal3 19584 38766 19584 38766 0 FrameData_O[13]
rlabel metal2 19776 39060 19776 39060 0 FrameData_O[14]
rlabel metal3 19152 38472 19152 38472 0 FrameData_O[15]
rlabel metal3 19776 39018 19776 39018 0 FrameData_O[16]
rlabel metal3 21090 33012 21090 33012 0 FrameData_O[17]
rlabel metal3 21138 33516 21138 33516 0 FrameData_O[18]
rlabel metal3 21138 34020 21138 34020 0 FrameData_O[19]
rlabel via2 21426 24948 21426 24948 0 FrameData_O[1]
rlabel metal4 8352 36330 8352 36330 0 FrameData_O[20]
rlabel metal3 16896 34188 16896 34188 0 FrameData_O[21]
rlabel metal3 21090 35532 21090 35532 0 FrameData_O[22]
rlabel metal2 11616 36246 11616 36246 0 FrameData_O[23]
rlabel metal2 19392 40446 19392 40446 0 FrameData_O[24]
rlabel metal4 12768 38346 12768 38346 0 FrameData_O[25]
rlabel metal3 21330 37548 21330 37548 0 FrameData_O[26]
rlabel metal4 19392 38766 19392 38766 0 FrameData_O[27]
rlabel metal2 13104 34608 13104 34608 0 FrameData_O[28]
rlabel metal3 18048 30492 18048 30492 0 FrameData_O[29]
rlabel metal2 19872 26292 19872 26292 0 FrameData_O[2]
rlabel metal3 16944 29232 16944 29232 0 FrameData_O[30]
rlabel metal2 17232 38976 17232 38976 0 FrameData_O[31]
rlabel metal3 20994 25956 20994 25956 0 FrameData_O[3]
rlabel via2 21426 26460 21426 26460 0 FrameData_O[4]
rlabel metal2 19968 27216 19968 27216 0 FrameData_O[5]
rlabel metal2 19968 27846 19968 27846 0 FrameData_O[6]
rlabel metal2 19392 28476 19392 28476 0 FrameData_O[7]
rlabel metal2 20400 31164 20400 31164 0 FrameData_O[8]
rlabel metal4 19968 30492 19968 30492 0 FrameData_O[9]
rlabel metal2 12672 28056 12672 28056 0 FrameStrobe[0]
rlabel metal2 17760 660 17760 660 0 FrameStrobe[10]
rlabel metal2 17952 240 17952 240 0 FrameStrobe[11]
rlabel metal2 18144 156 18144 156 0 FrameStrobe[12]
rlabel metal2 18336 660 18336 660 0 FrameStrobe[13]
rlabel metal2 18528 618 18528 618 0 FrameStrobe[14]
rlabel metal2 18720 450 18720 450 0 FrameStrobe[15]
rlabel metal2 18912 450 18912 450 0 FrameStrobe[16]
rlabel metal2 19104 450 19104 450 0 FrameStrobe[17]
rlabel metal2 19296 366 19296 366 0 FrameStrobe[18]
rlabel metal2 19488 282 19488 282 0 FrameStrobe[19]
rlabel metal2 12192 1974 12192 1974 0 FrameStrobe[1]
rlabel metal3 18912 30660 18912 30660 0 FrameStrobe[2]
rlabel metal2 2496 11550 2496 11550 0 FrameStrobe[3]
rlabel metal3 13728 18144 13728 18144 0 FrameStrobe[4]
rlabel metal2 14976 15414 14976 15414 0 FrameStrobe[5]
rlabel metal2 19248 1932 19248 1932 0 FrameStrobe[6]
rlabel metal2 16992 1386 16992 1386 0 FrameStrobe[7]
rlabel metal2 2400 35994 2400 35994 0 FrameStrobe[8]
rlabel metal2 2496 29484 2496 29484 0 FrameStrobe[9]
rlabel metal3 17328 40656 17328 40656 0 FrameStrobe_O[0]
rlabel metal2 18432 41454 18432 41454 0 FrameStrobe_O[10]
rlabel metal2 12672 34146 12672 34146 0 FrameStrobe_O[11]
rlabel metal2 18144 42264 18144 42264 0 FrameStrobe_O[12]
rlabel metal2 18336 42348 18336 42348 0 FrameStrobe_O[13]
rlabel metal2 18528 42474 18528 42474 0 FrameStrobe_O[14]
rlabel metal2 13248 38430 13248 38430 0 FrameStrobe_O[15]
rlabel metal3 15744 34944 15744 34944 0 FrameStrobe_O[16]
rlabel metal2 13632 38556 13632 38556 0 FrameStrobe_O[17]
rlabel metal2 14400 36414 14400 36414 0 FrameStrobe_O[18]
rlabel metal2 14064 35028 14064 35028 0 FrameStrobe_O[19]
rlabel metal2 19584 41790 19584 41790 0 FrameStrobe_O[1]
rlabel metal2 18048 39942 18048 39942 0 FrameStrobe_O[2]
rlabel metal3 15648 33012 15648 33012 0 FrameStrobe_O[3]
rlabel metal2 19968 40698 19968 40698 0 FrameStrobe_O[4]
rlabel metal4 16656 31920 16656 31920 0 FrameStrobe_O[5]
rlabel metal2 14976 18816 14976 18816 0 FrameStrobe_O[6]
rlabel metal2 17184 42138 17184 42138 0 FrameStrobe_O[7]
rlabel metal2 17376 42390 17376 42390 0 FrameStrobe_O[8]
rlabel metal2 13680 34944 13680 34944 0 FrameStrobe_O[9]
rlabel metal3 9600 1008 9600 1008 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit0.Q
rlabel metal2 12864 1218 12864 1218 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit1.Q
rlabel metal2 3408 36876 3408 36876 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit10.Q
rlabel metal2 5808 36540 5808 36540 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit11.Q
rlabel metal3 9936 37884 9936 37884 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit12.Q
rlabel metal2 8544 36960 8544 36960 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit13.Q
rlabel metal2 8832 36211 8832 36211 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit14.Q
rlabel metal2 7296 36834 7296 36834 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit15.Q
rlabel metal3 7200 33096 7200 33096 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit16.Q
rlabel metal2 4872 37394 4872 37394 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit17.Q
rlabel metal3 7824 38892 7824 38892 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit18.Q
rlabel metal2 9696 39109 9696 39109 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit19.Q
rlabel metal2 12192 25830 12192 25830 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit2.Q
rlabel metal3 8208 40404 8208 40404 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit20.Q
rlabel metal2 11520 40705 11520 40705 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit21.Q
rlabel metal2 5616 34608 5616 34608 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit22.Q
rlabel via2 7200 39729 7200 39729 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit23.Q
rlabel metal3 3312 2604 3312 2604 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit24.Q
rlabel metal2 3984 1932 3984 1932 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit25.Q
rlabel metal2 13152 29316 13152 29316 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit26.Q
rlabel metal3 13008 28560 13008 28560 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit27.Q
rlabel via1 14208 40407 14208 40407 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit28.Q
rlabel metal2 14400 39774 14400 39774 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit29.Q
rlabel metal2 13728 25585 13728 25585 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit3.Q
rlabel metal2 9408 31500 9408 31500 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit30.Q
rlabel metal2 9888 31122 9888 31122 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit31.Q
rlabel metal2 11472 35196 11472 35196 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit4.Q
rlabel metal2 13056 35445 13056 35445 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit5.Q
rlabel metal2 9264 18732 9264 18732 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit6.Q
rlabel metal2 10848 20325 10848 20325 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit7.Q
rlabel metal3 12054 38724 12054 38724 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit8.Q
rlabel metal3 12672 40908 12672 40908 0 Inst_E_TT_IF_ConfigMem.Inst_frame0_bit9.Q
rlabel metal2 5856 27384 5856 27384 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit0.Q
rlabel metal2 5808 25284 5808 25284 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit1.Q
rlabel metal2 14592 23142 14592 23142 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit10.Q
rlabel via1 16176 23094 16176 23094 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit11.Q
rlabel metal2 11376 37380 11376 37380 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit12.Q
rlabel metal2 13200 36876 13200 36876 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit13.Q
rlabel metal2 7680 12180 7680 12180 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit14.Q
rlabel metal3 9360 14196 9360 14196 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit15.Q
rlabel metal3 9456 8988 9456 8988 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit16.Q
rlabel metal2 10848 8701 10848 8701 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit17.Q
rlabel metal2 14496 24066 14496 24066 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit18.Q
rlabel metal2 16080 23835 16080 23835 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit19.Q
rlabel metal3 17184 21000 17184 21000 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit2.Q
rlabel metal2 10848 39144 10848 39144 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit20.Q
rlabel metal2 12384 39529 12384 39529 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit21.Q
rlabel metal2 7488 16716 7488 16716 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit22.Q
rlabel metal2 9744 15708 9744 15708 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit23.Q
rlabel metal2 9024 2142 9024 2142 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit24.Q
rlabel metal2 12000 2310 12000 2310 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit25.Q
rlabel metal3 14784 21000 14784 21000 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit26.Q
rlabel via1 16272 21583 16272 21583 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit27.Q
rlabel metal2 11136 38808 11136 38808 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit28.Q
rlabel metal2 12672 38847 12672 38847 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit29.Q
rlabel metal2 18048 21042 18048 21042 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit3.Q
rlabel metal2 8064 17556 8064 17556 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit30.Q
rlabel metal2 10800 18732 10800 18732 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit31.Q
rlabel metal2 7776 34230 7776 34230 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit4.Q
rlabel metal3 8352 37632 8352 37632 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit5.Q
rlabel metal2 3936 32844 3936 32844 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit6.Q
rlabel metal3 6432 35028 6432 35028 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit7.Q
rlabel metal2 9264 2856 9264 2856 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit8.Q
rlabel metal2 10272 4620 10272 4620 0 Inst_E_TT_IF_ConfigMem.Inst_frame1_bit9.Q
rlabel metal2 6720 25116 6720 25116 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit0.Q
rlabel metal2 19488 25788 19488 25788 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit1.Q
rlabel metal2 7584 19236 7584 19236 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit10.Q
rlabel metal2 1920 16842 1920 16842 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit11.Q
rlabel metal2 2880 19614 2880 19614 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit12.Q
rlabel metal2 17184 26250 17184 26250 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit13.Q
rlabel metal2 15744 26082 15744 26082 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit14.Q
rlabel metal2 17280 26166 17280 26166 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit15.Q
rlabel metal3 16944 35196 16944 35196 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit16.Q
rlabel metal2 14880 36918 14880 36918 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit17.Q
rlabel metal2 14784 35658 14784 35658 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit18.Q
rlabel metal2 4128 26082 4128 26082 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit19.Q
rlabel metal2 18960 26796 18960 26796 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit2.Q
rlabel metal3 4464 27636 4464 27636 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit20.Q
rlabel metal2 1344 26754 1344 26754 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit21.Q
rlabel metal2 10752 22050 10752 22050 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit22.Q
rlabel metal3 10368 22260 10368 22260 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit23.Q
rlabel metal2 11520 23226 11520 23226 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit24.Q
rlabel metal2 19824 22932 19824 22932 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit25.Q
rlabel metal2 20064 22890 20064 22890 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit26.Q
rlabel metal2 20147 22212 20147 22212 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit27.Q
rlabel metal2 19584 31668 19584 31668 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit28.Q
rlabel metal2 17664 33348 17664 33348 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit29.Q
rlabel metal2 17328 25200 17328 25200 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit3.Q
rlabel metal2 19584 30702 19584 30702 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit30.Q
rlabel metal3 6912 28392 6912 28392 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit31.Q
rlabel metal2 19488 34650 19488 34650 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit4.Q
rlabel metal3 19536 35868 19536 35868 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit5.Q
rlabel metal2 16752 33852 16752 33852 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit6.Q
rlabel metal2 7584 27090 7584 27090 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit7.Q
rlabel metal2 8352 27972 8352 27972 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit8.Q
rlabel metal2 8256 25830 8256 25830 0 Inst_E_TT_IF_ConfigMem.Inst_frame2_bit9.Q
rlabel metal2 9552 13440 9552 13440 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit0.Q
rlabel metal2 11328 13727 11328 13727 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit1.Q
rlabel metal2 4176 15708 4176 15708 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit10.Q
rlabel metal3 4080 17052 4080 17052 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit11.Q
rlabel metal2 14736 17220 14736 17220 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit12.Q
rlabel metal2 13104 17220 13104 17220 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit13.Q
rlabel metal2 15648 15960 15648 15960 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit14.Q
rlabel metal2 17280 16506 17280 16506 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit15.Q
rlabel metal2 2784 16513 2784 16513 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit16.Q
rlabel metal3 3504 14952 3504 14952 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit17.Q
rlabel metal2 3264 22050 3264 22050 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit18.Q
rlabel metal2 3024 18564 3024 18564 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit19.Q
rlabel metal2 3168 13986 3168 13986 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit2.Q
rlabel metal2 4416 20706 4416 20706 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit20.Q
rlabel metal2 15504 29652 15504 29652 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit21.Q
rlabel metal3 16800 27594 16800 27594 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit22.Q
rlabel metal2 14688 27888 14688 27888 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit23.Q
rlabel metal2 14208 33642 14208 33642 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit24.Q
rlabel metal3 14640 32844 14640 32844 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit25.Q
rlabel metal2 12672 33138 12672 33138 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit26.Q
rlabel metal2 1728 29568 1728 29568 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit27.Q
rlabel metal2 2304 30828 2304 30828 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit28.Q
rlabel metal2 2256 31332 2256 31332 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit29.Q
rlabel metal3 3312 11424 3312 11424 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit3.Q
rlabel metal2 8352 23898 8352 23898 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit30.Q
rlabel metal2 8544 24192 8544 24192 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit31.Q
rlabel metal3 13536 13440 13536 13440 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit4.Q
rlabel metal2 12048 14700 12048 14700 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit5.Q
rlabel metal2 16224 14364 16224 14364 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit6.Q
rlabel metal3 16608 14112 16608 14112 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit7.Q
rlabel metal2 2688 13020 2688 13020 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit8.Q
rlabel metal2 2736 11928 2736 11928 0 Inst_E_TT_IF_ConfigMem.Inst_frame3_bit9.Q
rlabel metal2 11088 1260 11088 1260 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit0.Q
rlabel metal2 9408 714 9408 714 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit1.Q
rlabel metal2 3456 10119 3456 10119 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit10.Q
rlabel metal2 2784 5334 2784 5334 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit11.Q
rlabel metal3 13920 13104 13920 13104 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit12.Q
rlabel metal2 12576 13314 12576 13314 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit13.Q
rlabel metal2 16656 11739 16656 11739 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit14.Q
rlabel metal2 15072 11508 15072 11508 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit15.Q
rlabel metal2 2784 7644 2784 7644 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit16.Q
rlabel metal2 2496 7224 2496 7224 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit17.Q
rlabel metal2 6912 11048 6912 11048 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit18.Q
rlabel metal2 5328 11172 5328 11172 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit19.Q
rlabel metal3 4416 6636 4416 6636 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit2.Q
rlabel metal2 13728 11977 13728 11977 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit20.Q
rlabel metal2 12192 11634 12192 11634 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit21.Q
rlabel metal2 15456 12555 15456 12555 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit22.Q
rlabel metal2 16944 11928 16944 11928 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit23.Q
rlabel via2 2208 3441 2208 3441 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit24.Q
rlabel metal2 3744 3486 3744 3486 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit25.Q
rlabel metal2 10176 7434 10176 7434 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit26.Q
rlabel metal2 11856 6636 11856 6636 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit27.Q
rlabel metal2 12288 21630 12288 21630 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit28.Q
rlabel metal2 13824 21837 13824 21837 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit29.Q
rlabel metal2 2880 3822 2880 3822 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit3.Q
rlabel metal2 12192 30702 12192 30702 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit30.Q
rlabel via1 13776 30655 13776 30655 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit31.Q
rlabel metal2 13920 6888 13920 6888 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit4.Q
rlabel metal2 12288 7434 12288 7434 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit5.Q
rlabel metal2 13440 9660 13440 9660 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit6.Q
rlabel metal2 15072 11046 15072 11046 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit7.Q
rlabel metal2 8880 3612 8880 3612 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit8.Q
rlabel metal2 2592 4998 2592 4998 0 Inst_E_TT_IF_ConfigMem.Inst_frame4_bit9.Q
rlabel metal2 7584 1512 7584 1512 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit0.Q
rlabel metal2 4464 4620 4464 4620 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit1.Q
rlabel metal2 19872 3402 19872 3402 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit10.Q
rlabel metal3 2928 8148 2928 8148 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit11.Q
rlabel metal2 3072 11459 3072 11459 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit12.Q
rlabel metal2 3072 9744 3072 9744 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit13.Q
rlabel metal2 7296 14109 7296 14109 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit14.Q
rlabel metal2 5760 13734 5760 13734 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit15.Q
rlabel metal2 4656 11844 4656 11844 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit16.Q
rlabel metal2 16656 8904 16656 8904 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit17.Q
rlabel metal2 15072 9198 15072 9198 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit18.Q
rlabel metal3 16944 9492 16944 9492 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit19.Q
rlabel metal2 4416 4410 4416 4410 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit2.Q
rlabel metal2 17664 19278 17664 19278 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit20.Q
rlabel via2 17652 18564 17652 18564 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit21.Q
rlabel metal2 15168 18732 15168 18732 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit22.Q
rlabel metal3 5760 9492 5760 9492 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit23.Q
rlabel metal2 6816 8946 6816 8946 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit24.Q
rlabel metal2 7008 8148 7008 8148 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit25.Q
rlabel metal2 7008 7441 7008 7441 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit26.Q
rlabel metal2 5280 6006 5280 6006 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit27.Q
rlabel metal2 15168 15960 15168 15960 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit28.Q
rlabel metal2 13488 15372 13488 15372 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit29.Q
rlabel metal2 5616 2436 5616 2436 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit3.Q
rlabel metal2 14784 7434 14784 7434 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit30.Q
rlabel metal2 16704 8022 16704 8022 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit31.Q
rlabel metal2 3456 5376 3456 5376 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit4.Q
rlabel metal2 18336 18144 18336 18144 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit5.Q
rlabel metal2 19714 19824 19714 19824 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit6.Q
rlabel metal2 19680 19572 19680 19572 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit7.Q
rlabel metal2 18048 6510 18048 6510 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit8.Q
rlabel metal2 17856 3864 17856 3864 0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit9.Q
rlabel metal2 16704 1680 16704 1680 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit0.Q
rlabel metal2 17664 1470 17664 1470 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit1.Q
rlabel metal2 9024 7056 9024 7056 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit10.Q
rlabel metal2 7392 6846 7392 6846 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit11.Q
rlabel metal2 9792 7434 9792 7434 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit12.Q
rlabel metal2 17760 14910 17760 14910 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit13.Q
rlabel metal3 18624 13860 18624 13860 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit14.Q
rlabel metal2 19968 12894 19968 12894 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit15.Q
rlabel metal2 19776 9786 19776 9786 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit16.Q
rlabel metal2 18864 10416 18864 10416 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit17.Q
rlabel metal2 20147 8562 20147 8562 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit18.Q
rlabel metal2 9072 11928 9072 11928 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit19.Q
rlabel via1 19344 3439 19344 3439 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit2.Q
rlabel metal3 7680 11970 7680 11970 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit20.Q
rlabel metal2 7824 12348 7824 12348 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit21.Q
rlabel metal2 11904 8694 11904 8694 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit22.Q
rlabel metal2 12864 8316 12864 8316 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit23.Q
rlabel metal2 13008 8652 13008 8652 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit24.Q
rlabel metal2 16416 6426 16416 6426 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit25.Q
rlabel metal3 19968 2100 19968 2100 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit26.Q
rlabel metal2 20448 1932 20448 1932 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit27.Q
rlabel metal2 19152 16212 19152 16212 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit28.Q
rlabel metal2 19872 16296 19872 16296 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit29.Q
rlabel metal2 19392 1386 19392 1386 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit3.Q
rlabel metal2 19008 15792 19008 15792 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit30.Q
rlabel metal2 7248 1764 7248 1764 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit31.Q
rlabel metal2 13536 5586 13536 5586 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit4.Q
rlabel metal2 15072 5929 15072 5929 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit5.Q
rlabel metal2 15552 4872 15552 4872 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit6.Q
rlabel metal2 11904 5082 11904 5082 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit7.Q
rlabel via1 13008 4120 13008 4120 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit8.Q
rlabel metal2 14208 2940 14208 2940 0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit9.Q
rlabel metal2 6144 21294 6144 21294 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit0.Q
rlabel metal2 7824 21000 7824 21000 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit1.Q
rlabel via2 7104 16214 7104 16214 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit10.Q
rlabel metal3 7248 15708 7248 15708 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit11.Q
rlabel metal2 7680 15036 7680 15036 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit12.Q
rlabel metal2 11664 15708 11664 15708 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit13.Q
rlabel metal3 10272 17220 10272 17220 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit14.Q
rlabel metal2 12432 17787 12432 17787 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit15.Q
rlabel metal2 7392 15584 7392 15584 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit16.Q
rlabel metal2 5856 17682 5856 17682 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit17.Q
rlabel metal2 11904 24353 11904 24353 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit18.Q
rlabel metal2 12048 23100 12048 23100 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit19.Q
rlabel metal3 5808 19488 5808 19488 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit2.Q
rlabel metal2 12000 24157 12000 24157 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit20.Q
rlabel metal2 18576 28980 18576 28980 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit21.Q
rlabel metal2 19584 29778 19584 29778 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit22.Q
rlabel metal2 17952 28098 17952 28098 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit23.Q
rlabel metal2 18816 37170 18816 37170 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit24.Q
rlabel metal2 20592 37464 20592 37464 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit25.Q
rlabel metal2 18048 35658 18048 35658 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit26.Q
rlabel metal2 9216 29400 9216 29400 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit27.Q
rlabel metal3 9888 29064 9888 29064 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit28.Q
rlabel metal2 8736 29232 8736 29232 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit29.Q
rlabel metal2 7776 18732 7776 18732 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit3.Q
rlabel metal2 15264 2310 15264 2310 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit30.Q
rlabel via1 16560 2634 16560 2634 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit31.Q
rlabel metal2 10560 32214 10560 32214 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit4.Q
rlabel metal2 12096 32421 12096 32421 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit5.Q
rlabel metal3 13920 18732 13920 18732 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit6.Q
rlabel metal2 12384 19824 12384 19824 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit7.Q
rlabel metal2 8064 22561 8064 22561 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit8.Q
rlabel metal3 6288 21756 6288 21756 0 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit9.Q
rlabel metal2 6144 33180 6144 33180 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit0.Q
rlabel metal3 5952 33054 5952 33054 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit1.Q
rlabel via1 12240 33679 12240 33679 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit10.Q
rlabel metal2 10656 33936 10656 33936 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit11.Q
rlabel metal2 3648 29694 3648 29694 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit12.Q
rlabel metal2 2112 37471 2112 37471 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit13.Q
rlabel metal2 2496 24192 2496 24192 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit14.Q
rlabel metal3 4560 25200 4560 25200 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit15.Q
rlabel metal2 3456 24234 3456 24234 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit16.Q
rlabel metal2 14112 30954 14112 30954 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit17.Q
rlabel metal3 17472 29778 17472 29778 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit18.Q
rlabel metal2 17856 30450 17856 30450 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit19.Q
rlabel metal2 2880 30156 2880 30156 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit2.Q
rlabel metal2 15888 38220 15888 38220 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit20.Q
rlabel metal2 16128 37926 16128 37926 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit21.Q
rlabel metal2 14880 37842 14880 37842 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit22.Q
rlabel metal2 6336 30492 6336 30492 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit23.Q
rlabel metal2 6240 32382 6240 32382 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit24.Q
rlabel metal2 5664 30324 5664 30324 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit25.Q
rlabel metal2 5616 18732 5616 18732 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit26.Q
rlabel metal2 7104 19537 7104 19537 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit27.Q
rlabel metal2 11712 26847 11712 26847 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit28.Q
rlabel via1 13307 26805 13307 26805 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit29.Q
rlabel metal2 2016 33054 2016 33054 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit3.Q
rlabel metal2 13344 19194 13344 19194 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit30.Q
rlabel metal2 14880 19537 14880 19537 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit31.Q
rlabel metal3 5712 33768 5712 33768 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit4.Q
rlabel metal2 1344 34986 1344 34986 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit5.Q
rlabel metal4 3600 36120 3600 36120 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit6.Q
rlabel metal2 3552 35952 3552 35952 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit7.Q
rlabel metal2 1632 39557 1632 39557 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit8.Q
rlabel metal3 12288 40950 12288 40950 0 Inst_E_TT_IF_ConfigMem.Inst_frame8_bit9.Q
rlabel metal2 3360 23520 3360 23520 0 Inst_E_TT_IF_ConfigMem.Inst_frame9_bit22.Q
rlabel metal2 6240 23268 6240 23268 0 Inst_E_TT_IF_ConfigMem.Inst_frame9_bit23.Q
rlabel metal2 11568 29820 11568 29820 0 Inst_E_TT_IF_ConfigMem.Inst_frame9_bit24.Q
rlabel metal2 13152 30499 13152 30499 0 Inst_E_TT_IF_ConfigMem.Inst_frame9_bit25.Q
rlabel metal2 16128 39984 16128 39984 0 Inst_E_TT_IF_ConfigMem.Inst_frame9_bit26.Q
rlabel metal2 17760 39396 17760 39396 0 Inst_E_TT_IF_ConfigMem.Inst_frame9_bit27.Q
rlabel metal2 6144 31500 6144 31500 0 Inst_E_TT_IF_ConfigMem.Inst_frame9_bit28.Q
rlabel via1 7680 31360 7680 31360 0 Inst_E_TT_IF_ConfigMem.Inst_frame9_bit29.Q
rlabel metal2 2016 28644 2016 28644 0 Inst_E_TT_IF_ConfigMem.Inst_frame9_bit30.Q
rlabel metal2 3552 28609 3552 28609 0 Inst_E_TT_IF_ConfigMem.Inst_frame9_bit31.Q
rlabel metal3 8016 29820 8016 29820 0 Inst_E_TT_IF_switch_matrix.N1BEG0
rlabel metal4 1248 32214 1248 32214 0 Inst_E_TT_IF_switch_matrix.N1BEG1
rlabel metal3 18576 39900 18576 39900 0 Inst_E_TT_IF_switch_matrix.N1BEG2
rlabel metal3 1536 38178 1536 38178 0 Inst_E_TT_IF_switch_matrix.N1BEG3
rlabel metal3 1248 34440 1248 34440 0 Inst_E_TT_IF_switch_matrix.N2BEG0
rlabel metal2 2304 33978 2304 33978 0 Inst_E_TT_IF_switch_matrix.N2BEG1
rlabel metal3 3456 32340 3456 32340 0 Inst_E_TT_IF_switch_matrix.N2BEG2
rlabel metal3 3408 35112 3408 35112 0 Inst_E_TT_IF_switch_matrix.N2BEG3
rlabel metal2 1536 35112 1536 35112 0 Inst_E_TT_IF_switch_matrix.N2BEG4
rlabel metal2 1536 37632 1536 37632 0 Inst_E_TT_IF_switch_matrix.N2BEG5
rlabel metal2 12384 34566 12384 34566 0 Inst_E_TT_IF_switch_matrix.N2BEG6
rlabel metal3 1584 37716 1584 37716 0 Inst_E_TT_IF_switch_matrix.N2BEG7
rlabel metal5 4656 31332 4656 31332 0 Inst_E_TT_IF_switch_matrix.N4BEG0
rlabel metal3 12432 31920 12432 31920 0 Inst_E_TT_IF_switch_matrix.N4BEG1
rlabel metal2 18144 38682 18144 38682 0 Inst_E_TT_IF_switch_matrix.N4BEG2
rlabel via1 4037 34944 4037 34944 0 Inst_E_TT_IF_switch_matrix.N4BEG3
rlabel metal5 11088 12096 11088 12096 0 Inst_E_TT_IF_switch_matrix.S1BEG0
rlabel metal3 15648 1008 15648 1008 0 Inst_E_TT_IF_switch_matrix.S1BEG1
rlabel metal4 17232 15288 17232 15288 0 Inst_E_TT_IF_switch_matrix.S1BEG2
rlabel metal3 13536 3780 13536 3780 0 Inst_E_TT_IF_switch_matrix.S1BEG3
rlabel metal3 5376 1848 5376 1848 0 Inst_E_TT_IF_switch_matrix.S2BEG0
rlabel metal5 12184 31416 12184 31416 0 Inst_E_TT_IF_switch_matrix.S2BEG1
rlabel metal3 14352 17052 14352 17052 0 Inst_E_TT_IF_switch_matrix.S2BEG2
rlabel metal4 10560 11424 10560 11424 0 Inst_E_TT_IF_switch_matrix.S2BEG3
rlabel metal3 6960 2688 6960 2688 0 Inst_E_TT_IF_switch_matrix.S2BEG4
rlabel metal4 11760 13608 11760 13608 0 Inst_E_TT_IF_switch_matrix.S2BEG5
rlabel metal2 14784 11718 14784 11718 0 Inst_E_TT_IF_switch_matrix.S2BEG6
rlabel metal4 1296 16716 1296 16716 0 Inst_E_TT_IF_switch_matrix.S2BEG7
rlabel metal5 13392 5040 13392 5040 0 Inst_E_TT_IF_switch_matrix.S4BEG0
rlabel metal3 20496 29988 20496 29988 0 Inst_E_TT_IF_switch_matrix.S4BEG1
rlabel metal3 19008 13692 19008 13692 0 Inst_E_TT_IF_switch_matrix.S4BEG2
rlabel metal3 1056 1848 1056 1848 0 Inst_E_TT_IF_switch_matrix.S4BEG3
rlabel metal2 17664 7014 17664 7014 0 Inst_E_TT_IF_switch_matrix.W1BEG0
rlabel metal3 20544 2268 20544 2268 0 Inst_E_TT_IF_switch_matrix.W1BEG1
rlabel metal2 13920 4242 13920 4242 0 Inst_E_TT_IF_switch_matrix.W1BEG2
rlabel metal3 16656 10584 16656 10584 0 Inst_E_TT_IF_switch_matrix.W1BEG3
rlabel metal4 12384 11130 12384 11130 0 Inst_E_TT_IF_switch_matrix.W2BEG0
rlabel metal2 14304 11718 14304 11718 0 Inst_E_TT_IF_switch_matrix.W2BEG1
rlabel metal3 19584 12264 19584 12264 0 Inst_E_TT_IF_switch_matrix.W2BEG2
rlabel metal2 10032 11760 10032 11760 0 Inst_E_TT_IF_switch_matrix.W2BEG3
rlabel metal4 1632 22344 1632 22344 0 Inst_E_TT_IF_switch_matrix.W2BEG4
rlabel metal3 13968 14196 13968 14196 0 Inst_E_TT_IF_switch_matrix.W2BEG5
rlabel metal3 14256 13272 14256 13272 0 Inst_E_TT_IF_switch_matrix.W2BEG6
rlabel metal2 9168 8666 9168 8666 0 Inst_E_TT_IF_switch_matrix.W2BEG7
rlabel metal3 2160 6636 2160 6636 0 Inst_E_TT_IF_switch_matrix.W2BEGb0
rlabel metal2 1536 19824 1536 19824 0 Inst_E_TT_IF_switch_matrix.W2BEGb1
rlabel metal2 13776 7056 13776 7056 0 Inst_E_TT_IF_switch_matrix.W2BEGb2
rlabel metal2 10656 3528 10656 3528 0 Inst_E_TT_IF_switch_matrix.W2BEGb3
rlabel metal3 6192 12432 6192 12432 0 Inst_E_TT_IF_switch_matrix.W2BEGb4
rlabel metal2 15840 8232 15840 8232 0 Inst_E_TT_IF_switch_matrix.W2BEGb5
rlabel metal2 2208 15960 2208 15960 0 Inst_E_TT_IF_switch_matrix.W2BEGb6
rlabel metal3 4080 12264 4080 12264 0 Inst_E_TT_IF_switch_matrix.W2BEGb7
rlabel metal2 2208 8309 2208 8309 0 Inst_E_TT_IF_switch_matrix.W6BEG0
rlabel metal2 1440 21588 1440 21588 0 Inst_E_TT_IF_switch_matrix.W6BEG1
rlabel metal2 15552 15750 15552 15750 0 Inst_E_TT_IF_switch_matrix.W6BEG10
rlabel metal2 1824 16254 1824 16254 0 Inst_E_TT_IF_switch_matrix.W6BEG11
rlabel metal2 14256 27552 14256 27552 0 Inst_E_TT_IF_switch_matrix.W6BEG2
rlabel metal2 2304 9366 2304 9366 0 Inst_E_TT_IF_switch_matrix.W6BEG3
rlabel metal2 4800 16002 4800 16002 0 Inst_E_TT_IF_switch_matrix.W6BEG4
rlabel metal2 12624 12432 12624 12432 0 Inst_E_TT_IF_switch_matrix.W6BEG5
rlabel metal2 1440 13482 1440 13482 0 Inst_E_TT_IF_switch_matrix.W6BEG6
rlabel metal2 2592 14028 2592 14028 0 Inst_E_TT_IF_switch_matrix.W6BEG7
rlabel metal3 1440 16422 1440 16422 0 Inst_E_TT_IF_switch_matrix.W6BEG8
rlabel metal3 14976 17808 14976 17808 0 Inst_E_TT_IF_switch_matrix.W6BEG9
rlabel metal3 6096 10248 6096 10248 0 Inst_E_TT_IF_switch_matrix.WW4BEG0
rlabel metal3 15792 16044 15792 16044 0 Inst_E_TT_IF_switch_matrix.WW4BEG1
rlabel metal3 16896 11424 16896 11424 0 Inst_E_TT_IF_switch_matrix.WW4BEG10
rlabel metal2 4597 8702 4597 8702 0 Inst_E_TT_IF_switch_matrix.WW4BEG11
rlabel metal3 5952 10500 5952 10500 0 Inst_E_TT_IF_switch_matrix.WW4BEG12
rlabel metal2 1440 6930 1440 6930 0 Inst_E_TT_IF_switch_matrix.WW4BEG13
rlabel metal4 13920 8652 13920 8652 0 Inst_E_TT_IF_switch_matrix.WW4BEG14
rlabel metal3 1392 11592 1392 11592 0 Inst_E_TT_IF_switch_matrix.WW4BEG15
rlabel metal2 15024 8148 15024 8148 0 Inst_E_TT_IF_switch_matrix.WW4BEG2
rlabel metal3 8400 16380 8400 16380 0 Inst_E_TT_IF_switch_matrix.WW4BEG3
rlabel metal2 1920 5838 1920 5838 0 Inst_E_TT_IF_switch_matrix.WW4BEG4
rlabel metal2 1824 6636 1824 6636 0 Inst_E_TT_IF_switch_matrix.WW4BEG5
rlabel metal2 13344 11004 13344 11004 0 Inst_E_TT_IF_switch_matrix.WW4BEG6
rlabel metal2 12288 6132 12288 6132 0 Inst_E_TT_IF_switch_matrix.WW4BEG7
rlabel metal4 1536 7686 1536 7686 0 Inst_E_TT_IF_switch_matrix.WW4BEG8
rlabel metal3 14016 14112 14016 14112 0 Inst_E_TT_IF_switch_matrix.WW4BEG9
rlabel metal2 1824 42600 1824 42600 0 N1BEG[0]
rlabel metal2 2016 41550 2016 41550 0 N1BEG[1]
rlabel via2 2208 42936 2208 42936 0 N1BEG[2]
rlabel metal2 1728 38514 1728 38514 0 N1BEG[3]
rlabel metal2 1824 576 1824 576 0 N1END[0]
rlabel metal2 2016 534 2016 534 0 N1END[1]
rlabel metal2 2208 744 2208 744 0 N1END[2]
rlabel metal2 2400 240 2400 240 0 N1END[3]
rlabel metal3 2208 34608 2208 34608 0 N2BEG[0]
rlabel metal2 2016 35280 2016 35280 0 N2BEG[1]
rlabel metal2 4608 37296 4608 37296 0 N2BEG[2]
rlabel metal3 3456 34944 3456 34944 0 N2BEG[3]
rlabel metal3 1872 36120 1872 36120 0 N2BEG[4]
rlabel metal2 1776 37632 1776 37632 0 N2BEG[5]
rlabel metal2 3744 42642 3744 42642 0 N2BEG[6]
rlabel metal2 1488 39060 1488 39060 0 N2BEG[7]
rlabel metal2 1536 36876 1536 36876 0 N2BEGb[0]
rlabel metal2 4416 37338 4416 37338 0 N2BEGb[1]
rlabel metal2 1536 41496 1536 41496 0 N2BEGb[2]
rlabel metal2 4080 36120 4080 36120 0 N2BEGb[3]
rlabel metal2 4032 37254 4032 37254 0 N2BEGb[4]
rlabel metal2 1632 41622 1632 41622 0 N2BEGb[5]
rlabel metal4 2112 38808 2112 38808 0 N2BEGb[6]
rlabel metal2 1728 32382 1728 32382 0 N2BEGb[7]
rlabel metal2 4128 576 4128 576 0 N2END[0]
rlabel metal3 672 29064 672 29064 0 N2END[1]
rlabel metal4 1152 15162 1152 15162 0 N2END[2]
rlabel metal6 2152 14238 2152 14238 0 N2END[3]
rlabel metal5 1148 5376 1148 5376 0 N2END[4]
rlabel metal2 5088 324 5088 324 0 N2END[5]
rlabel metal2 5280 114 5280 114 0 N2END[6]
rlabel metal2 384 11466 384 11466 0 N2END[7]
rlabel metal2 1248 37128 1248 37128 0 N2MID[0]
rlabel metal3 1056 29064 1056 29064 0 N2MID[1]
rlabel metal5 5376 12600 5376 12600 0 N2MID[2]
rlabel metal4 912 29148 912 29148 0 N2MID[3]
rlabel metal2 1344 35658 1344 35658 0 N2MID[4]
rlabel metal4 1440 40404 1440 40404 0 N2MID[5]
rlabel metal2 1632 38724 1632 38724 0 N2MID[6]
rlabel metal2 3936 324 3936 324 0 N2MID[7]
rlabel metal3 5184 37632 5184 37632 0 N4BEG[0]
rlabel metal2 7584 41802 7584 41802 0 N4BEG[10]
rlabel metal2 2208 40530 2208 40530 0 N4BEG[11]
rlabel metal2 3456 33474 3456 33474 0 N4BEG[12]
rlabel metal2 5856 41118 5856 41118 0 N4BEG[13]
rlabel metal2 19968 42084 19968 42084 0 N4BEG[14]
rlabel metal3 3120 38724 3120 38724 0 N4BEG[15]
rlabel metal2 2592 38094 2592 38094 0 N4BEG[1]
rlabel metal2 2976 38472 2976 38472 0 N4BEG[2]
rlabel metal2 6240 42264 6240 42264 0 N4BEG[3]
rlabel metal3 6192 36876 6192 36876 0 N4BEG[4]
rlabel metal2 7680 41034 7680 41034 0 N4BEG[5]
rlabel metal2 5280 39900 5280 39900 0 N4BEG[6]
rlabel metal3 7728 38724 7728 38724 0 N4BEG[7]
rlabel metal2 7104 39354 7104 39354 0 N4BEG[8]
rlabel metal2 4704 40068 4704 40068 0 N4BEG[9]
rlabel metal2 10464 1806 10464 1806 0 N4END[0]
rlabel metal2 7584 576 7584 576 0 N4END[10]
rlabel metal2 7776 492 7776 492 0 N4END[11]
rlabel metal2 7968 366 7968 366 0 N4END[12]
rlabel metal2 8160 660 8160 660 0 N4END[13]
rlabel metal3 1488 40320 1488 40320 0 N4END[14]
rlabel metal3 1296 38976 1296 38976 0 N4END[15]
rlabel metal2 11664 6300 11664 6300 0 N4END[1]
rlabel metal2 12288 30618 12288 30618 0 N4END[2]
rlabel metal2 8448 14616 8448 14616 0 N4END[3]
rlabel metal4 192 32760 192 32760 0 N4END[4]
rlabel metal4 2400 38220 2400 38220 0 N4END[5]
rlabel metal2 6816 660 6816 660 0 N4END[6]
rlabel metal2 7008 660 7008 660 0 N4END[7]
rlabel metal2 7200 660 7200 660 0 N4END[8]
rlabel metal2 7392 492 7392 492 0 N4END[9]
rlabel metal2 13824 32592 13824 32592 0 RST_N_TT_PROJECT
rlabel metal3 9360 2772 9360 2772 0 S1BEG[0]
rlabel metal2 16896 798 16896 798 0 S1BEG[1]
rlabel metal2 17280 2184 17280 2184 0 S1BEG[2]
rlabel metal2 14784 3066 14784 3066 0 S1BEG[3]
rlabel metal3 8544 11928 8544 11928 0 S1END[0]
rlabel metal3 17568 3444 17568 3444 0 S1END[1]
rlabel metal2 14111 19656 14111 19656 0 S1END[2]
rlabel metal2 11904 4494 11904 4494 0 S1END[3]
rlabel metal2 9504 618 9504 618 0 S2BEG[0]
rlabel metal2 9696 660 9696 660 0 S2BEG[1]
rlabel metal2 9888 1164 9888 1164 0 S2BEG[2]
rlabel metal2 10368 1848 10368 1848 0 S2BEG[3]
rlabel metal3 7344 2436 7344 2436 0 S2BEG[4]
rlabel metal3 2208 1638 2208 1638 0 S2BEG[5]
rlabel metal3 14688 11508 14688 11508 0 S2BEG[6]
rlabel metal2 10848 492 10848 492 0 S2BEG[7]
rlabel metal2 1824 1512 1824 1512 0 S2BEGb[0]
rlabel metal2 7584 2352 7584 2352 0 S2BEGb[1]
rlabel metal2 11424 450 11424 450 0 S2BEGb[2]
rlabel metal3 14256 2436 14256 2436 0 S2BEGb[3]
rlabel metal2 11808 870 11808 870 0 S2BEGb[4]
rlabel metal2 12000 870 12000 870 0 S2BEGb[5]
rlabel metal2 12192 912 12192 912 0 S2BEGb[6]
rlabel metal2 12384 282 12384 282 0 S2BEGb[7]
rlabel metal2 11040 42348 11040 42348 0 S2END[0]
rlabel metal2 5376 36162 5376 36162 0 S2END[1]
rlabel metal2 11424 41424 11424 41424 0 S2END[2]
rlabel metal2 11616 40794 11616 40794 0 S2END[3]
rlabel metal2 11808 41676 11808 41676 0 S2END[4]
rlabel metal2 12000 42516 12000 42516 0 S2END[5]
rlabel metal2 12192 42054 12192 42054 0 S2END[6]
rlabel metal2 12384 42726 12384 42726 0 S2END[7]
rlabel metal2 1632 1638 1632 1638 0 S2MID[0]
rlabel metal3 13680 2100 13680 2100 0 S2MID[1]
rlabel metal2 5088 1092 5088 1092 0 S2MID[2]
rlabel metal5 14784 3192 14784 3192 0 S2MID[3]
rlabel metal5 9380 2100 9380 2100 0 S2MID[4]
rlabel metal2 17568 2184 17568 2184 0 S2MID[5]
rlabel metal2 1824 3066 1824 3066 0 S2MID[6]
rlabel metal2 10752 41076 10752 41076 0 S2MID[7]
rlabel metal2 12576 660 12576 660 0 S4BEG[0]
rlabel metal3 16752 35784 16752 35784 0 S4BEG[10]
rlabel metal2 14688 660 14688 660 0 S4BEG[11]
rlabel metal2 14880 744 14880 744 0 S4BEG[12]
rlabel metal3 20592 2436 20592 2436 0 S4BEG[13]
rlabel metal2 15264 324 15264 324 0 S4BEG[14]
rlabel metal2 15456 660 15456 660 0 S4BEG[15]
rlabel metal2 12768 660 12768 660 0 S4BEG[1]
rlabel metal2 12960 660 12960 660 0 S4BEG[2]
rlabel metal2 13296 2940 13296 2940 0 S4BEG[3]
rlabel metal2 13344 534 13344 534 0 S4BEG[4]
rlabel metal2 13536 660 13536 660 0 S4BEG[5]
rlabel metal2 13728 660 13728 660 0 S4BEG[6]
rlabel metal2 13920 786 13920 786 0 S4BEG[7]
rlabel metal3 16416 10836 16416 10836 0 S4BEG[8]
rlabel metal2 14304 492 14304 492 0 S4BEG[9]
rlabel metal2 12576 42264 12576 42264 0 S4END[0]
rlabel metal2 14496 42306 14496 42306 0 S4END[10]
rlabel metal2 14688 42474 14688 42474 0 S4END[11]
rlabel metal2 14880 42054 14880 42054 0 S4END[12]
rlabel metal2 15072 42516 15072 42516 0 S4END[13]
rlabel metal2 15264 42726 15264 42726 0 S4END[14]
rlabel metal2 15456 42180 15456 42180 0 S4END[15]
rlabel metal2 15552 23184 15552 23184 0 S4END[1]
rlabel metal2 12576 36288 12576 36288 0 S4END[2]
rlabel metal2 13152 42306 13152 42306 0 S4END[3]
rlabel metal2 13344 42264 13344 42264 0 S4END[4]
rlabel metal2 13536 42222 13536 42222 0 S4END[5]
rlabel metal2 13728 42432 13728 42432 0 S4END[6]
rlabel metal2 13920 42180 13920 42180 0 S4END[7]
rlabel metal2 14112 42348 14112 42348 0 S4END[8]
rlabel metal2 14304 42642 14304 42642 0 S4END[9]
rlabel metal2 7680 19572 7680 19572 0 UIO_IN_TT_PROJECT0
rlabel metal2 17376 19866 17376 19866 0 UIO_IN_TT_PROJECT1
rlabel metal2 17856 34524 17856 34524 0 UIO_IN_TT_PROJECT2
rlabel metal4 15744 23310 15744 23310 0 UIO_IN_TT_PROJECT3
rlabel metal2 10176 21168 10176 21168 0 UIO_IN_TT_PROJECT4
rlabel metal3 20466 21420 20466 21420 0 UIO_IN_TT_PROJECT5
rlabel metal2 19488 29568 19488 29568 0 UIO_IN_TT_PROJECT6
rlabel metal4 14976 26418 14976 26418 0 UIO_IN_TT_PROJECT7
rlabel metal2 15360 3570 15360 3570 0 UIO_OE_TT_PROJECT0
rlabel metal3 19488 15582 19488 15582 0 UIO_OE_TT_PROJECT1
rlabel metal3 19344 11424 19344 11424 0 UIO_OE_TT_PROJECT2
rlabel metal2 2400 4746 2400 4746 0 UIO_OE_TT_PROJECT3
rlabel metal3 14208 12810 14208 12810 0 UIO_OE_TT_PROJECT4
rlabel metal3 15936 13020 15936 13020 0 UIO_OE_TT_PROJECT5
rlabel metal2 19584 13440 19584 13440 0 UIO_OE_TT_PROJECT6
rlabel metal4 16320 4158 16320 4158 0 UIO_OE_TT_PROJECT7
rlabel metal4 15744 6762 15744 6762 0 UIO_OUT_TT_PROJECT0
rlabel metal3 19440 13188 19440 13188 0 UIO_OUT_TT_PROJECT1
rlabel metal2 17184 16254 17184 16254 0 UIO_OUT_TT_PROJECT2
rlabel metal3 6528 13944 6528 13944 0 UIO_OUT_TT_PROJECT3
rlabel metal2 12192 8778 12192 8778 0 UIO_OUT_TT_PROJECT4
rlabel metal2 17568 7182 17568 7182 0 UIO_OUT_TT_PROJECT5
rlabel metal2 19392 16002 19392 16002 0 UIO_OUT_TT_PROJECT6
rlabel metal3 13824 10374 13824 10374 0 UIO_OUT_TT_PROJECT7
rlabel metal3 21330 14868 21330 14868 0 UI_IN_TT_PROJECT0
rlabel metal3 18096 29064 18096 29064 0 UI_IN_TT_PROJECT1
rlabel metal3 19296 30240 19296 30240 0 UI_IN_TT_PROJECT2
rlabel metal3 1824 29148 1824 29148 0 UI_IN_TT_PROJECT3
rlabel metal4 16320 19908 16320 19908 0 UI_IN_TT_PROJECT4
rlabel metal2 19584 25830 19584 25830 0 UI_IN_TT_PROJECT5
rlabel metal4 19488 25704 19488 25704 0 UI_IN_TT_PROJECT6
rlabel metal4 16704 22050 16704 22050 0 UI_IN_TT_PROJECT7
rlabel metal2 5568 6972 5568 6972 0 UO_OUT_TT_PROJECT0
rlabel metal2 12000 4074 12000 4074 0 UO_OUT_TT_PROJECT1
rlabel metal3 16752 11676 16752 11676 0 UO_OUT_TT_PROJECT2
rlabel metal2 18336 3654 18336 3654 0 UO_OUT_TT_PROJECT3
rlabel metal3 20946 4788 20946 4788 0 UO_OUT_TT_PROJECT4
rlabel metal2 12768 14364 12768 14364 0 UO_OUT_TT_PROJECT5
rlabel metal2 15072 10668 15072 10668 0 UO_OUT_TT_PROJECT6
rlabel metal3 15696 2604 15696 2604 0 UO_OUT_TT_PROJECT7
rlabel metal2 15648 660 15648 660 0 UserCLK
rlabel metal2 15072 34062 15072 34062 0 UserCLKo
rlabel metal3 174 84 174 84 0 W1BEG[0]
rlabel metal3 366 420 366 420 0 W1BEG[1]
rlabel metal3 126 756 126 756 0 W1BEG[2]
rlabel metal3 78 1092 78 1092 0 W1BEG[3]
rlabel metal3 558 1428 558 1428 0 W2BEG[0]
rlabel metal3 1230 1764 1230 1764 0 W2BEG[1]
rlabel metal3 414 2100 414 2100 0 W2BEG[2]
rlabel metal3 654 2436 654 2436 0 W2BEG[3]
rlabel metal3 462 2772 462 2772 0 W2BEG[4]
rlabel metal3 174 3108 174 3108 0 W2BEG[5]
rlabel metal4 11424 12474 11424 12474 0 W2BEG[6]
rlabel metal3 960 12432 960 12432 0 W2BEG[7]
rlabel metal3 768 15036 768 15036 0 W2BEGb[0]
rlabel metal5 1440 16212 1440 16212 0 W2BEGb[1]
rlabel metal3 654 4788 654 4788 0 W2BEGb[2]
rlabel metal3 1290 5124 1290 5124 0 W2BEGb[3]
rlabel metal3 3360 5544 3360 5544 0 W2BEGb[4]
rlabel metal3 174 5796 174 5796 0 W2BEGb[5]
rlabel metal3 990 6132 990 6132 0 W2BEGb[6]
rlabel metal3 366 6468 366 6468 0 W2BEGb[7]
rlabel metal3 1086 12180 1086 12180 0 W6BEG[0]
rlabel metal3 798 15540 798 15540 0 W6BEG[10]
rlabel metal3 798 15876 798 15876 0 W6BEG[11]
rlabel metal3 126 12516 126 12516 0 W6BEG[1]
rlabel metal3 126 12852 126 12852 0 W6BEG[2]
rlabel metal3 510 13188 510 13188 0 W6BEG[3]
rlabel metal4 4608 14322 4608 14322 0 W6BEG[4]
rlabel metal3 270 13860 270 13860 0 W6BEG[5]
rlabel metal2 1248 13734 1248 13734 0 W6BEG[6]
rlabel metal2 1248 14364 1248 14364 0 W6BEG[7]
rlabel metal3 654 14868 654 14868 0 W6BEG[8]
rlabel metal4 14976 16590 14976 16590 0 W6BEG[9]
rlabel metal3 78 6804 78 6804 0 WW4BEG[0]
rlabel metal2 240 924 240 924 0 WW4BEG[10]
rlabel metal2 4368 8820 4368 8820 0 WW4BEG[11]
rlabel metal3 318 10836 318 10836 0 WW4BEG[12]
rlabel metal2 1248 7308 1248 7308 0 WW4BEG[13]
rlabel metal3 990 11508 990 11508 0 WW4BEG[14]
rlabel metal3 318 11844 318 11844 0 WW4BEG[15]
rlabel metal3 126 7140 126 7140 0 WW4BEG[1]
rlabel metal3 414 7476 414 7476 0 WW4BEG[2]
rlabel metal3 1344 17640 1344 17640 0 WW4BEG[3]
rlabel metal2 1728 5544 1728 5544 0 WW4BEG[4]
rlabel metal2 1584 6636 1584 6636 0 WW4BEG[5]
rlabel metal3 126 8820 126 8820 0 WW4BEG[6]
rlabel metal4 10080 7896 10080 7896 0 WW4BEG[7]
rlabel metal2 1200 4788 1200 4788 0 WW4BEG[8]
rlabel metal2 1392 3612 1392 3612 0 WW4BEG[9]
rlabel metal2 1344 32466 1344 32466 0 _0000_
rlabel metal2 10560 28434 10560 28434 0 _0001_
rlabel metal2 9072 29484 9072 29484 0 _0002_
rlabel metal2 5664 25998 5664 25998 0 _0003_
rlabel metal2 17280 38430 17280 38430 0 _0004_
rlabel metal3 12720 36540 12720 36540 0 _0005_
rlabel metal2 18576 35364 18576 35364 0 _0006_
rlabel metal2 13440 28602 13440 28602 0 _0007_
rlabel metal2 19200 23436 19200 23436 0 _0008_
rlabel metal2 12144 7728 12144 7728 0 _0009_
rlabel metal2 11904 22470 11904 22470 0 _0010_
rlabel metal2 3648 26067 3648 26067 0 _0011_
rlabel metal2 15168 36897 15168 36897 0 _0012_
rlabel metal2 17376 26544 17376 26544 0 _0013_
rlabel metal2 5568 17472 5568 17472 0 _0014_
rlabel metal2 19104 34398 19104 34398 0 _0015_
rlabel metal3 19632 24612 19632 24612 0 _0016_
rlabel metal2 9600 24486 9600 24486 0 _0017_
rlabel metal2 3072 30744 3072 30744 0 _0018_
rlabel metal2 14592 34188 14592 34188 0 _0019_
rlabel metal2 16320 27384 16320 27384 0 _0020_
rlabel metal2 4416 21672 4416 21672 0 _0021_
rlabel metal3 14112 10164 14112 10164 0 _0022_
rlabel metal3 19920 14700 19920 14700 0 _0023_
rlabel metal2 14592 6510 14592 6510 0 _0024_
rlabel metal2 13152 8400 13152 8400 0 _0025_
rlabel metal2 11520 5964 11520 5964 0 _0026_
rlabel metal2 10512 12516 10512 12516 0 _0027_
rlabel metal2 18048 10122 18048 10122 0 _0028_
rlabel metal2 18336 4284 18336 4284 0 _0029_
rlabel metal2 10272 6509 10272 6509 0 _0030_
rlabel metal2 9456 29400 9456 29400 0 _0031_
rlabel metal2 19008 37464 19008 37464 0 _0032_
rlabel metal2 6720 29946 6720 29946 0 _0033_
rlabel metal2 16608 36624 16608 36624 0 _0034_
rlabel metal2 17376 33138 17376 33138 0 _0035_
rlabel metal2 4398 24661 4398 24661 0 _0036_
rlabel metal2 14496 39396 14496 39396 0 _0037_
rlabel metal3 6336 35448 6336 35448 0 _0038_
rlabel metal2 9024 33810 9024 33810 0 _0039_
rlabel metal2 6048 34776 6048 34776 0 _0040_
rlabel metal2 4608 35574 4608 35574 0 _0041_
rlabel metal2 10272 32886 10272 32886 0 _0042_
rlabel metal2 4320 32886 4320 32886 0 _0043_
rlabel metal3 9888 36036 9888 36036 0 _0044_
rlabel metal2 8256 32382 8256 32382 0 _0045_
rlabel metal2 8640 38724 8640 38724 0 _0046_
rlabel metal2 6432 35784 6432 35784 0 _0047_
rlabel metal2 6528 36204 6528 36204 0 _0048_
rlabel metal2 10032 32844 10032 32844 0 _0049_
rlabel metal3 9168 31416 9168 31416 0 _0050_
rlabel metal2 6720 6888 6720 6888 0 _0051_
rlabel metal3 5856 14700 5856 14700 0 _0052_
rlabel metal3 7104 14952 7104 14952 0 _0053_
rlabel metal2 6144 26628 6144 26628 0 _0054_
rlabel metal2 6946 26032 6946 26032 0 _0055_
rlabel metal2 6528 26880 6528 26880 0 _0056_
rlabel metal2 7008 26670 7008 26670 0 _0057_
rlabel metal3 6000 27132 6000 27132 0 _0058_
rlabel metal2 6336 27678 6336 27678 0 _0059_
rlabel metal2 17760 19362 17760 19362 0 _0060_
rlabel metal2 11904 18564 11904 18564 0 _0061_
rlabel metal2 17280 17766 17280 17766 0 _0062_
rlabel metal2 19872 31080 19872 31080 0 _0063_
rlabel metal2 18754 31507 18754 31507 0 _0064_
rlabel metal2 19296 32172 19296 32172 0 _0065_
rlabel metal2 19488 31248 19488 31248 0 _0066_
rlabel metal2 19872 32634 19872 32634 0 _0067_
rlabel metal2 19968 32634 19968 32634 0 _0068_
rlabel metal3 18288 17640 18288 17640 0 _0069_
rlabel metal2 14160 17724 14160 17724 0 _0070_
rlabel metal2 18048 7560 18048 7560 0 _0071_
rlabel metal2 19680 21504 19680 21504 0 _0072_
rlabel metal2 19042 23863 19042 23863 0 _0073_
rlabel metal3 19344 23772 19344 23772 0 _0074_
rlabel metal2 19296 22260 19296 22260 0 _0075_
rlabel metal2 18816 21966 18816 21966 0 _0076_
rlabel metal2 19584 21546 19584 21546 0 _0077_
rlabel metal3 7584 2016 7584 2016 0 _0078_
rlabel metal2 7584 15918 7584 15918 0 _0079_
rlabel metal2 4704 15036 4704 15036 0 _0080_
rlabel metal2 9984 21630 9984 21630 0 _0081_
rlabel metal2 11293 23050 11293 23050 0 _0082_
rlabel metal2 12000 22470 12000 22470 0 _0083_
rlabel metal2 10368 21756 10368 21756 0 _0084_
rlabel metal2 8832 22596 8832 22596 0 _0085_
rlabel metal3 9504 21504 9504 21504 0 _0086_
rlabel metal3 3312 7224 3312 7224 0 _0087_
rlabel metal2 12480 10416 12480 10416 0 _0088_
rlabel metal2 4416 26376 4416 26376 0 _0089_
rlabel via1 3796 26124 3796 26124 0 _0090_
rlabel via1 3526 26124 3526 26124 0 _0091_
rlabel metal2 4032 26208 4032 26208 0 _0092_
rlabel metal2 3173 26208 3173 26208 0 _0093_
rlabel metal2 4320 25746 4320 25746 0 _0094_
rlabel metal2 12576 14952 12576 14952 0 _0095_
rlabel metal2 13488 17892 13488 17892 0 _0096_
rlabel metal2 18048 35238 18048 35238 0 _0097_
rlabel metal2 16930 35104 16930 35104 0 _0098_
rlabel metal2 17184 35742 17184 35742 0 _0099_
rlabel metal2 17664 35364 17664 35364 0 _0100_
rlabel metal2 15936 35112 15936 35112 0 _0101_
rlabel metal2 15264 35826 15264 35826 0 _0102_
rlabel metal3 19392 19992 19392 19992 0 _0103_
rlabel metal3 13776 12180 13776 12180 0 _0104_
rlabel metal2 16704 25494 16704 25494 0 _0105_
rlabel metal2 16642 25948 16642 25948 0 _0106_
rlabel metal2 16896 26208 16896 26208 0 _0107_
rlabel metal2 17136 25284 17136 25284 0 _0108_
rlabel metal2 16320 26418 16320 26418 0 _0109_
rlabel metal2 16416 26586 16416 26586 0 _0110_
rlabel metal2 12624 2520 12624 2520 0 _0111_
rlabel metal2 4512 13860 4512 13860 0 _0112_
rlabel metal2 7872 19320 7872 19320 0 _0113_
rlabel metal2 5509 17094 5509 17094 0 _0114_
rlabel metal3 4656 18732 4656 18732 0 _0115_
rlabel metal2 7488 18648 7488 18648 0 _0116_
rlabel metal2 2400 19404 2400 19404 0 _0117_
rlabel metal2 7776 19740 7776 19740 0 _0118_
rlabel metal3 9792 27636 9792 27636 0 _0119_
rlabel metal2 10080 17262 10080 17262 0 _0120_
rlabel metal2 9168 26796 9168 26796 0 _0121_
rlabel metal2 9696 26880 9696 26880 0 _0122_
rlabel metal2 9504 27552 9504 27552 0 _0123_
rlabel metal2 9792 27048 9792 27048 0 _0124_
rlabel metal2 6528 24696 6528 24696 0 _0125_
rlabel metal3 8160 24444 8160 24444 0 _0126_
rlabel metal2 13536 17052 13536 17052 0 _0127_
rlabel metal2 19680 33936 19680 33936 0 _0128_
rlabel via1 19005 34356 19005 34356 0 _0129_
rlabel metal2 19248 34356 19248 34356 0 _0130_
rlabel metal2 19296 33936 19296 33936 0 _0131_
rlabel metal2 19968 34482 19968 34482 0 _0132_
rlabel metal2 19584 33558 19584 33558 0 _0133_
rlabel metal2 18240 9660 18240 9660 0 _0134_
rlabel metal2 19776 26208 19776 26208 0 _0135_
rlabel metal2 19138 24520 19138 24520 0 _0136_
rlabel metal2 19872 25368 19872 25368 0 _0137_
rlabel metal2 19488 25074 19488 25074 0 _0138_
rlabel metal2 20150 25452 20150 25452 0 _0139_
rlabel metal2 19680 25914 19680 25914 0 _0140_
rlabel metal3 7008 8484 7008 8484 0 _0141_
rlabel metal3 8304 23100 8304 23100 0 _0142_
rlabel metal2 9442 24520 9442 24520 0 _0143_
rlabel metal2 9696 24276 9696 24276 0 _0144_
rlabel metal2 8928 23394 8928 23394 0 _0145_
rlabel metal2 9312 25410 9312 25410 0 _0146_
rlabel metal2 8640 23982 8640 23982 0 _0147_
rlabel metal2 4608 17262 4608 17262 0 _0148_
rlabel metal2 1440 30324 1440 30324 0 _0149_
rlabel via1 4418 32172 4418 32172 0 _0150_
rlabel metal2 3072 30366 3072 30366 0 _0151_
rlabel metal2 1824 29652 1824 29652 0 _0152_
rlabel metal3 4752 28392 4752 28392 0 _0153_
rlabel metal3 2832 29064 2832 29064 0 _0154_
rlabel metal2 12672 11802 12672 11802 0 _0155_
rlabel metal3 15744 30660 15744 30660 0 _0156_
rlabel metal2 14693 33516 14693 33516 0 _0157_
rlabel metal3 14976 33096 14976 33096 0 _0158_
rlabel metal2 15072 31332 15072 31332 0 _0159_
rlabel metal2 15648 32298 15648 32298 0 _0160_
rlabel metal2 15360 30954 15360 30954 0 _0161_
rlabel metal2 19776 12474 19776 12474 0 _0162_
rlabel metal3 15888 29316 15888 29316 0 _0163_
rlabel metal2 15997 28441 15997 28441 0 _0164_
rlabel metal2 16416 27972 16416 27972 0 _0165_
rlabel metal3 15936 29064 15936 29064 0 _0166_
rlabel metal2 16128 27678 16128 27678 0 _0167_
rlabel metal3 16464 28140 16464 28140 0 _0168_
rlabel metal2 3744 16002 3744 16002 0 _0169_
rlabel metal2 2976 22554 2976 22554 0 _0170_
rlabel via1 4109 22260 4109 22260 0 _0171_
rlabel metal3 4128 21420 4128 21420 0 _0172_
rlabel metal2 3360 22050 3360 22050 0 _0173_
rlabel metal3 4032 19908 4032 19908 0 _0174_
rlabel metal2 3072 22134 3072 22134 0 _0175_
rlabel metal2 6720 5880 6720 5880 0 _0176_
rlabel metal2 5184 8946 5184 8946 0 _0177_
rlabel metal2 6288 5880 6288 5880 0 _0178_
rlabel metal2 7104 6636 7104 6636 0 _0179_
rlabel metal3 5808 6552 5808 6552 0 _0180_
rlabel metal3 5184 7140 5184 7140 0 _0181_
rlabel metal2 7872 9534 7872 9534 0 _0182_
rlabel metal2 5184 7182 5184 7182 0 _0183_
rlabel metal2 17568 18144 17568 18144 0 _0184_
rlabel metal2 17472 17304 17472 17304 0 _0185_
rlabel metal2 17136 16884 17136 16884 0 _0186_
rlabel via1 17184 19244 17184 19244 0 _0187_
rlabel metal2 17280 17220 17280 17220 0 _0188_
rlabel metal2 17856 17094 17856 17094 0 _0189_
rlabel metal2 15360 18522 15360 18522 0 _0190_
rlabel metal2 17664 17682 17664 17682 0 _0191_
rlabel metal2 17472 8148 17472 8148 0 _0192_
rlabel metal3 17808 8148 17808 8148 0 _0193_
rlabel metal2 17328 7980 17328 7980 0 _0194_
rlabel metal2 17088 9156 17088 9156 0 _0195_
rlabel metal2 17856 8736 17856 8736 0 _0196_
rlabel metal2 15936 7476 15936 7476 0 _0197_
rlabel metal2 17472 9576 17472 9576 0 _0198_
rlabel metal2 15744 7854 15744 7854 0 _0199_
rlabel metal2 4992 14112 4992 14112 0 _0200_
rlabel metal2 4848 12516 4848 12516 0 _0201_
rlabel metal2 5616 12516 5616 12516 0 _0202_
rlabel metal2 5472 12852 5472 12852 0 _0203_
rlabel metal2 5088 12605 5088 12605 0 _0204_
rlabel metal2 5136 12264 5136 12264 0 _0205_
rlabel metal2 7440 11676 7440 11676 0 _0206_
rlabel metal2 7488 11970 7488 11970 0 _0207_
rlabel metal2 4800 12012 4800 12012 0 _0208_
rlabel metal2 4848 11508 4848 11508 0 _0209_
rlabel metal2 1536 12600 1536 12600 0 _0210_
rlabel metal2 1728 14196 1728 14196 0 _0211_
rlabel metal2 2496 14028 2496 14028 0 _0212_
rlabel metal2 3648 8442 3648 8442 0 _0213_
rlabel metal2 1632 10836 1632 10836 0 _0214_
rlabel metal2 3456 8610 3456 8610 0 _0215_
rlabel metal2 18336 5796 18336 5796 0 _0216_
rlabel metal2 20256 6552 20256 6552 0 _0217_
rlabel metal2 17424 3612 17424 3612 0 _0218_
rlabel metal2 19776 3486 19776 3486 0 _0219_
rlabel metal2 19920 3612 19920 3612 0 _0220_
rlabel metal3 15120 11844 15120 11844 0 _0221_
rlabel metal2 19580 2436 19580 2436 0 _0222_
rlabel metal3 19632 2100 19632 2100 0 _0223_
rlabel metal2 19584 19698 19584 19698 0 _0224_
rlabel metal2 20016 17724 20016 17724 0 _0225_
rlabel metal2 18144 18522 18144 18522 0 _0226_
rlabel metal2 19968 20412 19968 20412 0 _0227_
rlabel metal2 20400 17724 20400 17724 0 _0228_
rlabel metal3 19968 18858 19968 18858 0 _0229_
rlabel metal3 19680 18732 19680 18732 0 _0230_
rlabel metal2 17952 20916 17952 20916 0 _0231_
rlabel metal2 5472 3864 5472 3864 0 _0232_
rlabel metal2 3264 2688 3264 2688 0 _0233_
rlabel metal2 6336 3696 6336 3696 0 _0234_
rlabel metal2 6576 3612 6576 3612 0 _0235_
rlabel metal2 3072 3318 3072 3318 0 _0236_
rlabel metal2 2112 3234 2112 3234 0 _0237_
rlabel metal3 2460 6468 2460 6468 0 _0238_
rlabel metal2 2208 6384 2208 6384 0 _0239_
rlabel metal2 9696 3108 9696 3108 0 _0240_
rlabel metal2 11328 3234 11328 3234 0 _0241_
rlabel metal3 6576 19236 6576 19236 0 _0242_
rlabel metal2 8544 4788 8544 4788 0 _0243_
rlabel metal2 8640 3696 8640 3696 0 _0244_
rlabel metal3 19776 15708 19776 15708 0 _0245_
rlabel metal2 19680 14574 19680 14574 0 _0246_
rlabel metal2 18144 15498 18144 15498 0 _0247_
rlabel metal2 13056 28644 13056 28644 0 _0248_
rlabel metal2 13824 27888 13824 27888 0 _0249_
rlabel metal2 12624 29064 12624 29064 0 _0250_
rlabel metal2 18816 15584 18816 15584 0 _0251_
rlabel metal3 18960 14700 18960 14700 0 _0252_
rlabel metal2 18720 14994 18720 14994 0 _0253_
rlabel metal2 19104 14742 19104 14742 0 _0254_
rlabel metal2 18432 14658 18432 14658 0 _0255_
rlabel metal2 18672 14532 18672 14532 0 _0256_
rlabel metal2 19968 16002 19968 16002 0 _0257_
rlabel metal2 19008 14868 19008 14868 0 _0258_
rlabel metal2 16032 6174 16032 6174 0 _0259_
rlabel metal2 16224 5082 16224 5082 0 _0260_
rlabel metal2 14016 40152 14016 40152 0 _0261_
rlabel metal2 14304 40320 14304 40320 0 _0262_
rlabel metal2 14400 19320 14400 19320 0 _0263_
rlabel via2 14305 7141 14305 7141 0 _0264_
rlabel metal2 19584 7098 19584 7098 0 _0265_
rlabel metal2 20064 2688 20064 2688 0 _0266_
rlabel metal2 19968 3024 19968 3024 0 _0267_
rlabel metal3 19920 6300 19920 6300 0 _0268_
rlabel metal2 20304 1764 20304 1764 0 _0269_
rlabel metal2 12720 7980 12720 7980 0 _0270_
rlabel metal2 10944 8820 10944 8820 0 _0271_
rlabel metal2 9840 32676 9840 32676 0 _0272_
rlabel metal2 9600 31332 9600 31332 0 _0273_
rlabel metal3 9072 17892 9072 17892 0 _0274_
rlabel metal2 10320 11172 10320 11172 0 _0275_
rlabel metal2 11616 9030 11616 9030 0 _0276_
rlabel via1 8928 8659 8928 8659 0 _0277_
rlabel via1 9024 8659 9024 8659 0 _0278_
rlabel metal2 12768 8610 12768 8610 0 _0279_
rlabel metal2 11184 8820 11184 8820 0 _0280_
rlabel metal2 10752 12222 10752 12222 0 _0281_
rlabel metal2 7776 9954 7776 9954 0 _0282_
rlabel metal2 7968 10080 7968 10080 0 _0283_
rlabel metal3 10320 12264 10320 12264 0 _0284_
rlabel metal2 7344 8148 7344 8148 0 _0285_
rlabel metal2 7488 10206 7488 10206 0 _0286_
rlabel metal2 7872 12852 7872 12852 0 _0287_
rlabel metal3 9264 13020 9264 13020 0 _0288_
rlabel metal3 18624 4620 18624 4620 0 _0289_
rlabel metal2 19968 8106 19968 8106 0 _0290_
rlabel metal4 19968 8316 19968 8316 0 _0291_
rlabel metal2 18240 4494 18240 4494 0 _0292_
rlabel metal2 19872 8694 19872 8694 0 _0293_
rlabel metal2 19968 8946 19968 8946 0 _0294_
rlabel metal3 18576 11844 18576 11844 0 _0295_
rlabel metal3 18528 4788 18528 4788 0 _0296_
rlabel metal2 19104 12558 19104 12558 0 _0297_
rlabel metal2 19392 13188 19392 13188 0 _0298_
rlabel metal2 19584 12012 19584 12012 0 _0299_
rlabel metal4 19488 10878 19488 10878 0 _0300_
rlabel metal3 19584 8358 19584 8358 0 _0301_
rlabel metal3 19824 14028 19824 14028 0 _0302_
rlabel metal3 17760 9660 17760 9660 0 _0303_
rlabel metal2 19584 14238 19584 14238 0 _0304_
rlabel metal3 19920 13356 19920 13356 0 _0305_
rlabel metal2 19728 12684 19728 12684 0 _0306_
rlabel metal2 11184 4284 11184 4284 0 _0307_
rlabel metal2 9792 5922 9792 5922 0 _0308_
rlabel metal2 9696 6132 9696 6132 0 _0309_
rlabel metal2 6528 4242 6528 4242 0 _0310_
rlabel metal2 7392 6510 7392 6510 0 _0311_
rlabel metal2 7872 6384 7872 6384 0 _0312_
rlabel metal3 9840 4116 9840 4116 0 _0313_
rlabel metal2 10464 5208 10464 5208 0 _0314_
rlabel metal2 9504 6972 9504 6972 0 _0315_
rlabel metal2 9696 7140 9696 7140 0 _0316_
rlabel metal2 13920 3780 13920 3780 0 _0317_
rlabel metal2 13824 3486 13824 3486 0 _0318_
rlabel metal2 15696 5124 15696 5124 0 _0319_
rlabel metal2 15264 5586 15264 5586 0 _0320_
rlabel metal2 19824 1092 19824 1092 0 _0321_
rlabel metal2 19584 1092 19584 1092 0 _0322_
rlabel metal2 16992 4368 16992 4368 0 _0323_
rlabel metal2 16704 4494 16704 4494 0 _0324_
rlabel metal3 9792 29148 9792 29148 0 _0325_
rlabel metal3 13110 30660 13110 30660 0 _0326_
rlabel metal3 7728 28308 7728 28308 0 _0327_
rlabel metal3 8592 28224 8592 28224 0 _0328_
rlabel metal2 14592 30450 14592 30450 0 _0329_
rlabel metal2 10176 30114 10176 30114 0 _0330_
rlabel metal2 9648 29400 9648 29400 0 _0331_
rlabel metal2 9840 29652 9840 29652 0 _0332_
rlabel metal2 9456 28560 9456 28560 0 _0333_
rlabel metal2 9312 29652 9312 29652 0 _0334_
rlabel metal3 18576 36876 18576 36876 0 _0335_
rlabel metal3 19152 37296 19152 37296 0 _0336_
rlabel metal2 19968 36162 19968 36162 0 _0337_
rlabel metal2 19584 36918 19584 36918 0 _0338_
rlabel metal2 19488 38640 19488 38640 0 _0339_
rlabel metal2 19968 37464 19968 37464 0 _0340_
rlabel metal2 19200 37464 19200 37464 0 _0341_
rlabel metal3 19488 37380 19488 37380 0 _0342_
rlabel metal3 19296 36708 19296 36708 0 _0343_
rlabel metal2 20352 36876 20352 36876 0 _0344_
rlabel metal2 19824 28224 19824 28224 0 _0345_
rlabel metal2 19824 29820 19824 29820 0 _0346_
rlabel metal2 12384 23226 12384 23226 0 _0347_
rlabel metal2 12240 23100 12240 23100 0 _0348_
rlabel metal2 7440 28308 7440 28308 0 _0349_
rlabel metal3 9648 34524 9648 34524 0 _0350_
rlabel metal2 7680 30828 7680 30828 0 _0351_
rlabel metal2 7632 29988 7632 29988 0 _0352_
rlabel metal3 8304 29652 8304 29652 0 _0353_
rlabel metal3 4032 32844 4032 32844 0 _0354_
rlabel metal2 3456 33180 3456 33180 0 _0355_
rlabel via1 16704 38217 16704 38217 0 _0356_
rlabel metal3 16032 36708 16032 36708 0 _0357_
rlabel metal2 16320 37044 16320 37044 0 _0358_
rlabel metal2 16320 38220 16320 38220 0 _0359_
rlabel metal3 17328 38052 17328 38052 0 _0360_
rlabel metal3 17088 37254 17088 37254 0 _0361_
rlabel metal2 19104 36918 19104 36918 0 _0362_
rlabel metal2 16800 36792 16800 36792 0 _0363_
rlabel metal2 16992 36918 16992 36918 0 _0364_
rlabel metal3 15456 31332 15456 31332 0 _0365_
rlabel metal2 17664 31038 17664 31038 0 _0366_
rlabel metal3 13680 29820 13680 29820 0 _0367_
rlabel metal2 13728 30156 13728 30156 0 _0368_
rlabel metal2 14016 31332 14016 31332 0 _0369_
rlabel metal2 17664 30030 17664 30030 0 _0370_
rlabel metal2 17568 29988 17568 29988 0 _0371_
rlabel metal2 5280 24528 5280 24528 0 _0372_
rlabel metal2 4416 23730 4416 23730 0 _0373_
rlabel metal2 4320 23814 4320 23814 0 _0374_
rlabel metal3 4848 24612 4848 24612 0 _0375_
rlabel metal2 5952 24486 5952 24486 0 _0376_
rlabel metal2 5472 25116 5472 25116 0 _0377_
rlabel metal2 5712 24612 5712 24612 0 _0378_
rlabel metal2 17472 21168 17472 21168 0 _0379_
rlabel metal3 17856 22092 17856 22092 0 _0380_
rlabel metal2 19440 32760 19440 32760 0 clknet_0_UserCLK
rlabel metal3 19824 23856 19824 23856 0 clknet_1_0__leaf_UserCLK
rlabel metal2 14880 33390 14880 33390 0 clknet_1_1__leaf_UserCLK
<< properties >>
string FIXED_BBOX 0 0 21504 43008
<< end >>
