 // NumberOfConfigBits: 298
module W_TT_IF_switch_matrix
    #(
        parameter NoConfigBits=298
    )
    (
        input  N1END0,
        input  N1END1,
        input  N1END2,
        input  N1END3,
        input  N2MID0,
        input  N2MID1,
        input  N2MID2,
        input  N2MID3,
        input  N2MID4,
        input  N2MID5,
        input  N2MID6,
        input  N2MID7,
        input  N2END0,
        input  N2END1,
        input  N2END2,
        input  N2END3,
        input  N2END4,
        input  N2END5,
        input  N2END6,
        input  N2END7,
        input  N4END0,
        input  N4END1,
        input  N4END2,
        input  N4END3,
        input  W1END0,
        input  W1END1,
        input  W1END2,
        input  W1END3,
        input  W2MID0,
        input  W2MID1,
        input  W2MID2,
        input  W2MID3,
        input  W2MID4,
        input  W2MID5,
        input  W2MID6,
        input  W2MID7,
        input  W2END0,
        input  W2END1,
        input  W2END2,
        input  W2END3,
        input  W2END4,
        input  W2END5,
        input  W2END6,
        input  W2END7,
        input  WW4END0,
        input  WW4END1,
        input  WW4END2,
        input  WW4END3,
        input  WW4END4,
        input  WW4END5,
        input  WW4END6,
        input  WW4END7,
        input  WW4END8,
        input  WW4END9,
        input  WW4END10,
        input  WW4END11,
        input  WW4END12,
        input  WW4END13,
        input  WW4END14,
        input  WW4END15,
        input  W6END0,
        input  W6END1,
        input  W6END2,
        input  W6END3,
        input  W6END4,
        input  W6END5,
        input  W6END6,
        input  W6END7,
        input  W6END8,
        input  W6END9,
        input  W6END10,
        input  W6END11,
        input  S1END0,
        input  S1END1,
        input  S1END2,
        input  S1END3,
        input  S2MID0,
        input  S2MID1,
        input  S2MID2,
        input  S2MID3,
        input  S2MID4,
        input  S2MID5,
        input  S2MID6,
        input  S2MID7,
        input  S2END0,
        input  S2END1,
        input  S2END2,
        input  S2END3,
        input  S2END4,
        input  S2END5,
        input  S2END6,
        input  S2END7,
        input  S4END0,
        input  S4END1,
        input  S4END2,
        input  S4END3,
        input  UO_OUT0,
        input  UO_OUT1,
        input  UO_OUT2,
        input  UO_OUT3,
        input  UO_OUT4,
        input  UO_OUT5,
        input  UO_OUT6,
        input  UO_OUT7,
        input  UIO_OUT0,
        input  UIO_OUT1,
        input  UIO_OUT2,
        input  UIO_OUT3,
        input  UIO_OUT4,
        input  UIO_OUT5,
        input  UIO_OUT6,
        input  UIO_OUT7,
        input  UIO_OE0,
        input  UIO_OE1,
        input  UIO_OE2,
        input  UIO_OE3,
        input  UIO_OE4,
        input  UIO_OE5,
        input  UIO_OE6,
        input  UIO_OE7,
        input  J_NS4_END0,
        input  J_NS4_END1,
        input  J_NS4_END2,
        input  J_NS4_END3,
        input  J_NS4_END4,
        input  J_NS4_END5,
        input  J_NS4_END6,
        input  J_NS4_END7,
        input  J_NS4_END8,
        input  J_NS4_END9,
        input  J_NS4_END10,
        input  J_NS4_END11,
        input  J_NS4_END12,
        input  J_NS4_END13,
        input  J_NS4_END14,
        input  J_NS4_END15,
        input  J_NS2_END0,
        input  J_NS2_END1,
        input  J_NS2_END2,
        input  J_NS2_END3,
        input  J_NS2_END4,
        input  J_NS2_END5,
        input  J_NS2_END6,
        input  J_NS2_END7,
        input  J_NS1_END0,
        input  J_NS1_END1,
        input  J_NS1_END2,
        input  J_NS1_END3,
        output  N1BEG0,
        output  N1BEG1,
        output  N1BEG2,
        output  N1BEG3,
        output  N2BEG0,
        output  N2BEG1,
        output  N2BEG2,
        output  N2BEG3,
        output  N2BEG4,
        output  N2BEG5,
        output  N2BEG6,
        output  N2BEG7,
        output  N2BEGb0,
        output  N2BEGb1,
        output  N2BEGb2,
        output  N2BEGb3,
        output  N2BEGb4,
        output  N2BEGb5,
        output  N2BEGb6,
        output  N2BEGb7,
        output  N4BEG0,
        output  N4BEG1,
        output  N4BEG2,
        output  N4BEG3,
        output  S1BEG0,
        output  S1BEG1,
        output  S1BEG2,
        output  S1BEG3,
        output  S2BEG0,
        output  S2BEG1,
        output  S2BEG2,
        output  S2BEG3,
        output  S2BEG4,
        output  S2BEG5,
        output  S2BEG6,
        output  S2BEG7,
        output  S2BEGb0,
        output  S2BEGb1,
        output  S2BEGb2,
        output  S2BEGb3,
        output  S2BEGb4,
        output  S2BEGb5,
        output  S2BEGb6,
        output  S2BEGb7,
        output  S4BEG0,
        output  S4BEG1,
        output  S4BEG2,
        output  S4BEG3,
        output  E1BEG0,
        output  E1BEG1,
        output  E1BEG2,
        output  E1BEG3,
        output  E2BEG0,
        output  E2BEG1,
        output  E2BEG2,
        output  E2BEG3,
        output  E2BEG4,
        output  E2BEG5,
        output  E2BEG6,
        output  E2BEG7,
        output  E2BEGb0,
        output  E2BEGb1,
        output  E2BEGb2,
        output  E2BEGb3,
        output  E2BEGb4,
        output  E2BEGb5,
        output  E2BEGb6,
        output  E2BEGb7,
        output  EE4BEG0,
        output  EE4BEG1,
        output  EE4BEG2,
        output  EE4BEG3,
        output  EE4BEG4,
        output  EE4BEG5,
        output  EE4BEG6,
        output  EE4BEG7,
        output  EE4BEG8,
        output  EE4BEG9,
        output  EE4BEG10,
        output  EE4BEG11,
        output  EE4BEG12,
        output  EE4BEG13,
        output  EE4BEG14,
        output  EE4BEG15,
        output  E6BEG0,
        output  E6BEG1,
        output  E6BEG2,
        output  E6BEG3,
        output  E6BEG4,
        output  E6BEG5,
        output  E6BEG6,
        output  E6BEG7,
        output  E6BEG8,
        output  E6BEG9,
        output  E6BEG10,
        output  E6BEG11,
        output  UI_IN0,
        output  UI_IN1,
        output  UI_IN2,
        output  UI_IN3,
        output  UI_IN4,
        output  UI_IN5,
        output  UI_IN6,
        output  UI_IN7,
        output  UIO_IN0,
        output  UIO_IN1,
        output  UIO_IN2,
        output  UIO_IN3,
        output  UIO_IN4,
        output  UIO_IN5,
        output  UIO_IN6,
        output  UIO_IN7,
        output  ENA,
        output  RST_N,
        output  J_NS4_BEG0,
        output  J_NS4_BEG1,
        output  J_NS4_BEG2,
        output  J_NS4_BEG3,
        output  J_NS4_BEG4,
        output  J_NS4_BEG5,
        output  J_NS4_BEG6,
        output  J_NS4_BEG7,
        output  J_NS4_BEG8,
        output  J_NS4_BEG9,
        output  J_NS4_BEG10,
        output  J_NS4_BEG11,
        output  J_NS4_BEG12,
        output  J_NS4_BEG13,
        output  J_NS4_BEG14,
        output  J_NS4_BEG15,
        output  J_NS2_BEG0,
        output  J_NS2_BEG1,
        output  J_NS2_BEG2,
        output  J_NS2_BEG3,
        output  J_NS2_BEG4,
        output  J_NS2_BEG5,
        output  J_NS2_BEG6,
        output  J_NS2_BEG7,
        output  J_NS1_BEG0,
        output  J_NS1_BEG1,
        output  J_NS1_BEG2,
        output  J_NS1_BEG3,
 //global
        input  [NoConfigBits-1:0] ConfigBits,
        input  [NoConfigBits-1:0] ConfigBits_N
);
parameter GND0 = 1'b0;
parameter GND = 1'b0;
parameter VCC0 = 1'b1;
parameter VCC = 1'b1;
parameter VDD0 = 1'b1;
parameter VDD = 1'b1;

wire[4-1:0] N1BEG0_input;
wire[4-1:0] N1BEG1_input;
wire[4-1:0] N1BEG2_input;
wire[4-1:0] N1BEG3_input;
wire[4-1:0] N2BEG0_input;
wire[4-1:0] N2BEG1_input;
wire[4-1:0] N2BEG2_input;
wire[4-1:0] N2BEG3_input;
wire[4-1:0] N2BEG4_input;
wire[4-1:0] N2BEG5_input;
wire[4-1:0] N2BEG6_input;
wire[4-1:0] N2BEG7_input;
wire[8-1:0] N4BEG0_input;
wire[8-1:0] N4BEG1_input;
wire[8-1:0] N4BEG2_input;
wire[8-1:0] N4BEG3_input;
wire[4-1:0] S1BEG0_input;
wire[4-1:0] S1BEG1_input;
wire[4-1:0] S1BEG2_input;
wire[4-1:0] S1BEG3_input;
wire[4-1:0] S2BEG0_input;
wire[4-1:0] S2BEG1_input;
wire[4-1:0] S2BEG2_input;
wire[4-1:0] S2BEG3_input;
wire[4-1:0] S2BEG4_input;
wire[4-1:0] S2BEG5_input;
wire[4-1:0] S2BEG6_input;
wire[4-1:0] S2BEG7_input;
wire[8-1:0] S4BEG0_input;
wire[8-1:0] S4BEG1_input;
wire[8-1:0] S4BEG2_input;
wire[8-1:0] S4BEG3_input;
wire[8-1:0] E1BEG0_input;
wire[8-1:0] E1BEG1_input;
wire[8-1:0] E1BEG2_input;
wire[8-1:0] E1BEG3_input;
wire[8-1:0] E2BEG0_input;
wire[8-1:0] E2BEG1_input;
wire[8-1:0] E2BEG2_input;
wire[8-1:0] E2BEG3_input;
wire[8-1:0] E2BEG4_input;
wire[8-1:0] E2BEG5_input;
wire[8-1:0] E2BEG6_input;
wire[8-1:0] E2BEG7_input;
wire[8-1:0] E2BEGb0_input;
wire[8-1:0] E2BEGb1_input;
wire[8-1:0] E2BEGb2_input;
wire[8-1:0] E2BEGb3_input;
wire[8-1:0] E2BEGb4_input;
wire[8-1:0] E2BEGb5_input;
wire[8-1:0] E2BEGb6_input;
wire[8-1:0] E2BEGb7_input;
wire[4-1:0] EE4BEG0_input;
wire[4-1:0] EE4BEG1_input;
wire[4-1:0] EE4BEG2_input;
wire[4-1:0] EE4BEG3_input;
wire[4-1:0] EE4BEG4_input;
wire[4-1:0] EE4BEG5_input;
wire[4-1:0] EE4BEG6_input;
wire[4-1:0] EE4BEG7_input;
wire[4-1:0] EE4BEG8_input;
wire[4-1:0] EE4BEG9_input;
wire[4-1:0] EE4BEG10_input;
wire[4-1:0] EE4BEG11_input;
wire[4-1:0] EE4BEG12_input;
wire[4-1:0] EE4BEG13_input;
wire[4-1:0] EE4BEG14_input;
wire[4-1:0] EE4BEG15_input;
wire[4-1:0] E6BEG0_input;
wire[4-1:0] E6BEG1_input;
wire[4-1:0] E6BEG2_input;
wire[4-1:0] E6BEG3_input;
wire[4-1:0] E6BEG4_input;
wire[4-1:0] E6BEG5_input;
wire[4-1:0] E6BEG6_input;
wire[4-1:0] E6BEG7_input;
wire[4-1:0] E6BEG8_input;
wire[4-1:0] E6BEG9_input;
wire[4-1:0] E6BEG10_input;
wire[4-1:0] E6BEG11_input;
wire[8-1:0] UI_IN0_input;
wire[8-1:0] UI_IN1_input;
wire[8-1:0] UI_IN2_input;
wire[8-1:0] UI_IN3_input;
wire[8-1:0] UI_IN4_input;
wire[8-1:0] UI_IN5_input;
wire[8-1:0] UI_IN6_input;
wire[8-1:0] UI_IN7_input;
wire[8-1:0] UIO_IN0_input;
wire[8-1:0] UIO_IN1_input;
wire[8-1:0] UIO_IN2_input;
wire[8-1:0] UIO_IN3_input;
wire[8-1:0] UIO_IN4_input;
wire[8-1:0] UIO_IN5_input;
wire[8-1:0] UIO_IN6_input;
wire[8-1:0] UIO_IN7_input;
wire[4-1:0] ENA_input;
wire[16-1:0] RST_N_input;
wire[4-1:0] J_NS4_BEG0_input;
wire[4-1:0] J_NS4_BEG1_input;
wire[4-1:0] J_NS4_BEG2_input;
wire[4-1:0] J_NS4_BEG3_input;
wire[4-1:0] J_NS4_BEG4_input;
wire[4-1:0] J_NS4_BEG5_input;
wire[4-1:0] J_NS4_BEG6_input;
wire[4-1:0] J_NS4_BEG7_input;
wire[4-1:0] J_NS4_BEG8_input;
wire[4-1:0] J_NS4_BEG9_input;
wire[4-1:0] J_NS4_BEG10_input;
wire[4-1:0] J_NS4_BEG11_input;
wire[4-1:0] J_NS4_BEG12_input;
wire[4-1:0] J_NS4_BEG13_input;
wire[4-1:0] J_NS4_BEG14_input;
wire[4-1:0] J_NS4_BEG15_input;
wire[4-1:0] J_NS2_BEG0_input;
wire[4-1:0] J_NS2_BEG1_input;
wire[4-1:0] J_NS2_BEG2_input;
wire[4-1:0] J_NS2_BEG3_input;
wire[4-1:0] J_NS2_BEG4_input;
wire[4-1:0] J_NS2_BEG5_input;
wire[4-1:0] J_NS2_BEG6_input;
wire[4-1:0] J_NS2_BEG7_input;
wire[4-1:0] J_NS1_BEG0_input;
wire[4-1:0] J_NS1_BEG1_input;
wire[4-1:0] J_NS1_BEG2_input;
wire[4-1:0] J_NS1_BEG3_input;
 //The configuration bits (if any) are just a long shift register
 //This shift register is padded to an even number of flops/latches
 //switch matrix multiplexer N1BEG0 MUX-4
assign N1BEG0_input = {J_NS1_END0,J_NS4_END12,W6END4,W1END0};
cus_mux41_buf inst_cus_mux41_buf_N1BEG0 (
    .A0(N1BEG0_input[0]),
    .A1(N1BEG0_input[1]),
    .A2(N1BEG0_input[2]),
    .A3(N1BEG0_input[3]),
    .S0(ConfigBits[0+0]),
    .S0N(ConfigBits_N[0+0]),
    .S1(ConfigBits[0+1]),
    .S1N(ConfigBits_N[0+1]),
    .X(N1BEG0)
);

 //switch matrix multiplexer N1BEG1 MUX-4
assign N1BEG1_input = {J_NS1_END1,J_NS4_END13,W6END5,W1END1};
cus_mux41_buf inst_cus_mux41_buf_N1BEG1 (
    .A0(N1BEG1_input[0]),
    .A1(N1BEG1_input[1]),
    .A2(N1BEG1_input[2]),
    .A3(N1BEG1_input[3]),
    .S0(ConfigBits[2+0]),
    .S0N(ConfigBits_N[2+0]),
    .S1(ConfigBits[2+1]),
    .S1N(ConfigBits_N[2+1]),
    .X(N1BEG1)
);

 //switch matrix multiplexer N1BEG2 MUX-4
assign N1BEG2_input = {J_NS1_END2,J_NS4_END14,W6END6,W1END2};
cus_mux41_buf inst_cus_mux41_buf_N1BEG2 (
    .A0(N1BEG2_input[0]),
    .A1(N1BEG2_input[1]),
    .A2(N1BEG2_input[2]),
    .A3(N1BEG2_input[3]),
    .S0(ConfigBits[4+0]),
    .S0N(ConfigBits_N[4+0]),
    .S1(ConfigBits[4+1]),
    .S1N(ConfigBits_N[4+1]),
    .X(N1BEG2)
);

 //switch matrix multiplexer N1BEG3 MUX-4
assign N1BEG3_input = {J_NS1_END3,J_NS4_END15,W6END7,W1END3};
cus_mux41_buf inst_cus_mux41_buf_N1BEG3 (
    .A0(N1BEG3_input[0]),
    .A1(N1BEG3_input[1]),
    .A2(N1BEG3_input[2]),
    .A3(N1BEG3_input[3]),
    .S0(ConfigBits[6+0]),
    .S0N(ConfigBits_N[6+0]),
    .S1(ConfigBits[6+1]),
    .S1N(ConfigBits_N[6+1]),
    .X(N1BEG3)
);

 //switch matrix multiplexer N2BEG0 MUX-4
assign N2BEG0_input = {J_NS2_END0,W6END7,W2END7,W2MID7};
cus_mux41_buf inst_cus_mux41_buf_N2BEG0 (
    .A0(N2BEG0_input[0]),
    .A1(N2BEG0_input[1]),
    .A2(N2BEG0_input[2]),
    .A3(N2BEG0_input[3]),
    .S0(ConfigBits[8+0]),
    .S0N(ConfigBits_N[8+0]),
    .S1(ConfigBits[8+1]),
    .S1N(ConfigBits_N[8+1]),
    .X(N2BEG0)
);

 //switch matrix multiplexer N2BEG1 MUX-4
assign N2BEG1_input = {J_NS2_END1,W6END6,W2END6,W2MID6};
cus_mux41_buf inst_cus_mux41_buf_N2BEG1 (
    .A0(N2BEG1_input[0]),
    .A1(N2BEG1_input[1]),
    .A2(N2BEG1_input[2]),
    .A3(N2BEG1_input[3]),
    .S0(ConfigBits[10+0]),
    .S0N(ConfigBits_N[10+0]),
    .S1(ConfigBits[10+1]),
    .S1N(ConfigBits_N[10+1]),
    .X(N2BEG1)
);

 //switch matrix multiplexer N2BEG2 MUX-4
assign N2BEG2_input = {J_NS2_END2,W6END5,W2END5,W2MID5};
cus_mux41_buf inst_cus_mux41_buf_N2BEG2 (
    .A0(N2BEG2_input[0]),
    .A1(N2BEG2_input[1]),
    .A2(N2BEG2_input[2]),
    .A3(N2BEG2_input[3]),
    .S0(ConfigBits[12+0]),
    .S0N(ConfigBits_N[12+0]),
    .S1(ConfigBits[12+1]),
    .S1N(ConfigBits_N[12+1]),
    .X(N2BEG2)
);

 //switch matrix multiplexer N2BEG3 MUX-4
assign N2BEG3_input = {J_NS2_END3,W6END4,W2END4,W2MID4};
cus_mux41_buf inst_cus_mux41_buf_N2BEG3 (
    .A0(N2BEG3_input[0]),
    .A1(N2BEG3_input[1]),
    .A2(N2BEG3_input[2]),
    .A3(N2BEG3_input[3]),
    .S0(ConfigBits[14+0]),
    .S0N(ConfigBits_N[14+0]),
    .S1(ConfigBits[14+1]),
    .S1N(ConfigBits_N[14+1]),
    .X(N2BEG3)
);

 //switch matrix multiplexer N2BEG4 MUX-4
assign N2BEG4_input = {J_NS2_END4,W6END3,W2END3,W2MID3};
cus_mux41_buf inst_cus_mux41_buf_N2BEG4 (
    .A0(N2BEG4_input[0]),
    .A1(N2BEG4_input[1]),
    .A2(N2BEG4_input[2]),
    .A3(N2BEG4_input[3]),
    .S0(ConfigBits[16+0]),
    .S0N(ConfigBits_N[16+0]),
    .S1(ConfigBits[16+1]),
    .S1N(ConfigBits_N[16+1]),
    .X(N2BEG4)
);

 //switch matrix multiplexer N2BEG5 MUX-4
assign N2BEG5_input = {J_NS2_END5,W6END2,W2END2,W2MID2};
cus_mux41_buf inst_cus_mux41_buf_N2BEG5 (
    .A0(N2BEG5_input[0]),
    .A1(N2BEG5_input[1]),
    .A2(N2BEG5_input[2]),
    .A3(N2BEG5_input[3]),
    .S0(ConfigBits[18+0]),
    .S0N(ConfigBits_N[18+0]),
    .S1(ConfigBits[18+1]),
    .S1N(ConfigBits_N[18+1]),
    .X(N2BEG5)
);

 //switch matrix multiplexer N2BEG6 MUX-4
assign N2BEG6_input = {J_NS2_END6,W6END1,W2END1,W2MID1};
cus_mux41_buf inst_cus_mux41_buf_N2BEG6 (
    .A0(N2BEG6_input[0]),
    .A1(N2BEG6_input[1]),
    .A2(N2BEG6_input[2]),
    .A3(N2BEG6_input[3]),
    .S0(ConfigBits[20+0]),
    .S0N(ConfigBits_N[20+0]),
    .S1(ConfigBits[20+1]),
    .S1N(ConfigBits_N[20+1]),
    .X(N2BEG6)
);

 //switch matrix multiplexer N2BEG7 MUX-4
assign N2BEG7_input = {J_NS2_END7,W6END0,W2END0,W2MID0};
cus_mux41_buf inst_cus_mux41_buf_N2BEG7 (
    .A0(N2BEG7_input[0]),
    .A1(N2BEG7_input[1]),
    .A2(N2BEG7_input[2]),
    .A3(N2BEG7_input[3]),
    .S0(ConfigBits[22+0]),
    .S0N(ConfigBits_N[22+0]),
    .S1(ConfigBits[22+1]),
    .S1N(ConfigBits_N[22+1]),
    .X(N2BEG7)
);

 //switch matrix multiplexer N2BEGb0 MUX-1
assign N2BEGb0 = N2MID0;

 //switch matrix multiplexer N2BEGb1 MUX-1
assign N2BEGb1 = N2MID1;

 //switch matrix multiplexer N2BEGb2 MUX-1
assign N2BEGb2 = N2MID2;

 //switch matrix multiplexer N2BEGb3 MUX-1
assign N2BEGb3 = N2MID3;

 //switch matrix multiplexer N2BEGb4 MUX-1
assign N2BEGb4 = N2MID4;

 //switch matrix multiplexer N2BEGb5 MUX-1
assign N2BEGb5 = N2MID5;

 //switch matrix multiplexer N2BEGb6 MUX-1
assign N2BEGb6 = N2MID6;

 //switch matrix multiplexer N2BEGb7 MUX-1
assign N2BEGb7 = N2MID7;

 //switch matrix multiplexer N4BEG0 MUX-8
assign N4BEG0_input = {J_NS2_END0,J_NS4_END12,J_NS4_END8,J_NS4_END4,J_NS4_END0,W6END8,WW4END0,W1END0};
cus_mux81_buf inst_cus_mux81_buf_N4BEG0 (
    .A0(N4BEG0_input[0]),
    .A1(N4BEG0_input[1]),
    .A2(N4BEG0_input[2]),
    .A3(N4BEG0_input[3]),
    .A4(N4BEG0_input[4]),
    .A5(N4BEG0_input[5]),
    .A6(N4BEG0_input[6]),
    .A7(N4BEG0_input[7]),
    .S0(ConfigBits[24+0]),
    .S0N(ConfigBits_N[24+0]),
    .S1(ConfigBits[24+1]),
    .S1N(ConfigBits_N[24+1]),
    .S2(ConfigBits[24+2]),
    .S2N(ConfigBits_N[24+2]),
    .X(N4BEG0)
);

 //switch matrix multiplexer N4BEG1 MUX-8
assign N4BEG1_input = {J_NS2_END1,J_NS4_END13,J_NS4_END9,J_NS4_END5,J_NS4_END1,W6END9,WW4END1,W1END1};
cus_mux81_buf inst_cus_mux81_buf_N4BEG1 (
    .A0(N4BEG1_input[0]),
    .A1(N4BEG1_input[1]),
    .A2(N4BEG1_input[2]),
    .A3(N4BEG1_input[3]),
    .A4(N4BEG1_input[4]),
    .A5(N4BEG1_input[5]),
    .A6(N4BEG1_input[6]),
    .A7(N4BEG1_input[7]),
    .S0(ConfigBits[27+0]),
    .S0N(ConfigBits_N[27+0]),
    .S1(ConfigBits[27+1]),
    .S1N(ConfigBits_N[27+1]),
    .S2(ConfigBits[27+2]),
    .S2N(ConfigBits_N[27+2]),
    .X(N4BEG1)
);

 //switch matrix multiplexer N4BEG2 MUX-8
assign N4BEG2_input = {J_NS2_END2,J_NS4_END14,J_NS4_END10,J_NS4_END6,J_NS4_END2,W6END10,WW4END2,W1END2};
cus_mux81_buf inst_cus_mux81_buf_N4BEG2 (
    .A0(N4BEG2_input[0]),
    .A1(N4BEG2_input[1]),
    .A2(N4BEG2_input[2]),
    .A3(N4BEG2_input[3]),
    .A4(N4BEG2_input[4]),
    .A5(N4BEG2_input[5]),
    .A6(N4BEG2_input[6]),
    .A7(N4BEG2_input[7]),
    .S0(ConfigBits[30+0]),
    .S0N(ConfigBits_N[30+0]),
    .S1(ConfigBits[30+1]),
    .S1N(ConfigBits_N[30+1]),
    .S2(ConfigBits[30+2]),
    .S2N(ConfigBits_N[30+2]),
    .X(N4BEG2)
);

 //switch matrix multiplexer N4BEG3 MUX-8
assign N4BEG3_input = {J_NS2_END3,J_NS4_END15,J_NS4_END11,J_NS4_END7,J_NS4_END3,W6END11,WW4END3,W1END3};
cus_mux81_buf inst_cus_mux81_buf_N4BEG3 (
    .A0(N4BEG3_input[0]),
    .A1(N4BEG3_input[1]),
    .A2(N4BEG3_input[2]),
    .A3(N4BEG3_input[3]),
    .A4(N4BEG3_input[4]),
    .A5(N4BEG3_input[5]),
    .A6(N4BEG3_input[6]),
    .A7(N4BEG3_input[7]),
    .S0(ConfigBits[33+0]),
    .S0N(ConfigBits_N[33+0]),
    .S1(ConfigBits[33+1]),
    .S1N(ConfigBits_N[33+1]),
    .S2(ConfigBits[33+2]),
    .S2N(ConfigBits_N[33+2]),
    .X(N4BEG3)
);

 //switch matrix multiplexer S1BEG0 MUX-4
assign S1BEG0_input = {J_NS1_END0,J_NS4_END12,W6END8,W1END0};
cus_mux41_buf inst_cus_mux41_buf_S1BEG0 (
    .A0(S1BEG0_input[0]),
    .A1(S1BEG0_input[1]),
    .A2(S1BEG0_input[2]),
    .A3(S1BEG0_input[3]),
    .S0(ConfigBits[36+0]),
    .S0N(ConfigBits_N[36+0]),
    .S1(ConfigBits[36+1]),
    .S1N(ConfigBits_N[36+1]),
    .X(S1BEG0)
);

 //switch matrix multiplexer S1BEG1 MUX-4
assign S1BEG1_input = {J_NS1_END1,J_NS4_END13,W6END9,W1END1};
cus_mux41_buf inst_cus_mux41_buf_S1BEG1 (
    .A0(S1BEG1_input[0]),
    .A1(S1BEG1_input[1]),
    .A2(S1BEG1_input[2]),
    .A3(S1BEG1_input[3]),
    .S0(ConfigBits[38+0]),
    .S0N(ConfigBits_N[38+0]),
    .S1(ConfigBits[38+1]),
    .S1N(ConfigBits_N[38+1]),
    .X(S1BEG1)
);

 //switch matrix multiplexer S1BEG2 MUX-4
assign S1BEG2_input = {J_NS1_END2,J_NS4_END14,W6END10,W1END2};
cus_mux41_buf inst_cus_mux41_buf_S1BEG2 (
    .A0(S1BEG2_input[0]),
    .A1(S1BEG2_input[1]),
    .A2(S1BEG2_input[2]),
    .A3(S1BEG2_input[3]),
    .S0(ConfigBits[40+0]),
    .S0N(ConfigBits_N[40+0]),
    .S1(ConfigBits[40+1]),
    .S1N(ConfigBits_N[40+1]),
    .X(S1BEG2)
);

 //switch matrix multiplexer S1BEG3 MUX-4
assign S1BEG3_input = {J_NS1_END3,J_NS4_END15,W6END11,W1END3};
cus_mux41_buf inst_cus_mux41_buf_S1BEG3 (
    .A0(S1BEG3_input[0]),
    .A1(S1BEG3_input[1]),
    .A2(S1BEG3_input[2]),
    .A3(S1BEG3_input[3]),
    .S0(ConfigBits[42+0]),
    .S0N(ConfigBits_N[42+0]),
    .S1(ConfigBits[42+1]),
    .S1N(ConfigBits_N[42+1]),
    .X(S1BEG3)
);

 //switch matrix multiplexer S2BEG0 MUX-4
assign S2BEG0_input = {J_NS2_END0,W6END8,W2END7,W2MID7};
cus_mux41_buf inst_cus_mux41_buf_S2BEG0 (
    .A0(S2BEG0_input[0]),
    .A1(S2BEG0_input[1]),
    .A2(S2BEG0_input[2]),
    .A3(S2BEG0_input[3]),
    .S0(ConfigBits[44+0]),
    .S0N(ConfigBits_N[44+0]),
    .S1(ConfigBits[44+1]),
    .S1N(ConfigBits_N[44+1]),
    .X(S2BEG0)
);

 //switch matrix multiplexer S2BEG1 MUX-4
assign S2BEG1_input = {J_NS2_END1,W6END9,W2END6,W2MID6};
cus_mux41_buf inst_cus_mux41_buf_S2BEG1 (
    .A0(S2BEG1_input[0]),
    .A1(S2BEG1_input[1]),
    .A2(S2BEG1_input[2]),
    .A3(S2BEG1_input[3]),
    .S0(ConfigBits[46+0]),
    .S0N(ConfigBits_N[46+0]),
    .S1(ConfigBits[46+1]),
    .S1N(ConfigBits_N[46+1]),
    .X(S2BEG1)
);

 //switch matrix multiplexer S2BEG2 MUX-4
assign S2BEG2_input = {J_NS2_END2,W6END10,W2END5,W2MID5};
cus_mux41_buf inst_cus_mux41_buf_S2BEG2 (
    .A0(S2BEG2_input[0]),
    .A1(S2BEG2_input[1]),
    .A2(S2BEG2_input[2]),
    .A3(S2BEG2_input[3]),
    .S0(ConfigBits[48+0]),
    .S0N(ConfigBits_N[48+0]),
    .S1(ConfigBits[48+1]),
    .S1N(ConfigBits_N[48+1]),
    .X(S2BEG2)
);

 //switch matrix multiplexer S2BEG3 MUX-4
assign S2BEG3_input = {J_NS2_END3,W6END11,W2END4,W2MID4};
cus_mux41_buf inst_cus_mux41_buf_S2BEG3 (
    .A0(S2BEG3_input[0]),
    .A1(S2BEG3_input[1]),
    .A2(S2BEG3_input[2]),
    .A3(S2BEG3_input[3]),
    .S0(ConfigBits[50+0]),
    .S0N(ConfigBits_N[50+0]),
    .S1(ConfigBits[50+1]),
    .S1N(ConfigBits_N[50+1]),
    .X(S2BEG3)
);

 //switch matrix multiplexer S2BEG4 MUX-4
assign S2BEG4_input = {J_NS2_END4,W2END3,W2MID3,W1END0};
cus_mux41_buf inst_cus_mux41_buf_S2BEG4 (
    .A0(S2BEG4_input[0]),
    .A1(S2BEG4_input[1]),
    .A2(S2BEG4_input[2]),
    .A3(S2BEG4_input[3]),
    .S0(ConfigBits[52+0]),
    .S0N(ConfigBits_N[52+0]),
    .S1(ConfigBits[52+1]),
    .S1N(ConfigBits_N[52+1]),
    .X(S2BEG4)
);

 //switch matrix multiplexer S2BEG5 MUX-4
assign S2BEG5_input = {J_NS2_END5,W2END2,W2MID2,W1END1};
cus_mux41_buf inst_cus_mux41_buf_S2BEG5 (
    .A0(S2BEG5_input[0]),
    .A1(S2BEG5_input[1]),
    .A2(S2BEG5_input[2]),
    .A3(S2BEG5_input[3]),
    .S0(ConfigBits[54+0]),
    .S0N(ConfigBits_N[54+0]),
    .S1(ConfigBits[54+1]),
    .S1N(ConfigBits_N[54+1]),
    .X(S2BEG5)
);

 //switch matrix multiplexer S2BEG6 MUX-4
assign S2BEG6_input = {J_NS2_END6,W2END1,W2MID1,W1END2};
cus_mux41_buf inst_cus_mux41_buf_S2BEG6 (
    .A0(S2BEG6_input[0]),
    .A1(S2BEG6_input[1]),
    .A2(S2BEG6_input[2]),
    .A3(S2BEG6_input[3]),
    .S0(ConfigBits[56+0]),
    .S0N(ConfigBits_N[56+0]),
    .S1(ConfigBits[56+1]),
    .S1N(ConfigBits_N[56+1]),
    .X(S2BEG6)
);

 //switch matrix multiplexer S2BEG7 MUX-4
assign S2BEG7_input = {J_NS2_END7,W2END0,W2MID0,W1END3};
cus_mux41_buf inst_cus_mux41_buf_S2BEG7 (
    .A0(S2BEG7_input[0]),
    .A1(S2BEG7_input[1]),
    .A2(S2BEG7_input[2]),
    .A3(S2BEG7_input[3]),
    .S0(ConfigBits[58+0]),
    .S0N(ConfigBits_N[58+0]),
    .S1(ConfigBits[58+1]),
    .S1N(ConfigBits_N[58+1]),
    .X(S2BEG7)
);

 //switch matrix multiplexer S2BEGb0 MUX-1
assign S2BEGb0 = S2MID0;

 //switch matrix multiplexer S2BEGb1 MUX-1
assign S2BEGb1 = S2MID1;

 //switch matrix multiplexer S2BEGb2 MUX-1
assign S2BEGb2 = S2MID2;

 //switch matrix multiplexer S2BEGb3 MUX-1
assign S2BEGb3 = S2MID3;

 //switch matrix multiplexer S2BEGb4 MUX-1
assign S2BEGb4 = S2MID4;

 //switch matrix multiplexer S2BEGb5 MUX-1
assign S2BEGb5 = S2MID5;

 //switch matrix multiplexer S2BEGb6 MUX-1
assign S2BEGb6 = S2MID6;

 //switch matrix multiplexer S2BEGb7 MUX-1
assign S2BEGb7 = S2MID7;

 //switch matrix multiplexer S4BEG0 MUX-8
assign S4BEG0_input = {J_NS2_END4,J_NS4_END12,J_NS4_END8,J_NS4_END4,J_NS4_END0,W6END4,WW4END12,W1END0};
cus_mux81_buf inst_cus_mux81_buf_S4BEG0 (
    .A0(S4BEG0_input[0]),
    .A1(S4BEG0_input[1]),
    .A2(S4BEG0_input[2]),
    .A3(S4BEG0_input[3]),
    .A4(S4BEG0_input[4]),
    .A5(S4BEG0_input[5]),
    .A6(S4BEG0_input[6]),
    .A7(S4BEG0_input[7]),
    .S0(ConfigBits[60+0]),
    .S0N(ConfigBits_N[60+0]),
    .S1(ConfigBits[60+1]),
    .S1N(ConfigBits_N[60+1]),
    .S2(ConfigBits[60+2]),
    .S2N(ConfigBits_N[60+2]),
    .X(S4BEG0)
);

 //switch matrix multiplexer S4BEG1 MUX-8
assign S4BEG1_input = {J_NS2_END5,J_NS4_END13,J_NS4_END9,J_NS4_END5,J_NS4_END1,W6END5,WW4END13,W1END1};
cus_mux81_buf inst_cus_mux81_buf_S4BEG1 (
    .A0(S4BEG1_input[0]),
    .A1(S4BEG1_input[1]),
    .A2(S4BEG1_input[2]),
    .A3(S4BEG1_input[3]),
    .A4(S4BEG1_input[4]),
    .A5(S4BEG1_input[5]),
    .A6(S4BEG1_input[6]),
    .A7(S4BEG1_input[7]),
    .S0(ConfigBits[63+0]),
    .S0N(ConfigBits_N[63+0]),
    .S1(ConfigBits[63+1]),
    .S1N(ConfigBits_N[63+1]),
    .S2(ConfigBits[63+2]),
    .S2N(ConfigBits_N[63+2]),
    .X(S4BEG1)
);

 //switch matrix multiplexer S4BEG2 MUX-8
assign S4BEG2_input = {J_NS2_END6,J_NS4_END14,J_NS4_END10,J_NS4_END6,J_NS4_END2,W6END6,WW4END14,W1END2};
cus_mux81_buf inst_cus_mux81_buf_S4BEG2 (
    .A0(S4BEG2_input[0]),
    .A1(S4BEG2_input[1]),
    .A2(S4BEG2_input[2]),
    .A3(S4BEG2_input[3]),
    .A4(S4BEG2_input[4]),
    .A5(S4BEG2_input[5]),
    .A6(S4BEG2_input[6]),
    .A7(S4BEG2_input[7]),
    .S0(ConfigBits[66+0]),
    .S0N(ConfigBits_N[66+0]),
    .S1(ConfigBits[66+1]),
    .S1N(ConfigBits_N[66+1]),
    .S2(ConfigBits[66+2]),
    .S2N(ConfigBits_N[66+2]),
    .X(S4BEG2)
);

 //switch matrix multiplexer S4BEG3 MUX-8
assign S4BEG3_input = {J_NS2_END7,J_NS4_END15,J_NS4_END11,J_NS4_END7,J_NS4_END3,W6END7,WW4END15,W1END3};
cus_mux81_buf inst_cus_mux81_buf_S4BEG3 (
    .A0(S4BEG3_input[0]),
    .A1(S4BEG3_input[1]),
    .A2(S4BEG3_input[2]),
    .A3(S4BEG3_input[3]),
    .A4(S4BEG3_input[4]),
    .A5(S4BEG3_input[5]),
    .A6(S4BEG3_input[6]),
    .A7(S4BEG3_input[7]),
    .S0(ConfigBits[69+0]),
    .S0N(ConfigBits_N[69+0]),
    .S1(ConfigBits[69+1]),
    .S1N(ConfigBits_N[69+1]),
    .S2(ConfigBits[69+2]),
    .S2N(ConfigBits_N[69+2]),
    .X(S4BEG3)
);

 //switch matrix multiplexer E1BEG0 MUX-8
assign E1BEG0_input = {UIO_OE7,UIO_OE6,UIO_OE2,UIO_OE0,UO_OUT7,UO_OUT2,S1END0,N1END0};
cus_mux81_buf inst_cus_mux81_buf_E1BEG0 (
    .A0(E1BEG0_input[0]),
    .A1(E1BEG0_input[1]),
    .A2(E1BEG0_input[2]),
    .A3(E1BEG0_input[3]),
    .A4(E1BEG0_input[4]),
    .A5(E1BEG0_input[5]),
    .A6(E1BEG0_input[6]),
    .A7(E1BEG0_input[7]),
    .S0(ConfigBits[72+0]),
    .S0N(ConfigBits_N[72+0]),
    .S1(ConfigBits[72+1]),
    .S1N(ConfigBits_N[72+1]),
    .S2(ConfigBits[72+2]),
    .S2N(ConfigBits_N[72+2]),
    .X(E1BEG0)
);

 //switch matrix multiplexer E1BEG1 MUX-8
assign E1BEG1_input = {UIO_OE6,UIO_OE5,UIO_OE1,UIO_OE0,UO_OUT6,UO_OUT3,S1END1,N1END1};
cus_mux81_buf inst_cus_mux81_buf_E1BEG1 (
    .A0(E1BEG1_input[0]),
    .A1(E1BEG1_input[1]),
    .A2(E1BEG1_input[2]),
    .A3(E1BEG1_input[3]),
    .A4(E1BEG1_input[4]),
    .A5(E1BEG1_input[5]),
    .A6(E1BEG1_input[6]),
    .A7(E1BEG1_input[7]),
    .S0(ConfigBits[75+0]),
    .S0N(ConfigBits_N[75+0]),
    .S1(ConfigBits[75+1]),
    .S1N(ConfigBits_N[75+1]),
    .S2(ConfigBits[75+2]),
    .S2N(ConfigBits_N[75+2]),
    .X(E1BEG1)
);

 //switch matrix multiplexer E1BEG2 MUX-8
assign E1BEG2_input = {UIO_OE5,UIO_OE4,UIO_OE3,UIO_OE2,UO_OUT5,UO_OUT0,S1END2,N1END2};
cus_mux81_buf inst_cus_mux81_buf_E1BEG2 (
    .A0(E1BEG2_input[0]),
    .A1(E1BEG2_input[1]),
    .A2(E1BEG2_input[2]),
    .A3(E1BEG2_input[3]),
    .A4(E1BEG2_input[4]),
    .A5(E1BEG2_input[5]),
    .A6(E1BEG2_input[6]),
    .A7(E1BEG2_input[7]),
    .S0(ConfigBits[78+0]),
    .S0N(ConfigBits_N[78+0]),
    .S1(ConfigBits[78+1]),
    .S1N(ConfigBits_N[78+1]),
    .S2(ConfigBits[78+2]),
    .S2N(ConfigBits_N[78+2]),
    .X(E1BEG2)
);

 //switch matrix multiplexer E1BEG3 MUX-8
assign E1BEG3_input = {UIO_OE7,UIO_OE4,UIO_OE3,UIO_OE1,UO_OUT4,UO_OUT1,S1END3,N1END3};
cus_mux81_buf inst_cus_mux81_buf_E1BEG3 (
    .A0(E1BEG3_input[0]),
    .A1(E1BEG3_input[1]),
    .A2(E1BEG3_input[2]),
    .A3(E1BEG3_input[3]),
    .A4(E1BEG3_input[4]),
    .A5(E1BEG3_input[5]),
    .A6(E1BEG3_input[6]),
    .A7(E1BEG3_input[7]),
    .S0(ConfigBits[81+0]),
    .S0N(ConfigBits_N[81+0]),
    .S1(ConfigBits[81+1]),
    .S1N(ConfigBits_N[81+1]),
    .S2(ConfigBits[81+2]),
    .S2N(ConfigBits_N[81+2]),
    .X(E1BEG3)
);

 //switch matrix multiplexer E2BEG0 MUX-8
assign E2BEG0_input = {J_NS1_END0,J_NS2_END7,J_NS2_END0,J_NS4_END0,UIO_OE7,UIO_OUT0,UO_OUT3,UO_OUT0};
cus_mux81_buf inst_cus_mux81_buf_E2BEG0 (
    .A0(E2BEG0_input[0]),
    .A1(E2BEG0_input[1]),
    .A2(E2BEG0_input[2]),
    .A3(E2BEG0_input[3]),
    .A4(E2BEG0_input[4]),
    .A5(E2BEG0_input[5]),
    .A6(E2BEG0_input[6]),
    .A7(E2BEG0_input[7]),
    .S0(ConfigBits[84+0]),
    .S0N(ConfigBits_N[84+0]),
    .S1(ConfigBits[84+1]),
    .S1N(ConfigBits_N[84+1]),
    .S2(ConfigBits[84+2]),
    .S2N(ConfigBits_N[84+2]),
    .X(E2BEG0)
);

 //switch matrix multiplexer E2BEG1 MUX-8
assign E2BEG1_input = {J_NS1_END1,J_NS2_END6,J_NS2_END1,J_NS4_END1,UIO_OE6,UIO_OUT1,UO_OUT2,UO_OUT1};
cus_mux81_buf inst_cus_mux81_buf_E2BEG1 (
    .A0(E2BEG1_input[0]),
    .A1(E2BEG1_input[1]),
    .A2(E2BEG1_input[2]),
    .A3(E2BEG1_input[3]),
    .A4(E2BEG1_input[4]),
    .A5(E2BEG1_input[5]),
    .A6(E2BEG1_input[6]),
    .A7(E2BEG1_input[7]),
    .S0(ConfigBits[87+0]),
    .S0N(ConfigBits_N[87+0]),
    .S1(ConfigBits[87+1]),
    .S1N(ConfigBits_N[87+1]),
    .S2(ConfigBits[87+2]),
    .S2N(ConfigBits_N[87+2]),
    .X(E2BEG1)
);

 //switch matrix multiplexer E2BEG2 MUX-8
assign E2BEG2_input = {J_NS1_END2,J_NS2_END5,J_NS2_END2,J_NS4_END2,UIO_OE5,UIO_OUT2,UO_OUT2,UO_OUT1};
cus_mux81_buf inst_cus_mux81_buf_E2BEG2 (
    .A0(E2BEG2_input[0]),
    .A1(E2BEG2_input[1]),
    .A2(E2BEG2_input[2]),
    .A3(E2BEG2_input[3]),
    .A4(E2BEG2_input[4]),
    .A5(E2BEG2_input[5]),
    .A6(E2BEG2_input[6]),
    .A7(E2BEG2_input[7]),
    .S0(ConfigBits[90+0]),
    .S0N(ConfigBits_N[90+0]),
    .S1(ConfigBits[90+1]),
    .S1N(ConfigBits_N[90+1]),
    .S2(ConfigBits[90+2]),
    .S2N(ConfigBits_N[90+2]),
    .X(E2BEG2)
);

 //switch matrix multiplexer E2BEG3 MUX-8
assign E2BEG3_input = {J_NS1_END3,J_NS2_END4,J_NS2_END3,J_NS4_END3,UIO_OE4,UIO_OUT3,UO_OUT3,UO_OUT0};
cus_mux81_buf inst_cus_mux81_buf_E2BEG3 (
    .A0(E2BEG3_input[0]),
    .A1(E2BEG3_input[1]),
    .A2(E2BEG3_input[2]),
    .A3(E2BEG3_input[3]),
    .A4(E2BEG3_input[4]),
    .A5(E2BEG3_input[5]),
    .A6(E2BEG3_input[6]),
    .A7(E2BEG3_input[7]),
    .S0(ConfigBits[93+0]),
    .S0N(ConfigBits_N[93+0]),
    .S1(ConfigBits[93+1]),
    .S1N(ConfigBits_N[93+1]),
    .S2(ConfigBits[93+2]),
    .S2N(ConfigBits_N[93+2]),
    .X(E2BEG3)
);

 //switch matrix multiplexer E2BEG4 MUX-8
assign E2BEG4_input = {J_NS1_END3,J_NS2_END4,J_NS2_END3,J_NS4_END4,UIO_OE3,UIO_OUT4,UO_OUT7,UO_OUT4};
cus_mux81_buf inst_cus_mux81_buf_E2BEG4 (
    .A0(E2BEG4_input[0]),
    .A1(E2BEG4_input[1]),
    .A2(E2BEG4_input[2]),
    .A3(E2BEG4_input[3]),
    .A4(E2BEG4_input[4]),
    .A5(E2BEG4_input[5]),
    .A6(E2BEG4_input[6]),
    .A7(E2BEG4_input[7]),
    .S0(ConfigBits[96+0]),
    .S0N(ConfigBits_N[96+0]),
    .S1(ConfigBits[96+1]),
    .S1N(ConfigBits_N[96+1]),
    .S2(ConfigBits[96+2]),
    .S2N(ConfigBits_N[96+2]),
    .X(E2BEG4)
);

 //switch matrix multiplexer E2BEG5 MUX-8
assign E2BEG5_input = {J_NS1_END2,J_NS2_END5,J_NS2_END2,J_NS4_END5,UIO_OE2,UIO_OUT5,UO_OUT6,UO_OUT5};
cus_mux81_buf inst_cus_mux81_buf_E2BEG5 (
    .A0(E2BEG5_input[0]),
    .A1(E2BEG5_input[1]),
    .A2(E2BEG5_input[2]),
    .A3(E2BEG5_input[3]),
    .A4(E2BEG5_input[4]),
    .A5(E2BEG5_input[5]),
    .A6(E2BEG5_input[6]),
    .A7(E2BEG5_input[7]),
    .S0(ConfigBits[99+0]),
    .S0N(ConfigBits_N[99+0]),
    .S1(ConfigBits[99+1]),
    .S1N(ConfigBits_N[99+1]),
    .S2(ConfigBits[99+2]),
    .S2N(ConfigBits_N[99+2]),
    .X(E2BEG5)
);

 //switch matrix multiplexer E2BEG6 MUX-8
assign E2BEG6_input = {J_NS1_END1,J_NS2_END6,J_NS2_END1,J_NS4_END6,UIO_OE1,UIO_OUT6,UO_OUT6,UO_OUT5};
cus_mux81_buf inst_cus_mux81_buf_E2BEG6 (
    .A0(E2BEG6_input[0]),
    .A1(E2BEG6_input[1]),
    .A2(E2BEG6_input[2]),
    .A3(E2BEG6_input[3]),
    .A4(E2BEG6_input[4]),
    .A5(E2BEG6_input[5]),
    .A6(E2BEG6_input[6]),
    .A7(E2BEG6_input[7]),
    .S0(ConfigBits[102+0]),
    .S0N(ConfigBits_N[102+0]),
    .S1(ConfigBits[102+1]),
    .S1N(ConfigBits_N[102+1]),
    .S2(ConfigBits[102+2]),
    .S2N(ConfigBits_N[102+2]),
    .X(E2BEG6)
);

 //switch matrix multiplexer E2BEG7 MUX-8
assign E2BEG7_input = {J_NS1_END0,J_NS2_END7,J_NS2_END0,J_NS4_END7,UIO_OE0,UIO_OUT7,UO_OUT7,UO_OUT4};
cus_mux81_buf inst_cus_mux81_buf_E2BEG7 (
    .A0(E2BEG7_input[0]),
    .A1(E2BEG7_input[1]),
    .A2(E2BEG7_input[2]),
    .A3(E2BEG7_input[3]),
    .A4(E2BEG7_input[4]),
    .A5(E2BEG7_input[5]),
    .A6(E2BEG7_input[6]),
    .A7(E2BEG7_input[7]),
    .S0(ConfigBits[105+0]),
    .S0N(ConfigBits_N[105+0]),
    .S1(ConfigBits[105+1]),
    .S1N(ConfigBits_N[105+1]),
    .S2(ConfigBits[105+2]),
    .S2N(ConfigBits_N[105+2]),
    .X(E2BEG7)
);

 //switch matrix multiplexer E2BEGb0 MUX-8
assign E2BEGb0_input = {J_NS2_END7,J_NS2_END0,J_NS4_END8,UIO_OE0,UIO_OUT7,UIO_OUT3,UIO_OUT0,W2END7};
cus_mux81_buf inst_cus_mux81_buf_E2BEGb0 (
    .A0(E2BEGb0_input[0]),
    .A1(E2BEGb0_input[1]),
    .A2(E2BEGb0_input[2]),
    .A3(E2BEGb0_input[3]),
    .A4(E2BEGb0_input[4]),
    .A5(E2BEGb0_input[5]),
    .A6(E2BEGb0_input[6]),
    .A7(E2BEGb0_input[7]),
    .S0(ConfigBits[108+0]),
    .S0N(ConfigBits_N[108+0]),
    .S1(ConfigBits[108+1]),
    .S1N(ConfigBits_N[108+1]),
    .S2(ConfigBits[108+2]),
    .S2N(ConfigBits_N[108+2]),
    .X(E2BEGb0)
);

 //switch matrix multiplexer E2BEGb1 MUX-8
assign E2BEGb1_input = {J_NS2_END6,J_NS2_END1,J_NS4_END9,UIO_OE1,UIO_OUT6,UIO_OUT2,UIO_OUT1,W2END6};
cus_mux81_buf inst_cus_mux81_buf_E2BEGb1 (
    .A0(E2BEGb1_input[0]),
    .A1(E2BEGb1_input[1]),
    .A2(E2BEGb1_input[2]),
    .A3(E2BEGb1_input[3]),
    .A4(E2BEGb1_input[4]),
    .A5(E2BEGb1_input[5]),
    .A6(E2BEGb1_input[6]),
    .A7(E2BEGb1_input[7]),
    .S0(ConfigBits[111+0]),
    .S0N(ConfigBits_N[111+0]),
    .S1(ConfigBits[111+1]),
    .S1N(ConfigBits_N[111+1]),
    .S2(ConfigBits[111+2]),
    .S2N(ConfigBits_N[111+2]),
    .X(E2BEGb1)
);

 //switch matrix multiplexer E2BEGb2 MUX-8
assign E2BEGb2_input = {J_NS2_END5,J_NS2_END2,J_NS4_END10,UIO_OE2,UIO_OUT5,UIO_OUT2,UIO_OUT1,W2END5};
cus_mux81_buf inst_cus_mux81_buf_E2BEGb2 (
    .A0(E2BEGb2_input[0]),
    .A1(E2BEGb2_input[1]),
    .A2(E2BEGb2_input[2]),
    .A3(E2BEGb2_input[3]),
    .A4(E2BEGb2_input[4]),
    .A5(E2BEGb2_input[5]),
    .A6(E2BEGb2_input[6]),
    .A7(E2BEGb2_input[7]),
    .S0(ConfigBits[114+0]),
    .S0N(ConfigBits_N[114+0]),
    .S1(ConfigBits[114+1]),
    .S1N(ConfigBits_N[114+1]),
    .S2(ConfigBits[114+2]),
    .S2N(ConfigBits_N[114+2]),
    .X(E2BEGb2)
);

 //switch matrix multiplexer E2BEGb3 MUX-8
assign E2BEGb3_input = {J_NS2_END4,J_NS2_END3,J_NS4_END11,UIO_OE3,UIO_OUT4,UIO_OUT3,UIO_OUT0,W2END4};
cus_mux81_buf inst_cus_mux81_buf_E2BEGb3 (
    .A0(E2BEGb3_input[0]),
    .A1(E2BEGb3_input[1]),
    .A2(E2BEGb3_input[2]),
    .A3(E2BEGb3_input[3]),
    .A4(E2BEGb3_input[4]),
    .A5(E2BEGb3_input[5]),
    .A6(E2BEGb3_input[6]),
    .A7(E2BEGb3_input[7]),
    .S0(ConfigBits[117+0]),
    .S0N(ConfigBits_N[117+0]),
    .S1(ConfigBits[117+1]),
    .S1N(ConfigBits_N[117+1]),
    .S2(ConfigBits[117+2]),
    .S2N(ConfigBits_N[117+2]),
    .X(E2BEGb3)
);

 //switch matrix multiplexer E2BEGb4 MUX-8
assign E2BEGb4_input = {J_NS2_END4,J_NS2_END3,J_NS4_END12,UIO_OE4,UIO_OUT7,UIO_OUT4,UIO_OUT3,W2END3};
cus_mux81_buf inst_cus_mux81_buf_E2BEGb4 (
    .A0(E2BEGb4_input[0]),
    .A1(E2BEGb4_input[1]),
    .A2(E2BEGb4_input[2]),
    .A3(E2BEGb4_input[3]),
    .A4(E2BEGb4_input[4]),
    .A5(E2BEGb4_input[5]),
    .A6(E2BEGb4_input[6]),
    .A7(E2BEGb4_input[7]),
    .S0(ConfigBits[120+0]),
    .S0N(ConfigBits_N[120+0]),
    .S1(ConfigBits[120+1]),
    .S1N(ConfigBits_N[120+1]),
    .S2(ConfigBits[120+2]),
    .S2N(ConfigBits_N[120+2]),
    .X(E2BEGb4)
);

 //switch matrix multiplexer E2BEGb5 MUX-8
assign E2BEGb5_input = {J_NS2_END5,J_NS2_END2,J_NS4_END13,UIO_OE5,UIO_OUT6,UIO_OUT5,UIO_OUT2,W2END2};
cus_mux81_buf inst_cus_mux81_buf_E2BEGb5 (
    .A0(E2BEGb5_input[0]),
    .A1(E2BEGb5_input[1]),
    .A2(E2BEGb5_input[2]),
    .A3(E2BEGb5_input[3]),
    .A4(E2BEGb5_input[4]),
    .A5(E2BEGb5_input[5]),
    .A6(E2BEGb5_input[6]),
    .A7(E2BEGb5_input[7]),
    .S0(ConfigBits[123+0]),
    .S0N(ConfigBits_N[123+0]),
    .S1(ConfigBits[123+1]),
    .S1N(ConfigBits_N[123+1]),
    .S2(ConfigBits[123+2]),
    .S2N(ConfigBits_N[123+2]),
    .X(E2BEGb5)
);

 //switch matrix multiplexer E2BEGb6 MUX-8
assign E2BEGb6_input = {J_NS2_END6,J_NS2_END1,J_NS4_END14,UIO_OE6,UIO_OUT6,UIO_OUT5,UIO_OUT1,W2END1};
cus_mux81_buf inst_cus_mux81_buf_E2BEGb6 (
    .A0(E2BEGb6_input[0]),
    .A1(E2BEGb6_input[1]),
    .A2(E2BEGb6_input[2]),
    .A3(E2BEGb6_input[3]),
    .A4(E2BEGb6_input[4]),
    .A5(E2BEGb6_input[5]),
    .A6(E2BEGb6_input[6]),
    .A7(E2BEGb6_input[7]),
    .S0(ConfigBits[126+0]),
    .S0N(ConfigBits_N[126+0]),
    .S1(ConfigBits[126+1]),
    .S1N(ConfigBits_N[126+1]),
    .S2(ConfigBits[126+2]),
    .S2N(ConfigBits_N[126+2]),
    .X(E2BEGb6)
);

 //switch matrix multiplexer E2BEGb7 MUX-8
assign E2BEGb7_input = {J_NS2_END7,J_NS2_END0,J_NS4_END15,UIO_OE7,UIO_OUT7,UIO_OUT4,UIO_OUT0,W2END0};
cus_mux81_buf inst_cus_mux81_buf_E2BEGb7 (
    .A0(E2BEGb7_input[0]),
    .A1(E2BEGb7_input[1]),
    .A2(E2BEGb7_input[2]),
    .A3(E2BEGb7_input[3]),
    .A4(E2BEGb7_input[4]),
    .A5(E2BEGb7_input[5]),
    .A6(E2BEGb7_input[6]),
    .A7(E2BEGb7_input[7]),
    .S0(ConfigBits[129+0]),
    .S0N(ConfigBits_N[129+0]),
    .S1(ConfigBits[129+1]),
    .S1N(ConfigBits_N[129+1]),
    .S2(ConfigBits[129+2]),
    .S2N(ConfigBits_N[129+2]),
    .X(E2BEGb7)
);

 //switch matrix multiplexer EE4BEG0 MUX-4
assign EE4BEG0_input = {J_NS2_END7,J_NS4_END15,UIO_OE4,UO_OUT0};
cus_mux41_buf inst_cus_mux41_buf_EE4BEG0 (
    .A0(EE4BEG0_input[0]),
    .A1(EE4BEG0_input[1]),
    .A2(EE4BEG0_input[2]),
    .A3(EE4BEG0_input[3]),
    .S0(ConfigBits[132+0]),
    .S0N(ConfigBits_N[132+0]),
    .S1(ConfigBits[132+1]),
    .S1N(ConfigBits_N[132+1]),
    .X(EE4BEG0)
);

 //switch matrix multiplexer EE4BEG1 MUX-4
assign EE4BEG1_input = {J_NS2_END6,J_NS4_END14,UIO_OE5,UO_OUT1};
cus_mux41_buf inst_cus_mux41_buf_EE4BEG1 (
    .A0(EE4BEG1_input[0]),
    .A1(EE4BEG1_input[1]),
    .A2(EE4BEG1_input[2]),
    .A3(EE4BEG1_input[3]),
    .S0(ConfigBits[134+0]),
    .S0N(ConfigBits_N[134+0]),
    .S1(ConfigBits[134+1]),
    .S1N(ConfigBits_N[134+1]),
    .X(EE4BEG1)
);

 //switch matrix multiplexer EE4BEG2 MUX-4
assign EE4BEG2_input = {J_NS2_END5,J_NS4_END13,UIO_OE6,UO_OUT2};
cus_mux41_buf inst_cus_mux41_buf_EE4BEG2 (
    .A0(EE4BEG2_input[0]),
    .A1(EE4BEG2_input[1]),
    .A2(EE4BEG2_input[2]),
    .A3(EE4BEG2_input[3]),
    .S0(ConfigBits[136+0]),
    .S0N(ConfigBits_N[136+0]),
    .S1(ConfigBits[136+1]),
    .S1N(ConfigBits_N[136+1]),
    .X(EE4BEG2)
);

 //switch matrix multiplexer EE4BEG3 MUX-4
assign EE4BEG3_input = {J_NS2_END4,J_NS4_END12,UIO_OE7,UO_OUT3};
cus_mux41_buf inst_cus_mux41_buf_EE4BEG3 (
    .A0(EE4BEG3_input[0]),
    .A1(EE4BEG3_input[1]),
    .A2(EE4BEG3_input[2]),
    .A3(EE4BEG3_input[3]),
    .S0(ConfigBits[138+0]),
    .S0N(ConfigBits_N[138+0]),
    .S1(ConfigBits[138+1]),
    .S1N(ConfigBits_N[138+1]),
    .X(EE4BEG3)
);

 //switch matrix multiplexer EE4BEG4 MUX-4
assign EE4BEG4_input = {J_NS2_END3,J_NS4_END11,UIO_OE0,UO_OUT4};
cus_mux41_buf inst_cus_mux41_buf_EE4BEG4 (
    .A0(EE4BEG4_input[0]),
    .A1(EE4BEG4_input[1]),
    .A2(EE4BEG4_input[2]),
    .A3(EE4BEG4_input[3]),
    .S0(ConfigBits[140+0]),
    .S0N(ConfigBits_N[140+0]),
    .S1(ConfigBits[140+1]),
    .S1N(ConfigBits_N[140+1]),
    .X(EE4BEG4)
);

 //switch matrix multiplexer EE4BEG5 MUX-4
assign EE4BEG5_input = {J_NS2_END2,J_NS4_END10,UIO_OE1,UO_OUT5};
cus_mux41_buf inst_cus_mux41_buf_EE4BEG5 (
    .A0(EE4BEG5_input[0]),
    .A1(EE4BEG5_input[1]),
    .A2(EE4BEG5_input[2]),
    .A3(EE4BEG5_input[3]),
    .S0(ConfigBits[142+0]),
    .S0N(ConfigBits_N[142+0]),
    .S1(ConfigBits[142+1]),
    .S1N(ConfigBits_N[142+1]),
    .X(EE4BEG5)
);

 //switch matrix multiplexer EE4BEG6 MUX-4
assign EE4BEG6_input = {J_NS2_END1,J_NS4_END9,UIO_OE2,UO_OUT6};
cus_mux41_buf inst_cus_mux41_buf_EE4BEG6 (
    .A0(EE4BEG6_input[0]),
    .A1(EE4BEG6_input[1]),
    .A2(EE4BEG6_input[2]),
    .A3(EE4BEG6_input[3]),
    .S0(ConfigBits[144+0]),
    .S0N(ConfigBits_N[144+0]),
    .S1(ConfigBits[144+1]),
    .S1N(ConfigBits_N[144+1]),
    .X(EE4BEG6)
);

 //switch matrix multiplexer EE4BEG7 MUX-4
assign EE4BEG7_input = {J_NS2_END0,J_NS4_END8,UIO_OE3,UO_OUT7};
cus_mux41_buf inst_cus_mux41_buf_EE4BEG7 (
    .A0(EE4BEG7_input[0]),
    .A1(EE4BEG7_input[1]),
    .A2(EE4BEG7_input[2]),
    .A3(EE4BEG7_input[3]),
    .S0(ConfigBits[146+0]),
    .S0N(ConfigBits_N[146+0]),
    .S1(ConfigBits[146+1]),
    .S1N(ConfigBits_N[146+1]),
    .X(EE4BEG7)
);

 //switch matrix multiplexer EE4BEG8 MUX-4
assign EE4BEG8_input = {J_NS2_END7,J_NS4_END7,UIO_OUT0,UO_OUT4};
cus_mux41_buf inst_cus_mux41_buf_EE4BEG8 (
    .A0(EE4BEG8_input[0]),
    .A1(EE4BEG8_input[1]),
    .A2(EE4BEG8_input[2]),
    .A3(EE4BEG8_input[3]),
    .S0(ConfigBits[148+0]),
    .S0N(ConfigBits_N[148+0]),
    .S1(ConfigBits[148+1]),
    .S1N(ConfigBits_N[148+1]),
    .X(EE4BEG8)
);

 //switch matrix multiplexer EE4BEG9 MUX-4
assign EE4BEG9_input = {J_NS2_END6,J_NS4_END6,UIO_OUT1,UO_OUT5};
cus_mux41_buf inst_cus_mux41_buf_EE4BEG9 (
    .A0(EE4BEG9_input[0]),
    .A1(EE4BEG9_input[1]),
    .A2(EE4BEG9_input[2]),
    .A3(EE4BEG9_input[3]),
    .S0(ConfigBits[150+0]),
    .S0N(ConfigBits_N[150+0]),
    .S1(ConfigBits[150+1]),
    .S1N(ConfigBits_N[150+1]),
    .X(EE4BEG9)
);

 //switch matrix multiplexer EE4BEG10 MUX-4
assign EE4BEG10_input = {J_NS2_END5,J_NS4_END5,UIO_OUT2,UO_OUT6};
cus_mux41_buf inst_cus_mux41_buf_EE4BEG10 (
    .A0(EE4BEG10_input[0]),
    .A1(EE4BEG10_input[1]),
    .A2(EE4BEG10_input[2]),
    .A3(EE4BEG10_input[3]),
    .S0(ConfigBits[152+0]),
    .S0N(ConfigBits_N[152+0]),
    .S1(ConfigBits[152+1]),
    .S1N(ConfigBits_N[152+1]),
    .X(EE4BEG10)
);

 //switch matrix multiplexer EE4BEG11 MUX-4
assign EE4BEG11_input = {J_NS2_END4,J_NS4_END4,UIO_OUT3,UO_OUT7};
cus_mux41_buf inst_cus_mux41_buf_EE4BEG11 (
    .A0(EE4BEG11_input[0]),
    .A1(EE4BEG11_input[1]),
    .A2(EE4BEG11_input[2]),
    .A3(EE4BEG11_input[3]),
    .S0(ConfigBits[154+0]),
    .S0N(ConfigBits_N[154+0]),
    .S1(ConfigBits[154+1]),
    .S1N(ConfigBits_N[154+1]),
    .X(EE4BEG11)
);

 //switch matrix multiplexer EE4BEG12 MUX-4
assign EE4BEG12_input = {J_NS2_END3,J_NS4_END3,UIO_OUT4,UO_OUT0};
cus_mux41_buf inst_cus_mux41_buf_EE4BEG12 (
    .A0(EE4BEG12_input[0]),
    .A1(EE4BEG12_input[1]),
    .A2(EE4BEG12_input[2]),
    .A3(EE4BEG12_input[3]),
    .S0(ConfigBits[156+0]),
    .S0N(ConfigBits_N[156+0]),
    .S1(ConfigBits[156+1]),
    .S1N(ConfigBits_N[156+1]),
    .X(EE4BEG12)
);

 //switch matrix multiplexer EE4BEG13 MUX-4
assign EE4BEG13_input = {J_NS2_END2,J_NS4_END2,UIO_OUT5,UO_OUT1};
cus_mux41_buf inst_cus_mux41_buf_EE4BEG13 (
    .A0(EE4BEG13_input[0]),
    .A1(EE4BEG13_input[1]),
    .A2(EE4BEG13_input[2]),
    .A3(EE4BEG13_input[3]),
    .S0(ConfigBits[158+0]),
    .S0N(ConfigBits_N[158+0]),
    .S1(ConfigBits[158+1]),
    .S1N(ConfigBits_N[158+1]),
    .X(EE4BEG13)
);

 //switch matrix multiplexer EE4BEG14 MUX-4
assign EE4BEG14_input = {J_NS2_END1,J_NS4_END1,UIO_OUT6,UO_OUT2};
cus_mux41_buf inst_cus_mux41_buf_EE4BEG14 (
    .A0(EE4BEG14_input[0]),
    .A1(EE4BEG14_input[1]),
    .A2(EE4BEG14_input[2]),
    .A3(EE4BEG14_input[3]),
    .S0(ConfigBits[160+0]),
    .S0N(ConfigBits_N[160+0]),
    .S1(ConfigBits[160+1]),
    .S1N(ConfigBits_N[160+1]),
    .X(EE4BEG14)
);

 //switch matrix multiplexer EE4BEG15 MUX-4
assign EE4BEG15_input = {J_NS2_END0,J_NS4_END0,UIO_OUT7,UO_OUT3};
cus_mux41_buf inst_cus_mux41_buf_EE4BEG15 (
    .A0(EE4BEG15_input[0]),
    .A1(EE4BEG15_input[1]),
    .A2(EE4BEG15_input[2]),
    .A3(EE4BEG15_input[3]),
    .S0(ConfigBits[162+0]),
    .S0N(ConfigBits_N[162+0]),
    .S1(ConfigBits[162+1]),
    .S1N(ConfigBits_N[162+1]),
    .X(EE4BEG15)
);

 //switch matrix multiplexer E6BEG0 MUX-4
assign E6BEG0_input = {J_NS4_END15,J_NS4_END11,S4END0,N4END0};
cus_mux41_buf inst_cus_mux41_buf_E6BEG0 (
    .A0(E6BEG0_input[0]),
    .A1(E6BEG0_input[1]),
    .A2(E6BEG0_input[2]),
    .A3(E6BEG0_input[3]),
    .S0(ConfigBits[164+0]),
    .S0N(ConfigBits_N[164+0]),
    .S1(ConfigBits[164+1]),
    .S1N(ConfigBits_N[164+1]),
    .X(E6BEG0)
);

 //switch matrix multiplexer E6BEG1 MUX-4
assign E6BEG1_input = {J_NS4_END14,J_NS4_END10,S4END1,N4END1};
cus_mux41_buf inst_cus_mux41_buf_E6BEG1 (
    .A0(E6BEG1_input[0]),
    .A1(E6BEG1_input[1]),
    .A2(E6BEG1_input[2]),
    .A3(E6BEG1_input[3]),
    .S0(ConfigBits[166+0]),
    .S0N(ConfigBits_N[166+0]),
    .S1(ConfigBits[166+1]),
    .S1N(ConfigBits_N[166+1]),
    .X(E6BEG1)
);

 //switch matrix multiplexer E6BEG2 MUX-4
assign E6BEG2_input = {J_NS4_END13,J_NS4_END9,S4END2,N4END2};
cus_mux41_buf inst_cus_mux41_buf_E6BEG2 (
    .A0(E6BEG2_input[0]),
    .A1(E6BEG2_input[1]),
    .A2(E6BEG2_input[2]),
    .A3(E6BEG2_input[3]),
    .S0(ConfigBits[168+0]),
    .S0N(ConfigBits_N[168+0]),
    .S1(ConfigBits[168+1]),
    .S1N(ConfigBits_N[168+1]),
    .X(E6BEG2)
);

 //switch matrix multiplexer E6BEG3 MUX-4
assign E6BEG3_input = {J_NS4_END12,J_NS4_END8,S4END3,N4END3};
cus_mux41_buf inst_cus_mux41_buf_E6BEG3 (
    .A0(E6BEG3_input[0]),
    .A1(E6BEG3_input[1]),
    .A2(E6BEG3_input[2]),
    .A3(E6BEG3_input[3]),
    .S0(ConfigBits[170+0]),
    .S0N(ConfigBits_N[170+0]),
    .S1(ConfigBits[170+1]),
    .S1N(ConfigBits_N[170+1]),
    .X(E6BEG3)
);

 //switch matrix multiplexer E6BEG4 MUX-4
assign E6BEG4_input = {J_NS2_END0,J_NS4_END11,J_NS4_END7,UIO_OUT4};
cus_mux41_buf inst_cus_mux41_buf_E6BEG4 (
    .A0(E6BEG4_input[0]),
    .A1(E6BEG4_input[1]),
    .A2(E6BEG4_input[2]),
    .A3(E6BEG4_input[3]),
    .S0(ConfigBits[172+0]),
    .S0N(ConfigBits_N[172+0]),
    .S1(ConfigBits[172+1]),
    .S1N(ConfigBits_N[172+1]),
    .X(E6BEG4)
);

 //switch matrix multiplexer E6BEG5 MUX-4
assign E6BEG5_input = {J_NS2_END1,J_NS4_END10,J_NS4_END6,UIO_OUT5};
cus_mux41_buf inst_cus_mux41_buf_E6BEG5 (
    .A0(E6BEG5_input[0]),
    .A1(E6BEG5_input[1]),
    .A2(E6BEG5_input[2]),
    .A3(E6BEG5_input[3]),
    .S0(ConfigBits[174+0]),
    .S0N(ConfigBits_N[174+0]),
    .S1(ConfigBits[174+1]),
    .S1N(ConfigBits_N[174+1]),
    .X(E6BEG5)
);

 //switch matrix multiplexer E6BEG6 MUX-4
assign E6BEG6_input = {J_NS2_END2,J_NS4_END9,J_NS4_END5,UIO_OUT6};
cus_mux41_buf inst_cus_mux41_buf_E6BEG6 (
    .A0(E6BEG6_input[0]),
    .A1(E6BEG6_input[1]),
    .A2(E6BEG6_input[2]),
    .A3(E6BEG6_input[3]),
    .S0(ConfigBits[176+0]),
    .S0N(ConfigBits_N[176+0]),
    .S1(ConfigBits[176+1]),
    .S1N(ConfigBits_N[176+1]),
    .X(E6BEG6)
);

 //switch matrix multiplexer E6BEG7 MUX-4
assign E6BEG7_input = {J_NS2_END3,J_NS4_END8,J_NS4_END4,UIO_OUT7};
cus_mux41_buf inst_cus_mux41_buf_E6BEG7 (
    .A0(E6BEG7_input[0]),
    .A1(E6BEG7_input[1]),
    .A2(E6BEG7_input[2]),
    .A3(E6BEG7_input[3]),
    .S0(ConfigBits[178+0]),
    .S0N(ConfigBits_N[178+0]),
    .S1(ConfigBits[178+1]),
    .S1N(ConfigBits_N[178+1]),
    .X(E6BEG7)
);

 //switch matrix multiplexer E6BEG8 MUX-4
assign E6BEG8_input = {J_NS2_END4,J_NS4_END7,J_NS4_END3,UIO_OUT0};
cus_mux41_buf inst_cus_mux41_buf_E6BEG8 (
    .A0(E6BEG8_input[0]),
    .A1(E6BEG8_input[1]),
    .A2(E6BEG8_input[2]),
    .A3(E6BEG8_input[3]),
    .S0(ConfigBits[180+0]),
    .S0N(ConfigBits_N[180+0]),
    .S1(ConfigBits[180+1]),
    .S1N(ConfigBits_N[180+1]),
    .X(E6BEG8)
);

 //switch matrix multiplexer E6BEG9 MUX-4
assign E6BEG9_input = {J_NS2_END5,J_NS4_END6,J_NS4_END2,UIO_OUT1};
cus_mux41_buf inst_cus_mux41_buf_E6BEG9 (
    .A0(E6BEG9_input[0]),
    .A1(E6BEG9_input[1]),
    .A2(E6BEG9_input[2]),
    .A3(E6BEG9_input[3]),
    .S0(ConfigBits[182+0]),
    .S0N(ConfigBits_N[182+0]),
    .S1(ConfigBits[182+1]),
    .S1N(ConfigBits_N[182+1]),
    .X(E6BEG9)
);

 //switch matrix multiplexer E6BEG10 MUX-4
assign E6BEG10_input = {J_NS2_END6,J_NS4_END5,J_NS4_END1,UIO_OUT2};
cus_mux41_buf inst_cus_mux41_buf_E6BEG10 (
    .A0(E6BEG10_input[0]),
    .A1(E6BEG10_input[1]),
    .A2(E6BEG10_input[2]),
    .A3(E6BEG10_input[3]),
    .S0(ConfigBits[184+0]),
    .S0N(ConfigBits_N[184+0]),
    .S1(ConfigBits[184+1]),
    .S1N(ConfigBits_N[184+1]),
    .X(E6BEG10)
);

 //switch matrix multiplexer E6BEG11 MUX-4
assign E6BEG11_input = {J_NS2_END7,J_NS4_END4,J_NS4_END0,UIO_OUT3};
cus_mux41_buf inst_cus_mux41_buf_E6BEG11 (
    .A0(E6BEG11_input[0]),
    .A1(E6BEG11_input[1]),
    .A2(E6BEG11_input[2]),
    .A3(E6BEG11_input[3]),
    .S0(ConfigBits[186+0]),
    .S0N(ConfigBits_N[186+0]),
    .S1(ConfigBits[186+1]),
    .S1N(ConfigBits_N[186+1]),
    .X(E6BEG11)
);

 //switch matrix multiplexer UI_IN0 MUX-8
assign UI_IN0_input = {GND0,J_NS2_END0,J_NS4_END0,W6END0,WW4END8,WW4END0,W2END0,W2MID0};
cus_mux81_buf inst_cus_mux81_buf_UI_IN0 (
    .A0(UI_IN0_input[0]),
    .A1(UI_IN0_input[1]),
    .A2(UI_IN0_input[2]),
    .A3(UI_IN0_input[3]),
    .A4(UI_IN0_input[4]),
    .A5(UI_IN0_input[5]),
    .A6(UI_IN0_input[6]),
    .A7(UI_IN0_input[7]),
    .S0(ConfigBits[188+0]),
    .S0N(ConfigBits_N[188+0]),
    .S1(ConfigBits[188+1]),
    .S1N(ConfigBits_N[188+1]),
    .S2(ConfigBits[188+2]),
    .S2N(ConfigBits_N[188+2]),
    .X(UI_IN0)
);

 //switch matrix multiplexer UI_IN1 MUX-8
assign UI_IN1_input = {GND0,J_NS2_END1,J_NS4_END1,W6END1,WW4END9,WW4END1,W2END1,W2MID1};
cus_mux81_buf inst_cus_mux81_buf_UI_IN1 (
    .A0(UI_IN1_input[0]),
    .A1(UI_IN1_input[1]),
    .A2(UI_IN1_input[2]),
    .A3(UI_IN1_input[3]),
    .A4(UI_IN1_input[4]),
    .A5(UI_IN1_input[5]),
    .A6(UI_IN1_input[6]),
    .A7(UI_IN1_input[7]),
    .S0(ConfigBits[191+0]),
    .S0N(ConfigBits_N[191+0]),
    .S1(ConfigBits[191+1]),
    .S1N(ConfigBits_N[191+1]),
    .S2(ConfigBits[191+2]),
    .S2N(ConfigBits_N[191+2]),
    .X(UI_IN1)
);

 //switch matrix multiplexer UI_IN2 MUX-8
assign UI_IN2_input = {GND0,J_NS2_END2,J_NS4_END2,W6END2,WW4END10,WW4END2,W2END2,W2MID2};
cus_mux81_buf inst_cus_mux81_buf_UI_IN2 (
    .A0(UI_IN2_input[0]),
    .A1(UI_IN2_input[1]),
    .A2(UI_IN2_input[2]),
    .A3(UI_IN2_input[3]),
    .A4(UI_IN2_input[4]),
    .A5(UI_IN2_input[5]),
    .A6(UI_IN2_input[6]),
    .A7(UI_IN2_input[7]),
    .S0(ConfigBits[194+0]),
    .S0N(ConfigBits_N[194+0]),
    .S1(ConfigBits[194+1]),
    .S1N(ConfigBits_N[194+1]),
    .S2(ConfigBits[194+2]),
    .S2N(ConfigBits_N[194+2]),
    .X(UI_IN2)
);

 //switch matrix multiplexer UI_IN3 MUX-8
assign UI_IN3_input = {GND0,J_NS2_END3,J_NS4_END3,W6END3,WW4END11,WW4END3,W2END3,W2MID3};
cus_mux81_buf inst_cus_mux81_buf_UI_IN3 (
    .A0(UI_IN3_input[0]),
    .A1(UI_IN3_input[1]),
    .A2(UI_IN3_input[2]),
    .A3(UI_IN3_input[3]),
    .A4(UI_IN3_input[4]),
    .A5(UI_IN3_input[5]),
    .A6(UI_IN3_input[6]),
    .A7(UI_IN3_input[7]),
    .S0(ConfigBits[197+0]),
    .S0N(ConfigBits_N[197+0]),
    .S1(ConfigBits[197+1]),
    .S1N(ConfigBits_N[197+1]),
    .S2(ConfigBits[197+2]),
    .S2N(ConfigBits_N[197+2]),
    .X(UI_IN3)
);

 //switch matrix multiplexer UI_IN4 MUX-8
assign UI_IN4_input = {GND0,J_NS2_END4,J_NS4_END4,W6END4,WW4END12,WW4END4,W2END4,W2MID4};
cus_mux81_buf inst_cus_mux81_buf_UI_IN4 (
    .A0(UI_IN4_input[0]),
    .A1(UI_IN4_input[1]),
    .A2(UI_IN4_input[2]),
    .A3(UI_IN4_input[3]),
    .A4(UI_IN4_input[4]),
    .A5(UI_IN4_input[5]),
    .A6(UI_IN4_input[6]),
    .A7(UI_IN4_input[7]),
    .S0(ConfigBits[200+0]),
    .S0N(ConfigBits_N[200+0]),
    .S1(ConfigBits[200+1]),
    .S1N(ConfigBits_N[200+1]),
    .S2(ConfigBits[200+2]),
    .S2N(ConfigBits_N[200+2]),
    .X(UI_IN4)
);

 //switch matrix multiplexer UI_IN5 MUX-8
assign UI_IN5_input = {GND0,J_NS2_END5,J_NS4_END5,W6END5,WW4END13,WW4END5,W2END5,W2MID5};
cus_mux81_buf inst_cus_mux81_buf_UI_IN5 (
    .A0(UI_IN5_input[0]),
    .A1(UI_IN5_input[1]),
    .A2(UI_IN5_input[2]),
    .A3(UI_IN5_input[3]),
    .A4(UI_IN5_input[4]),
    .A5(UI_IN5_input[5]),
    .A6(UI_IN5_input[6]),
    .A7(UI_IN5_input[7]),
    .S0(ConfigBits[203+0]),
    .S0N(ConfigBits_N[203+0]),
    .S1(ConfigBits[203+1]),
    .S1N(ConfigBits_N[203+1]),
    .S2(ConfigBits[203+2]),
    .S2N(ConfigBits_N[203+2]),
    .X(UI_IN5)
);

 //switch matrix multiplexer UI_IN6 MUX-8
assign UI_IN6_input = {GND0,J_NS2_END6,J_NS4_END6,W6END6,WW4END14,WW4END6,W2END6,W2MID6};
cus_mux81_buf inst_cus_mux81_buf_UI_IN6 (
    .A0(UI_IN6_input[0]),
    .A1(UI_IN6_input[1]),
    .A2(UI_IN6_input[2]),
    .A3(UI_IN6_input[3]),
    .A4(UI_IN6_input[4]),
    .A5(UI_IN6_input[5]),
    .A6(UI_IN6_input[6]),
    .A7(UI_IN6_input[7]),
    .S0(ConfigBits[206+0]),
    .S0N(ConfigBits_N[206+0]),
    .S1(ConfigBits[206+1]),
    .S1N(ConfigBits_N[206+1]),
    .S2(ConfigBits[206+2]),
    .S2N(ConfigBits_N[206+2]),
    .X(UI_IN6)
);

 //switch matrix multiplexer UI_IN7 MUX-8
assign UI_IN7_input = {GND0,J_NS2_END7,J_NS4_END7,W6END7,WW4END15,WW4END7,W2END7,W2MID7};
cus_mux81_buf inst_cus_mux81_buf_UI_IN7 (
    .A0(UI_IN7_input[0]),
    .A1(UI_IN7_input[1]),
    .A2(UI_IN7_input[2]),
    .A3(UI_IN7_input[3]),
    .A4(UI_IN7_input[4]),
    .A5(UI_IN7_input[5]),
    .A6(UI_IN7_input[6]),
    .A7(UI_IN7_input[7]),
    .S0(ConfigBits[209+0]),
    .S0N(ConfigBits_N[209+0]),
    .S1(ConfigBits[209+1]),
    .S1N(ConfigBits_N[209+1]),
    .S2(ConfigBits[209+2]),
    .S2N(ConfigBits_N[209+2]),
    .X(UI_IN7)
);

 //switch matrix multiplexer UIO_IN0 MUX-8
assign UIO_IN0_input = {GND0,J_NS2_END0,J_NS4_END8,W6END8,WW4END8,WW4END0,W2END0,W2MID0};
cus_mux81_buf inst_cus_mux81_buf_UIO_IN0 (
    .A0(UIO_IN0_input[0]),
    .A1(UIO_IN0_input[1]),
    .A2(UIO_IN0_input[2]),
    .A3(UIO_IN0_input[3]),
    .A4(UIO_IN0_input[4]),
    .A5(UIO_IN0_input[5]),
    .A6(UIO_IN0_input[6]),
    .A7(UIO_IN0_input[7]),
    .S0(ConfigBits[212+0]),
    .S0N(ConfigBits_N[212+0]),
    .S1(ConfigBits[212+1]),
    .S1N(ConfigBits_N[212+1]),
    .S2(ConfigBits[212+2]),
    .S2N(ConfigBits_N[212+2]),
    .X(UIO_IN0)
);

 //switch matrix multiplexer UIO_IN1 MUX-8
assign UIO_IN1_input = {GND0,J_NS2_END1,J_NS4_END9,W6END9,WW4END9,WW4END1,W2END1,W2MID1};
cus_mux81_buf inst_cus_mux81_buf_UIO_IN1 (
    .A0(UIO_IN1_input[0]),
    .A1(UIO_IN1_input[1]),
    .A2(UIO_IN1_input[2]),
    .A3(UIO_IN1_input[3]),
    .A4(UIO_IN1_input[4]),
    .A5(UIO_IN1_input[5]),
    .A6(UIO_IN1_input[6]),
    .A7(UIO_IN1_input[7]),
    .S0(ConfigBits[215+0]),
    .S0N(ConfigBits_N[215+0]),
    .S1(ConfigBits[215+1]),
    .S1N(ConfigBits_N[215+1]),
    .S2(ConfigBits[215+2]),
    .S2N(ConfigBits_N[215+2]),
    .X(UIO_IN1)
);

 //switch matrix multiplexer UIO_IN2 MUX-8
assign UIO_IN2_input = {GND0,J_NS2_END2,J_NS4_END10,W6END10,WW4END10,WW4END2,W2END2,W2MID2};
cus_mux81_buf inst_cus_mux81_buf_UIO_IN2 (
    .A0(UIO_IN2_input[0]),
    .A1(UIO_IN2_input[1]),
    .A2(UIO_IN2_input[2]),
    .A3(UIO_IN2_input[3]),
    .A4(UIO_IN2_input[4]),
    .A5(UIO_IN2_input[5]),
    .A6(UIO_IN2_input[6]),
    .A7(UIO_IN2_input[7]),
    .S0(ConfigBits[218+0]),
    .S0N(ConfigBits_N[218+0]),
    .S1(ConfigBits[218+1]),
    .S1N(ConfigBits_N[218+1]),
    .S2(ConfigBits[218+2]),
    .S2N(ConfigBits_N[218+2]),
    .X(UIO_IN2)
);

 //switch matrix multiplexer UIO_IN3 MUX-8
assign UIO_IN3_input = {GND0,J_NS2_END3,J_NS4_END11,W6END11,WW4END11,WW4END3,W2END3,W2MID3};
cus_mux81_buf inst_cus_mux81_buf_UIO_IN3 (
    .A0(UIO_IN3_input[0]),
    .A1(UIO_IN3_input[1]),
    .A2(UIO_IN3_input[2]),
    .A3(UIO_IN3_input[3]),
    .A4(UIO_IN3_input[4]),
    .A5(UIO_IN3_input[5]),
    .A6(UIO_IN3_input[6]),
    .A7(UIO_IN3_input[7]),
    .S0(ConfigBits[221+0]),
    .S0N(ConfigBits_N[221+0]),
    .S1(ConfigBits[221+1]),
    .S1N(ConfigBits_N[221+1]),
    .S2(ConfigBits[221+2]),
    .S2N(ConfigBits_N[221+2]),
    .X(UIO_IN3)
);

 //switch matrix multiplexer UIO_IN4 MUX-8
assign UIO_IN4_input = {GND0,J_NS2_END4,J_NS4_END12,WW4END12,WW4END4,W2END4,W2MID4,W1END0};
cus_mux81_buf inst_cus_mux81_buf_UIO_IN4 (
    .A0(UIO_IN4_input[0]),
    .A1(UIO_IN4_input[1]),
    .A2(UIO_IN4_input[2]),
    .A3(UIO_IN4_input[3]),
    .A4(UIO_IN4_input[4]),
    .A5(UIO_IN4_input[5]),
    .A6(UIO_IN4_input[6]),
    .A7(UIO_IN4_input[7]),
    .S0(ConfigBits[224+0]),
    .S0N(ConfigBits_N[224+0]),
    .S1(ConfigBits[224+1]),
    .S1N(ConfigBits_N[224+1]),
    .S2(ConfigBits[224+2]),
    .S2N(ConfigBits_N[224+2]),
    .X(UIO_IN4)
);

 //switch matrix multiplexer UIO_IN5 MUX-8
assign UIO_IN5_input = {GND0,J_NS2_END5,J_NS4_END13,WW4END13,WW4END5,W2END5,W2MID5,W1END1};
cus_mux81_buf inst_cus_mux81_buf_UIO_IN5 (
    .A0(UIO_IN5_input[0]),
    .A1(UIO_IN5_input[1]),
    .A2(UIO_IN5_input[2]),
    .A3(UIO_IN5_input[3]),
    .A4(UIO_IN5_input[4]),
    .A5(UIO_IN5_input[5]),
    .A6(UIO_IN5_input[6]),
    .A7(UIO_IN5_input[7]),
    .S0(ConfigBits[227+0]),
    .S0N(ConfigBits_N[227+0]),
    .S1(ConfigBits[227+1]),
    .S1N(ConfigBits_N[227+1]),
    .S2(ConfigBits[227+2]),
    .S2N(ConfigBits_N[227+2]),
    .X(UIO_IN5)
);

 //switch matrix multiplexer UIO_IN6 MUX-8
assign UIO_IN6_input = {GND0,J_NS2_END6,J_NS4_END14,WW4END14,WW4END6,W2END6,W2MID6,W1END2};
cus_mux81_buf inst_cus_mux81_buf_UIO_IN6 (
    .A0(UIO_IN6_input[0]),
    .A1(UIO_IN6_input[1]),
    .A2(UIO_IN6_input[2]),
    .A3(UIO_IN6_input[3]),
    .A4(UIO_IN6_input[4]),
    .A5(UIO_IN6_input[5]),
    .A6(UIO_IN6_input[6]),
    .A7(UIO_IN6_input[7]),
    .S0(ConfigBits[230+0]),
    .S0N(ConfigBits_N[230+0]),
    .S1(ConfigBits[230+1]),
    .S1N(ConfigBits_N[230+1]),
    .S2(ConfigBits[230+2]),
    .S2N(ConfigBits_N[230+2]),
    .X(UIO_IN6)
);

 //switch matrix multiplexer UIO_IN7 MUX-8
assign UIO_IN7_input = {GND0,J_NS2_END7,J_NS4_END15,WW4END15,WW4END7,W2END7,W2MID7,W1END3};
cus_mux81_buf inst_cus_mux81_buf_UIO_IN7 (
    .A0(UIO_IN7_input[0]),
    .A1(UIO_IN7_input[1]),
    .A2(UIO_IN7_input[2]),
    .A3(UIO_IN7_input[3]),
    .A4(UIO_IN7_input[4]),
    .A5(UIO_IN7_input[5]),
    .A6(UIO_IN7_input[6]),
    .A7(UIO_IN7_input[7]),
    .S0(ConfigBits[233+0]),
    .S0N(ConfigBits_N[233+0]),
    .S1(ConfigBits[233+1]),
    .S1N(ConfigBits_N[233+1]),
    .S2(ConfigBits[233+2]),
    .S2N(ConfigBits_N[233+2]),
    .X(UIO_IN7)
);

 //switch matrix multiplexer ENA MUX-4
assign ENA_input = {VCC0,GND0,W2MID6,N2MID6};
cus_mux41_buf inst_cus_mux41_buf_ENA (
    .A0(ENA_input[0]),
    .A1(ENA_input[1]),
    .A2(ENA_input[2]),
    .A3(ENA_input[3]),
    .S0(ConfigBits[236+0]),
    .S0N(ConfigBits_N[236+0]),
    .S1(ConfigBits[236+1]),
    .S1N(ConfigBits_N[236+1]),
    .X(ENA)
);

 //switch matrix multiplexer RST_N MUX-16
assign RST_N_input = {VCC0,GND0,S2END3,S2END2,S2MID0,W2END5,W2END4,W2END3,W2END2,W2END1,W2MID6,W2MID3,W2MID0,N2END3,N2END2,N2MID6};
cus_mux161_buf inst_cus_mux161_buf_RST_N (
    .A0(RST_N_input[0]),
    .A1(RST_N_input[1]),
    .A2(RST_N_input[2]),
    .A3(RST_N_input[3]),
    .A4(RST_N_input[4]),
    .A5(RST_N_input[5]),
    .A6(RST_N_input[6]),
    .A7(RST_N_input[7]),
    .A8(RST_N_input[8]),
    .A9(RST_N_input[9]),
    .A10(RST_N_input[10]),
    .A11(RST_N_input[11]),
    .A12(RST_N_input[12]),
    .A13(RST_N_input[13]),
    .A14(RST_N_input[14]),
    .A15(RST_N_input[15]),
    .S0(ConfigBits[238+0]),
    .S0N(ConfigBits_N[238+0]),
    .S1(ConfigBits[238+1]),
    .S1N(ConfigBits_N[238+1]),
    .S2(ConfigBits[238+2]),
    .S2N(ConfigBits_N[238+2]),
    .S3(ConfigBits[238+3]),
    .S3N(ConfigBits_N[238+3]),
    .X(RST_N)
);

 //switch matrix multiplexer J_NS4_BEG0 MUX-4
assign J_NS4_BEG0_input = {S4END0,S1END0,N4END0,N1END0};
cus_mux41_buf inst_cus_mux41_buf_J_NS4_BEG0 (
    .A0(J_NS4_BEG0_input[0]),
    .A1(J_NS4_BEG0_input[1]),
    .A2(J_NS4_BEG0_input[2]),
    .A3(J_NS4_BEG0_input[3]),
    .S0(ConfigBits[242+0]),
    .S0N(ConfigBits_N[242+0]),
    .S1(ConfigBits[242+1]),
    .S1N(ConfigBits_N[242+1]),
    .X(J_NS4_BEG0)
);

 //switch matrix multiplexer J_NS4_BEG1 MUX-4
assign J_NS4_BEG1_input = {S4END1,S1END1,N4END1,N1END1};
cus_mux41_buf inst_cus_mux41_buf_J_NS4_BEG1 (
    .A0(J_NS4_BEG1_input[0]),
    .A1(J_NS4_BEG1_input[1]),
    .A2(J_NS4_BEG1_input[2]),
    .A3(J_NS4_BEG1_input[3]),
    .S0(ConfigBits[244+0]),
    .S0N(ConfigBits_N[244+0]),
    .S1(ConfigBits[244+1]),
    .S1N(ConfigBits_N[244+1]),
    .X(J_NS4_BEG1)
);

 //switch matrix multiplexer J_NS4_BEG2 MUX-4
assign J_NS4_BEG2_input = {S4END2,S1END2,N4END2,N1END2};
cus_mux41_buf inst_cus_mux41_buf_J_NS4_BEG2 (
    .A0(J_NS4_BEG2_input[0]),
    .A1(J_NS4_BEG2_input[1]),
    .A2(J_NS4_BEG2_input[2]),
    .A3(J_NS4_BEG2_input[3]),
    .S0(ConfigBits[246+0]),
    .S0N(ConfigBits_N[246+0]),
    .S1(ConfigBits[246+1]),
    .S1N(ConfigBits_N[246+1]),
    .X(J_NS4_BEG2)
);

 //switch matrix multiplexer J_NS4_BEG3 MUX-4
assign J_NS4_BEG3_input = {S4END3,S1END3,N4END3,N1END3};
cus_mux41_buf inst_cus_mux41_buf_J_NS4_BEG3 (
    .A0(J_NS4_BEG3_input[0]),
    .A1(J_NS4_BEG3_input[1]),
    .A2(J_NS4_BEG3_input[2]),
    .A3(J_NS4_BEG3_input[3]),
    .S0(ConfigBits[248+0]),
    .S0N(ConfigBits_N[248+0]),
    .S1(ConfigBits[248+1]),
    .S1N(ConfigBits_N[248+1]),
    .X(J_NS4_BEG3)
);

 //switch matrix multiplexer J_NS4_BEG4 MUX-4
assign J_NS4_BEG4_input = {S4END0,S1END0,N4END0,N1END0};
cus_mux41_buf inst_cus_mux41_buf_J_NS4_BEG4 (
    .A0(J_NS4_BEG4_input[0]),
    .A1(J_NS4_BEG4_input[1]),
    .A2(J_NS4_BEG4_input[2]),
    .A3(J_NS4_BEG4_input[3]),
    .S0(ConfigBits[250+0]),
    .S0N(ConfigBits_N[250+0]),
    .S1(ConfigBits[250+1]),
    .S1N(ConfigBits_N[250+1]),
    .X(J_NS4_BEG4)
);

 //switch matrix multiplexer J_NS4_BEG5 MUX-4
assign J_NS4_BEG5_input = {S4END1,S1END1,N4END1,N1END1};
cus_mux41_buf inst_cus_mux41_buf_J_NS4_BEG5 (
    .A0(J_NS4_BEG5_input[0]),
    .A1(J_NS4_BEG5_input[1]),
    .A2(J_NS4_BEG5_input[2]),
    .A3(J_NS4_BEG5_input[3]),
    .S0(ConfigBits[252+0]),
    .S0N(ConfigBits_N[252+0]),
    .S1(ConfigBits[252+1]),
    .S1N(ConfigBits_N[252+1]),
    .X(J_NS4_BEG5)
);

 //switch matrix multiplexer J_NS4_BEG6 MUX-4
assign J_NS4_BEG6_input = {S4END2,S1END2,N4END2,N1END2};
cus_mux41_buf inst_cus_mux41_buf_J_NS4_BEG6 (
    .A0(J_NS4_BEG6_input[0]),
    .A1(J_NS4_BEG6_input[1]),
    .A2(J_NS4_BEG6_input[2]),
    .A3(J_NS4_BEG6_input[3]),
    .S0(ConfigBits[254+0]),
    .S0N(ConfigBits_N[254+0]),
    .S1(ConfigBits[254+1]),
    .S1N(ConfigBits_N[254+1]),
    .X(J_NS4_BEG6)
);

 //switch matrix multiplexer J_NS4_BEG7 MUX-4
assign J_NS4_BEG7_input = {S4END3,S1END3,N4END3,N1END3};
cus_mux41_buf inst_cus_mux41_buf_J_NS4_BEG7 (
    .A0(J_NS4_BEG7_input[0]),
    .A1(J_NS4_BEG7_input[1]),
    .A2(J_NS4_BEG7_input[2]),
    .A3(J_NS4_BEG7_input[3]),
    .S0(ConfigBits[256+0]),
    .S0N(ConfigBits_N[256+0]),
    .S1(ConfigBits[256+1]),
    .S1N(ConfigBits_N[256+1]),
    .X(J_NS4_BEG7)
);

 //switch matrix multiplexer J_NS4_BEG8 MUX-4
assign J_NS4_BEG8_input = {S4END0,S1END0,N4END0,N1END0};
cus_mux41_buf inst_cus_mux41_buf_J_NS4_BEG8 (
    .A0(J_NS4_BEG8_input[0]),
    .A1(J_NS4_BEG8_input[1]),
    .A2(J_NS4_BEG8_input[2]),
    .A3(J_NS4_BEG8_input[3]),
    .S0(ConfigBits[258+0]),
    .S0N(ConfigBits_N[258+0]),
    .S1(ConfigBits[258+1]),
    .S1N(ConfigBits_N[258+1]),
    .X(J_NS4_BEG8)
);

 //switch matrix multiplexer J_NS4_BEG9 MUX-4
assign J_NS4_BEG9_input = {S4END1,S1END1,N4END1,N1END1};
cus_mux41_buf inst_cus_mux41_buf_J_NS4_BEG9 (
    .A0(J_NS4_BEG9_input[0]),
    .A1(J_NS4_BEG9_input[1]),
    .A2(J_NS4_BEG9_input[2]),
    .A3(J_NS4_BEG9_input[3]),
    .S0(ConfigBits[260+0]),
    .S0N(ConfigBits_N[260+0]),
    .S1(ConfigBits[260+1]),
    .S1N(ConfigBits_N[260+1]),
    .X(J_NS4_BEG9)
);

 //switch matrix multiplexer J_NS4_BEG10 MUX-4
assign J_NS4_BEG10_input = {S4END2,S1END2,N4END2,N1END2};
cus_mux41_buf inst_cus_mux41_buf_J_NS4_BEG10 (
    .A0(J_NS4_BEG10_input[0]),
    .A1(J_NS4_BEG10_input[1]),
    .A2(J_NS4_BEG10_input[2]),
    .A3(J_NS4_BEG10_input[3]),
    .S0(ConfigBits[262+0]),
    .S0N(ConfigBits_N[262+0]),
    .S1(ConfigBits[262+1]),
    .S1N(ConfigBits_N[262+1]),
    .X(J_NS4_BEG10)
);

 //switch matrix multiplexer J_NS4_BEG11 MUX-4
assign J_NS4_BEG11_input = {S4END3,S1END3,N4END3,N1END3};
cus_mux41_buf inst_cus_mux41_buf_J_NS4_BEG11 (
    .A0(J_NS4_BEG11_input[0]),
    .A1(J_NS4_BEG11_input[1]),
    .A2(J_NS4_BEG11_input[2]),
    .A3(J_NS4_BEG11_input[3]),
    .S0(ConfigBits[264+0]),
    .S0N(ConfigBits_N[264+0]),
    .S1(ConfigBits[264+1]),
    .S1N(ConfigBits_N[264+1]),
    .X(J_NS4_BEG11)
);

 //switch matrix multiplexer J_NS4_BEG12 MUX-4
assign J_NS4_BEG12_input = {S4END0,S1END0,N4END0,N1END0};
cus_mux41_buf inst_cus_mux41_buf_J_NS4_BEG12 (
    .A0(J_NS4_BEG12_input[0]),
    .A1(J_NS4_BEG12_input[1]),
    .A2(J_NS4_BEG12_input[2]),
    .A3(J_NS4_BEG12_input[3]),
    .S0(ConfigBits[266+0]),
    .S0N(ConfigBits_N[266+0]),
    .S1(ConfigBits[266+1]),
    .S1N(ConfigBits_N[266+1]),
    .X(J_NS4_BEG12)
);

 //switch matrix multiplexer J_NS4_BEG13 MUX-4
assign J_NS4_BEG13_input = {S4END1,S1END1,N4END1,N1END1};
cus_mux41_buf inst_cus_mux41_buf_J_NS4_BEG13 (
    .A0(J_NS4_BEG13_input[0]),
    .A1(J_NS4_BEG13_input[1]),
    .A2(J_NS4_BEG13_input[2]),
    .A3(J_NS4_BEG13_input[3]),
    .S0(ConfigBits[268+0]),
    .S0N(ConfigBits_N[268+0]),
    .S1(ConfigBits[268+1]),
    .S1N(ConfigBits_N[268+1]),
    .X(J_NS4_BEG13)
);

 //switch matrix multiplexer J_NS4_BEG14 MUX-4
assign J_NS4_BEG14_input = {S4END2,S1END2,N4END2,N1END2};
cus_mux41_buf inst_cus_mux41_buf_J_NS4_BEG14 (
    .A0(J_NS4_BEG14_input[0]),
    .A1(J_NS4_BEG14_input[1]),
    .A2(J_NS4_BEG14_input[2]),
    .A3(J_NS4_BEG14_input[3]),
    .S0(ConfigBits[270+0]),
    .S0N(ConfigBits_N[270+0]),
    .S1(ConfigBits[270+1]),
    .S1N(ConfigBits_N[270+1]),
    .X(J_NS4_BEG14)
);

 //switch matrix multiplexer J_NS4_BEG15 MUX-4
assign J_NS4_BEG15_input = {S4END3,S1END3,N4END3,N1END3};
cus_mux41_buf inst_cus_mux41_buf_J_NS4_BEG15 (
    .A0(J_NS4_BEG15_input[0]),
    .A1(J_NS4_BEG15_input[1]),
    .A2(J_NS4_BEG15_input[2]),
    .A3(J_NS4_BEG15_input[3]),
    .S0(ConfigBits[272+0]),
    .S0N(ConfigBits_N[272+0]),
    .S1(ConfigBits[272+1]),
    .S1N(ConfigBits_N[272+1]),
    .X(J_NS4_BEG15)
);

 //switch matrix multiplexer J_NS2_BEG0 MUX-4
assign J_NS2_BEG0_input = {S2END0,S2MID0,N2END0,N2MID0};
cus_mux41_buf inst_cus_mux41_buf_J_NS2_BEG0 (
    .A0(J_NS2_BEG0_input[0]),
    .A1(J_NS2_BEG0_input[1]),
    .A2(J_NS2_BEG0_input[2]),
    .A3(J_NS2_BEG0_input[3]),
    .S0(ConfigBits[274+0]),
    .S0N(ConfigBits_N[274+0]),
    .S1(ConfigBits[274+1]),
    .S1N(ConfigBits_N[274+1]),
    .X(J_NS2_BEG0)
);

 //switch matrix multiplexer J_NS2_BEG1 MUX-4
assign J_NS2_BEG1_input = {S2END1,S2MID1,N2END1,N2MID1};
cus_mux41_buf inst_cus_mux41_buf_J_NS2_BEG1 (
    .A0(J_NS2_BEG1_input[0]),
    .A1(J_NS2_BEG1_input[1]),
    .A2(J_NS2_BEG1_input[2]),
    .A3(J_NS2_BEG1_input[3]),
    .S0(ConfigBits[276+0]),
    .S0N(ConfigBits_N[276+0]),
    .S1(ConfigBits[276+1]),
    .S1N(ConfigBits_N[276+1]),
    .X(J_NS2_BEG1)
);

 //switch matrix multiplexer J_NS2_BEG2 MUX-4
assign J_NS2_BEG2_input = {S2END2,S2MID2,N2END2,N2MID2};
cus_mux41_buf inst_cus_mux41_buf_J_NS2_BEG2 (
    .A0(J_NS2_BEG2_input[0]),
    .A1(J_NS2_BEG2_input[1]),
    .A2(J_NS2_BEG2_input[2]),
    .A3(J_NS2_BEG2_input[3]),
    .S0(ConfigBits[278+0]),
    .S0N(ConfigBits_N[278+0]),
    .S1(ConfigBits[278+1]),
    .S1N(ConfigBits_N[278+1]),
    .X(J_NS2_BEG2)
);

 //switch matrix multiplexer J_NS2_BEG3 MUX-4
assign J_NS2_BEG3_input = {S2END3,S2MID3,N2END3,N2MID3};
cus_mux41_buf inst_cus_mux41_buf_J_NS2_BEG3 (
    .A0(J_NS2_BEG3_input[0]),
    .A1(J_NS2_BEG3_input[1]),
    .A2(J_NS2_BEG3_input[2]),
    .A3(J_NS2_BEG3_input[3]),
    .S0(ConfigBits[280+0]),
    .S0N(ConfigBits_N[280+0]),
    .S1(ConfigBits[280+1]),
    .S1N(ConfigBits_N[280+1]),
    .X(J_NS2_BEG3)
);

 //switch matrix multiplexer J_NS2_BEG4 MUX-4
assign J_NS2_BEG4_input = {S2END4,S2MID4,N2END4,N2MID4};
cus_mux41_buf inst_cus_mux41_buf_J_NS2_BEG4 (
    .A0(J_NS2_BEG4_input[0]),
    .A1(J_NS2_BEG4_input[1]),
    .A2(J_NS2_BEG4_input[2]),
    .A3(J_NS2_BEG4_input[3]),
    .S0(ConfigBits[282+0]),
    .S0N(ConfigBits_N[282+0]),
    .S1(ConfigBits[282+1]),
    .S1N(ConfigBits_N[282+1]),
    .X(J_NS2_BEG4)
);

 //switch matrix multiplexer J_NS2_BEG5 MUX-4
assign J_NS2_BEG5_input = {S2END5,S2MID5,N2END5,N2MID5};
cus_mux41_buf inst_cus_mux41_buf_J_NS2_BEG5 (
    .A0(J_NS2_BEG5_input[0]),
    .A1(J_NS2_BEG5_input[1]),
    .A2(J_NS2_BEG5_input[2]),
    .A3(J_NS2_BEG5_input[3]),
    .S0(ConfigBits[284+0]),
    .S0N(ConfigBits_N[284+0]),
    .S1(ConfigBits[284+1]),
    .S1N(ConfigBits_N[284+1]),
    .X(J_NS2_BEG5)
);

 //switch matrix multiplexer J_NS2_BEG6 MUX-4
assign J_NS2_BEG6_input = {S2END6,S2MID6,N2END6,N2MID6};
cus_mux41_buf inst_cus_mux41_buf_J_NS2_BEG6 (
    .A0(J_NS2_BEG6_input[0]),
    .A1(J_NS2_BEG6_input[1]),
    .A2(J_NS2_BEG6_input[2]),
    .A3(J_NS2_BEG6_input[3]),
    .S0(ConfigBits[286+0]),
    .S0N(ConfigBits_N[286+0]),
    .S1(ConfigBits[286+1]),
    .S1N(ConfigBits_N[286+1]),
    .X(J_NS2_BEG6)
);

 //switch matrix multiplexer J_NS2_BEG7 MUX-4
assign J_NS2_BEG7_input = {S2END7,S2MID7,N2END7,N2MID7};
cus_mux41_buf inst_cus_mux41_buf_J_NS2_BEG7 (
    .A0(J_NS2_BEG7_input[0]),
    .A1(J_NS2_BEG7_input[1]),
    .A2(J_NS2_BEG7_input[2]),
    .A3(J_NS2_BEG7_input[3]),
    .S0(ConfigBits[288+0]),
    .S0N(ConfigBits_N[288+0]),
    .S1(ConfigBits[288+1]),
    .S1N(ConfigBits_N[288+1]),
    .X(J_NS2_BEG7)
);

 //switch matrix multiplexer J_NS1_BEG0 MUX-4
assign J_NS1_BEG0_input = {GND0,S1END0,W6END0,N1END0};
cus_mux41_buf inst_cus_mux41_buf_J_NS1_BEG0 (
    .A0(J_NS1_BEG0_input[0]),
    .A1(J_NS1_BEG0_input[1]),
    .A2(J_NS1_BEG0_input[2]),
    .A3(J_NS1_BEG0_input[3]),
    .S0(ConfigBits[290+0]),
    .S0N(ConfigBits_N[290+0]),
    .S1(ConfigBits[290+1]),
    .S1N(ConfigBits_N[290+1]),
    .X(J_NS1_BEG0)
);

 //switch matrix multiplexer J_NS1_BEG1 MUX-4
assign J_NS1_BEG1_input = {GND0,S1END1,W6END1,N1END1};
cus_mux41_buf inst_cus_mux41_buf_J_NS1_BEG1 (
    .A0(J_NS1_BEG1_input[0]),
    .A1(J_NS1_BEG1_input[1]),
    .A2(J_NS1_BEG1_input[2]),
    .A3(J_NS1_BEG1_input[3]),
    .S0(ConfigBits[292+0]),
    .S0N(ConfigBits_N[292+0]),
    .S1(ConfigBits[292+1]),
    .S1N(ConfigBits_N[292+1]),
    .X(J_NS1_BEG1)
);

 //switch matrix multiplexer J_NS1_BEG2 MUX-4
assign J_NS1_BEG2_input = {GND0,S1END2,W6END2,N1END2};
cus_mux41_buf inst_cus_mux41_buf_J_NS1_BEG2 (
    .A0(J_NS1_BEG2_input[0]),
    .A1(J_NS1_BEG2_input[1]),
    .A2(J_NS1_BEG2_input[2]),
    .A3(J_NS1_BEG2_input[3]),
    .S0(ConfigBits[294+0]),
    .S0N(ConfigBits_N[294+0]),
    .S1(ConfigBits[294+1]),
    .S1N(ConfigBits_N[294+1]),
    .X(J_NS1_BEG2)
);

 //switch matrix multiplexer J_NS1_BEG3 MUX-4
assign J_NS1_BEG3_input = {GND0,S1END3,W6END3,N1END3};
cus_mux41_buf inst_cus_mux41_buf_J_NS1_BEG3 (
    .A0(J_NS1_BEG3_input[0]),
    .A1(J_NS1_BEG3_input[1]),
    .A2(J_NS1_BEG3_input[2]),
    .A3(J_NS1_BEG3_input[3]),
    .S0(ConfigBits[296+0]),
    .S0N(ConfigBits_N[296+0]),
    .S1(ConfigBits[296+1]),
    .S1N(ConfigBits_N[296+1]),
    .X(J_NS1_BEG3)
);

endmodule