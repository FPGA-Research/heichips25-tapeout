module heichips25_example_small (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net25;

 sg13g2_and2_1 _29_ (.A(net1),
    .B(net9),
    .X(_00_));
 sg13g2_and2_1 _30_ (.A(net2),
    .B(net10),
    .X(_01_));
 sg13g2_xor2_1 _31_ (.B(net10),
    .A(net2),
    .X(_02_));
 sg13g2_xor2_1 _32_ (.B(_02_),
    .A(_00_),
    .X(net18));
 sg13g2_a21oi_2 _33_ (.B1(_01_),
    .Y(_03_),
    .A2(_02_),
    .A1(_00_));
 sg13g2_and2_1 _34_ (.A(net3),
    .B(net11),
    .X(_04_));
 sg13g2_xnor2_1 _35_ (.Y(_05_),
    .A(net3),
    .B(net11));
 sg13g2_nor2_1 _36_ (.A(_03_),
    .B(_05_),
    .Y(_06_));
 sg13g2_xor2_1 _37_ (.B(_05_),
    .A(_03_),
    .X(net19));
 sg13g2_or2_1 _38_ (.X(_07_),
    .B(net12),
    .A(net4));
 sg13g2_and2_1 _39_ (.A(net4),
    .B(net12),
    .X(_08_));
 sg13g2_xor2_1 _40_ (.B(net12),
    .A(net4),
    .X(_09_));
 sg13g2_nor2_1 _41_ (.A(_04_),
    .B(_06_),
    .Y(_10_));
 sg13g2_xnor2_1 _42_ (.Y(net20),
    .A(_09_),
    .B(_10_));
 sg13g2_nand2b_1 _43_ (.Y(_11_),
    .B(_09_),
    .A_N(_05_));
 sg13g2_a21oi_1 _44_ (.A1(_04_),
    .A2(_07_),
    .Y(_12_),
    .B1(_08_));
 sg13g2_o21ai_1 _45_ (.B1(_12_),
    .Y(_13_),
    .A1(_03_),
    .A2(_11_));
 sg13g2_nand2_1 _46_ (.Y(_14_),
    .A(net5),
    .B(net13));
 sg13g2_xor2_1 _47_ (.B(net13),
    .A(net5),
    .X(_15_));
 sg13g2_inv_1 _48_ (.Y(_16_),
    .A(_15_));
 sg13g2_nand2_1 _49_ (.Y(_17_),
    .A(_13_),
    .B(_15_));
 sg13g2_xnor2_1 _50_ (.Y(net21),
    .A(_13_),
    .B(_16_));
 sg13g2_nor2_1 _51_ (.A(net6),
    .B(net14),
    .Y(_18_));
 sg13g2_xnor2_1 _52_ (.Y(_19_),
    .A(net6),
    .B(net14));
 sg13g2_nand2_1 _53_ (.Y(_20_),
    .A(_14_),
    .B(_17_));
 sg13g2_xnor2_1 _54_ (.Y(net22),
    .A(_19_),
    .B(_20_));
 sg13g2_nor2_1 _55_ (.A(_16_),
    .B(_19_),
    .Y(_21_));
 sg13g2_nor2_1 _56_ (.A(_14_),
    .B(_18_),
    .Y(_22_));
 sg13g2_a221oi_1 _57_ (.B2(_21_),
    .C1(_22_),
    .B1(_13_),
    .A1(net6),
    .Y(_23_),
    .A2(net14));
 sg13g2_nand2_1 _58_ (.Y(_24_),
    .A(net7),
    .B(net15));
 sg13g2_nor2_1 _59_ (.A(net7),
    .B(net15),
    .Y(_25_));
 sg13g2_xor2_1 _60_ (.B(net15),
    .A(net7),
    .X(_26_));
 sg13g2_xnor2_1 _61_ (.Y(net23),
    .A(_23_),
    .B(_26_));
 sg13g2_o21ai_1 _62_ (.B1(_24_),
    .Y(_27_),
    .A1(_23_),
    .A2(_25_));
 sg13g2_xnor2_1 _63_ (.Y(_28_),
    .A(net8),
    .B(net16));
 sg13g2_xnor2_1 _64_ (.Y(net24),
    .A(_27_),
    .B(_28_));
 sg13g2_xor2_1 _65_ (.B(net9),
    .A(net1),
    .X(net17));
 sg13g2_tielo heichips25_example_small_26 (.L_LO(net26));
 sg13g2_tielo heichips25_example_small_27 (.L_LO(net27));
 sg13g2_tielo heichips25_example_small_28 (.L_LO(net28));
 sg13g2_tielo heichips25_example_small_29 (.L_LO(net29));
 sg13g2_tielo heichips25_example_small_30 (.L_LO(net30));
 sg13g2_tielo heichips25_example_small_31 (.L_LO(net31));
 sg13g2_tielo heichips25_example_small_32 (.L_LO(net32));
 sg13g2_tielo heichips25_example_small_33 (.L_LO(net33));
 sg13g2_tielo heichips25_example_small_34 (.L_LO(net34));
 sg13g2_tielo heichips25_example_small_35 (.L_LO(net35));
 sg13g2_tielo heichips25_example_small_36 (.L_LO(net36));
 sg13g2_tielo heichips25_example_small_37 (.L_LO(net37));
 sg13g2_tielo heichips25_example_small_38 (.L_LO(net38));
 sg13g2_tielo heichips25_example_small_39 (.L_LO(net39));
 sg13g2_tielo heichips25_example_small_40 (.L_LO(net40));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[4]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[5]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(uio_in[6]),
    .X(net15));
 sg13g2_buf_1 input16 (.A(uio_in[7]),
    .X(net16));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[0]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[1]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[2]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[3]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[4]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[5]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[6]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[7]));
 sg13g2_tielo heichips25_example_small_25 (.L_LO(net25));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_decap_8 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_0_868 ();
 sg13g2_decap_8 FILLER_0_875 ();
 sg13g2_decap_8 FILLER_0_882 ();
 sg13g2_decap_8 FILLER_0_889 ();
 sg13g2_decap_8 FILLER_0_896 ();
 sg13g2_decap_8 FILLER_0_903 ();
 sg13g2_decap_8 FILLER_0_910 ();
 sg13g2_decap_8 FILLER_0_917 ();
 sg13g2_decap_8 FILLER_0_924 ();
 sg13g2_decap_8 FILLER_0_931 ();
 sg13g2_decap_8 FILLER_0_938 ();
 sg13g2_decap_8 FILLER_0_945 ();
 sg13g2_decap_8 FILLER_0_952 ();
 sg13g2_decap_8 FILLER_0_959 ();
 sg13g2_decap_8 FILLER_0_966 ();
 sg13g2_decap_8 FILLER_0_973 ();
 sg13g2_decap_8 FILLER_0_980 ();
 sg13g2_decap_8 FILLER_0_987 ();
 sg13g2_decap_8 FILLER_0_994 ();
 sg13g2_decap_8 FILLER_0_1001 ();
 sg13g2_decap_8 FILLER_0_1008 ();
 sg13g2_decap_8 FILLER_0_1015 ();
 sg13g2_decap_8 FILLER_0_1022 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_decap_8 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_1_868 ();
 sg13g2_decap_8 FILLER_1_875 ();
 sg13g2_decap_8 FILLER_1_882 ();
 sg13g2_decap_8 FILLER_1_889 ();
 sg13g2_decap_8 FILLER_1_896 ();
 sg13g2_decap_8 FILLER_1_903 ();
 sg13g2_decap_8 FILLER_1_910 ();
 sg13g2_decap_8 FILLER_1_917 ();
 sg13g2_decap_8 FILLER_1_924 ();
 sg13g2_decap_8 FILLER_1_931 ();
 sg13g2_decap_8 FILLER_1_938 ();
 sg13g2_decap_8 FILLER_1_945 ();
 sg13g2_decap_8 FILLER_1_952 ();
 sg13g2_decap_8 FILLER_1_959 ();
 sg13g2_decap_8 FILLER_1_966 ();
 sg13g2_decap_8 FILLER_1_973 ();
 sg13g2_decap_8 FILLER_1_980 ();
 sg13g2_decap_8 FILLER_1_987 ();
 sg13g2_decap_8 FILLER_1_994 ();
 sg13g2_decap_8 FILLER_1_1001 ();
 sg13g2_decap_8 FILLER_1_1008 ();
 sg13g2_decap_8 FILLER_1_1015 ();
 sg13g2_decap_8 FILLER_1_1022 ();
 sg13g2_decap_8 FILLER_2_4 ();
 sg13g2_decap_8 FILLER_2_11 ();
 sg13g2_decap_8 FILLER_2_18 ();
 sg13g2_decap_8 FILLER_2_25 ();
 sg13g2_decap_8 FILLER_2_32 ();
 sg13g2_decap_8 FILLER_2_39 ();
 sg13g2_decap_8 FILLER_2_46 ();
 sg13g2_decap_8 FILLER_2_53 ();
 sg13g2_decap_8 FILLER_2_60 ();
 sg13g2_decap_8 FILLER_2_67 ();
 sg13g2_decap_8 FILLER_2_74 ();
 sg13g2_decap_8 FILLER_2_81 ();
 sg13g2_decap_8 FILLER_2_88 ();
 sg13g2_decap_8 FILLER_2_95 ();
 sg13g2_decap_8 FILLER_2_102 ();
 sg13g2_decap_8 FILLER_2_109 ();
 sg13g2_decap_8 FILLER_2_116 ();
 sg13g2_decap_8 FILLER_2_123 ();
 sg13g2_decap_8 FILLER_2_130 ();
 sg13g2_decap_8 FILLER_2_137 ();
 sg13g2_decap_8 FILLER_2_144 ();
 sg13g2_decap_8 FILLER_2_151 ();
 sg13g2_decap_8 FILLER_2_158 ();
 sg13g2_decap_8 FILLER_2_165 ();
 sg13g2_decap_8 FILLER_2_172 ();
 sg13g2_decap_8 FILLER_2_179 ();
 sg13g2_decap_8 FILLER_2_186 ();
 sg13g2_decap_8 FILLER_2_193 ();
 sg13g2_decap_8 FILLER_2_200 ();
 sg13g2_decap_8 FILLER_2_207 ();
 sg13g2_decap_8 FILLER_2_214 ();
 sg13g2_decap_8 FILLER_2_221 ();
 sg13g2_decap_8 FILLER_2_228 ();
 sg13g2_decap_8 FILLER_2_235 ();
 sg13g2_decap_8 FILLER_2_242 ();
 sg13g2_decap_8 FILLER_2_249 ();
 sg13g2_decap_8 FILLER_2_256 ();
 sg13g2_decap_8 FILLER_2_263 ();
 sg13g2_decap_8 FILLER_2_270 ();
 sg13g2_decap_8 FILLER_2_277 ();
 sg13g2_decap_8 FILLER_2_284 ();
 sg13g2_decap_8 FILLER_2_291 ();
 sg13g2_decap_8 FILLER_2_298 ();
 sg13g2_decap_8 FILLER_2_305 ();
 sg13g2_decap_8 FILLER_2_312 ();
 sg13g2_decap_8 FILLER_2_319 ();
 sg13g2_decap_8 FILLER_2_326 ();
 sg13g2_decap_8 FILLER_2_333 ();
 sg13g2_decap_8 FILLER_2_340 ();
 sg13g2_decap_8 FILLER_2_347 ();
 sg13g2_decap_8 FILLER_2_354 ();
 sg13g2_decap_8 FILLER_2_361 ();
 sg13g2_decap_8 FILLER_2_368 ();
 sg13g2_decap_8 FILLER_2_375 ();
 sg13g2_decap_8 FILLER_2_382 ();
 sg13g2_decap_8 FILLER_2_389 ();
 sg13g2_decap_8 FILLER_2_396 ();
 sg13g2_decap_8 FILLER_2_403 ();
 sg13g2_decap_8 FILLER_2_410 ();
 sg13g2_decap_8 FILLER_2_417 ();
 sg13g2_decap_8 FILLER_2_424 ();
 sg13g2_decap_8 FILLER_2_431 ();
 sg13g2_decap_8 FILLER_2_438 ();
 sg13g2_decap_8 FILLER_2_445 ();
 sg13g2_decap_8 FILLER_2_452 ();
 sg13g2_decap_8 FILLER_2_459 ();
 sg13g2_decap_8 FILLER_2_466 ();
 sg13g2_decap_8 FILLER_2_473 ();
 sg13g2_decap_8 FILLER_2_480 ();
 sg13g2_decap_8 FILLER_2_487 ();
 sg13g2_decap_8 FILLER_2_494 ();
 sg13g2_decap_8 FILLER_2_501 ();
 sg13g2_decap_8 FILLER_2_508 ();
 sg13g2_decap_8 FILLER_2_515 ();
 sg13g2_decap_8 FILLER_2_522 ();
 sg13g2_decap_8 FILLER_2_529 ();
 sg13g2_decap_8 FILLER_2_536 ();
 sg13g2_decap_8 FILLER_2_543 ();
 sg13g2_decap_8 FILLER_2_550 ();
 sg13g2_decap_8 FILLER_2_557 ();
 sg13g2_decap_8 FILLER_2_564 ();
 sg13g2_decap_8 FILLER_2_571 ();
 sg13g2_decap_8 FILLER_2_578 ();
 sg13g2_decap_8 FILLER_2_585 ();
 sg13g2_decap_8 FILLER_2_592 ();
 sg13g2_decap_8 FILLER_2_599 ();
 sg13g2_decap_8 FILLER_2_606 ();
 sg13g2_decap_8 FILLER_2_613 ();
 sg13g2_decap_8 FILLER_2_620 ();
 sg13g2_decap_8 FILLER_2_627 ();
 sg13g2_decap_8 FILLER_2_634 ();
 sg13g2_decap_8 FILLER_2_641 ();
 sg13g2_decap_8 FILLER_2_648 ();
 sg13g2_decap_8 FILLER_2_655 ();
 sg13g2_decap_8 FILLER_2_662 ();
 sg13g2_decap_8 FILLER_2_669 ();
 sg13g2_decap_8 FILLER_2_676 ();
 sg13g2_decap_8 FILLER_2_683 ();
 sg13g2_decap_8 FILLER_2_690 ();
 sg13g2_decap_8 FILLER_2_697 ();
 sg13g2_decap_8 FILLER_2_704 ();
 sg13g2_decap_8 FILLER_2_711 ();
 sg13g2_decap_8 FILLER_2_718 ();
 sg13g2_decap_8 FILLER_2_725 ();
 sg13g2_decap_8 FILLER_2_732 ();
 sg13g2_decap_8 FILLER_2_739 ();
 sg13g2_decap_8 FILLER_2_746 ();
 sg13g2_decap_8 FILLER_2_753 ();
 sg13g2_decap_8 FILLER_2_760 ();
 sg13g2_decap_8 FILLER_2_767 ();
 sg13g2_decap_8 FILLER_2_774 ();
 sg13g2_decap_8 FILLER_2_781 ();
 sg13g2_decap_8 FILLER_2_788 ();
 sg13g2_decap_8 FILLER_2_795 ();
 sg13g2_decap_8 FILLER_2_802 ();
 sg13g2_decap_8 FILLER_2_809 ();
 sg13g2_decap_8 FILLER_2_816 ();
 sg13g2_decap_8 FILLER_2_823 ();
 sg13g2_decap_8 FILLER_2_830 ();
 sg13g2_decap_8 FILLER_2_837 ();
 sg13g2_decap_8 FILLER_2_844 ();
 sg13g2_decap_8 FILLER_2_851 ();
 sg13g2_decap_8 FILLER_2_858 ();
 sg13g2_decap_8 FILLER_2_865 ();
 sg13g2_decap_8 FILLER_2_872 ();
 sg13g2_decap_8 FILLER_2_879 ();
 sg13g2_decap_8 FILLER_2_886 ();
 sg13g2_decap_8 FILLER_2_893 ();
 sg13g2_decap_8 FILLER_2_900 ();
 sg13g2_decap_8 FILLER_2_907 ();
 sg13g2_decap_8 FILLER_2_914 ();
 sg13g2_decap_8 FILLER_2_921 ();
 sg13g2_decap_8 FILLER_2_928 ();
 sg13g2_decap_8 FILLER_2_935 ();
 sg13g2_decap_8 FILLER_2_942 ();
 sg13g2_decap_8 FILLER_2_949 ();
 sg13g2_decap_8 FILLER_2_956 ();
 sg13g2_decap_8 FILLER_2_963 ();
 sg13g2_decap_8 FILLER_2_970 ();
 sg13g2_decap_8 FILLER_2_977 ();
 sg13g2_decap_8 FILLER_2_984 ();
 sg13g2_decap_8 FILLER_2_991 ();
 sg13g2_decap_8 FILLER_2_998 ();
 sg13g2_decap_8 FILLER_2_1005 ();
 sg13g2_decap_8 FILLER_2_1012 ();
 sg13g2_decap_8 FILLER_2_1019 ();
 sg13g2_fill_2 FILLER_2_1026 ();
 sg13g2_fill_1 FILLER_2_1028 ();
 sg13g2_decap_8 FILLER_3_4 ();
 sg13g2_decap_8 FILLER_3_11 ();
 sg13g2_decap_8 FILLER_3_18 ();
 sg13g2_decap_8 FILLER_3_25 ();
 sg13g2_decap_8 FILLER_3_32 ();
 sg13g2_decap_8 FILLER_3_39 ();
 sg13g2_decap_8 FILLER_3_46 ();
 sg13g2_decap_8 FILLER_3_53 ();
 sg13g2_decap_8 FILLER_3_60 ();
 sg13g2_decap_8 FILLER_3_67 ();
 sg13g2_decap_8 FILLER_3_74 ();
 sg13g2_decap_8 FILLER_3_81 ();
 sg13g2_decap_8 FILLER_3_88 ();
 sg13g2_decap_8 FILLER_3_95 ();
 sg13g2_decap_8 FILLER_3_102 ();
 sg13g2_decap_8 FILLER_3_109 ();
 sg13g2_decap_8 FILLER_3_116 ();
 sg13g2_decap_8 FILLER_3_123 ();
 sg13g2_decap_8 FILLER_3_130 ();
 sg13g2_decap_8 FILLER_3_137 ();
 sg13g2_decap_8 FILLER_3_144 ();
 sg13g2_decap_8 FILLER_3_151 ();
 sg13g2_decap_8 FILLER_3_158 ();
 sg13g2_decap_8 FILLER_3_165 ();
 sg13g2_decap_8 FILLER_3_172 ();
 sg13g2_decap_8 FILLER_3_179 ();
 sg13g2_decap_8 FILLER_3_186 ();
 sg13g2_decap_8 FILLER_3_193 ();
 sg13g2_decap_8 FILLER_3_200 ();
 sg13g2_decap_8 FILLER_3_207 ();
 sg13g2_decap_8 FILLER_3_214 ();
 sg13g2_decap_8 FILLER_3_221 ();
 sg13g2_decap_8 FILLER_3_228 ();
 sg13g2_decap_8 FILLER_3_235 ();
 sg13g2_decap_8 FILLER_3_242 ();
 sg13g2_decap_8 FILLER_3_249 ();
 sg13g2_decap_8 FILLER_3_256 ();
 sg13g2_decap_8 FILLER_3_263 ();
 sg13g2_decap_8 FILLER_3_270 ();
 sg13g2_decap_8 FILLER_3_277 ();
 sg13g2_decap_8 FILLER_3_284 ();
 sg13g2_decap_8 FILLER_3_291 ();
 sg13g2_decap_8 FILLER_3_298 ();
 sg13g2_decap_8 FILLER_3_305 ();
 sg13g2_decap_8 FILLER_3_312 ();
 sg13g2_decap_8 FILLER_3_319 ();
 sg13g2_decap_8 FILLER_3_326 ();
 sg13g2_decap_8 FILLER_3_333 ();
 sg13g2_decap_8 FILLER_3_340 ();
 sg13g2_decap_8 FILLER_3_347 ();
 sg13g2_decap_8 FILLER_3_354 ();
 sg13g2_decap_8 FILLER_3_361 ();
 sg13g2_decap_8 FILLER_3_368 ();
 sg13g2_decap_8 FILLER_3_375 ();
 sg13g2_decap_8 FILLER_3_382 ();
 sg13g2_decap_8 FILLER_3_389 ();
 sg13g2_decap_8 FILLER_3_396 ();
 sg13g2_decap_8 FILLER_3_403 ();
 sg13g2_decap_8 FILLER_3_410 ();
 sg13g2_decap_8 FILLER_3_417 ();
 sg13g2_decap_8 FILLER_3_424 ();
 sg13g2_decap_8 FILLER_3_431 ();
 sg13g2_decap_8 FILLER_3_438 ();
 sg13g2_decap_8 FILLER_3_445 ();
 sg13g2_decap_8 FILLER_3_452 ();
 sg13g2_decap_8 FILLER_3_459 ();
 sg13g2_decap_8 FILLER_3_466 ();
 sg13g2_decap_8 FILLER_3_473 ();
 sg13g2_decap_8 FILLER_3_480 ();
 sg13g2_decap_8 FILLER_3_487 ();
 sg13g2_decap_8 FILLER_3_494 ();
 sg13g2_decap_8 FILLER_3_501 ();
 sg13g2_decap_8 FILLER_3_508 ();
 sg13g2_decap_8 FILLER_3_515 ();
 sg13g2_decap_8 FILLER_3_522 ();
 sg13g2_decap_8 FILLER_3_529 ();
 sg13g2_decap_8 FILLER_3_536 ();
 sg13g2_decap_8 FILLER_3_543 ();
 sg13g2_decap_8 FILLER_3_550 ();
 sg13g2_decap_8 FILLER_3_557 ();
 sg13g2_decap_8 FILLER_3_564 ();
 sg13g2_decap_8 FILLER_3_571 ();
 sg13g2_decap_8 FILLER_3_578 ();
 sg13g2_decap_8 FILLER_3_585 ();
 sg13g2_decap_8 FILLER_3_592 ();
 sg13g2_decap_8 FILLER_3_599 ();
 sg13g2_decap_8 FILLER_3_606 ();
 sg13g2_decap_8 FILLER_3_613 ();
 sg13g2_decap_8 FILLER_3_620 ();
 sg13g2_decap_8 FILLER_3_627 ();
 sg13g2_decap_8 FILLER_3_634 ();
 sg13g2_decap_8 FILLER_3_641 ();
 sg13g2_decap_8 FILLER_3_648 ();
 sg13g2_decap_8 FILLER_3_655 ();
 sg13g2_decap_8 FILLER_3_662 ();
 sg13g2_decap_8 FILLER_3_669 ();
 sg13g2_decap_8 FILLER_3_676 ();
 sg13g2_decap_8 FILLER_3_683 ();
 sg13g2_decap_8 FILLER_3_690 ();
 sg13g2_decap_8 FILLER_3_697 ();
 sg13g2_decap_8 FILLER_3_704 ();
 sg13g2_decap_8 FILLER_3_711 ();
 sg13g2_decap_8 FILLER_3_718 ();
 sg13g2_decap_8 FILLER_3_725 ();
 sg13g2_decap_8 FILLER_3_732 ();
 sg13g2_decap_8 FILLER_3_739 ();
 sg13g2_decap_8 FILLER_3_746 ();
 sg13g2_decap_8 FILLER_3_753 ();
 sg13g2_decap_8 FILLER_3_760 ();
 sg13g2_decap_8 FILLER_3_767 ();
 sg13g2_decap_8 FILLER_3_774 ();
 sg13g2_decap_8 FILLER_3_781 ();
 sg13g2_decap_8 FILLER_3_788 ();
 sg13g2_decap_8 FILLER_3_795 ();
 sg13g2_decap_8 FILLER_3_802 ();
 sg13g2_decap_8 FILLER_3_809 ();
 sg13g2_decap_8 FILLER_3_816 ();
 sg13g2_decap_8 FILLER_3_823 ();
 sg13g2_decap_8 FILLER_3_830 ();
 sg13g2_decap_8 FILLER_3_837 ();
 sg13g2_decap_8 FILLER_3_844 ();
 sg13g2_decap_8 FILLER_3_851 ();
 sg13g2_decap_8 FILLER_3_858 ();
 sg13g2_decap_8 FILLER_3_865 ();
 sg13g2_decap_8 FILLER_3_872 ();
 sg13g2_decap_8 FILLER_3_879 ();
 sg13g2_decap_8 FILLER_3_886 ();
 sg13g2_decap_8 FILLER_3_893 ();
 sg13g2_decap_8 FILLER_3_900 ();
 sg13g2_decap_8 FILLER_3_907 ();
 sg13g2_decap_8 FILLER_3_914 ();
 sg13g2_decap_8 FILLER_3_921 ();
 sg13g2_decap_8 FILLER_3_928 ();
 sg13g2_decap_8 FILLER_3_935 ();
 sg13g2_decap_8 FILLER_3_942 ();
 sg13g2_decap_8 FILLER_3_949 ();
 sg13g2_decap_8 FILLER_3_956 ();
 sg13g2_decap_8 FILLER_3_963 ();
 sg13g2_decap_8 FILLER_3_970 ();
 sg13g2_decap_8 FILLER_3_977 ();
 sg13g2_decap_8 FILLER_3_984 ();
 sg13g2_decap_8 FILLER_3_991 ();
 sg13g2_decap_8 FILLER_3_998 ();
 sg13g2_decap_8 FILLER_3_1005 ();
 sg13g2_decap_8 FILLER_3_1012 ();
 sg13g2_decap_8 FILLER_3_1019 ();
 sg13g2_fill_2 FILLER_3_1026 ();
 sg13g2_fill_1 FILLER_3_1028 ();
 sg13g2_decap_8 FILLER_4_4 ();
 sg13g2_decap_8 FILLER_4_11 ();
 sg13g2_decap_8 FILLER_4_18 ();
 sg13g2_decap_8 FILLER_4_25 ();
 sg13g2_decap_8 FILLER_4_32 ();
 sg13g2_decap_8 FILLER_4_39 ();
 sg13g2_decap_8 FILLER_4_46 ();
 sg13g2_decap_8 FILLER_4_53 ();
 sg13g2_decap_8 FILLER_4_60 ();
 sg13g2_decap_8 FILLER_4_67 ();
 sg13g2_decap_8 FILLER_4_74 ();
 sg13g2_decap_8 FILLER_4_81 ();
 sg13g2_decap_8 FILLER_4_88 ();
 sg13g2_decap_8 FILLER_4_95 ();
 sg13g2_decap_8 FILLER_4_102 ();
 sg13g2_decap_8 FILLER_4_109 ();
 sg13g2_decap_8 FILLER_4_116 ();
 sg13g2_decap_8 FILLER_4_123 ();
 sg13g2_decap_8 FILLER_4_130 ();
 sg13g2_decap_8 FILLER_4_137 ();
 sg13g2_decap_8 FILLER_4_144 ();
 sg13g2_decap_8 FILLER_4_151 ();
 sg13g2_decap_8 FILLER_4_158 ();
 sg13g2_decap_8 FILLER_4_165 ();
 sg13g2_decap_8 FILLER_4_172 ();
 sg13g2_decap_8 FILLER_4_179 ();
 sg13g2_decap_8 FILLER_4_186 ();
 sg13g2_decap_8 FILLER_4_193 ();
 sg13g2_decap_8 FILLER_4_200 ();
 sg13g2_decap_8 FILLER_4_207 ();
 sg13g2_decap_8 FILLER_4_214 ();
 sg13g2_decap_8 FILLER_4_221 ();
 sg13g2_decap_8 FILLER_4_228 ();
 sg13g2_decap_8 FILLER_4_235 ();
 sg13g2_decap_8 FILLER_4_242 ();
 sg13g2_decap_8 FILLER_4_249 ();
 sg13g2_decap_8 FILLER_4_256 ();
 sg13g2_decap_8 FILLER_4_263 ();
 sg13g2_decap_8 FILLER_4_270 ();
 sg13g2_decap_8 FILLER_4_277 ();
 sg13g2_decap_8 FILLER_4_284 ();
 sg13g2_decap_8 FILLER_4_291 ();
 sg13g2_decap_8 FILLER_4_298 ();
 sg13g2_decap_8 FILLER_4_305 ();
 sg13g2_decap_8 FILLER_4_312 ();
 sg13g2_decap_8 FILLER_4_319 ();
 sg13g2_decap_8 FILLER_4_326 ();
 sg13g2_decap_8 FILLER_4_333 ();
 sg13g2_decap_8 FILLER_4_340 ();
 sg13g2_decap_8 FILLER_4_347 ();
 sg13g2_decap_8 FILLER_4_354 ();
 sg13g2_decap_8 FILLER_4_361 ();
 sg13g2_decap_8 FILLER_4_368 ();
 sg13g2_decap_8 FILLER_4_375 ();
 sg13g2_decap_8 FILLER_4_382 ();
 sg13g2_decap_8 FILLER_4_389 ();
 sg13g2_decap_8 FILLER_4_396 ();
 sg13g2_decap_8 FILLER_4_403 ();
 sg13g2_decap_8 FILLER_4_410 ();
 sg13g2_decap_8 FILLER_4_417 ();
 sg13g2_decap_8 FILLER_4_424 ();
 sg13g2_decap_8 FILLER_4_431 ();
 sg13g2_decap_8 FILLER_4_438 ();
 sg13g2_decap_8 FILLER_4_445 ();
 sg13g2_decap_8 FILLER_4_452 ();
 sg13g2_decap_8 FILLER_4_459 ();
 sg13g2_decap_8 FILLER_4_466 ();
 sg13g2_decap_8 FILLER_4_473 ();
 sg13g2_decap_8 FILLER_4_480 ();
 sg13g2_decap_8 FILLER_4_487 ();
 sg13g2_decap_8 FILLER_4_494 ();
 sg13g2_decap_8 FILLER_4_501 ();
 sg13g2_decap_8 FILLER_4_508 ();
 sg13g2_decap_8 FILLER_4_515 ();
 sg13g2_decap_8 FILLER_4_522 ();
 sg13g2_decap_8 FILLER_4_529 ();
 sg13g2_decap_8 FILLER_4_536 ();
 sg13g2_decap_8 FILLER_4_543 ();
 sg13g2_decap_8 FILLER_4_550 ();
 sg13g2_decap_8 FILLER_4_557 ();
 sg13g2_decap_8 FILLER_4_564 ();
 sg13g2_decap_8 FILLER_4_571 ();
 sg13g2_decap_8 FILLER_4_578 ();
 sg13g2_decap_8 FILLER_4_585 ();
 sg13g2_decap_8 FILLER_4_592 ();
 sg13g2_decap_8 FILLER_4_599 ();
 sg13g2_decap_8 FILLER_4_606 ();
 sg13g2_decap_8 FILLER_4_613 ();
 sg13g2_decap_8 FILLER_4_620 ();
 sg13g2_decap_8 FILLER_4_627 ();
 sg13g2_decap_8 FILLER_4_634 ();
 sg13g2_decap_8 FILLER_4_641 ();
 sg13g2_decap_8 FILLER_4_648 ();
 sg13g2_decap_8 FILLER_4_655 ();
 sg13g2_decap_8 FILLER_4_662 ();
 sg13g2_decap_8 FILLER_4_669 ();
 sg13g2_decap_8 FILLER_4_676 ();
 sg13g2_decap_8 FILLER_4_683 ();
 sg13g2_decap_8 FILLER_4_690 ();
 sg13g2_decap_8 FILLER_4_697 ();
 sg13g2_decap_8 FILLER_4_704 ();
 sg13g2_decap_8 FILLER_4_711 ();
 sg13g2_decap_8 FILLER_4_718 ();
 sg13g2_decap_8 FILLER_4_725 ();
 sg13g2_decap_8 FILLER_4_732 ();
 sg13g2_decap_8 FILLER_4_739 ();
 sg13g2_decap_8 FILLER_4_746 ();
 sg13g2_decap_8 FILLER_4_753 ();
 sg13g2_decap_8 FILLER_4_760 ();
 sg13g2_decap_8 FILLER_4_767 ();
 sg13g2_decap_8 FILLER_4_774 ();
 sg13g2_decap_8 FILLER_4_781 ();
 sg13g2_decap_8 FILLER_4_788 ();
 sg13g2_decap_8 FILLER_4_795 ();
 sg13g2_decap_8 FILLER_4_802 ();
 sg13g2_decap_8 FILLER_4_809 ();
 sg13g2_decap_8 FILLER_4_816 ();
 sg13g2_decap_8 FILLER_4_823 ();
 sg13g2_decap_8 FILLER_4_830 ();
 sg13g2_decap_8 FILLER_4_837 ();
 sg13g2_decap_8 FILLER_4_844 ();
 sg13g2_decap_8 FILLER_4_851 ();
 sg13g2_decap_8 FILLER_4_858 ();
 sg13g2_decap_8 FILLER_4_865 ();
 sg13g2_decap_8 FILLER_4_872 ();
 sg13g2_decap_8 FILLER_4_879 ();
 sg13g2_decap_8 FILLER_4_886 ();
 sg13g2_decap_8 FILLER_4_893 ();
 sg13g2_decap_8 FILLER_4_900 ();
 sg13g2_decap_8 FILLER_4_907 ();
 sg13g2_decap_8 FILLER_4_914 ();
 sg13g2_decap_8 FILLER_4_921 ();
 sg13g2_decap_8 FILLER_4_928 ();
 sg13g2_decap_8 FILLER_4_935 ();
 sg13g2_decap_8 FILLER_4_942 ();
 sg13g2_decap_8 FILLER_4_949 ();
 sg13g2_decap_8 FILLER_4_956 ();
 sg13g2_decap_8 FILLER_4_963 ();
 sg13g2_decap_8 FILLER_4_970 ();
 sg13g2_decap_8 FILLER_4_977 ();
 sg13g2_decap_8 FILLER_4_984 ();
 sg13g2_decap_8 FILLER_4_991 ();
 sg13g2_decap_8 FILLER_4_998 ();
 sg13g2_decap_8 FILLER_4_1005 ();
 sg13g2_decap_8 FILLER_4_1012 ();
 sg13g2_decap_8 FILLER_4_1019 ();
 sg13g2_fill_2 FILLER_4_1026 ();
 sg13g2_fill_1 FILLER_4_1028 ();
 sg13g2_decap_8 FILLER_5_4 ();
 sg13g2_decap_8 FILLER_5_11 ();
 sg13g2_decap_8 FILLER_5_18 ();
 sg13g2_decap_8 FILLER_5_25 ();
 sg13g2_decap_8 FILLER_5_32 ();
 sg13g2_decap_8 FILLER_5_39 ();
 sg13g2_decap_8 FILLER_5_46 ();
 sg13g2_decap_8 FILLER_5_53 ();
 sg13g2_decap_8 FILLER_5_60 ();
 sg13g2_decap_8 FILLER_5_67 ();
 sg13g2_decap_8 FILLER_5_74 ();
 sg13g2_decap_8 FILLER_5_81 ();
 sg13g2_decap_8 FILLER_5_88 ();
 sg13g2_decap_8 FILLER_5_95 ();
 sg13g2_decap_8 FILLER_5_102 ();
 sg13g2_decap_8 FILLER_5_109 ();
 sg13g2_decap_8 FILLER_5_116 ();
 sg13g2_decap_8 FILLER_5_123 ();
 sg13g2_decap_8 FILLER_5_130 ();
 sg13g2_decap_8 FILLER_5_137 ();
 sg13g2_decap_8 FILLER_5_144 ();
 sg13g2_decap_8 FILLER_5_151 ();
 sg13g2_decap_8 FILLER_5_158 ();
 sg13g2_decap_8 FILLER_5_165 ();
 sg13g2_decap_8 FILLER_5_172 ();
 sg13g2_decap_8 FILLER_5_179 ();
 sg13g2_decap_8 FILLER_5_186 ();
 sg13g2_decap_8 FILLER_5_193 ();
 sg13g2_decap_8 FILLER_5_200 ();
 sg13g2_decap_8 FILLER_5_207 ();
 sg13g2_decap_8 FILLER_5_214 ();
 sg13g2_decap_8 FILLER_5_221 ();
 sg13g2_decap_8 FILLER_5_228 ();
 sg13g2_decap_8 FILLER_5_235 ();
 sg13g2_decap_8 FILLER_5_242 ();
 sg13g2_decap_8 FILLER_5_249 ();
 sg13g2_decap_8 FILLER_5_256 ();
 sg13g2_decap_8 FILLER_5_263 ();
 sg13g2_decap_8 FILLER_5_270 ();
 sg13g2_decap_8 FILLER_5_277 ();
 sg13g2_decap_8 FILLER_5_284 ();
 sg13g2_decap_8 FILLER_5_291 ();
 sg13g2_decap_8 FILLER_5_298 ();
 sg13g2_decap_8 FILLER_5_305 ();
 sg13g2_decap_8 FILLER_5_312 ();
 sg13g2_decap_8 FILLER_5_319 ();
 sg13g2_decap_8 FILLER_5_326 ();
 sg13g2_decap_8 FILLER_5_333 ();
 sg13g2_decap_8 FILLER_5_340 ();
 sg13g2_decap_8 FILLER_5_347 ();
 sg13g2_decap_8 FILLER_5_354 ();
 sg13g2_decap_8 FILLER_5_361 ();
 sg13g2_decap_8 FILLER_5_368 ();
 sg13g2_decap_8 FILLER_5_375 ();
 sg13g2_decap_8 FILLER_5_382 ();
 sg13g2_decap_8 FILLER_5_389 ();
 sg13g2_decap_8 FILLER_5_396 ();
 sg13g2_decap_8 FILLER_5_403 ();
 sg13g2_decap_8 FILLER_5_410 ();
 sg13g2_decap_8 FILLER_5_417 ();
 sg13g2_decap_8 FILLER_5_424 ();
 sg13g2_decap_8 FILLER_5_431 ();
 sg13g2_decap_8 FILLER_5_438 ();
 sg13g2_decap_8 FILLER_5_445 ();
 sg13g2_decap_8 FILLER_5_452 ();
 sg13g2_decap_8 FILLER_5_459 ();
 sg13g2_decap_8 FILLER_5_466 ();
 sg13g2_decap_8 FILLER_5_473 ();
 sg13g2_decap_8 FILLER_5_480 ();
 sg13g2_decap_8 FILLER_5_487 ();
 sg13g2_decap_8 FILLER_5_494 ();
 sg13g2_decap_8 FILLER_5_501 ();
 sg13g2_decap_8 FILLER_5_508 ();
 sg13g2_decap_8 FILLER_5_515 ();
 sg13g2_decap_8 FILLER_5_522 ();
 sg13g2_decap_8 FILLER_5_529 ();
 sg13g2_decap_8 FILLER_5_536 ();
 sg13g2_decap_8 FILLER_5_543 ();
 sg13g2_decap_8 FILLER_5_550 ();
 sg13g2_decap_8 FILLER_5_557 ();
 sg13g2_decap_8 FILLER_5_564 ();
 sg13g2_decap_8 FILLER_5_571 ();
 sg13g2_decap_8 FILLER_5_578 ();
 sg13g2_decap_8 FILLER_5_585 ();
 sg13g2_decap_8 FILLER_5_592 ();
 sg13g2_decap_8 FILLER_5_599 ();
 sg13g2_decap_8 FILLER_5_606 ();
 sg13g2_decap_8 FILLER_5_613 ();
 sg13g2_decap_8 FILLER_5_620 ();
 sg13g2_decap_8 FILLER_5_627 ();
 sg13g2_decap_8 FILLER_5_634 ();
 sg13g2_decap_8 FILLER_5_641 ();
 sg13g2_decap_8 FILLER_5_648 ();
 sg13g2_decap_8 FILLER_5_655 ();
 sg13g2_decap_8 FILLER_5_662 ();
 sg13g2_decap_8 FILLER_5_669 ();
 sg13g2_decap_8 FILLER_5_676 ();
 sg13g2_decap_8 FILLER_5_683 ();
 sg13g2_decap_8 FILLER_5_690 ();
 sg13g2_decap_8 FILLER_5_697 ();
 sg13g2_decap_8 FILLER_5_704 ();
 sg13g2_decap_8 FILLER_5_711 ();
 sg13g2_decap_8 FILLER_5_718 ();
 sg13g2_decap_8 FILLER_5_725 ();
 sg13g2_decap_8 FILLER_5_732 ();
 sg13g2_decap_8 FILLER_5_739 ();
 sg13g2_decap_8 FILLER_5_746 ();
 sg13g2_decap_8 FILLER_5_753 ();
 sg13g2_decap_8 FILLER_5_760 ();
 sg13g2_decap_8 FILLER_5_767 ();
 sg13g2_decap_8 FILLER_5_774 ();
 sg13g2_decap_8 FILLER_5_781 ();
 sg13g2_decap_8 FILLER_5_788 ();
 sg13g2_decap_8 FILLER_5_795 ();
 sg13g2_decap_8 FILLER_5_802 ();
 sg13g2_decap_8 FILLER_5_809 ();
 sg13g2_decap_8 FILLER_5_816 ();
 sg13g2_decap_8 FILLER_5_823 ();
 sg13g2_decap_8 FILLER_5_830 ();
 sg13g2_decap_8 FILLER_5_837 ();
 sg13g2_decap_8 FILLER_5_844 ();
 sg13g2_decap_8 FILLER_5_851 ();
 sg13g2_decap_8 FILLER_5_858 ();
 sg13g2_decap_8 FILLER_5_865 ();
 sg13g2_decap_8 FILLER_5_872 ();
 sg13g2_decap_8 FILLER_5_879 ();
 sg13g2_decap_8 FILLER_5_886 ();
 sg13g2_decap_8 FILLER_5_893 ();
 sg13g2_decap_8 FILLER_5_900 ();
 sg13g2_decap_8 FILLER_5_907 ();
 sg13g2_decap_8 FILLER_5_914 ();
 sg13g2_decap_8 FILLER_5_921 ();
 sg13g2_decap_8 FILLER_5_928 ();
 sg13g2_decap_8 FILLER_5_935 ();
 sg13g2_decap_8 FILLER_5_942 ();
 sg13g2_decap_8 FILLER_5_949 ();
 sg13g2_decap_8 FILLER_5_956 ();
 sg13g2_decap_8 FILLER_5_963 ();
 sg13g2_decap_8 FILLER_5_970 ();
 sg13g2_decap_8 FILLER_5_977 ();
 sg13g2_decap_8 FILLER_5_984 ();
 sg13g2_decap_8 FILLER_5_991 ();
 sg13g2_decap_8 FILLER_5_998 ();
 sg13g2_decap_8 FILLER_5_1005 ();
 sg13g2_decap_8 FILLER_5_1012 ();
 sg13g2_decap_8 FILLER_5_1019 ();
 sg13g2_fill_2 FILLER_5_1026 ();
 sg13g2_fill_1 FILLER_5_1028 ();
 sg13g2_decap_8 FILLER_6_4 ();
 sg13g2_decap_8 FILLER_6_11 ();
 sg13g2_decap_8 FILLER_6_18 ();
 sg13g2_decap_8 FILLER_6_25 ();
 sg13g2_decap_8 FILLER_6_32 ();
 sg13g2_decap_8 FILLER_6_39 ();
 sg13g2_decap_8 FILLER_6_46 ();
 sg13g2_decap_8 FILLER_6_53 ();
 sg13g2_decap_8 FILLER_6_60 ();
 sg13g2_decap_8 FILLER_6_67 ();
 sg13g2_decap_8 FILLER_6_74 ();
 sg13g2_decap_8 FILLER_6_81 ();
 sg13g2_decap_8 FILLER_6_88 ();
 sg13g2_decap_8 FILLER_6_95 ();
 sg13g2_decap_8 FILLER_6_102 ();
 sg13g2_decap_8 FILLER_6_109 ();
 sg13g2_decap_8 FILLER_6_116 ();
 sg13g2_decap_8 FILLER_6_123 ();
 sg13g2_decap_8 FILLER_6_130 ();
 sg13g2_decap_8 FILLER_6_137 ();
 sg13g2_decap_8 FILLER_6_144 ();
 sg13g2_decap_8 FILLER_6_151 ();
 sg13g2_decap_8 FILLER_6_158 ();
 sg13g2_decap_8 FILLER_6_165 ();
 sg13g2_decap_8 FILLER_6_172 ();
 sg13g2_decap_8 FILLER_6_179 ();
 sg13g2_decap_8 FILLER_6_186 ();
 sg13g2_decap_8 FILLER_6_193 ();
 sg13g2_decap_8 FILLER_6_200 ();
 sg13g2_decap_8 FILLER_6_207 ();
 sg13g2_decap_8 FILLER_6_214 ();
 sg13g2_decap_8 FILLER_6_221 ();
 sg13g2_decap_8 FILLER_6_228 ();
 sg13g2_decap_8 FILLER_6_235 ();
 sg13g2_decap_8 FILLER_6_242 ();
 sg13g2_decap_8 FILLER_6_249 ();
 sg13g2_decap_8 FILLER_6_256 ();
 sg13g2_decap_8 FILLER_6_263 ();
 sg13g2_decap_8 FILLER_6_270 ();
 sg13g2_decap_8 FILLER_6_277 ();
 sg13g2_decap_8 FILLER_6_284 ();
 sg13g2_decap_8 FILLER_6_291 ();
 sg13g2_decap_8 FILLER_6_298 ();
 sg13g2_decap_8 FILLER_6_305 ();
 sg13g2_decap_8 FILLER_6_312 ();
 sg13g2_decap_8 FILLER_6_319 ();
 sg13g2_decap_8 FILLER_6_326 ();
 sg13g2_decap_8 FILLER_6_333 ();
 sg13g2_decap_8 FILLER_6_340 ();
 sg13g2_decap_8 FILLER_6_347 ();
 sg13g2_decap_8 FILLER_6_354 ();
 sg13g2_decap_8 FILLER_6_361 ();
 sg13g2_decap_8 FILLER_6_368 ();
 sg13g2_decap_8 FILLER_6_375 ();
 sg13g2_decap_8 FILLER_6_382 ();
 sg13g2_decap_8 FILLER_6_389 ();
 sg13g2_decap_8 FILLER_6_396 ();
 sg13g2_decap_8 FILLER_6_403 ();
 sg13g2_decap_8 FILLER_6_410 ();
 sg13g2_decap_8 FILLER_6_417 ();
 sg13g2_decap_8 FILLER_6_424 ();
 sg13g2_decap_8 FILLER_6_431 ();
 sg13g2_decap_8 FILLER_6_438 ();
 sg13g2_decap_8 FILLER_6_445 ();
 sg13g2_decap_8 FILLER_6_452 ();
 sg13g2_decap_8 FILLER_6_459 ();
 sg13g2_decap_8 FILLER_6_466 ();
 sg13g2_decap_8 FILLER_6_473 ();
 sg13g2_decap_8 FILLER_6_480 ();
 sg13g2_decap_8 FILLER_6_487 ();
 sg13g2_decap_8 FILLER_6_494 ();
 sg13g2_decap_8 FILLER_6_501 ();
 sg13g2_decap_8 FILLER_6_508 ();
 sg13g2_decap_8 FILLER_6_515 ();
 sg13g2_decap_8 FILLER_6_522 ();
 sg13g2_decap_8 FILLER_6_529 ();
 sg13g2_decap_8 FILLER_6_536 ();
 sg13g2_decap_8 FILLER_6_543 ();
 sg13g2_decap_8 FILLER_6_550 ();
 sg13g2_decap_8 FILLER_6_557 ();
 sg13g2_decap_8 FILLER_6_564 ();
 sg13g2_decap_8 FILLER_6_571 ();
 sg13g2_decap_8 FILLER_6_578 ();
 sg13g2_decap_8 FILLER_6_585 ();
 sg13g2_decap_8 FILLER_6_592 ();
 sg13g2_decap_8 FILLER_6_599 ();
 sg13g2_decap_8 FILLER_6_606 ();
 sg13g2_decap_8 FILLER_6_613 ();
 sg13g2_decap_8 FILLER_6_620 ();
 sg13g2_decap_8 FILLER_6_627 ();
 sg13g2_decap_8 FILLER_6_634 ();
 sg13g2_decap_8 FILLER_6_641 ();
 sg13g2_decap_8 FILLER_6_648 ();
 sg13g2_decap_8 FILLER_6_655 ();
 sg13g2_decap_8 FILLER_6_662 ();
 sg13g2_decap_8 FILLER_6_669 ();
 sg13g2_decap_8 FILLER_6_676 ();
 sg13g2_decap_8 FILLER_6_683 ();
 sg13g2_decap_8 FILLER_6_690 ();
 sg13g2_decap_8 FILLER_6_697 ();
 sg13g2_decap_8 FILLER_6_704 ();
 sg13g2_decap_8 FILLER_6_711 ();
 sg13g2_decap_8 FILLER_6_718 ();
 sg13g2_decap_8 FILLER_6_725 ();
 sg13g2_decap_8 FILLER_6_732 ();
 sg13g2_decap_8 FILLER_6_739 ();
 sg13g2_decap_8 FILLER_6_746 ();
 sg13g2_decap_8 FILLER_6_753 ();
 sg13g2_decap_8 FILLER_6_760 ();
 sg13g2_decap_8 FILLER_6_767 ();
 sg13g2_decap_8 FILLER_6_774 ();
 sg13g2_decap_8 FILLER_6_781 ();
 sg13g2_decap_8 FILLER_6_788 ();
 sg13g2_decap_8 FILLER_6_795 ();
 sg13g2_decap_8 FILLER_6_802 ();
 sg13g2_decap_8 FILLER_6_809 ();
 sg13g2_decap_8 FILLER_6_816 ();
 sg13g2_decap_8 FILLER_6_823 ();
 sg13g2_decap_8 FILLER_6_830 ();
 sg13g2_decap_8 FILLER_6_837 ();
 sg13g2_decap_8 FILLER_6_844 ();
 sg13g2_decap_8 FILLER_6_851 ();
 sg13g2_decap_8 FILLER_6_858 ();
 sg13g2_decap_8 FILLER_6_865 ();
 sg13g2_decap_8 FILLER_6_872 ();
 sg13g2_decap_8 FILLER_6_879 ();
 sg13g2_decap_8 FILLER_6_886 ();
 sg13g2_decap_8 FILLER_6_893 ();
 sg13g2_decap_8 FILLER_6_900 ();
 sg13g2_decap_8 FILLER_6_907 ();
 sg13g2_decap_8 FILLER_6_914 ();
 sg13g2_decap_8 FILLER_6_921 ();
 sg13g2_decap_8 FILLER_6_928 ();
 sg13g2_decap_8 FILLER_6_935 ();
 sg13g2_decap_8 FILLER_6_942 ();
 sg13g2_decap_8 FILLER_6_949 ();
 sg13g2_decap_8 FILLER_6_956 ();
 sg13g2_decap_8 FILLER_6_963 ();
 sg13g2_decap_8 FILLER_6_970 ();
 sg13g2_decap_8 FILLER_6_977 ();
 sg13g2_decap_8 FILLER_6_984 ();
 sg13g2_decap_8 FILLER_6_991 ();
 sg13g2_decap_8 FILLER_6_998 ();
 sg13g2_decap_8 FILLER_6_1005 ();
 sg13g2_decap_8 FILLER_6_1012 ();
 sg13g2_decap_8 FILLER_6_1019 ();
 sg13g2_fill_2 FILLER_6_1026 ();
 sg13g2_fill_1 FILLER_6_1028 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_decap_8 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_7_868 ();
 sg13g2_decap_8 FILLER_7_875 ();
 sg13g2_decap_8 FILLER_7_882 ();
 sg13g2_decap_8 FILLER_7_889 ();
 sg13g2_decap_8 FILLER_7_896 ();
 sg13g2_decap_8 FILLER_7_903 ();
 sg13g2_decap_8 FILLER_7_910 ();
 sg13g2_decap_8 FILLER_7_917 ();
 sg13g2_decap_8 FILLER_7_924 ();
 sg13g2_decap_8 FILLER_7_931 ();
 sg13g2_decap_8 FILLER_7_938 ();
 sg13g2_decap_8 FILLER_7_945 ();
 sg13g2_decap_8 FILLER_7_952 ();
 sg13g2_decap_8 FILLER_7_959 ();
 sg13g2_decap_8 FILLER_7_966 ();
 sg13g2_decap_8 FILLER_7_973 ();
 sg13g2_decap_8 FILLER_7_980 ();
 sg13g2_decap_8 FILLER_7_987 ();
 sg13g2_decap_8 FILLER_7_994 ();
 sg13g2_decap_8 FILLER_7_1001 ();
 sg13g2_decap_8 FILLER_7_1008 ();
 sg13g2_decap_8 FILLER_7_1015 ();
 sg13g2_decap_8 FILLER_7_1022 ();
 sg13g2_decap_8 FILLER_8_4 ();
 sg13g2_decap_8 FILLER_8_11 ();
 sg13g2_decap_8 FILLER_8_18 ();
 sg13g2_decap_8 FILLER_8_25 ();
 sg13g2_decap_8 FILLER_8_32 ();
 sg13g2_decap_8 FILLER_8_39 ();
 sg13g2_decap_8 FILLER_8_46 ();
 sg13g2_decap_8 FILLER_8_53 ();
 sg13g2_decap_8 FILLER_8_60 ();
 sg13g2_decap_8 FILLER_8_67 ();
 sg13g2_decap_8 FILLER_8_74 ();
 sg13g2_decap_8 FILLER_8_81 ();
 sg13g2_decap_8 FILLER_8_88 ();
 sg13g2_decap_8 FILLER_8_95 ();
 sg13g2_decap_8 FILLER_8_102 ();
 sg13g2_decap_8 FILLER_8_109 ();
 sg13g2_decap_8 FILLER_8_116 ();
 sg13g2_decap_8 FILLER_8_123 ();
 sg13g2_decap_8 FILLER_8_130 ();
 sg13g2_decap_8 FILLER_8_137 ();
 sg13g2_decap_8 FILLER_8_144 ();
 sg13g2_decap_8 FILLER_8_151 ();
 sg13g2_decap_8 FILLER_8_158 ();
 sg13g2_decap_8 FILLER_8_165 ();
 sg13g2_decap_8 FILLER_8_172 ();
 sg13g2_decap_8 FILLER_8_179 ();
 sg13g2_decap_8 FILLER_8_186 ();
 sg13g2_decap_8 FILLER_8_193 ();
 sg13g2_decap_8 FILLER_8_200 ();
 sg13g2_decap_8 FILLER_8_207 ();
 sg13g2_decap_8 FILLER_8_214 ();
 sg13g2_decap_8 FILLER_8_221 ();
 sg13g2_decap_8 FILLER_8_228 ();
 sg13g2_decap_8 FILLER_8_235 ();
 sg13g2_decap_8 FILLER_8_242 ();
 sg13g2_decap_8 FILLER_8_249 ();
 sg13g2_decap_8 FILLER_8_256 ();
 sg13g2_decap_8 FILLER_8_263 ();
 sg13g2_decap_8 FILLER_8_270 ();
 sg13g2_decap_8 FILLER_8_277 ();
 sg13g2_decap_8 FILLER_8_284 ();
 sg13g2_decap_8 FILLER_8_291 ();
 sg13g2_decap_8 FILLER_8_298 ();
 sg13g2_decap_8 FILLER_8_305 ();
 sg13g2_decap_8 FILLER_8_312 ();
 sg13g2_decap_8 FILLER_8_319 ();
 sg13g2_decap_8 FILLER_8_326 ();
 sg13g2_decap_8 FILLER_8_333 ();
 sg13g2_decap_8 FILLER_8_340 ();
 sg13g2_decap_8 FILLER_8_347 ();
 sg13g2_decap_8 FILLER_8_354 ();
 sg13g2_decap_8 FILLER_8_361 ();
 sg13g2_decap_8 FILLER_8_368 ();
 sg13g2_decap_8 FILLER_8_375 ();
 sg13g2_decap_8 FILLER_8_382 ();
 sg13g2_decap_8 FILLER_8_389 ();
 sg13g2_decap_8 FILLER_8_396 ();
 sg13g2_decap_8 FILLER_8_403 ();
 sg13g2_decap_8 FILLER_8_410 ();
 sg13g2_decap_8 FILLER_8_417 ();
 sg13g2_decap_8 FILLER_8_424 ();
 sg13g2_decap_8 FILLER_8_431 ();
 sg13g2_decap_8 FILLER_8_438 ();
 sg13g2_decap_8 FILLER_8_445 ();
 sg13g2_decap_8 FILLER_8_452 ();
 sg13g2_decap_8 FILLER_8_459 ();
 sg13g2_decap_8 FILLER_8_466 ();
 sg13g2_decap_8 FILLER_8_473 ();
 sg13g2_decap_8 FILLER_8_480 ();
 sg13g2_decap_8 FILLER_8_487 ();
 sg13g2_decap_8 FILLER_8_494 ();
 sg13g2_decap_8 FILLER_8_501 ();
 sg13g2_decap_8 FILLER_8_508 ();
 sg13g2_decap_8 FILLER_8_515 ();
 sg13g2_decap_8 FILLER_8_522 ();
 sg13g2_decap_8 FILLER_8_529 ();
 sg13g2_decap_8 FILLER_8_536 ();
 sg13g2_decap_8 FILLER_8_543 ();
 sg13g2_decap_8 FILLER_8_550 ();
 sg13g2_decap_8 FILLER_8_557 ();
 sg13g2_decap_8 FILLER_8_564 ();
 sg13g2_decap_8 FILLER_8_571 ();
 sg13g2_decap_8 FILLER_8_578 ();
 sg13g2_decap_8 FILLER_8_585 ();
 sg13g2_decap_8 FILLER_8_592 ();
 sg13g2_decap_8 FILLER_8_599 ();
 sg13g2_decap_8 FILLER_8_606 ();
 sg13g2_decap_8 FILLER_8_613 ();
 sg13g2_decap_8 FILLER_8_620 ();
 sg13g2_decap_8 FILLER_8_627 ();
 sg13g2_decap_8 FILLER_8_634 ();
 sg13g2_decap_8 FILLER_8_641 ();
 sg13g2_decap_8 FILLER_8_648 ();
 sg13g2_decap_8 FILLER_8_655 ();
 sg13g2_decap_8 FILLER_8_662 ();
 sg13g2_decap_8 FILLER_8_669 ();
 sg13g2_decap_8 FILLER_8_676 ();
 sg13g2_decap_8 FILLER_8_683 ();
 sg13g2_decap_8 FILLER_8_690 ();
 sg13g2_decap_8 FILLER_8_697 ();
 sg13g2_decap_8 FILLER_8_704 ();
 sg13g2_decap_8 FILLER_8_711 ();
 sg13g2_decap_8 FILLER_8_718 ();
 sg13g2_decap_8 FILLER_8_725 ();
 sg13g2_decap_8 FILLER_8_732 ();
 sg13g2_decap_8 FILLER_8_739 ();
 sg13g2_decap_8 FILLER_8_746 ();
 sg13g2_decap_8 FILLER_8_753 ();
 sg13g2_decap_8 FILLER_8_760 ();
 sg13g2_decap_8 FILLER_8_767 ();
 sg13g2_decap_8 FILLER_8_774 ();
 sg13g2_decap_8 FILLER_8_781 ();
 sg13g2_decap_8 FILLER_8_788 ();
 sg13g2_decap_8 FILLER_8_795 ();
 sg13g2_decap_8 FILLER_8_802 ();
 sg13g2_decap_8 FILLER_8_809 ();
 sg13g2_decap_8 FILLER_8_816 ();
 sg13g2_decap_8 FILLER_8_823 ();
 sg13g2_decap_8 FILLER_8_830 ();
 sg13g2_decap_8 FILLER_8_837 ();
 sg13g2_decap_8 FILLER_8_844 ();
 sg13g2_decap_8 FILLER_8_851 ();
 sg13g2_decap_8 FILLER_8_858 ();
 sg13g2_decap_8 FILLER_8_865 ();
 sg13g2_decap_8 FILLER_8_872 ();
 sg13g2_decap_8 FILLER_8_879 ();
 sg13g2_decap_8 FILLER_8_886 ();
 sg13g2_decap_8 FILLER_8_893 ();
 sg13g2_decap_8 FILLER_8_900 ();
 sg13g2_decap_8 FILLER_8_907 ();
 sg13g2_decap_8 FILLER_8_914 ();
 sg13g2_decap_8 FILLER_8_921 ();
 sg13g2_decap_8 FILLER_8_928 ();
 sg13g2_decap_8 FILLER_8_935 ();
 sg13g2_decap_8 FILLER_8_942 ();
 sg13g2_decap_8 FILLER_8_949 ();
 sg13g2_decap_8 FILLER_8_956 ();
 sg13g2_decap_8 FILLER_8_963 ();
 sg13g2_decap_8 FILLER_8_970 ();
 sg13g2_decap_8 FILLER_8_977 ();
 sg13g2_decap_8 FILLER_8_984 ();
 sg13g2_decap_8 FILLER_8_991 ();
 sg13g2_decap_8 FILLER_8_998 ();
 sg13g2_decap_8 FILLER_8_1005 ();
 sg13g2_decap_8 FILLER_8_1012 ();
 sg13g2_decap_8 FILLER_8_1019 ();
 sg13g2_fill_2 FILLER_8_1026 ();
 sg13g2_fill_1 FILLER_8_1028 ();
 sg13g2_decap_8 FILLER_9_4 ();
 sg13g2_decap_8 FILLER_9_11 ();
 sg13g2_decap_8 FILLER_9_18 ();
 sg13g2_decap_8 FILLER_9_25 ();
 sg13g2_decap_8 FILLER_9_32 ();
 sg13g2_decap_8 FILLER_9_39 ();
 sg13g2_decap_8 FILLER_9_46 ();
 sg13g2_decap_8 FILLER_9_53 ();
 sg13g2_decap_8 FILLER_9_60 ();
 sg13g2_decap_8 FILLER_9_67 ();
 sg13g2_decap_8 FILLER_9_74 ();
 sg13g2_decap_8 FILLER_9_81 ();
 sg13g2_decap_8 FILLER_9_88 ();
 sg13g2_decap_8 FILLER_9_95 ();
 sg13g2_decap_8 FILLER_9_102 ();
 sg13g2_decap_8 FILLER_9_109 ();
 sg13g2_decap_8 FILLER_9_116 ();
 sg13g2_decap_8 FILLER_9_123 ();
 sg13g2_decap_8 FILLER_9_130 ();
 sg13g2_decap_8 FILLER_9_137 ();
 sg13g2_decap_8 FILLER_9_144 ();
 sg13g2_decap_8 FILLER_9_151 ();
 sg13g2_decap_8 FILLER_9_158 ();
 sg13g2_decap_8 FILLER_9_165 ();
 sg13g2_decap_8 FILLER_9_172 ();
 sg13g2_decap_8 FILLER_9_179 ();
 sg13g2_decap_8 FILLER_9_186 ();
 sg13g2_decap_8 FILLER_9_193 ();
 sg13g2_decap_8 FILLER_9_200 ();
 sg13g2_decap_8 FILLER_9_207 ();
 sg13g2_decap_8 FILLER_9_214 ();
 sg13g2_decap_8 FILLER_9_221 ();
 sg13g2_decap_8 FILLER_9_228 ();
 sg13g2_decap_8 FILLER_9_235 ();
 sg13g2_decap_8 FILLER_9_242 ();
 sg13g2_decap_8 FILLER_9_249 ();
 sg13g2_decap_8 FILLER_9_256 ();
 sg13g2_decap_8 FILLER_9_263 ();
 sg13g2_decap_8 FILLER_9_270 ();
 sg13g2_decap_8 FILLER_9_277 ();
 sg13g2_decap_8 FILLER_9_284 ();
 sg13g2_decap_8 FILLER_9_291 ();
 sg13g2_decap_8 FILLER_9_298 ();
 sg13g2_decap_8 FILLER_9_305 ();
 sg13g2_decap_8 FILLER_9_312 ();
 sg13g2_decap_8 FILLER_9_319 ();
 sg13g2_decap_8 FILLER_9_326 ();
 sg13g2_decap_8 FILLER_9_333 ();
 sg13g2_decap_8 FILLER_9_340 ();
 sg13g2_decap_8 FILLER_9_347 ();
 sg13g2_decap_8 FILLER_9_354 ();
 sg13g2_decap_8 FILLER_9_361 ();
 sg13g2_decap_8 FILLER_9_368 ();
 sg13g2_decap_8 FILLER_9_375 ();
 sg13g2_decap_8 FILLER_9_382 ();
 sg13g2_decap_8 FILLER_9_389 ();
 sg13g2_decap_8 FILLER_9_396 ();
 sg13g2_decap_8 FILLER_9_403 ();
 sg13g2_decap_8 FILLER_9_410 ();
 sg13g2_decap_8 FILLER_9_417 ();
 sg13g2_decap_8 FILLER_9_424 ();
 sg13g2_decap_8 FILLER_9_431 ();
 sg13g2_decap_8 FILLER_9_438 ();
 sg13g2_decap_8 FILLER_9_445 ();
 sg13g2_decap_8 FILLER_9_452 ();
 sg13g2_decap_8 FILLER_9_459 ();
 sg13g2_decap_8 FILLER_9_466 ();
 sg13g2_decap_8 FILLER_9_473 ();
 sg13g2_decap_8 FILLER_9_480 ();
 sg13g2_decap_8 FILLER_9_487 ();
 sg13g2_decap_8 FILLER_9_494 ();
 sg13g2_decap_8 FILLER_9_501 ();
 sg13g2_decap_8 FILLER_9_508 ();
 sg13g2_decap_8 FILLER_9_515 ();
 sg13g2_decap_8 FILLER_9_522 ();
 sg13g2_decap_8 FILLER_9_529 ();
 sg13g2_decap_8 FILLER_9_536 ();
 sg13g2_decap_8 FILLER_9_543 ();
 sg13g2_decap_8 FILLER_9_550 ();
 sg13g2_decap_8 FILLER_9_557 ();
 sg13g2_decap_8 FILLER_9_564 ();
 sg13g2_decap_8 FILLER_9_571 ();
 sg13g2_decap_8 FILLER_9_578 ();
 sg13g2_decap_8 FILLER_9_585 ();
 sg13g2_decap_8 FILLER_9_592 ();
 sg13g2_decap_8 FILLER_9_599 ();
 sg13g2_decap_8 FILLER_9_606 ();
 sg13g2_decap_8 FILLER_9_613 ();
 sg13g2_decap_8 FILLER_9_620 ();
 sg13g2_decap_8 FILLER_9_627 ();
 sg13g2_decap_8 FILLER_9_634 ();
 sg13g2_decap_8 FILLER_9_641 ();
 sg13g2_decap_8 FILLER_9_648 ();
 sg13g2_decap_8 FILLER_9_655 ();
 sg13g2_decap_8 FILLER_9_662 ();
 sg13g2_decap_8 FILLER_9_669 ();
 sg13g2_decap_8 FILLER_9_676 ();
 sg13g2_decap_8 FILLER_9_683 ();
 sg13g2_decap_8 FILLER_9_690 ();
 sg13g2_decap_8 FILLER_9_697 ();
 sg13g2_decap_8 FILLER_9_704 ();
 sg13g2_decap_8 FILLER_9_711 ();
 sg13g2_decap_8 FILLER_9_718 ();
 sg13g2_decap_8 FILLER_9_725 ();
 sg13g2_decap_8 FILLER_9_732 ();
 sg13g2_decap_8 FILLER_9_739 ();
 sg13g2_decap_8 FILLER_9_746 ();
 sg13g2_decap_8 FILLER_9_753 ();
 sg13g2_decap_8 FILLER_9_760 ();
 sg13g2_decap_8 FILLER_9_767 ();
 sg13g2_decap_8 FILLER_9_774 ();
 sg13g2_decap_8 FILLER_9_781 ();
 sg13g2_decap_8 FILLER_9_788 ();
 sg13g2_decap_8 FILLER_9_795 ();
 sg13g2_decap_8 FILLER_9_802 ();
 sg13g2_decap_8 FILLER_9_809 ();
 sg13g2_decap_8 FILLER_9_816 ();
 sg13g2_decap_8 FILLER_9_823 ();
 sg13g2_decap_8 FILLER_9_830 ();
 sg13g2_decap_8 FILLER_9_837 ();
 sg13g2_decap_8 FILLER_9_844 ();
 sg13g2_decap_8 FILLER_9_851 ();
 sg13g2_decap_8 FILLER_9_858 ();
 sg13g2_decap_8 FILLER_9_865 ();
 sg13g2_decap_8 FILLER_9_872 ();
 sg13g2_decap_8 FILLER_9_879 ();
 sg13g2_decap_8 FILLER_9_886 ();
 sg13g2_decap_8 FILLER_9_893 ();
 sg13g2_decap_8 FILLER_9_900 ();
 sg13g2_decap_8 FILLER_9_907 ();
 sg13g2_decap_8 FILLER_9_914 ();
 sg13g2_decap_8 FILLER_9_921 ();
 sg13g2_decap_8 FILLER_9_928 ();
 sg13g2_decap_8 FILLER_9_935 ();
 sg13g2_decap_8 FILLER_9_942 ();
 sg13g2_decap_8 FILLER_9_949 ();
 sg13g2_decap_8 FILLER_9_956 ();
 sg13g2_decap_8 FILLER_9_963 ();
 sg13g2_decap_8 FILLER_9_970 ();
 sg13g2_decap_8 FILLER_9_977 ();
 sg13g2_decap_8 FILLER_9_984 ();
 sg13g2_decap_8 FILLER_9_991 ();
 sg13g2_decap_8 FILLER_9_998 ();
 sg13g2_decap_8 FILLER_9_1005 ();
 sg13g2_decap_8 FILLER_9_1012 ();
 sg13g2_decap_8 FILLER_9_1019 ();
 sg13g2_fill_2 FILLER_9_1026 ();
 sg13g2_fill_1 FILLER_9_1028 ();
 sg13g2_decap_8 FILLER_10_4 ();
 sg13g2_decap_8 FILLER_10_11 ();
 sg13g2_decap_8 FILLER_10_18 ();
 sg13g2_decap_8 FILLER_10_25 ();
 sg13g2_decap_8 FILLER_10_32 ();
 sg13g2_decap_8 FILLER_10_39 ();
 sg13g2_decap_8 FILLER_10_46 ();
 sg13g2_decap_8 FILLER_10_53 ();
 sg13g2_decap_8 FILLER_10_60 ();
 sg13g2_decap_8 FILLER_10_67 ();
 sg13g2_decap_8 FILLER_10_74 ();
 sg13g2_decap_8 FILLER_10_81 ();
 sg13g2_decap_8 FILLER_10_88 ();
 sg13g2_decap_8 FILLER_10_95 ();
 sg13g2_decap_8 FILLER_10_102 ();
 sg13g2_decap_8 FILLER_10_109 ();
 sg13g2_decap_8 FILLER_10_116 ();
 sg13g2_decap_8 FILLER_10_123 ();
 sg13g2_decap_8 FILLER_10_130 ();
 sg13g2_decap_8 FILLER_10_137 ();
 sg13g2_decap_8 FILLER_10_144 ();
 sg13g2_decap_8 FILLER_10_151 ();
 sg13g2_decap_8 FILLER_10_158 ();
 sg13g2_decap_8 FILLER_10_165 ();
 sg13g2_decap_8 FILLER_10_172 ();
 sg13g2_decap_8 FILLER_10_179 ();
 sg13g2_decap_8 FILLER_10_186 ();
 sg13g2_decap_8 FILLER_10_193 ();
 sg13g2_decap_8 FILLER_10_200 ();
 sg13g2_decap_8 FILLER_10_207 ();
 sg13g2_decap_8 FILLER_10_214 ();
 sg13g2_decap_8 FILLER_10_221 ();
 sg13g2_decap_8 FILLER_10_228 ();
 sg13g2_decap_8 FILLER_10_235 ();
 sg13g2_decap_8 FILLER_10_242 ();
 sg13g2_decap_8 FILLER_10_249 ();
 sg13g2_decap_8 FILLER_10_256 ();
 sg13g2_decap_8 FILLER_10_263 ();
 sg13g2_decap_8 FILLER_10_270 ();
 sg13g2_decap_8 FILLER_10_277 ();
 sg13g2_decap_8 FILLER_10_284 ();
 sg13g2_decap_8 FILLER_10_291 ();
 sg13g2_decap_8 FILLER_10_298 ();
 sg13g2_decap_8 FILLER_10_305 ();
 sg13g2_decap_8 FILLER_10_312 ();
 sg13g2_decap_8 FILLER_10_319 ();
 sg13g2_decap_8 FILLER_10_326 ();
 sg13g2_decap_8 FILLER_10_333 ();
 sg13g2_decap_8 FILLER_10_340 ();
 sg13g2_decap_8 FILLER_10_347 ();
 sg13g2_decap_8 FILLER_10_354 ();
 sg13g2_decap_8 FILLER_10_361 ();
 sg13g2_decap_8 FILLER_10_368 ();
 sg13g2_decap_8 FILLER_10_375 ();
 sg13g2_decap_8 FILLER_10_382 ();
 sg13g2_decap_8 FILLER_10_389 ();
 sg13g2_decap_8 FILLER_10_396 ();
 sg13g2_decap_8 FILLER_10_403 ();
 sg13g2_decap_8 FILLER_10_410 ();
 sg13g2_decap_8 FILLER_10_417 ();
 sg13g2_decap_8 FILLER_10_424 ();
 sg13g2_decap_8 FILLER_10_431 ();
 sg13g2_decap_8 FILLER_10_438 ();
 sg13g2_decap_8 FILLER_10_445 ();
 sg13g2_decap_8 FILLER_10_452 ();
 sg13g2_decap_8 FILLER_10_459 ();
 sg13g2_decap_8 FILLER_10_466 ();
 sg13g2_decap_8 FILLER_10_473 ();
 sg13g2_decap_8 FILLER_10_480 ();
 sg13g2_decap_8 FILLER_10_487 ();
 sg13g2_decap_8 FILLER_10_494 ();
 sg13g2_decap_8 FILLER_10_501 ();
 sg13g2_decap_8 FILLER_10_508 ();
 sg13g2_decap_8 FILLER_10_515 ();
 sg13g2_decap_8 FILLER_10_522 ();
 sg13g2_decap_8 FILLER_10_529 ();
 sg13g2_decap_8 FILLER_10_536 ();
 sg13g2_decap_8 FILLER_10_543 ();
 sg13g2_decap_8 FILLER_10_550 ();
 sg13g2_decap_8 FILLER_10_557 ();
 sg13g2_decap_8 FILLER_10_564 ();
 sg13g2_decap_8 FILLER_10_571 ();
 sg13g2_decap_8 FILLER_10_578 ();
 sg13g2_decap_8 FILLER_10_585 ();
 sg13g2_decap_8 FILLER_10_592 ();
 sg13g2_decap_8 FILLER_10_599 ();
 sg13g2_decap_8 FILLER_10_606 ();
 sg13g2_decap_8 FILLER_10_613 ();
 sg13g2_decap_8 FILLER_10_620 ();
 sg13g2_decap_8 FILLER_10_627 ();
 sg13g2_decap_8 FILLER_10_634 ();
 sg13g2_decap_8 FILLER_10_641 ();
 sg13g2_decap_8 FILLER_10_648 ();
 sg13g2_decap_8 FILLER_10_655 ();
 sg13g2_decap_8 FILLER_10_662 ();
 sg13g2_decap_8 FILLER_10_669 ();
 sg13g2_decap_8 FILLER_10_676 ();
 sg13g2_decap_8 FILLER_10_683 ();
 sg13g2_decap_8 FILLER_10_690 ();
 sg13g2_decap_8 FILLER_10_697 ();
 sg13g2_decap_8 FILLER_10_704 ();
 sg13g2_decap_8 FILLER_10_711 ();
 sg13g2_decap_8 FILLER_10_718 ();
 sg13g2_decap_8 FILLER_10_725 ();
 sg13g2_decap_8 FILLER_10_732 ();
 sg13g2_decap_8 FILLER_10_739 ();
 sg13g2_decap_8 FILLER_10_746 ();
 sg13g2_decap_8 FILLER_10_753 ();
 sg13g2_decap_8 FILLER_10_760 ();
 sg13g2_decap_8 FILLER_10_767 ();
 sg13g2_decap_8 FILLER_10_774 ();
 sg13g2_decap_8 FILLER_10_781 ();
 sg13g2_decap_8 FILLER_10_788 ();
 sg13g2_decap_8 FILLER_10_795 ();
 sg13g2_decap_8 FILLER_10_802 ();
 sg13g2_decap_8 FILLER_10_809 ();
 sg13g2_decap_8 FILLER_10_816 ();
 sg13g2_decap_8 FILLER_10_823 ();
 sg13g2_decap_8 FILLER_10_830 ();
 sg13g2_decap_8 FILLER_10_837 ();
 sg13g2_decap_8 FILLER_10_844 ();
 sg13g2_decap_8 FILLER_10_851 ();
 sg13g2_decap_8 FILLER_10_858 ();
 sg13g2_decap_8 FILLER_10_865 ();
 sg13g2_decap_8 FILLER_10_872 ();
 sg13g2_decap_8 FILLER_10_879 ();
 sg13g2_decap_8 FILLER_10_886 ();
 sg13g2_decap_8 FILLER_10_893 ();
 sg13g2_decap_8 FILLER_10_900 ();
 sg13g2_decap_8 FILLER_10_907 ();
 sg13g2_decap_8 FILLER_10_914 ();
 sg13g2_decap_8 FILLER_10_921 ();
 sg13g2_decap_8 FILLER_10_928 ();
 sg13g2_decap_8 FILLER_10_935 ();
 sg13g2_decap_8 FILLER_10_942 ();
 sg13g2_decap_8 FILLER_10_949 ();
 sg13g2_decap_8 FILLER_10_956 ();
 sg13g2_decap_8 FILLER_10_963 ();
 sg13g2_decap_8 FILLER_10_970 ();
 sg13g2_decap_8 FILLER_10_977 ();
 sg13g2_decap_8 FILLER_10_984 ();
 sg13g2_decap_8 FILLER_10_991 ();
 sg13g2_decap_8 FILLER_10_998 ();
 sg13g2_decap_8 FILLER_10_1005 ();
 sg13g2_decap_8 FILLER_10_1012 ();
 sg13g2_decap_8 FILLER_10_1019 ();
 sg13g2_fill_2 FILLER_10_1026 ();
 sg13g2_fill_1 FILLER_10_1028 ();
 sg13g2_decap_8 FILLER_11_4 ();
 sg13g2_decap_8 FILLER_11_11 ();
 sg13g2_decap_8 FILLER_11_18 ();
 sg13g2_decap_8 FILLER_11_25 ();
 sg13g2_decap_8 FILLER_11_32 ();
 sg13g2_decap_8 FILLER_11_39 ();
 sg13g2_decap_8 FILLER_11_46 ();
 sg13g2_decap_8 FILLER_11_53 ();
 sg13g2_decap_8 FILLER_11_60 ();
 sg13g2_decap_8 FILLER_11_67 ();
 sg13g2_decap_8 FILLER_11_74 ();
 sg13g2_decap_8 FILLER_11_81 ();
 sg13g2_decap_8 FILLER_11_88 ();
 sg13g2_decap_8 FILLER_11_95 ();
 sg13g2_decap_8 FILLER_11_102 ();
 sg13g2_decap_8 FILLER_11_109 ();
 sg13g2_decap_8 FILLER_11_116 ();
 sg13g2_decap_8 FILLER_11_123 ();
 sg13g2_decap_8 FILLER_11_130 ();
 sg13g2_decap_8 FILLER_11_137 ();
 sg13g2_decap_8 FILLER_11_144 ();
 sg13g2_decap_8 FILLER_11_151 ();
 sg13g2_decap_8 FILLER_11_158 ();
 sg13g2_decap_8 FILLER_11_165 ();
 sg13g2_decap_8 FILLER_11_172 ();
 sg13g2_decap_8 FILLER_11_179 ();
 sg13g2_decap_8 FILLER_11_186 ();
 sg13g2_decap_8 FILLER_11_193 ();
 sg13g2_decap_8 FILLER_11_200 ();
 sg13g2_decap_8 FILLER_11_207 ();
 sg13g2_decap_8 FILLER_11_214 ();
 sg13g2_decap_8 FILLER_11_221 ();
 sg13g2_decap_8 FILLER_11_228 ();
 sg13g2_decap_8 FILLER_11_235 ();
 sg13g2_decap_8 FILLER_11_242 ();
 sg13g2_decap_8 FILLER_11_249 ();
 sg13g2_decap_8 FILLER_11_256 ();
 sg13g2_decap_8 FILLER_11_263 ();
 sg13g2_decap_8 FILLER_11_270 ();
 sg13g2_decap_8 FILLER_11_277 ();
 sg13g2_decap_8 FILLER_11_284 ();
 sg13g2_decap_8 FILLER_11_291 ();
 sg13g2_decap_8 FILLER_11_298 ();
 sg13g2_decap_8 FILLER_11_305 ();
 sg13g2_decap_8 FILLER_11_312 ();
 sg13g2_decap_8 FILLER_11_319 ();
 sg13g2_decap_8 FILLER_11_326 ();
 sg13g2_decap_8 FILLER_11_333 ();
 sg13g2_decap_8 FILLER_11_340 ();
 sg13g2_decap_8 FILLER_11_347 ();
 sg13g2_decap_8 FILLER_11_354 ();
 sg13g2_decap_8 FILLER_11_361 ();
 sg13g2_decap_8 FILLER_11_368 ();
 sg13g2_decap_8 FILLER_11_375 ();
 sg13g2_decap_8 FILLER_11_382 ();
 sg13g2_decap_8 FILLER_11_389 ();
 sg13g2_decap_8 FILLER_11_396 ();
 sg13g2_decap_8 FILLER_11_403 ();
 sg13g2_decap_8 FILLER_11_410 ();
 sg13g2_decap_8 FILLER_11_417 ();
 sg13g2_decap_8 FILLER_11_424 ();
 sg13g2_decap_8 FILLER_11_431 ();
 sg13g2_decap_8 FILLER_11_438 ();
 sg13g2_decap_8 FILLER_11_445 ();
 sg13g2_decap_8 FILLER_11_452 ();
 sg13g2_decap_8 FILLER_11_459 ();
 sg13g2_decap_8 FILLER_11_466 ();
 sg13g2_decap_8 FILLER_11_473 ();
 sg13g2_decap_8 FILLER_11_480 ();
 sg13g2_decap_8 FILLER_11_487 ();
 sg13g2_decap_8 FILLER_11_494 ();
 sg13g2_decap_8 FILLER_11_501 ();
 sg13g2_decap_8 FILLER_11_508 ();
 sg13g2_decap_8 FILLER_11_515 ();
 sg13g2_decap_8 FILLER_11_522 ();
 sg13g2_decap_8 FILLER_11_529 ();
 sg13g2_decap_8 FILLER_11_536 ();
 sg13g2_decap_8 FILLER_11_543 ();
 sg13g2_decap_8 FILLER_11_550 ();
 sg13g2_decap_8 FILLER_11_557 ();
 sg13g2_decap_8 FILLER_11_564 ();
 sg13g2_decap_8 FILLER_11_571 ();
 sg13g2_decap_8 FILLER_11_578 ();
 sg13g2_decap_8 FILLER_11_585 ();
 sg13g2_decap_8 FILLER_11_592 ();
 sg13g2_decap_8 FILLER_11_599 ();
 sg13g2_decap_8 FILLER_11_606 ();
 sg13g2_decap_8 FILLER_11_613 ();
 sg13g2_decap_8 FILLER_11_620 ();
 sg13g2_decap_8 FILLER_11_627 ();
 sg13g2_decap_8 FILLER_11_634 ();
 sg13g2_decap_8 FILLER_11_641 ();
 sg13g2_decap_8 FILLER_11_648 ();
 sg13g2_decap_8 FILLER_11_655 ();
 sg13g2_decap_8 FILLER_11_662 ();
 sg13g2_decap_8 FILLER_11_669 ();
 sg13g2_decap_8 FILLER_11_676 ();
 sg13g2_decap_8 FILLER_11_683 ();
 sg13g2_decap_8 FILLER_11_690 ();
 sg13g2_decap_8 FILLER_11_697 ();
 sg13g2_decap_8 FILLER_11_704 ();
 sg13g2_decap_8 FILLER_11_711 ();
 sg13g2_decap_8 FILLER_11_718 ();
 sg13g2_decap_8 FILLER_11_725 ();
 sg13g2_decap_8 FILLER_11_732 ();
 sg13g2_decap_8 FILLER_11_739 ();
 sg13g2_decap_8 FILLER_11_746 ();
 sg13g2_decap_8 FILLER_11_753 ();
 sg13g2_decap_8 FILLER_11_760 ();
 sg13g2_decap_8 FILLER_11_767 ();
 sg13g2_decap_8 FILLER_11_774 ();
 sg13g2_decap_8 FILLER_11_781 ();
 sg13g2_decap_8 FILLER_11_788 ();
 sg13g2_decap_8 FILLER_11_795 ();
 sg13g2_decap_8 FILLER_11_802 ();
 sg13g2_decap_8 FILLER_11_809 ();
 sg13g2_decap_8 FILLER_11_816 ();
 sg13g2_decap_8 FILLER_11_823 ();
 sg13g2_decap_8 FILLER_11_830 ();
 sg13g2_decap_8 FILLER_11_837 ();
 sg13g2_decap_8 FILLER_11_844 ();
 sg13g2_decap_8 FILLER_11_851 ();
 sg13g2_decap_8 FILLER_11_858 ();
 sg13g2_decap_8 FILLER_11_865 ();
 sg13g2_decap_8 FILLER_11_872 ();
 sg13g2_decap_8 FILLER_11_879 ();
 sg13g2_decap_8 FILLER_11_886 ();
 sg13g2_decap_8 FILLER_11_893 ();
 sg13g2_decap_8 FILLER_11_900 ();
 sg13g2_decap_8 FILLER_11_907 ();
 sg13g2_decap_8 FILLER_11_914 ();
 sg13g2_decap_8 FILLER_11_921 ();
 sg13g2_decap_8 FILLER_11_928 ();
 sg13g2_decap_8 FILLER_11_935 ();
 sg13g2_decap_8 FILLER_11_942 ();
 sg13g2_decap_8 FILLER_11_949 ();
 sg13g2_decap_8 FILLER_11_956 ();
 sg13g2_decap_8 FILLER_11_963 ();
 sg13g2_decap_8 FILLER_11_970 ();
 sg13g2_decap_8 FILLER_11_977 ();
 sg13g2_decap_8 FILLER_11_984 ();
 sg13g2_decap_8 FILLER_11_991 ();
 sg13g2_decap_8 FILLER_11_998 ();
 sg13g2_decap_8 FILLER_11_1005 ();
 sg13g2_decap_8 FILLER_11_1012 ();
 sg13g2_decap_8 FILLER_11_1019 ();
 sg13g2_fill_2 FILLER_11_1026 ();
 sg13g2_fill_1 FILLER_11_1028 ();
 sg13g2_decap_8 FILLER_12_4 ();
 sg13g2_decap_8 FILLER_12_11 ();
 sg13g2_decap_8 FILLER_12_18 ();
 sg13g2_decap_8 FILLER_12_25 ();
 sg13g2_decap_8 FILLER_12_32 ();
 sg13g2_decap_8 FILLER_12_39 ();
 sg13g2_decap_8 FILLER_12_46 ();
 sg13g2_decap_8 FILLER_12_53 ();
 sg13g2_decap_8 FILLER_12_60 ();
 sg13g2_decap_8 FILLER_12_67 ();
 sg13g2_decap_8 FILLER_12_74 ();
 sg13g2_decap_8 FILLER_12_81 ();
 sg13g2_decap_8 FILLER_12_88 ();
 sg13g2_decap_8 FILLER_12_95 ();
 sg13g2_decap_8 FILLER_12_102 ();
 sg13g2_decap_8 FILLER_12_109 ();
 sg13g2_decap_8 FILLER_12_116 ();
 sg13g2_decap_8 FILLER_12_123 ();
 sg13g2_decap_8 FILLER_12_130 ();
 sg13g2_decap_8 FILLER_12_137 ();
 sg13g2_decap_8 FILLER_12_144 ();
 sg13g2_decap_8 FILLER_12_151 ();
 sg13g2_decap_8 FILLER_12_158 ();
 sg13g2_decap_8 FILLER_12_165 ();
 sg13g2_decap_8 FILLER_12_172 ();
 sg13g2_decap_8 FILLER_12_179 ();
 sg13g2_decap_8 FILLER_12_186 ();
 sg13g2_decap_8 FILLER_12_193 ();
 sg13g2_decap_8 FILLER_12_200 ();
 sg13g2_decap_8 FILLER_12_207 ();
 sg13g2_decap_8 FILLER_12_214 ();
 sg13g2_decap_8 FILLER_12_221 ();
 sg13g2_decap_8 FILLER_12_228 ();
 sg13g2_decap_8 FILLER_12_235 ();
 sg13g2_decap_8 FILLER_12_242 ();
 sg13g2_decap_8 FILLER_12_249 ();
 sg13g2_decap_8 FILLER_12_256 ();
 sg13g2_decap_8 FILLER_12_263 ();
 sg13g2_decap_8 FILLER_12_270 ();
 sg13g2_decap_8 FILLER_12_277 ();
 sg13g2_decap_8 FILLER_12_284 ();
 sg13g2_decap_8 FILLER_12_291 ();
 sg13g2_decap_8 FILLER_12_298 ();
 sg13g2_decap_8 FILLER_12_305 ();
 sg13g2_decap_8 FILLER_12_312 ();
 sg13g2_decap_8 FILLER_12_319 ();
 sg13g2_decap_8 FILLER_12_326 ();
 sg13g2_decap_8 FILLER_12_333 ();
 sg13g2_decap_8 FILLER_12_340 ();
 sg13g2_decap_8 FILLER_12_347 ();
 sg13g2_decap_8 FILLER_12_354 ();
 sg13g2_decap_8 FILLER_12_361 ();
 sg13g2_decap_8 FILLER_12_368 ();
 sg13g2_decap_8 FILLER_12_375 ();
 sg13g2_decap_8 FILLER_12_382 ();
 sg13g2_decap_8 FILLER_12_389 ();
 sg13g2_decap_8 FILLER_12_396 ();
 sg13g2_decap_8 FILLER_12_403 ();
 sg13g2_decap_8 FILLER_12_410 ();
 sg13g2_decap_8 FILLER_12_417 ();
 sg13g2_decap_8 FILLER_12_424 ();
 sg13g2_decap_8 FILLER_12_431 ();
 sg13g2_decap_8 FILLER_12_438 ();
 sg13g2_decap_8 FILLER_12_445 ();
 sg13g2_decap_8 FILLER_12_452 ();
 sg13g2_decap_8 FILLER_12_459 ();
 sg13g2_decap_8 FILLER_12_466 ();
 sg13g2_decap_8 FILLER_12_473 ();
 sg13g2_decap_8 FILLER_12_480 ();
 sg13g2_decap_8 FILLER_12_487 ();
 sg13g2_decap_8 FILLER_12_494 ();
 sg13g2_decap_8 FILLER_12_501 ();
 sg13g2_decap_8 FILLER_12_508 ();
 sg13g2_decap_8 FILLER_12_515 ();
 sg13g2_decap_8 FILLER_12_522 ();
 sg13g2_decap_8 FILLER_12_529 ();
 sg13g2_decap_8 FILLER_12_536 ();
 sg13g2_decap_8 FILLER_12_543 ();
 sg13g2_decap_8 FILLER_12_550 ();
 sg13g2_decap_8 FILLER_12_557 ();
 sg13g2_decap_8 FILLER_12_564 ();
 sg13g2_decap_8 FILLER_12_571 ();
 sg13g2_decap_8 FILLER_12_578 ();
 sg13g2_decap_8 FILLER_12_585 ();
 sg13g2_decap_8 FILLER_12_592 ();
 sg13g2_decap_8 FILLER_12_599 ();
 sg13g2_decap_8 FILLER_12_606 ();
 sg13g2_decap_8 FILLER_12_613 ();
 sg13g2_decap_8 FILLER_12_620 ();
 sg13g2_decap_8 FILLER_12_627 ();
 sg13g2_decap_8 FILLER_12_634 ();
 sg13g2_decap_8 FILLER_12_641 ();
 sg13g2_decap_8 FILLER_12_648 ();
 sg13g2_decap_8 FILLER_12_655 ();
 sg13g2_decap_8 FILLER_12_662 ();
 sg13g2_decap_8 FILLER_12_669 ();
 sg13g2_decap_8 FILLER_12_676 ();
 sg13g2_decap_8 FILLER_12_683 ();
 sg13g2_decap_8 FILLER_12_690 ();
 sg13g2_decap_8 FILLER_12_697 ();
 sg13g2_decap_8 FILLER_12_704 ();
 sg13g2_decap_8 FILLER_12_711 ();
 sg13g2_decap_8 FILLER_12_718 ();
 sg13g2_decap_8 FILLER_12_725 ();
 sg13g2_decap_8 FILLER_12_732 ();
 sg13g2_decap_8 FILLER_12_739 ();
 sg13g2_decap_8 FILLER_12_746 ();
 sg13g2_decap_8 FILLER_12_753 ();
 sg13g2_decap_8 FILLER_12_760 ();
 sg13g2_decap_8 FILLER_12_767 ();
 sg13g2_decap_8 FILLER_12_774 ();
 sg13g2_decap_8 FILLER_12_781 ();
 sg13g2_decap_8 FILLER_12_788 ();
 sg13g2_decap_8 FILLER_12_795 ();
 sg13g2_decap_8 FILLER_12_802 ();
 sg13g2_decap_8 FILLER_12_809 ();
 sg13g2_decap_8 FILLER_12_816 ();
 sg13g2_decap_8 FILLER_12_823 ();
 sg13g2_decap_8 FILLER_12_830 ();
 sg13g2_decap_8 FILLER_12_837 ();
 sg13g2_decap_8 FILLER_12_844 ();
 sg13g2_decap_8 FILLER_12_851 ();
 sg13g2_decap_8 FILLER_12_858 ();
 sg13g2_decap_8 FILLER_12_865 ();
 sg13g2_decap_8 FILLER_12_872 ();
 sg13g2_decap_8 FILLER_12_879 ();
 sg13g2_decap_8 FILLER_12_886 ();
 sg13g2_decap_8 FILLER_12_893 ();
 sg13g2_decap_8 FILLER_12_900 ();
 sg13g2_decap_8 FILLER_12_907 ();
 sg13g2_decap_8 FILLER_12_914 ();
 sg13g2_decap_8 FILLER_12_921 ();
 sg13g2_decap_8 FILLER_12_928 ();
 sg13g2_decap_8 FILLER_12_935 ();
 sg13g2_decap_8 FILLER_12_942 ();
 sg13g2_decap_8 FILLER_12_949 ();
 sg13g2_decap_8 FILLER_12_956 ();
 sg13g2_decap_8 FILLER_12_963 ();
 sg13g2_decap_8 FILLER_12_970 ();
 sg13g2_decap_8 FILLER_12_977 ();
 sg13g2_decap_8 FILLER_12_984 ();
 sg13g2_decap_8 FILLER_12_991 ();
 sg13g2_decap_8 FILLER_12_998 ();
 sg13g2_decap_8 FILLER_12_1005 ();
 sg13g2_decap_8 FILLER_12_1012 ();
 sg13g2_decap_8 FILLER_12_1019 ();
 sg13g2_fill_2 FILLER_12_1026 ();
 sg13g2_fill_1 FILLER_12_1028 ();
 sg13g2_decap_8 FILLER_13_4 ();
 sg13g2_decap_8 FILLER_13_11 ();
 sg13g2_decap_8 FILLER_13_18 ();
 sg13g2_decap_8 FILLER_13_25 ();
 sg13g2_decap_8 FILLER_13_32 ();
 sg13g2_decap_8 FILLER_13_39 ();
 sg13g2_decap_8 FILLER_13_46 ();
 sg13g2_decap_8 FILLER_13_53 ();
 sg13g2_decap_8 FILLER_13_60 ();
 sg13g2_decap_8 FILLER_13_67 ();
 sg13g2_decap_8 FILLER_13_74 ();
 sg13g2_decap_8 FILLER_13_81 ();
 sg13g2_decap_8 FILLER_13_88 ();
 sg13g2_decap_8 FILLER_13_95 ();
 sg13g2_decap_8 FILLER_13_102 ();
 sg13g2_decap_8 FILLER_13_109 ();
 sg13g2_decap_8 FILLER_13_116 ();
 sg13g2_decap_8 FILLER_13_123 ();
 sg13g2_decap_8 FILLER_13_130 ();
 sg13g2_decap_8 FILLER_13_137 ();
 sg13g2_decap_8 FILLER_13_144 ();
 sg13g2_decap_8 FILLER_13_151 ();
 sg13g2_decap_8 FILLER_13_158 ();
 sg13g2_decap_8 FILLER_13_165 ();
 sg13g2_decap_8 FILLER_13_172 ();
 sg13g2_decap_8 FILLER_13_179 ();
 sg13g2_decap_8 FILLER_13_186 ();
 sg13g2_decap_8 FILLER_13_193 ();
 sg13g2_decap_8 FILLER_13_200 ();
 sg13g2_decap_8 FILLER_13_207 ();
 sg13g2_decap_8 FILLER_13_214 ();
 sg13g2_decap_8 FILLER_13_221 ();
 sg13g2_decap_8 FILLER_13_228 ();
 sg13g2_decap_8 FILLER_13_235 ();
 sg13g2_decap_8 FILLER_13_242 ();
 sg13g2_decap_8 FILLER_13_249 ();
 sg13g2_decap_8 FILLER_13_256 ();
 sg13g2_decap_8 FILLER_13_263 ();
 sg13g2_decap_8 FILLER_13_270 ();
 sg13g2_decap_8 FILLER_13_277 ();
 sg13g2_decap_8 FILLER_13_284 ();
 sg13g2_decap_8 FILLER_13_291 ();
 sg13g2_decap_8 FILLER_13_298 ();
 sg13g2_decap_8 FILLER_13_305 ();
 sg13g2_decap_8 FILLER_13_312 ();
 sg13g2_decap_8 FILLER_13_319 ();
 sg13g2_decap_8 FILLER_13_326 ();
 sg13g2_decap_8 FILLER_13_333 ();
 sg13g2_decap_8 FILLER_13_340 ();
 sg13g2_decap_8 FILLER_13_347 ();
 sg13g2_decap_8 FILLER_13_354 ();
 sg13g2_decap_8 FILLER_13_361 ();
 sg13g2_decap_8 FILLER_13_368 ();
 sg13g2_decap_8 FILLER_13_375 ();
 sg13g2_decap_8 FILLER_13_382 ();
 sg13g2_decap_8 FILLER_13_389 ();
 sg13g2_decap_8 FILLER_13_396 ();
 sg13g2_decap_8 FILLER_13_403 ();
 sg13g2_decap_8 FILLER_13_410 ();
 sg13g2_decap_8 FILLER_13_417 ();
 sg13g2_decap_8 FILLER_13_424 ();
 sg13g2_decap_8 FILLER_13_431 ();
 sg13g2_decap_8 FILLER_13_438 ();
 sg13g2_decap_8 FILLER_13_445 ();
 sg13g2_decap_8 FILLER_13_452 ();
 sg13g2_decap_8 FILLER_13_459 ();
 sg13g2_decap_8 FILLER_13_466 ();
 sg13g2_decap_8 FILLER_13_473 ();
 sg13g2_decap_8 FILLER_13_480 ();
 sg13g2_decap_8 FILLER_13_487 ();
 sg13g2_decap_8 FILLER_13_494 ();
 sg13g2_decap_8 FILLER_13_501 ();
 sg13g2_decap_8 FILLER_13_508 ();
 sg13g2_decap_8 FILLER_13_515 ();
 sg13g2_decap_8 FILLER_13_522 ();
 sg13g2_decap_8 FILLER_13_529 ();
 sg13g2_decap_8 FILLER_13_536 ();
 sg13g2_decap_8 FILLER_13_543 ();
 sg13g2_decap_8 FILLER_13_550 ();
 sg13g2_decap_8 FILLER_13_557 ();
 sg13g2_decap_8 FILLER_13_564 ();
 sg13g2_decap_8 FILLER_13_571 ();
 sg13g2_decap_8 FILLER_13_578 ();
 sg13g2_decap_8 FILLER_13_585 ();
 sg13g2_decap_8 FILLER_13_592 ();
 sg13g2_decap_8 FILLER_13_599 ();
 sg13g2_decap_8 FILLER_13_606 ();
 sg13g2_decap_8 FILLER_13_613 ();
 sg13g2_decap_8 FILLER_13_620 ();
 sg13g2_decap_8 FILLER_13_627 ();
 sg13g2_decap_8 FILLER_13_634 ();
 sg13g2_decap_8 FILLER_13_641 ();
 sg13g2_decap_8 FILLER_13_648 ();
 sg13g2_decap_8 FILLER_13_655 ();
 sg13g2_decap_8 FILLER_13_662 ();
 sg13g2_decap_8 FILLER_13_669 ();
 sg13g2_decap_8 FILLER_13_676 ();
 sg13g2_decap_8 FILLER_13_683 ();
 sg13g2_decap_8 FILLER_13_690 ();
 sg13g2_decap_8 FILLER_13_697 ();
 sg13g2_decap_8 FILLER_13_704 ();
 sg13g2_decap_8 FILLER_13_711 ();
 sg13g2_decap_8 FILLER_13_718 ();
 sg13g2_decap_8 FILLER_13_725 ();
 sg13g2_decap_8 FILLER_13_732 ();
 sg13g2_decap_8 FILLER_13_739 ();
 sg13g2_decap_8 FILLER_13_746 ();
 sg13g2_decap_8 FILLER_13_753 ();
 sg13g2_decap_8 FILLER_13_760 ();
 sg13g2_decap_8 FILLER_13_767 ();
 sg13g2_decap_8 FILLER_13_774 ();
 sg13g2_decap_8 FILLER_13_781 ();
 sg13g2_decap_8 FILLER_13_788 ();
 sg13g2_decap_8 FILLER_13_795 ();
 sg13g2_decap_8 FILLER_13_802 ();
 sg13g2_decap_8 FILLER_13_809 ();
 sg13g2_decap_8 FILLER_13_816 ();
 sg13g2_decap_8 FILLER_13_823 ();
 sg13g2_decap_8 FILLER_13_830 ();
 sg13g2_decap_8 FILLER_13_837 ();
 sg13g2_decap_8 FILLER_13_844 ();
 sg13g2_decap_8 FILLER_13_851 ();
 sg13g2_decap_8 FILLER_13_858 ();
 sg13g2_decap_8 FILLER_13_865 ();
 sg13g2_decap_8 FILLER_13_872 ();
 sg13g2_decap_8 FILLER_13_879 ();
 sg13g2_decap_8 FILLER_13_886 ();
 sg13g2_decap_8 FILLER_13_893 ();
 sg13g2_decap_8 FILLER_13_900 ();
 sg13g2_decap_8 FILLER_13_907 ();
 sg13g2_decap_8 FILLER_13_914 ();
 sg13g2_decap_8 FILLER_13_921 ();
 sg13g2_decap_8 FILLER_13_928 ();
 sg13g2_decap_8 FILLER_13_935 ();
 sg13g2_decap_8 FILLER_13_942 ();
 sg13g2_decap_8 FILLER_13_949 ();
 sg13g2_decap_8 FILLER_13_956 ();
 sg13g2_decap_8 FILLER_13_963 ();
 sg13g2_decap_8 FILLER_13_970 ();
 sg13g2_decap_8 FILLER_13_977 ();
 sg13g2_decap_8 FILLER_13_984 ();
 sg13g2_decap_8 FILLER_13_991 ();
 sg13g2_decap_8 FILLER_13_998 ();
 sg13g2_decap_8 FILLER_13_1005 ();
 sg13g2_decap_8 FILLER_13_1012 ();
 sg13g2_decap_8 FILLER_13_1019 ();
 sg13g2_fill_2 FILLER_13_1026 ();
 sg13g2_fill_1 FILLER_13_1028 ();
 sg13g2_decap_8 FILLER_14_4 ();
 sg13g2_decap_8 FILLER_14_11 ();
 sg13g2_decap_8 FILLER_14_18 ();
 sg13g2_decap_8 FILLER_14_25 ();
 sg13g2_decap_8 FILLER_14_32 ();
 sg13g2_decap_8 FILLER_14_39 ();
 sg13g2_decap_8 FILLER_14_46 ();
 sg13g2_decap_8 FILLER_14_53 ();
 sg13g2_decap_8 FILLER_14_60 ();
 sg13g2_decap_8 FILLER_14_67 ();
 sg13g2_decap_8 FILLER_14_74 ();
 sg13g2_decap_8 FILLER_14_81 ();
 sg13g2_decap_8 FILLER_14_88 ();
 sg13g2_decap_8 FILLER_14_95 ();
 sg13g2_decap_8 FILLER_14_102 ();
 sg13g2_decap_8 FILLER_14_109 ();
 sg13g2_decap_8 FILLER_14_116 ();
 sg13g2_decap_8 FILLER_14_123 ();
 sg13g2_decap_8 FILLER_14_130 ();
 sg13g2_decap_8 FILLER_14_137 ();
 sg13g2_decap_8 FILLER_14_144 ();
 sg13g2_decap_8 FILLER_14_151 ();
 sg13g2_decap_8 FILLER_14_158 ();
 sg13g2_decap_8 FILLER_14_165 ();
 sg13g2_decap_8 FILLER_14_172 ();
 sg13g2_decap_8 FILLER_14_179 ();
 sg13g2_decap_8 FILLER_14_186 ();
 sg13g2_decap_8 FILLER_14_193 ();
 sg13g2_decap_8 FILLER_14_200 ();
 sg13g2_decap_8 FILLER_14_207 ();
 sg13g2_decap_8 FILLER_14_214 ();
 sg13g2_decap_8 FILLER_14_221 ();
 sg13g2_decap_8 FILLER_14_228 ();
 sg13g2_decap_8 FILLER_14_235 ();
 sg13g2_decap_8 FILLER_14_242 ();
 sg13g2_decap_8 FILLER_14_249 ();
 sg13g2_decap_8 FILLER_14_256 ();
 sg13g2_decap_8 FILLER_14_263 ();
 sg13g2_decap_8 FILLER_14_270 ();
 sg13g2_decap_8 FILLER_14_277 ();
 sg13g2_decap_8 FILLER_14_284 ();
 sg13g2_decap_8 FILLER_14_291 ();
 sg13g2_decap_8 FILLER_14_298 ();
 sg13g2_decap_8 FILLER_14_305 ();
 sg13g2_decap_8 FILLER_14_312 ();
 sg13g2_decap_8 FILLER_14_319 ();
 sg13g2_decap_8 FILLER_14_326 ();
 sg13g2_decap_8 FILLER_14_333 ();
 sg13g2_decap_8 FILLER_14_340 ();
 sg13g2_decap_8 FILLER_14_347 ();
 sg13g2_decap_8 FILLER_14_354 ();
 sg13g2_decap_8 FILLER_14_361 ();
 sg13g2_decap_8 FILLER_14_368 ();
 sg13g2_decap_8 FILLER_14_375 ();
 sg13g2_decap_8 FILLER_14_382 ();
 sg13g2_decap_8 FILLER_14_389 ();
 sg13g2_decap_8 FILLER_14_396 ();
 sg13g2_decap_8 FILLER_14_403 ();
 sg13g2_decap_8 FILLER_14_410 ();
 sg13g2_decap_8 FILLER_14_417 ();
 sg13g2_decap_8 FILLER_14_424 ();
 sg13g2_decap_8 FILLER_14_431 ();
 sg13g2_decap_8 FILLER_14_438 ();
 sg13g2_decap_8 FILLER_14_445 ();
 sg13g2_decap_8 FILLER_14_452 ();
 sg13g2_decap_8 FILLER_14_459 ();
 sg13g2_decap_8 FILLER_14_466 ();
 sg13g2_decap_8 FILLER_14_473 ();
 sg13g2_decap_8 FILLER_14_480 ();
 sg13g2_decap_8 FILLER_14_487 ();
 sg13g2_decap_8 FILLER_14_494 ();
 sg13g2_decap_8 FILLER_14_501 ();
 sg13g2_decap_8 FILLER_14_508 ();
 sg13g2_decap_8 FILLER_14_515 ();
 sg13g2_decap_8 FILLER_14_522 ();
 sg13g2_decap_8 FILLER_14_529 ();
 sg13g2_decap_8 FILLER_14_536 ();
 sg13g2_decap_8 FILLER_14_543 ();
 sg13g2_decap_8 FILLER_14_550 ();
 sg13g2_decap_8 FILLER_14_557 ();
 sg13g2_decap_8 FILLER_14_564 ();
 sg13g2_decap_8 FILLER_14_571 ();
 sg13g2_decap_8 FILLER_14_578 ();
 sg13g2_decap_8 FILLER_14_585 ();
 sg13g2_decap_8 FILLER_14_592 ();
 sg13g2_decap_8 FILLER_14_599 ();
 sg13g2_decap_8 FILLER_14_606 ();
 sg13g2_decap_8 FILLER_14_613 ();
 sg13g2_decap_8 FILLER_14_620 ();
 sg13g2_decap_8 FILLER_14_627 ();
 sg13g2_decap_8 FILLER_14_634 ();
 sg13g2_decap_8 FILLER_14_641 ();
 sg13g2_decap_8 FILLER_14_648 ();
 sg13g2_decap_8 FILLER_14_655 ();
 sg13g2_decap_8 FILLER_14_662 ();
 sg13g2_decap_8 FILLER_14_669 ();
 sg13g2_decap_8 FILLER_14_676 ();
 sg13g2_decap_8 FILLER_14_683 ();
 sg13g2_decap_8 FILLER_14_690 ();
 sg13g2_decap_8 FILLER_14_697 ();
 sg13g2_decap_8 FILLER_14_704 ();
 sg13g2_decap_8 FILLER_14_711 ();
 sg13g2_decap_8 FILLER_14_718 ();
 sg13g2_decap_8 FILLER_14_725 ();
 sg13g2_decap_8 FILLER_14_732 ();
 sg13g2_decap_8 FILLER_14_739 ();
 sg13g2_decap_8 FILLER_14_746 ();
 sg13g2_decap_8 FILLER_14_753 ();
 sg13g2_decap_8 FILLER_14_760 ();
 sg13g2_decap_8 FILLER_14_767 ();
 sg13g2_decap_8 FILLER_14_774 ();
 sg13g2_decap_8 FILLER_14_781 ();
 sg13g2_decap_8 FILLER_14_788 ();
 sg13g2_decap_8 FILLER_14_795 ();
 sg13g2_decap_8 FILLER_14_802 ();
 sg13g2_decap_8 FILLER_14_809 ();
 sg13g2_decap_8 FILLER_14_816 ();
 sg13g2_decap_8 FILLER_14_823 ();
 sg13g2_decap_8 FILLER_14_830 ();
 sg13g2_decap_8 FILLER_14_837 ();
 sg13g2_decap_8 FILLER_14_844 ();
 sg13g2_decap_8 FILLER_14_851 ();
 sg13g2_decap_8 FILLER_14_858 ();
 sg13g2_decap_8 FILLER_14_865 ();
 sg13g2_decap_8 FILLER_14_872 ();
 sg13g2_decap_8 FILLER_14_879 ();
 sg13g2_decap_8 FILLER_14_886 ();
 sg13g2_decap_8 FILLER_14_893 ();
 sg13g2_decap_8 FILLER_14_900 ();
 sg13g2_decap_8 FILLER_14_907 ();
 sg13g2_decap_8 FILLER_14_914 ();
 sg13g2_decap_8 FILLER_14_921 ();
 sg13g2_decap_8 FILLER_14_928 ();
 sg13g2_decap_8 FILLER_14_935 ();
 sg13g2_decap_8 FILLER_14_942 ();
 sg13g2_decap_8 FILLER_14_949 ();
 sg13g2_decap_8 FILLER_14_956 ();
 sg13g2_decap_8 FILLER_14_963 ();
 sg13g2_decap_8 FILLER_14_970 ();
 sg13g2_decap_8 FILLER_14_977 ();
 sg13g2_decap_8 FILLER_14_984 ();
 sg13g2_decap_8 FILLER_14_991 ();
 sg13g2_decap_8 FILLER_14_998 ();
 sg13g2_decap_8 FILLER_14_1005 ();
 sg13g2_decap_8 FILLER_14_1012 ();
 sg13g2_decap_8 FILLER_14_1019 ();
 sg13g2_fill_2 FILLER_14_1026 ();
 sg13g2_fill_1 FILLER_14_1028 ();
 sg13g2_decap_8 FILLER_15_4 ();
 sg13g2_decap_8 FILLER_15_11 ();
 sg13g2_decap_8 FILLER_15_18 ();
 sg13g2_decap_8 FILLER_15_25 ();
 sg13g2_decap_8 FILLER_15_32 ();
 sg13g2_decap_8 FILLER_15_39 ();
 sg13g2_decap_8 FILLER_15_46 ();
 sg13g2_decap_8 FILLER_15_53 ();
 sg13g2_decap_8 FILLER_15_60 ();
 sg13g2_decap_8 FILLER_15_67 ();
 sg13g2_decap_8 FILLER_15_74 ();
 sg13g2_decap_8 FILLER_15_81 ();
 sg13g2_decap_8 FILLER_15_88 ();
 sg13g2_decap_8 FILLER_15_95 ();
 sg13g2_decap_8 FILLER_15_102 ();
 sg13g2_decap_8 FILLER_15_109 ();
 sg13g2_decap_8 FILLER_15_116 ();
 sg13g2_decap_8 FILLER_15_123 ();
 sg13g2_decap_8 FILLER_15_130 ();
 sg13g2_decap_8 FILLER_15_137 ();
 sg13g2_decap_8 FILLER_15_144 ();
 sg13g2_decap_8 FILLER_15_151 ();
 sg13g2_decap_8 FILLER_15_158 ();
 sg13g2_decap_8 FILLER_15_165 ();
 sg13g2_decap_8 FILLER_15_172 ();
 sg13g2_decap_8 FILLER_15_179 ();
 sg13g2_decap_8 FILLER_15_186 ();
 sg13g2_decap_8 FILLER_15_193 ();
 sg13g2_decap_8 FILLER_15_200 ();
 sg13g2_decap_8 FILLER_15_207 ();
 sg13g2_decap_8 FILLER_15_214 ();
 sg13g2_decap_8 FILLER_15_221 ();
 sg13g2_decap_8 FILLER_15_228 ();
 sg13g2_decap_8 FILLER_15_235 ();
 sg13g2_decap_8 FILLER_15_242 ();
 sg13g2_decap_8 FILLER_15_249 ();
 sg13g2_decap_8 FILLER_15_256 ();
 sg13g2_decap_8 FILLER_15_263 ();
 sg13g2_decap_8 FILLER_15_270 ();
 sg13g2_decap_8 FILLER_15_277 ();
 sg13g2_decap_8 FILLER_15_284 ();
 sg13g2_decap_8 FILLER_15_291 ();
 sg13g2_decap_8 FILLER_15_298 ();
 sg13g2_decap_8 FILLER_15_305 ();
 sg13g2_decap_8 FILLER_15_312 ();
 sg13g2_decap_8 FILLER_15_319 ();
 sg13g2_decap_8 FILLER_15_326 ();
 sg13g2_decap_8 FILLER_15_333 ();
 sg13g2_decap_8 FILLER_15_340 ();
 sg13g2_decap_8 FILLER_15_347 ();
 sg13g2_decap_8 FILLER_15_354 ();
 sg13g2_decap_8 FILLER_15_361 ();
 sg13g2_decap_8 FILLER_15_368 ();
 sg13g2_decap_8 FILLER_15_375 ();
 sg13g2_decap_8 FILLER_15_382 ();
 sg13g2_decap_8 FILLER_15_389 ();
 sg13g2_decap_8 FILLER_15_396 ();
 sg13g2_decap_8 FILLER_15_403 ();
 sg13g2_decap_8 FILLER_15_410 ();
 sg13g2_decap_8 FILLER_15_417 ();
 sg13g2_decap_8 FILLER_15_424 ();
 sg13g2_decap_8 FILLER_15_431 ();
 sg13g2_decap_8 FILLER_15_438 ();
 sg13g2_decap_8 FILLER_15_445 ();
 sg13g2_decap_8 FILLER_15_452 ();
 sg13g2_decap_8 FILLER_15_459 ();
 sg13g2_decap_8 FILLER_15_466 ();
 sg13g2_decap_8 FILLER_15_473 ();
 sg13g2_decap_8 FILLER_15_480 ();
 sg13g2_decap_8 FILLER_15_487 ();
 sg13g2_decap_8 FILLER_15_494 ();
 sg13g2_decap_8 FILLER_15_501 ();
 sg13g2_decap_8 FILLER_15_508 ();
 sg13g2_decap_8 FILLER_15_515 ();
 sg13g2_decap_8 FILLER_15_522 ();
 sg13g2_decap_8 FILLER_15_529 ();
 sg13g2_decap_8 FILLER_15_536 ();
 sg13g2_decap_8 FILLER_15_543 ();
 sg13g2_decap_8 FILLER_15_550 ();
 sg13g2_decap_8 FILLER_15_557 ();
 sg13g2_decap_8 FILLER_15_564 ();
 sg13g2_decap_8 FILLER_15_571 ();
 sg13g2_decap_8 FILLER_15_578 ();
 sg13g2_decap_8 FILLER_15_585 ();
 sg13g2_decap_8 FILLER_15_592 ();
 sg13g2_decap_8 FILLER_15_599 ();
 sg13g2_decap_8 FILLER_15_606 ();
 sg13g2_decap_8 FILLER_15_613 ();
 sg13g2_decap_8 FILLER_15_620 ();
 sg13g2_decap_8 FILLER_15_627 ();
 sg13g2_decap_8 FILLER_15_634 ();
 sg13g2_decap_8 FILLER_15_641 ();
 sg13g2_decap_8 FILLER_15_648 ();
 sg13g2_decap_8 FILLER_15_655 ();
 sg13g2_decap_8 FILLER_15_662 ();
 sg13g2_decap_8 FILLER_15_669 ();
 sg13g2_decap_8 FILLER_15_676 ();
 sg13g2_decap_8 FILLER_15_683 ();
 sg13g2_decap_8 FILLER_15_690 ();
 sg13g2_decap_8 FILLER_15_697 ();
 sg13g2_decap_8 FILLER_15_704 ();
 sg13g2_decap_8 FILLER_15_711 ();
 sg13g2_decap_8 FILLER_15_718 ();
 sg13g2_decap_8 FILLER_15_725 ();
 sg13g2_decap_8 FILLER_15_732 ();
 sg13g2_decap_8 FILLER_15_739 ();
 sg13g2_decap_8 FILLER_15_746 ();
 sg13g2_decap_8 FILLER_15_753 ();
 sg13g2_decap_8 FILLER_15_760 ();
 sg13g2_decap_8 FILLER_15_767 ();
 sg13g2_decap_8 FILLER_15_774 ();
 sg13g2_decap_8 FILLER_15_781 ();
 sg13g2_decap_8 FILLER_15_788 ();
 sg13g2_decap_8 FILLER_15_795 ();
 sg13g2_decap_8 FILLER_15_802 ();
 sg13g2_decap_8 FILLER_15_809 ();
 sg13g2_decap_8 FILLER_15_816 ();
 sg13g2_decap_8 FILLER_15_823 ();
 sg13g2_decap_8 FILLER_15_830 ();
 sg13g2_decap_8 FILLER_15_837 ();
 sg13g2_decap_8 FILLER_15_844 ();
 sg13g2_decap_8 FILLER_15_851 ();
 sg13g2_decap_8 FILLER_15_858 ();
 sg13g2_decap_8 FILLER_15_865 ();
 sg13g2_decap_8 FILLER_15_872 ();
 sg13g2_decap_8 FILLER_15_879 ();
 sg13g2_decap_8 FILLER_15_886 ();
 sg13g2_decap_8 FILLER_15_893 ();
 sg13g2_decap_8 FILLER_15_900 ();
 sg13g2_decap_8 FILLER_15_907 ();
 sg13g2_decap_8 FILLER_15_914 ();
 sg13g2_decap_8 FILLER_15_921 ();
 sg13g2_decap_8 FILLER_15_928 ();
 sg13g2_decap_8 FILLER_15_935 ();
 sg13g2_decap_8 FILLER_15_942 ();
 sg13g2_decap_8 FILLER_15_949 ();
 sg13g2_decap_8 FILLER_15_956 ();
 sg13g2_decap_8 FILLER_15_963 ();
 sg13g2_decap_8 FILLER_15_970 ();
 sg13g2_decap_8 FILLER_15_977 ();
 sg13g2_decap_8 FILLER_15_984 ();
 sg13g2_decap_8 FILLER_15_991 ();
 sg13g2_decap_8 FILLER_15_998 ();
 sg13g2_decap_8 FILLER_15_1005 ();
 sg13g2_decap_8 FILLER_15_1012 ();
 sg13g2_decap_8 FILLER_15_1019 ();
 sg13g2_fill_2 FILLER_15_1026 ();
 sg13g2_fill_1 FILLER_15_1028 ();
 sg13g2_decap_8 FILLER_16_4 ();
 sg13g2_decap_8 FILLER_16_11 ();
 sg13g2_decap_8 FILLER_16_18 ();
 sg13g2_decap_8 FILLER_16_25 ();
 sg13g2_decap_8 FILLER_16_32 ();
 sg13g2_decap_8 FILLER_16_39 ();
 sg13g2_decap_8 FILLER_16_46 ();
 sg13g2_decap_8 FILLER_16_53 ();
 sg13g2_decap_8 FILLER_16_60 ();
 sg13g2_decap_8 FILLER_16_67 ();
 sg13g2_decap_8 FILLER_16_74 ();
 sg13g2_decap_8 FILLER_16_81 ();
 sg13g2_decap_8 FILLER_16_88 ();
 sg13g2_decap_8 FILLER_16_95 ();
 sg13g2_decap_8 FILLER_16_102 ();
 sg13g2_decap_8 FILLER_16_109 ();
 sg13g2_decap_8 FILLER_16_116 ();
 sg13g2_decap_8 FILLER_16_123 ();
 sg13g2_decap_8 FILLER_16_130 ();
 sg13g2_decap_8 FILLER_16_137 ();
 sg13g2_decap_8 FILLER_16_144 ();
 sg13g2_decap_8 FILLER_16_151 ();
 sg13g2_decap_8 FILLER_16_158 ();
 sg13g2_decap_8 FILLER_16_165 ();
 sg13g2_decap_8 FILLER_16_172 ();
 sg13g2_decap_8 FILLER_16_179 ();
 sg13g2_decap_8 FILLER_16_186 ();
 sg13g2_decap_8 FILLER_16_193 ();
 sg13g2_decap_8 FILLER_16_200 ();
 sg13g2_decap_8 FILLER_16_207 ();
 sg13g2_decap_8 FILLER_16_214 ();
 sg13g2_decap_8 FILLER_16_221 ();
 sg13g2_decap_8 FILLER_16_228 ();
 sg13g2_decap_8 FILLER_16_235 ();
 sg13g2_decap_8 FILLER_16_242 ();
 sg13g2_decap_8 FILLER_16_249 ();
 sg13g2_decap_8 FILLER_16_256 ();
 sg13g2_decap_8 FILLER_16_263 ();
 sg13g2_decap_8 FILLER_16_270 ();
 sg13g2_decap_8 FILLER_16_277 ();
 sg13g2_decap_8 FILLER_16_284 ();
 sg13g2_decap_8 FILLER_16_291 ();
 sg13g2_decap_8 FILLER_16_298 ();
 sg13g2_decap_8 FILLER_16_305 ();
 sg13g2_decap_8 FILLER_16_312 ();
 sg13g2_decap_8 FILLER_16_319 ();
 sg13g2_decap_8 FILLER_16_326 ();
 sg13g2_decap_8 FILLER_16_333 ();
 sg13g2_decap_8 FILLER_16_340 ();
 sg13g2_decap_8 FILLER_16_347 ();
 sg13g2_decap_8 FILLER_16_354 ();
 sg13g2_decap_8 FILLER_16_361 ();
 sg13g2_decap_8 FILLER_16_368 ();
 sg13g2_decap_8 FILLER_16_375 ();
 sg13g2_decap_8 FILLER_16_382 ();
 sg13g2_decap_8 FILLER_16_389 ();
 sg13g2_decap_8 FILLER_16_396 ();
 sg13g2_decap_8 FILLER_16_403 ();
 sg13g2_decap_8 FILLER_16_410 ();
 sg13g2_decap_8 FILLER_16_417 ();
 sg13g2_decap_8 FILLER_16_424 ();
 sg13g2_decap_8 FILLER_16_431 ();
 sg13g2_decap_8 FILLER_16_438 ();
 sg13g2_decap_8 FILLER_16_445 ();
 sg13g2_decap_8 FILLER_16_452 ();
 sg13g2_decap_8 FILLER_16_459 ();
 sg13g2_decap_8 FILLER_16_466 ();
 sg13g2_decap_8 FILLER_16_473 ();
 sg13g2_decap_8 FILLER_16_480 ();
 sg13g2_decap_8 FILLER_16_487 ();
 sg13g2_decap_8 FILLER_16_494 ();
 sg13g2_decap_8 FILLER_16_501 ();
 sg13g2_decap_8 FILLER_16_508 ();
 sg13g2_decap_8 FILLER_16_515 ();
 sg13g2_decap_8 FILLER_16_522 ();
 sg13g2_decap_8 FILLER_16_529 ();
 sg13g2_decap_8 FILLER_16_536 ();
 sg13g2_decap_8 FILLER_16_543 ();
 sg13g2_decap_8 FILLER_16_550 ();
 sg13g2_decap_8 FILLER_16_557 ();
 sg13g2_decap_8 FILLER_16_564 ();
 sg13g2_decap_8 FILLER_16_571 ();
 sg13g2_decap_8 FILLER_16_578 ();
 sg13g2_decap_8 FILLER_16_585 ();
 sg13g2_decap_8 FILLER_16_592 ();
 sg13g2_decap_8 FILLER_16_599 ();
 sg13g2_decap_8 FILLER_16_606 ();
 sg13g2_decap_8 FILLER_16_613 ();
 sg13g2_decap_8 FILLER_16_620 ();
 sg13g2_decap_8 FILLER_16_627 ();
 sg13g2_decap_8 FILLER_16_634 ();
 sg13g2_decap_8 FILLER_16_641 ();
 sg13g2_decap_8 FILLER_16_648 ();
 sg13g2_decap_8 FILLER_16_655 ();
 sg13g2_decap_8 FILLER_16_662 ();
 sg13g2_decap_8 FILLER_16_669 ();
 sg13g2_decap_8 FILLER_16_676 ();
 sg13g2_decap_8 FILLER_16_683 ();
 sg13g2_decap_8 FILLER_16_690 ();
 sg13g2_decap_8 FILLER_16_697 ();
 sg13g2_decap_8 FILLER_16_704 ();
 sg13g2_decap_8 FILLER_16_711 ();
 sg13g2_decap_8 FILLER_16_718 ();
 sg13g2_decap_8 FILLER_16_725 ();
 sg13g2_decap_8 FILLER_16_732 ();
 sg13g2_decap_8 FILLER_16_739 ();
 sg13g2_decap_8 FILLER_16_746 ();
 sg13g2_decap_8 FILLER_16_753 ();
 sg13g2_decap_8 FILLER_16_760 ();
 sg13g2_decap_8 FILLER_16_767 ();
 sg13g2_decap_8 FILLER_16_774 ();
 sg13g2_decap_8 FILLER_16_781 ();
 sg13g2_decap_8 FILLER_16_788 ();
 sg13g2_decap_8 FILLER_16_795 ();
 sg13g2_decap_8 FILLER_16_802 ();
 sg13g2_decap_8 FILLER_16_809 ();
 sg13g2_decap_8 FILLER_16_816 ();
 sg13g2_decap_8 FILLER_16_823 ();
 sg13g2_decap_8 FILLER_16_830 ();
 sg13g2_decap_8 FILLER_16_837 ();
 sg13g2_decap_8 FILLER_16_844 ();
 sg13g2_decap_8 FILLER_16_851 ();
 sg13g2_decap_8 FILLER_16_858 ();
 sg13g2_decap_8 FILLER_16_865 ();
 sg13g2_decap_8 FILLER_16_872 ();
 sg13g2_decap_8 FILLER_16_879 ();
 sg13g2_decap_8 FILLER_16_886 ();
 sg13g2_decap_8 FILLER_16_893 ();
 sg13g2_decap_8 FILLER_16_900 ();
 sg13g2_decap_8 FILLER_16_907 ();
 sg13g2_decap_8 FILLER_16_914 ();
 sg13g2_decap_8 FILLER_16_921 ();
 sg13g2_decap_8 FILLER_16_928 ();
 sg13g2_decap_8 FILLER_16_935 ();
 sg13g2_decap_8 FILLER_16_942 ();
 sg13g2_decap_8 FILLER_16_949 ();
 sg13g2_decap_8 FILLER_16_956 ();
 sg13g2_decap_8 FILLER_16_963 ();
 sg13g2_decap_8 FILLER_16_970 ();
 sg13g2_decap_8 FILLER_16_977 ();
 sg13g2_decap_8 FILLER_16_984 ();
 sg13g2_decap_8 FILLER_16_991 ();
 sg13g2_decap_8 FILLER_16_998 ();
 sg13g2_decap_8 FILLER_16_1005 ();
 sg13g2_decap_8 FILLER_16_1012 ();
 sg13g2_decap_8 FILLER_16_1019 ();
 sg13g2_fill_2 FILLER_16_1026 ();
 sg13g2_fill_1 FILLER_16_1028 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_decap_8 FILLER_17_427 ();
 sg13g2_decap_8 FILLER_17_434 ();
 sg13g2_decap_8 FILLER_17_441 ();
 sg13g2_decap_8 FILLER_17_448 ();
 sg13g2_decap_8 FILLER_17_455 ();
 sg13g2_decap_8 FILLER_17_462 ();
 sg13g2_decap_8 FILLER_17_469 ();
 sg13g2_decap_8 FILLER_17_476 ();
 sg13g2_decap_8 FILLER_17_483 ();
 sg13g2_decap_8 FILLER_17_490 ();
 sg13g2_decap_8 FILLER_17_497 ();
 sg13g2_decap_8 FILLER_17_504 ();
 sg13g2_decap_8 FILLER_17_511 ();
 sg13g2_decap_8 FILLER_17_518 ();
 sg13g2_decap_8 FILLER_17_525 ();
 sg13g2_decap_8 FILLER_17_532 ();
 sg13g2_decap_8 FILLER_17_539 ();
 sg13g2_decap_8 FILLER_17_546 ();
 sg13g2_decap_8 FILLER_17_553 ();
 sg13g2_decap_8 FILLER_17_560 ();
 sg13g2_decap_8 FILLER_17_567 ();
 sg13g2_decap_8 FILLER_17_574 ();
 sg13g2_decap_8 FILLER_17_581 ();
 sg13g2_decap_8 FILLER_17_588 ();
 sg13g2_decap_8 FILLER_17_595 ();
 sg13g2_decap_8 FILLER_17_602 ();
 sg13g2_decap_8 FILLER_17_609 ();
 sg13g2_decap_8 FILLER_17_616 ();
 sg13g2_decap_8 FILLER_17_623 ();
 sg13g2_decap_8 FILLER_17_630 ();
 sg13g2_decap_8 FILLER_17_637 ();
 sg13g2_decap_8 FILLER_17_644 ();
 sg13g2_decap_8 FILLER_17_651 ();
 sg13g2_decap_8 FILLER_17_658 ();
 sg13g2_decap_8 FILLER_17_665 ();
 sg13g2_decap_8 FILLER_17_672 ();
 sg13g2_decap_8 FILLER_17_679 ();
 sg13g2_decap_8 FILLER_17_686 ();
 sg13g2_decap_8 FILLER_17_693 ();
 sg13g2_decap_8 FILLER_17_700 ();
 sg13g2_decap_8 FILLER_17_707 ();
 sg13g2_decap_8 FILLER_17_714 ();
 sg13g2_decap_8 FILLER_17_721 ();
 sg13g2_decap_8 FILLER_17_728 ();
 sg13g2_decap_8 FILLER_17_735 ();
 sg13g2_decap_8 FILLER_17_742 ();
 sg13g2_decap_8 FILLER_17_749 ();
 sg13g2_decap_8 FILLER_17_756 ();
 sg13g2_decap_8 FILLER_17_763 ();
 sg13g2_decap_8 FILLER_17_770 ();
 sg13g2_decap_8 FILLER_17_777 ();
 sg13g2_decap_8 FILLER_17_784 ();
 sg13g2_decap_8 FILLER_17_791 ();
 sg13g2_decap_8 FILLER_17_798 ();
 sg13g2_decap_8 FILLER_17_805 ();
 sg13g2_decap_8 FILLER_17_812 ();
 sg13g2_decap_8 FILLER_17_819 ();
 sg13g2_decap_8 FILLER_17_826 ();
 sg13g2_decap_8 FILLER_17_833 ();
 sg13g2_decap_8 FILLER_17_840 ();
 sg13g2_decap_8 FILLER_17_847 ();
 sg13g2_decap_8 FILLER_17_854 ();
 sg13g2_decap_8 FILLER_17_861 ();
 sg13g2_decap_8 FILLER_17_868 ();
 sg13g2_decap_8 FILLER_17_875 ();
 sg13g2_decap_8 FILLER_17_882 ();
 sg13g2_decap_8 FILLER_17_889 ();
 sg13g2_decap_8 FILLER_17_896 ();
 sg13g2_decap_8 FILLER_17_903 ();
 sg13g2_decap_8 FILLER_17_910 ();
 sg13g2_decap_8 FILLER_17_917 ();
 sg13g2_decap_8 FILLER_17_924 ();
 sg13g2_decap_8 FILLER_17_931 ();
 sg13g2_decap_8 FILLER_17_938 ();
 sg13g2_decap_8 FILLER_17_945 ();
 sg13g2_decap_8 FILLER_17_952 ();
 sg13g2_decap_8 FILLER_17_959 ();
 sg13g2_decap_8 FILLER_17_966 ();
 sg13g2_decap_8 FILLER_17_973 ();
 sg13g2_decap_8 FILLER_17_980 ();
 sg13g2_decap_8 FILLER_17_987 ();
 sg13g2_decap_8 FILLER_17_994 ();
 sg13g2_decap_8 FILLER_17_1001 ();
 sg13g2_decap_8 FILLER_17_1008 ();
 sg13g2_decap_8 FILLER_17_1015 ();
 sg13g2_decap_8 FILLER_17_1022 ();
 sg13g2_decap_8 FILLER_18_4 ();
 sg13g2_decap_8 FILLER_18_11 ();
 sg13g2_decap_8 FILLER_18_18 ();
 sg13g2_decap_8 FILLER_18_25 ();
 sg13g2_decap_8 FILLER_18_32 ();
 sg13g2_decap_8 FILLER_18_39 ();
 sg13g2_decap_8 FILLER_18_46 ();
 sg13g2_decap_8 FILLER_18_53 ();
 sg13g2_decap_8 FILLER_18_60 ();
 sg13g2_decap_8 FILLER_18_67 ();
 sg13g2_decap_8 FILLER_18_74 ();
 sg13g2_decap_8 FILLER_18_81 ();
 sg13g2_decap_8 FILLER_18_88 ();
 sg13g2_decap_8 FILLER_18_95 ();
 sg13g2_decap_8 FILLER_18_102 ();
 sg13g2_decap_8 FILLER_18_109 ();
 sg13g2_decap_8 FILLER_18_116 ();
 sg13g2_decap_8 FILLER_18_123 ();
 sg13g2_decap_8 FILLER_18_130 ();
 sg13g2_decap_8 FILLER_18_137 ();
 sg13g2_decap_8 FILLER_18_144 ();
 sg13g2_decap_8 FILLER_18_151 ();
 sg13g2_decap_8 FILLER_18_158 ();
 sg13g2_decap_8 FILLER_18_165 ();
 sg13g2_decap_8 FILLER_18_172 ();
 sg13g2_decap_8 FILLER_18_179 ();
 sg13g2_decap_8 FILLER_18_186 ();
 sg13g2_decap_8 FILLER_18_193 ();
 sg13g2_decap_8 FILLER_18_200 ();
 sg13g2_decap_8 FILLER_18_207 ();
 sg13g2_decap_8 FILLER_18_214 ();
 sg13g2_decap_8 FILLER_18_221 ();
 sg13g2_decap_8 FILLER_18_228 ();
 sg13g2_decap_8 FILLER_18_235 ();
 sg13g2_decap_8 FILLER_18_242 ();
 sg13g2_decap_8 FILLER_18_249 ();
 sg13g2_decap_8 FILLER_18_256 ();
 sg13g2_decap_8 FILLER_18_263 ();
 sg13g2_decap_8 FILLER_18_270 ();
 sg13g2_decap_8 FILLER_18_277 ();
 sg13g2_decap_8 FILLER_18_284 ();
 sg13g2_decap_8 FILLER_18_291 ();
 sg13g2_decap_8 FILLER_18_298 ();
 sg13g2_decap_8 FILLER_18_305 ();
 sg13g2_decap_8 FILLER_18_312 ();
 sg13g2_decap_8 FILLER_18_319 ();
 sg13g2_decap_8 FILLER_18_326 ();
 sg13g2_decap_8 FILLER_18_333 ();
 sg13g2_decap_8 FILLER_18_340 ();
 sg13g2_decap_8 FILLER_18_347 ();
 sg13g2_decap_8 FILLER_18_354 ();
 sg13g2_decap_8 FILLER_18_361 ();
 sg13g2_decap_8 FILLER_18_368 ();
 sg13g2_decap_8 FILLER_18_375 ();
 sg13g2_decap_8 FILLER_18_382 ();
 sg13g2_decap_8 FILLER_18_389 ();
 sg13g2_decap_8 FILLER_18_396 ();
 sg13g2_decap_8 FILLER_18_403 ();
 sg13g2_decap_8 FILLER_18_410 ();
 sg13g2_decap_8 FILLER_18_417 ();
 sg13g2_decap_8 FILLER_18_424 ();
 sg13g2_decap_8 FILLER_18_431 ();
 sg13g2_decap_8 FILLER_18_438 ();
 sg13g2_decap_8 FILLER_18_445 ();
 sg13g2_decap_8 FILLER_18_452 ();
 sg13g2_decap_8 FILLER_18_459 ();
 sg13g2_decap_8 FILLER_18_466 ();
 sg13g2_decap_8 FILLER_18_473 ();
 sg13g2_decap_8 FILLER_18_480 ();
 sg13g2_decap_8 FILLER_18_487 ();
 sg13g2_decap_8 FILLER_18_494 ();
 sg13g2_decap_8 FILLER_18_501 ();
 sg13g2_decap_8 FILLER_18_508 ();
 sg13g2_decap_8 FILLER_18_515 ();
 sg13g2_decap_8 FILLER_18_522 ();
 sg13g2_decap_8 FILLER_18_529 ();
 sg13g2_decap_8 FILLER_18_536 ();
 sg13g2_decap_8 FILLER_18_543 ();
 sg13g2_decap_8 FILLER_18_550 ();
 sg13g2_decap_8 FILLER_18_557 ();
 sg13g2_decap_8 FILLER_18_564 ();
 sg13g2_decap_8 FILLER_18_571 ();
 sg13g2_decap_8 FILLER_18_578 ();
 sg13g2_decap_8 FILLER_18_585 ();
 sg13g2_decap_8 FILLER_18_592 ();
 sg13g2_decap_8 FILLER_18_599 ();
 sg13g2_decap_8 FILLER_18_606 ();
 sg13g2_decap_8 FILLER_18_613 ();
 sg13g2_decap_8 FILLER_18_620 ();
 sg13g2_decap_8 FILLER_18_627 ();
 sg13g2_decap_8 FILLER_18_634 ();
 sg13g2_decap_8 FILLER_18_641 ();
 sg13g2_decap_8 FILLER_18_648 ();
 sg13g2_decap_8 FILLER_18_655 ();
 sg13g2_decap_8 FILLER_18_662 ();
 sg13g2_decap_8 FILLER_18_669 ();
 sg13g2_decap_8 FILLER_18_676 ();
 sg13g2_decap_8 FILLER_18_683 ();
 sg13g2_decap_8 FILLER_18_690 ();
 sg13g2_decap_8 FILLER_18_697 ();
 sg13g2_decap_8 FILLER_18_704 ();
 sg13g2_decap_8 FILLER_18_711 ();
 sg13g2_decap_8 FILLER_18_718 ();
 sg13g2_decap_8 FILLER_18_725 ();
 sg13g2_decap_8 FILLER_18_732 ();
 sg13g2_decap_8 FILLER_18_739 ();
 sg13g2_decap_8 FILLER_18_746 ();
 sg13g2_decap_8 FILLER_18_753 ();
 sg13g2_decap_8 FILLER_18_760 ();
 sg13g2_decap_8 FILLER_18_767 ();
 sg13g2_decap_8 FILLER_18_774 ();
 sg13g2_decap_8 FILLER_18_781 ();
 sg13g2_decap_8 FILLER_18_788 ();
 sg13g2_decap_8 FILLER_18_795 ();
 sg13g2_decap_8 FILLER_18_802 ();
 sg13g2_decap_8 FILLER_18_809 ();
 sg13g2_decap_8 FILLER_18_816 ();
 sg13g2_decap_8 FILLER_18_823 ();
 sg13g2_decap_8 FILLER_18_830 ();
 sg13g2_decap_8 FILLER_18_837 ();
 sg13g2_decap_8 FILLER_18_844 ();
 sg13g2_decap_8 FILLER_18_851 ();
 sg13g2_decap_8 FILLER_18_858 ();
 sg13g2_decap_8 FILLER_18_865 ();
 sg13g2_decap_8 FILLER_18_872 ();
 sg13g2_decap_8 FILLER_18_879 ();
 sg13g2_decap_8 FILLER_18_886 ();
 sg13g2_decap_8 FILLER_18_893 ();
 sg13g2_decap_8 FILLER_18_900 ();
 sg13g2_decap_8 FILLER_18_907 ();
 sg13g2_decap_8 FILLER_18_914 ();
 sg13g2_decap_8 FILLER_18_921 ();
 sg13g2_decap_8 FILLER_18_928 ();
 sg13g2_decap_8 FILLER_18_935 ();
 sg13g2_decap_8 FILLER_18_942 ();
 sg13g2_decap_8 FILLER_18_949 ();
 sg13g2_decap_8 FILLER_18_956 ();
 sg13g2_decap_8 FILLER_18_963 ();
 sg13g2_decap_8 FILLER_18_970 ();
 sg13g2_decap_8 FILLER_18_977 ();
 sg13g2_decap_8 FILLER_18_984 ();
 sg13g2_decap_8 FILLER_18_991 ();
 sg13g2_decap_8 FILLER_18_998 ();
 sg13g2_decap_8 FILLER_18_1005 ();
 sg13g2_decap_8 FILLER_18_1012 ();
 sg13g2_decap_8 FILLER_18_1019 ();
 sg13g2_fill_2 FILLER_18_1026 ();
 sg13g2_fill_1 FILLER_18_1028 ();
 sg13g2_decap_8 FILLER_19_4 ();
 sg13g2_decap_8 FILLER_19_11 ();
 sg13g2_decap_8 FILLER_19_18 ();
 sg13g2_decap_8 FILLER_19_25 ();
 sg13g2_decap_8 FILLER_19_32 ();
 sg13g2_decap_8 FILLER_19_39 ();
 sg13g2_decap_8 FILLER_19_46 ();
 sg13g2_decap_8 FILLER_19_53 ();
 sg13g2_decap_8 FILLER_19_60 ();
 sg13g2_decap_8 FILLER_19_67 ();
 sg13g2_decap_8 FILLER_19_74 ();
 sg13g2_decap_8 FILLER_19_81 ();
 sg13g2_decap_8 FILLER_19_88 ();
 sg13g2_decap_8 FILLER_19_95 ();
 sg13g2_decap_8 FILLER_19_102 ();
 sg13g2_decap_8 FILLER_19_109 ();
 sg13g2_decap_8 FILLER_19_116 ();
 sg13g2_decap_8 FILLER_19_123 ();
 sg13g2_decap_8 FILLER_19_130 ();
 sg13g2_decap_8 FILLER_19_137 ();
 sg13g2_decap_8 FILLER_19_144 ();
 sg13g2_decap_8 FILLER_19_151 ();
 sg13g2_decap_8 FILLER_19_158 ();
 sg13g2_decap_8 FILLER_19_165 ();
 sg13g2_decap_8 FILLER_19_172 ();
 sg13g2_decap_8 FILLER_19_179 ();
 sg13g2_decap_8 FILLER_19_186 ();
 sg13g2_decap_8 FILLER_19_193 ();
 sg13g2_decap_8 FILLER_19_200 ();
 sg13g2_decap_8 FILLER_19_207 ();
 sg13g2_decap_8 FILLER_19_214 ();
 sg13g2_decap_8 FILLER_19_221 ();
 sg13g2_decap_8 FILLER_19_228 ();
 sg13g2_decap_8 FILLER_19_235 ();
 sg13g2_decap_8 FILLER_19_242 ();
 sg13g2_decap_8 FILLER_19_249 ();
 sg13g2_decap_8 FILLER_19_256 ();
 sg13g2_decap_8 FILLER_19_263 ();
 sg13g2_decap_8 FILLER_19_270 ();
 sg13g2_decap_8 FILLER_19_277 ();
 sg13g2_decap_8 FILLER_19_284 ();
 sg13g2_decap_8 FILLER_19_291 ();
 sg13g2_decap_8 FILLER_19_298 ();
 sg13g2_decap_8 FILLER_19_305 ();
 sg13g2_decap_8 FILLER_19_312 ();
 sg13g2_decap_8 FILLER_19_319 ();
 sg13g2_decap_8 FILLER_19_326 ();
 sg13g2_decap_8 FILLER_19_333 ();
 sg13g2_decap_8 FILLER_19_340 ();
 sg13g2_decap_8 FILLER_19_347 ();
 sg13g2_decap_8 FILLER_19_354 ();
 sg13g2_decap_8 FILLER_19_361 ();
 sg13g2_decap_8 FILLER_19_368 ();
 sg13g2_decap_8 FILLER_19_375 ();
 sg13g2_decap_8 FILLER_19_382 ();
 sg13g2_decap_8 FILLER_19_389 ();
 sg13g2_decap_8 FILLER_19_396 ();
 sg13g2_decap_8 FILLER_19_403 ();
 sg13g2_decap_8 FILLER_19_410 ();
 sg13g2_decap_8 FILLER_19_417 ();
 sg13g2_decap_8 FILLER_19_424 ();
 sg13g2_decap_8 FILLER_19_431 ();
 sg13g2_decap_8 FILLER_19_438 ();
 sg13g2_decap_8 FILLER_19_445 ();
 sg13g2_decap_8 FILLER_19_452 ();
 sg13g2_decap_8 FILLER_19_459 ();
 sg13g2_decap_8 FILLER_19_466 ();
 sg13g2_decap_8 FILLER_19_473 ();
 sg13g2_decap_8 FILLER_19_480 ();
 sg13g2_decap_8 FILLER_19_487 ();
 sg13g2_decap_8 FILLER_19_494 ();
 sg13g2_decap_8 FILLER_19_501 ();
 sg13g2_decap_8 FILLER_19_508 ();
 sg13g2_decap_8 FILLER_19_515 ();
 sg13g2_decap_8 FILLER_19_522 ();
 sg13g2_decap_8 FILLER_19_529 ();
 sg13g2_decap_8 FILLER_19_536 ();
 sg13g2_decap_8 FILLER_19_543 ();
 sg13g2_decap_8 FILLER_19_550 ();
 sg13g2_decap_8 FILLER_19_557 ();
 sg13g2_decap_8 FILLER_19_564 ();
 sg13g2_decap_8 FILLER_19_571 ();
 sg13g2_decap_8 FILLER_19_578 ();
 sg13g2_decap_8 FILLER_19_585 ();
 sg13g2_decap_8 FILLER_19_592 ();
 sg13g2_decap_8 FILLER_19_599 ();
 sg13g2_decap_8 FILLER_19_606 ();
 sg13g2_decap_8 FILLER_19_613 ();
 sg13g2_decap_8 FILLER_19_620 ();
 sg13g2_decap_8 FILLER_19_627 ();
 sg13g2_decap_8 FILLER_19_634 ();
 sg13g2_decap_8 FILLER_19_641 ();
 sg13g2_decap_8 FILLER_19_648 ();
 sg13g2_decap_8 FILLER_19_655 ();
 sg13g2_decap_8 FILLER_19_662 ();
 sg13g2_decap_8 FILLER_19_669 ();
 sg13g2_decap_8 FILLER_19_676 ();
 sg13g2_decap_8 FILLER_19_683 ();
 sg13g2_decap_8 FILLER_19_690 ();
 sg13g2_decap_8 FILLER_19_697 ();
 sg13g2_decap_8 FILLER_19_704 ();
 sg13g2_decap_8 FILLER_19_711 ();
 sg13g2_decap_8 FILLER_19_718 ();
 sg13g2_decap_8 FILLER_19_725 ();
 sg13g2_decap_8 FILLER_19_732 ();
 sg13g2_decap_8 FILLER_19_739 ();
 sg13g2_decap_8 FILLER_19_746 ();
 sg13g2_decap_8 FILLER_19_753 ();
 sg13g2_decap_8 FILLER_19_760 ();
 sg13g2_decap_8 FILLER_19_767 ();
 sg13g2_decap_8 FILLER_19_774 ();
 sg13g2_decap_8 FILLER_19_781 ();
 sg13g2_decap_8 FILLER_19_788 ();
 sg13g2_decap_8 FILLER_19_795 ();
 sg13g2_decap_8 FILLER_19_802 ();
 sg13g2_decap_8 FILLER_19_809 ();
 sg13g2_decap_8 FILLER_19_816 ();
 sg13g2_decap_8 FILLER_19_823 ();
 sg13g2_decap_8 FILLER_19_830 ();
 sg13g2_decap_8 FILLER_19_837 ();
 sg13g2_decap_8 FILLER_19_844 ();
 sg13g2_decap_8 FILLER_19_851 ();
 sg13g2_decap_8 FILLER_19_858 ();
 sg13g2_decap_8 FILLER_19_865 ();
 sg13g2_decap_8 FILLER_19_872 ();
 sg13g2_decap_8 FILLER_19_879 ();
 sg13g2_decap_8 FILLER_19_886 ();
 sg13g2_decap_8 FILLER_19_893 ();
 sg13g2_decap_8 FILLER_19_900 ();
 sg13g2_decap_8 FILLER_19_907 ();
 sg13g2_decap_8 FILLER_19_914 ();
 sg13g2_decap_8 FILLER_19_921 ();
 sg13g2_decap_8 FILLER_19_928 ();
 sg13g2_decap_8 FILLER_19_935 ();
 sg13g2_decap_8 FILLER_19_942 ();
 sg13g2_decap_8 FILLER_19_949 ();
 sg13g2_decap_8 FILLER_19_956 ();
 sg13g2_decap_8 FILLER_19_963 ();
 sg13g2_decap_8 FILLER_19_970 ();
 sg13g2_decap_8 FILLER_19_977 ();
 sg13g2_decap_8 FILLER_19_984 ();
 sg13g2_decap_8 FILLER_19_991 ();
 sg13g2_decap_8 FILLER_19_998 ();
 sg13g2_decap_8 FILLER_19_1005 ();
 sg13g2_decap_8 FILLER_19_1012 ();
 sg13g2_decap_8 FILLER_19_1019 ();
 sg13g2_fill_2 FILLER_19_1026 ();
 sg13g2_fill_1 FILLER_19_1028 ();
 sg13g2_decap_8 FILLER_20_4 ();
 sg13g2_decap_8 FILLER_20_11 ();
 sg13g2_decap_8 FILLER_20_18 ();
 sg13g2_decap_8 FILLER_20_25 ();
 sg13g2_decap_8 FILLER_20_32 ();
 sg13g2_decap_8 FILLER_20_39 ();
 sg13g2_decap_8 FILLER_20_46 ();
 sg13g2_decap_8 FILLER_20_53 ();
 sg13g2_decap_8 FILLER_20_60 ();
 sg13g2_decap_8 FILLER_20_67 ();
 sg13g2_decap_8 FILLER_20_74 ();
 sg13g2_decap_8 FILLER_20_81 ();
 sg13g2_decap_8 FILLER_20_88 ();
 sg13g2_decap_8 FILLER_20_95 ();
 sg13g2_decap_8 FILLER_20_102 ();
 sg13g2_decap_8 FILLER_20_109 ();
 sg13g2_decap_8 FILLER_20_116 ();
 sg13g2_decap_8 FILLER_20_123 ();
 sg13g2_decap_8 FILLER_20_130 ();
 sg13g2_decap_8 FILLER_20_137 ();
 sg13g2_decap_8 FILLER_20_144 ();
 sg13g2_decap_8 FILLER_20_151 ();
 sg13g2_decap_8 FILLER_20_158 ();
 sg13g2_decap_8 FILLER_20_165 ();
 sg13g2_decap_8 FILLER_20_172 ();
 sg13g2_decap_8 FILLER_20_179 ();
 sg13g2_decap_8 FILLER_20_186 ();
 sg13g2_decap_8 FILLER_20_193 ();
 sg13g2_decap_8 FILLER_20_200 ();
 sg13g2_decap_8 FILLER_20_207 ();
 sg13g2_decap_8 FILLER_20_214 ();
 sg13g2_decap_8 FILLER_20_221 ();
 sg13g2_decap_8 FILLER_20_228 ();
 sg13g2_decap_8 FILLER_20_235 ();
 sg13g2_decap_8 FILLER_20_242 ();
 sg13g2_decap_8 FILLER_20_249 ();
 sg13g2_decap_8 FILLER_20_256 ();
 sg13g2_decap_8 FILLER_20_263 ();
 sg13g2_decap_8 FILLER_20_270 ();
 sg13g2_decap_8 FILLER_20_277 ();
 sg13g2_decap_8 FILLER_20_284 ();
 sg13g2_decap_8 FILLER_20_291 ();
 sg13g2_decap_8 FILLER_20_298 ();
 sg13g2_decap_8 FILLER_20_305 ();
 sg13g2_decap_8 FILLER_20_312 ();
 sg13g2_decap_8 FILLER_20_319 ();
 sg13g2_decap_8 FILLER_20_326 ();
 sg13g2_decap_8 FILLER_20_333 ();
 sg13g2_decap_8 FILLER_20_340 ();
 sg13g2_decap_8 FILLER_20_347 ();
 sg13g2_decap_8 FILLER_20_354 ();
 sg13g2_decap_8 FILLER_20_361 ();
 sg13g2_decap_8 FILLER_20_368 ();
 sg13g2_decap_8 FILLER_20_375 ();
 sg13g2_decap_8 FILLER_20_382 ();
 sg13g2_decap_8 FILLER_20_389 ();
 sg13g2_decap_8 FILLER_20_396 ();
 sg13g2_decap_8 FILLER_20_403 ();
 sg13g2_decap_8 FILLER_20_410 ();
 sg13g2_decap_8 FILLER_20_417 ();
 sg13g2_decap_8 FILLER_20_424 ();
 sg13g2_decap_8 FILLER_20_431 ();
 sg13g2_decap_8 FILLER_20_438 ();
 sg13g2_decap_8 FILLER_20_445 ();
 sg13g2_decap_8 FILLER_20_452 ();
 sg13g2_decap_8 FILLER_20_459 ();
 sg13g2_decap_8 FILLER_20_466 ();
 sg13g2_decap_8 FILLER_20_473 ();
 sg13g2_decap_8 FILLER_20_480 ();
 sg13g2_decap_8 FILLER_20_487 ();
 sg13g2_decap_8 FILLER_20_494 ();
 sg13g2_decap_8 FILLER_20_501 ();
 sg13g2_decap_8 FILLER_20_508 ();
 sg13g2_decap_8 FILLER_20_515 ();
 sg13g2_decap_8 FILLER_20_522 ();
 sg13g2_decap_8 FILLER_20_529 ();
 sg13g2_decap_8 FILLER_20_536 ();
 sg13g2_decap_8 FILLER_20_543 ();
 sg13g2_decap_8 FILLER_20_550 ();
 sg13g2_decap_8 FILLER_20_557 ();
 sg13g2_decap_8 FILLER_20_564 ();
 sg13g2_decap_8 FILLER_20_571 ();
 sg13g2_decap_8 FILLER_20_578 ();
 sg13g2_decap_8 FILLER_20_585 ();
 sg13g2_decap_8 FILLER_20_592 ();
 sg13g2_decap_8 FILLER_20_599 ();
 sg13g2_decap_8 FILLER_20_606 ();
 sg13g2_decap_8 FILLER_20_613 ();
 sg13g2_decap_8 FILLER_20_620 ();
 sg13g2_decap_8 FILLER_20_627 ();
 sg13g2_decap_8 FILLER_20_634 ();
 sg13g2_decap_8 FILLER_20_641 ();
 sg13g2_decap_8 FILLER_20_648 ();
 sg13g2_decap_8 FILLER_20_655 ();
 sg13g2_decap_8 FILLER_20_662 ();
 sg13g2_decap_8 FILLER_20_669 ();
 sg13g2_decap_8 FILLER_20_676 ();
 sg13g2_decap_8 FILLER_20_683 ();
 sg13g2_decap_8 FILLER_20_690 ();
 sg13g2_decap_8 FILLER_20_697 ();
 sg13g2_decap_8 FILLER_20_704 ();
 sg13g2_decap_8 FILLER_20_711 ();
 sg13g2_decap_8 FILLER_20_718 ();
 sg13g2_decap_8 FILLER_20_725 ();
 sg13g2_decap_8 FILLER_20_732 ();
 sg13g2_decap_8 FILLER_20_739 ();
 sg13g2_decap_8 FILLER_20_746 ();
 sg13g2_decap_8 FILLER_20_753 ();
 sg13g2_decap_8 FILLER_20_760 ();
 sg13g2_decap_8 FILLER_20_767 ();
 sg13g2_decap_8 FILLER_20_774 ();
 sg13g2_decap_8 FILLER_20_781 ();
 sg13g2_decap_8 FILLER_20_788 ();
 sg13g2_decap_8 FILLER_20_795 ();
 sg13g2_decap_8 FILLER_20_802 ();
 sg13g2_decap_8 FILLER_20_809 ();
 sg13g2_decap_8 FILLER_20_816 ();
 sg13g2_decap_8 FILLER_20_823 ();
 sg13g2_decap_8 FILLER_20_830 ();
 sg13g2_decap_8 FILLER_20_837 ();
 sg13g2_decap_8 FILLER_20_844 ();
 sg13g2_decap_8 FILLER_20_851 ();
 sg13g2_decap_8 FILLER_20_858 ();
 sg13g2_decap_8 FILLER_20_865 ();
 sg13g2_decap_8 FILLER_20_872 ();
 sg13g2_decap_8 FILLER_20_879 ();
 sg13g2_decap_8 FILLER_20_886 ();
 sg13g2_decap_8 FILLER_20_893 ();
 sg13g2_decap_8 FILLER_20_900 ();
 sg13g2_decap_8 FILLER_20_907 ();
 sg13g2_decap_8 FILLER_20_914 ();
 sg13g2_decap_8 FILLER_20_921 ();
 sg13g2_decap_8 FILLER_20_928 ();
 sg13g2_decap_8 FILLER_20_935 ();
 sg13g2_decap_8 FILLER_20_942 ();
 sg13g2_decap_8 FILLER_20_949 ();
 sg13g2_decap_8 FILLER_20_956 ();
 sg13g2_decap_8 FILLER_20_963 ();
 sg13g2_decap_8 FILLER_20_970 ();
 sg13g2_decap_8 FILLER_20_977 ();
 sg13g2_decap_8 FILLER_20_984 ();
 sg13g2_decap_8 FILLER_20_991 ();
 sg13g2_decap_8 FILLER_20_998 ();
 sg13g2_decap_8 FILLER_20_1005 ();
 sg13g2_decap_8 FILLER_20_1012 ();
 sg13g2_decap_8 FILLER_20_1019 ();
 sg13g2_fill_2 FILLER_20_1026 ();
 sg13g2_fill_1 FILLER_20_1028 ();
 sg13g2_decap_8 FILLER_21_4 ();
 sg13g2_decap_8 FILLER_21_11 ();
 sg13g2_decap_8 FILLER_21_18 ();
 sg13g2_decap_8 FILLER_21_25 ();
 sg13g2_decap_8 FILLER_21_32 ();
 sg13g2_decap_8 FILLER_21_39 ();
 sg13g2_decap_8 FILLER_21_46 ();
 sg13g2_decap_8 FILLER_21_53 ();
 sg13g2_decap_8 FILLER_21_60 ();
 sg13g2_decap_8 FILLER_21_67 ();
 sg13g2_decap_8 FILLER_21_74 ();
 sg13g2_decap_8 FILLER_21_81 ();
 sg13g2_decap_8 FILLER_21_88 ();
 sg13g2_decap_8 FILLER_21_95 ();
 sg13g2_decap_8 FILLER_21_102 ();
 sg13g2_decap_8 FILLER_21_109 ();
 sg13g2_decap_8 FILLER_21_116 ();
 sg13g2_decap_8 FILLER_21_123 ();
 sg13g2_decap_8 FILLER_21_130 ();
 sg13g2_decap_8 FILLER_21_137 ();
 sg13g2_decap_8 FILLER_21_144 ();
 sg13g2_decap_8 FILLER_21_151 ();
 sg13g2_decap_8 FILLER_21_158 ();
 sg13g2_decap_8 FILLER_21_165 ();
 sg13g2_decap_8 FILLER_21_172 ();
 sg13g2_decap_8 FILLER_21_179 ();
 sg13g2_decap_8 FILLER_21_186 ();
 sg13g2_decap_8 FILLER_21_193 ();
 sg13g2_decap_8 FILLER_21_200 ();
 sg13g2_decap_8 FILLER_21_207 ();
 sg13g2_decap_8 FILLER_21_214 ();
 sg13g2_decap_8 FILLER_21_221 ();
 sg13g2_decap_8 FILLER_21_228 ();
 sg13g2_decap_8 FILLER_21_235 ();
 sg13g2_decap_8 FILLER_21_242 ();
 sg13g2_decap_8 FILLER_21_249 ();
 sg13g2_decap_8 FILLER_21_256 ();
 sg13g2_decap_8 FILLER_21_263 ();
 sg13g2_decap_8 FILLER_21_270 ();
 sg13g2_decap_8 FILLER_21_277 ();
 sg13g2_decap_8 FILLER_21_284 ();
 sg13g2_decap_8 FILLER_21_291 ();
 sg13g2_decap_8 FILLER_21_298 ();
 sg13g2_decap_8 FILLER_21_305 ();
 sg13g2_decap_8 FILLER_21_312 ();
 sg13g2_decap_8 FILLER_21_319 ();
 sg13g2_decap_8 FILLER_21_326 ();
 sg13g2_decap_8 FILLER_21_333 ();
 sg13g2_decap_8 FILLER_21_340 ();
 sg13g2_decap_8 FILLER_21_347 ();
 sg13g2_decap_8 FILLER_21_354 ();
 sg13g2_decap_8 FILLER_21_361 ();
 sg13g2_decap_8 FILLER_21_368 ();
 sg13g2_decap_8 FILLER_21_375 ();
 sg13g2_decap_8 FILLER_21_382 ();
 sg13g2_decap_8 FILLER_21_389 ();
 sg13g2_decap_8 FILLER_21_396 ();
 sg13g2_decap_8 FILLER_21_403 ();
 sg13g2_decap_8 FILLER_21_410 ();
 sg13g2_decap_8 FILLER_21_417 ();
 sg13g2_decap_8 FILLER_21_424 ();
 sg13g2_decap_8 FILLER_21_431 ();
 sg13g2_decap_8 FILLER_21_438 ();
 sg13g2_decap_8 FILLER_21_445 ();
 sg13g2_decap_8 FILLER_21_452 ();
 sg13g2_decap_8 FILLER_21_459 ();
 sg13g2_decap_8 FILLER_21_466 ();
 sg13g2_decap_8 FILLER_21_473 ();
 sg13g2_decap_8 FILLER_21_480 ();
 sg13g2_decap_8 FILLER_21_487 ();
 sg13g2_decap_8 FILLER_21_494 ();
 sg13g2_decap_8 FILLER_21_501 ();
 sg13g2_decap_8 FILLER_21_508 ();
 sg13g2_decap_8 FILLER_21_515 ();
 sg13g2_decap_8 FILLER_21_522 ();
 sg13g2_decap_8 FILLER_21_529 ();
 sg13g2_decap_8 FILLER_21_536 ();
 sg13g2_decap_8 FILLER_21_543 ();
 sg13g2_decap_8 FILLER_21_550 ();
 sg13g2_decap_8 FILLER_21_557 ();
 sg13g2_decap_8 FILLER_21_564 ();
 sg13g2_decap_8 FILLER_21_571 ();
 sg13g2_decap_8 FILLER_21_578 ();
 sg13g2_decap_8 FILLER_21_585 ();
 sg13g2_decap_8 FILLER_21_592 ();
 sg13g2_decap_8 FILLER_21_599 ();
 sg13g2_decap_8 FILLER_21_606 ();
 sg13g2_decap_8 FILLER_21_613 ();
 sg13g2_decap_8 FILLER_21_620 ();
 sg13g2_decap_8 FILLER_21_627 ();
 sg13g2_decap_8 FILLER_21_634 ();
 sg13g2_decap_8 FILLER_21_641 ();
 sg13g2_decap_8 FILLER_21_648 ();
 sg13g2_decap_8 FILLER_21_655 ();
 sg13g2_decap_8 FILLER_21_662 ();
 sg13g2_decap_8 FILLER_21_669 ();
 sg13g2_decap_8 FILLER_21_676 ();
 sg13g2_decap_8 FILLER_21_683 ();
 sg13g2_decap_8 FILLER_21_690 ();
 sg13g2_decap_8 FILLER_21_697 ();
 sg13g2_decap_8 FILLER_21_704 ();
 sg13g2_decap_8 FILLER_21_711 ();
 sg13g2_decap_8 FILLER_21_718 ();
 sg13g2_decap_8 FILLER_21_725 ();
 sg13g2_decap_8 FILLER_21_732 ();
 sg13g2_decap_8 FILLER_21_739 ();
 sg13g2_decap_8 FILLER_21_746 ();
 sg13g2_decap_8 FILLER_21_753 ();
 sg13g2_decap_8 FILLER_21_760 ();
 sg13g2_decap_8 FILLER_21_767 ();
 sg13g2_decap_8 FILLER_21_774 ();
 sg13g2_decap_8 FILLER_21_781 ();
 sg13g2_decap_8 FILLER_21_788 ();
 sg13g2_decap_8 FILLER_21_795 ();
 sg13g2_decap_8 FILLER_21_802 ();
 sg13g2_decap_8 FILLER_21_809 ();
 sg13g2_decap_8 FILLER_21_816 ();
 sg13g2_decap_8 FILLER_21_823 ();
 sg13g2_decap_8 FILLER_21_830 ();
 sg13g2_decap_8 FILLER_21_837 ();
 sg13g2_decap_8 FILLER_21_844 ();
 sg13g2_decap_8 FILLER_21_851 ();
 sg13g2_decap_8 FILLER_21_858 ();
 sg13g2_decap_8 FILLER_21_865 ();
 sg13g2_decap_8 FILLER_21_872 ();
 sg13g2_decap_8 FILLER_21_879 ();
 sg13g2_decap_8 FILLER_21_886 ();
 sg13g2_decap_8 FILLER_21_893 ();
 sg13g2_decap_8 FILLER_21_900 ();
 sg13g2_decap_8 FILLER_21_907 ();
 sg13g2_decap_8 FILLER_21_914 ();
 sg13g2_decap_8 FILLER_21_921 ();
 sg13g2_decap_8 FILLER_21_928 ();
 sg13g2_decap_8 FILLER_21_935 ();
 sg13g2_decap_8 FILLER_21_942 ();
 sg13g2_decap_8 FILLER_21_949 ();
 sg13g2_decap_8 FILLER_21_956 ();
 sg13g2_decap_8 FILLER_21_963 ();
 sg13g2_decap_8 FILLER_21_970 ();
 sg13g2_decap_8 FILLER_21_977 ();
 sg13g2_decap_8 FILLER_21_984 ();
 sg13g2_decap_8 FILLER_21_991 ();
 sg13g2_decap_8 FILLER_21_998 ();
 sg13g2_decap_8 FILLER_21_1005 ();
 sg13g2_decap_8 FILLER_21_1012 ();
 sg13g2_decap_8 FILLER_21_1019 ();
 sg13g2_fill_2 FILLER_21_1026 ();
 sg13g2_fill_1 FILLER_21_1028 ();
 sg13g2_decap_8 FILLER_22_4 ();
 sg13g2_decap_8 FILLER_22_11 ();
 sg13g2_decap_8 FILLER_22_18 ();
 sg13g2_decap_8 FILLER_22_25 ();
 sg13g2_decap_8 FILLER_22_32 ();
 sg13g2_decap_8 FILLER_22_39 ();
 sg13g2_decap_8 FILLER_22_46 ();
 sg13g2_decap_8 FILLER_22_53 ();
 sg13g2_decap_8 FILLER_22_60 ();
 sg13g2_decap_8 FILLER_22_67 ();
 sg13g2_decap_8 FILLER_22_74 ();
 sg13g2_decap_8 FILLER_22_81 ();
 sg13g2_decap_8 FILLER_22_88 ();
 sg13g2_decap_8 FILLER_22_95 ();
 sg13g2_decap_8 FILLER_22_102 ();
 sg13g2_decap_8 FILLER_22_109 ();
 sg13g2_decap_8 FILLER_22_116 ();
 sg13g2_decap_8 FILLER_22_123 ();
 sg13g2_decap_8 FILLER_22_130 ();
 sg13g2_decap_8 FILLER_22_137 ();
 sg13g2_decap_8 FILLER_22_144 ();
 sg13g2_decap_8 FILLER_22_151 ();
 sg13g2_decap_8 FILLER_22_158 ();
 sg13g2_decap_8 FILLER_22_165 ();
 sg13g2_decap_8 FILLER_22_172 ();
 sg13g2_decap_8 FILLER_22_179 ();
 sg13g2_decap_8 FILLER_22_186 ();
 sg13g2_decap_8 FILLER_22_193 ();
 sg13g2_decap_8 FILLER_22_200 ();
 sg13g2_decap_8 FILLER_22_207 ();
 sg13g2_decap_8 FILLER_22_214 ();
 sg13g2_decap_8 FILLER_22_221 ();
 sg13g2_decap_8 FILLER_22_228 ();
 sg13g2_decap_8 FILLER_22_235 ();
 sg13g2_decap_8 FILLER_22_242 ();
 sg13g2_decap_8 FILLER_22_249 ();
 sg13g2_decap_8 FILLER_22_256 ();
 sg13g2_decap_8 FILLER_22_263 ();
 sg13g2_decap_8 FILLER_22_270 ();
 sg13g2_decap_8 FILLER_22_277 ();
 sg13g2_decap_8 FILLER_22_284 ();
 sg13g2_decap_8 FILLER_22_291 ();
 sg13g2_decap_8 FILLER_22_298 ();
 sg13g2_decap_8 FILLER_22_305 ();
 sg13g2_decap_8 FILLER_22_312 ();
 sg13g2_decap_8 FILLER_22_319 ();
 sg13g2_decap_8 FILLER_22_326 ();
 sg13g2_decap_8 FILLER_22_333 ();
 sg13g2_decap_8 FILLER_22_340 ();
 sg13g2_decap_8 FILLER_22_347 ();
 sg13g2_decap_8 FILLER_22_354 ();
 sg13g2_decap_8 FILLER_22_361 ();
 sg13g2_decap_8 FILLER_22_368 ();
 sg13g2_decap_8 FILLER_22_375 ();
 sg13g2_decap_8 FILLER_22_382 ();
 sg13g2_decap_8 FILLER_22_389 ();
 sg13g2_decap_8 FILLER_22_396 ();
 sg13g2_decap_8 FILLER_22_403 ();
 sg13g2_decap_8 FILLER_22_410 ();
 sg13g2_decap_8 FILLER_22_417 ();
 sg13g2_decap_8 FILLER_22_424 ();
 sg13g2_decap_8 FILLER_22_431 ();
 sg13g2_decap_8 FILLER_22_438 ();
 sg13g2_decap_8 FILLER_22_445 ();
 sg13g2_decap_8 FILLER_22_452 ();
 sg13g2_decap_8 FILLER_22_459 ();
 sg13g2_decap_8 FILLER_22_466 ();
 sg13g2_decap_8 FILLER_22_473 ();
 sg13g2_decap_8 FILLER_22_480 ();
 sg13g2_decap_8 FILLER_22_487 ();
 sg13g2_decap_8 FILLER_22_494 ();
 sg13g2_decap_8 FILLER_22_501 ();
 sg13g2_decap_8 FILLER_22_508 ();
 sg13g2_decap_8 FILLER_22_515 ();
 sg13g2_decap_8 FILLER_22_522 ();
 sg13g2_decap_8 FILLER_22_529 ();
 sg13g2_decap_8 FILLER_22_536 ();
 sg13g2_decap_8 FILLER_22_543 ();
 sg13g2_decap_8 FILLER_22_550 ();
 sg13g2_decap_8 FILLER_22_557 ();
 sg13g2_decap_8 FILLER_22_564 ();
 sg13g2_decap_8 FILLER_22_571 ();
 sg13g2_decap_8 FILLER_22_578 ();
 sg13g2_decap_8 FILLER_22_585 ();
 sg13g2_decap_8 FILLER_22_592 ();
 sg13g2_decap_8 FILLER_22_599 ();
 sg13g2_decap_8 FILLER_22_606 ();
 sg13g2_decap_8 FILLER_22_613 ();
 sg13g2_decap_8 FILLER_22_620 ();
 sg13g2_decap_8 FILLER_22_627 ();
 sg13g2_decap_8 FILLER_22_634 ();
 sg13g2_decap_8 FILLER_22_641 ();
 sg13g2_decap_8 FILLER_22_648 ();
 sg13g2_decap_8 FILLER_22_655 ();
 sg13g2_decap_8 FILLER_22_662 ();
 sg13g2_decap_8 FILLER_22_669 ();
 sg13g2_decap_8 FILLER_22_676 ();
 sg13g2_decap_8 FILLER_22_683 ();
 sg13g2_decap_8 FILLER_22_690 ();
 sg13g2_decap_8 FILLER_22_697 ();
 sg13g2_decap_8 FILLER_22_704 ();
 sg13g2_decap_8 FILLER_22_711 ();
 sg13g2_decap_8 FILLER_22_718 ();
 sg13g2_decap_8 FILLER_22_725 ();
 sg13g2_decap_8 FILLER_22_732 ();
 sg13g2_decap_8 FILLER_22_739 ();
 sg13g2_decap_8 FILLER_22_746 ();
 sg13g2_decap_8 FILLER_22_753 ();
 sg13g2_decap_8 FILLER_22_760 ();
 sg13g2_decap_8 FILLER_22_767 ();
 sg13g2_decap_8 FILLER_22_774 ();
 sg13g2_decap_8 FILLER_22_781 ();
 sg13g2_decap_8 FILLER_22_788 ();
 sg13g2_decap_8 FILLER_22_795 ();
 sg13g2_decap_8 FILLER_22_802 ();
 sg13g2_decap_8 FILLER_22_809 ();
 sg13g2_decap_8 FILLER_22_816 ();
 sg13g2_decap_8 FILLER_22_823 ();
 sg13g2_decap_8 FILLER_22_830 ();
 sg13g2_decap_8 FILLER_22_837 ();
 sg13g2_decap_8 FILLER_22_844 ();
 sg13g2_decap_8 FILLER_22_851 ();
 sg13g2_decap_8 FILLER_22_858 ();
 sg13g2_decap_8 FILLER_22_865 ();
 sg13g2_decap_8 FILLER_22_872 ();
 sg13g2_decap_8 FILLER_22_879 ();
 sg13g2_decap_8 FILLER_22_886 ();
 sg13g2_decap_8 FILLER_22_893 ();
 sg13g2_decap_8 FILLER_22_900 ();
 sg13g2_decap_8 FILLER_22_907 ();
 sg13g2_decap_8 FILLER_22_914 ();
 sg13g2_decap_8 FILLER_22_921 ();
 sg13g2_decap_8 FILLER_22_928 ();
 sg13g2_decap_8 FILLER_22_935 ();
 sg13g2_decap_8 FILLER_22_942 ();
 sg13g2_decap_8 FILLER_22_949 ();
 sg13g2_decap_8 FILLER_22_956 ();
 sg13g2_decap_8 FILLER_22_963 ();
 sg13g2_decap_8 FILLER_22_970 ();
 sg13g2_decap_8 FILLER_22_977 ();
 sg13g2_decap_8 FILLER_22_984 ();
 sg13g2_decap_8 FILLER_22_991 ();
 sg13g2_decap_8 FILLER_22_998 ();
 sg13g2_decap_8 FILLER_22_1005 ();
 sg13g2_decap_8 FILLER_22_1012 ();
 sg13g2_decap_8 FILLER_22_1019 ();
 sg13g2_fill_2 FILLER_22_1026 ();
 sg13g2_fill_1 FILLER_22_1028 ();
 sg13g2_decap_8 FILLER_23_4 ();
 sg13g2_decap_8 FILLER_23_11 ();
 sg13g2_decap_8 FILLER_23_18 ();
 sg13g2_decap_8 FILLER_23_25 ();
 sg13g2_decap_8 FILLER_23_32 ();
 sg13g2_decap_8 FILLER_23_39 ();
 sg13g2_decap_8 FILLER_23_46 ();
 sg13g2_decap_8 FILLER_23_53 ();
 sg13g2_decap_8 FILLER_23_60 ();
 sg13g2_decap_8 FILLER_23_67 ();
 sg13g2_decap_8 FILLER_23_74 ();
 sg13g2_decap_8 FILLER_23_81 ();
 sg13g2_decap_8 FILLER_23_88 ();
 sg13g2_decap_8 FILLER_23_95 ();
 sg13g2_decap_8 FILLER_23_102 ();
 sg13g2_decap_8 FILLER_23_109 ();
 sg13g2_decap_8 FILLER_23_116 ();
 sg13g2_decap_8 FILLER_23_123 ();
 sg13g2_decap_8 FILLER_23_130 ();
 sg13g2_decap_8 FILLER_23_137 ();
 sg13g2_decap_8 FILLER_23_144 ();
 sg13g2_decap_8 FILLER_23_151 ();
 sg13g2_decap_8 FILLER_23_158 ();
 sg13g2_decap_8 FILLER_23_165 ();
 sg13g2_decap_8 FILLER_23_172 ();
 sg13g2_decap_8 FILLER_23_179 ();
 sg13g2_decap_8 FILLER_23_186 ();
 sg13g2_decap_8 FILLER_23_193 ();
 sg13g2_decap_8 FILLER_23_200 ();
 sg13g2_decap_8 FILLER_23_207 ();
 sg13g2_decap_8 FILLER_23_214 ();
 sg13g2_decap_8 FILLER_23_221 ();
 sg13g2_decap_8 FILLER_23_228 ();
 sg13g2_decap_8 FILLER_23_235 ();
 sg13g2_decap_8 FILLER_23_242 ();
 sg13g2_decap_8 FILLER_23_249 ();
 sg13g2_decap_8 FILLER_23_256 ();
 sg13g2_decap_8 FILLER_23_263 ();
 sg13g2_decap_8 FILLER_23_270 ();
 sg13g2_decap_8 FILLER_23_277 ();
 sg13g2_decap_8 FILLER_23_284 ();
 sg13g2_decap_8 FILLER_23_291 ();
 sg13g2_decap_8 FILLER_23_298 ();
 sg13g2_decap_8 FILLER_23_305 ();
 sg13g2_decap_8 FILLER_23_312 ();
 sg13g2_decap_8 FILLER_23_319 ();
 sg13g2_decap_8 FILLER_23_326 ();
 sg13g2_decap_8 FILLER_23_333 ();
 sg13g2_decap_8 FILLER_23_340 ();
 sg13g2_decap_8 FILLER_23_347 ();
 sg13g2_decap_8 FILLER_23_354 ();
 sg13g2_decap_8 FILLER_23_361 ();
 sg13g2_decap_8 FILLER_23_368 ();
 sg13g2_decap_8 FILLER_23_375 ();
 sg13g2_decap_8 FILLER_23_382 ();
 sg13g2_decap_8 FILLER_23_389 ();
 sg13g2_decap_8 FILLER_23_396 ();
 sg13g2_decap_8 FILLER_23_403 ();
 sg13g2_decap_8 FILLER_23_410 ();
 sg13g2_decap_8 FILLER_23_417 ();
 sg13g2_decap_8 FILLER_23_424 ();
 sg13g2_decap_8 FILLER_23_431 ();
 sg13g2_decap_8 FILLER_23_438 ();
 sg13g2_decap_8 FILLER_23_445 ();
 sg13g2_decap_8 FILLER_23_452 ();
 sg13g2_decap_8 FILLER_23_459 ();
 sg13g2_decap_8 FILLER_23_466 ();
 sg13g2_decap_8 FILLER_23_473 ();
 sg13g2_decap_8 FILLER_23_480 ();
 sg13g2_decap_8 FILLER_23_487 ();
 sg13g2_decap_8 FILLER_23_494 ();
 sg13g2_decap_8 FILLER_23_501 ();
 sg13g2_decap_8 FILLER_23_508 ();
 sg13g2_decap_8 FILLER_23_515 ();
 sg13g2_decap_8 FILLER_23_522 ();
 sg13g2_decap_8 FILLER_23_529 ();
 sg13g2_decap_8 FILLER_23_536 ();
 sg13g2_decap_8 FILLER_23_543 ();
 sg13g2_decap_8 FILLER_23_550 ();
 sg13g2_decap_8 FILLER_23_557 ();
 sg13g2_decap_8 FILLER_23_564 ();
 sg13g2_decap_8 FILLER_23_571 ();
 sg13g2_decap_8 FILLER_23_578 ();
 sg13g2_decap_8 FILLER_23_585 ();
 sg13g2_decap_8 FILLER_23_592 ();
 sg13g2_decap_8 FILLER_23_599 ();
 sg13g2_decap_8 FILLER_23_606 ();
 sg13g2_decap_8 FILLER_23_613 ();
 sg13g2_decap_8 FILLER_23_620 ();
 sg13g2_decap_8 FILLER_23_627 ();
 sg13g2_decap_8 FILLER_23_634 ();
 sg13g2_decap_8 FILLER_23_641 ();
 sg13g2_decap_8 FILLER_23_648 ();
 sg13g2_decap_8 FILLER_23_655 ();
 sg13g2_decap_8 FILLER_23_662 ();
 sg13g2_decap_8 FILLER_23_669 ();
 sg13g2_decap_8 FILLER_23_676 ();
 sg13g2_decap_8 FILLER_23_683 ();
 sg13g2_decap_8 FILLER_23_690 ();
 sg13g2_decap_8 FILLER_23_697 ();
 sg13g2_decap_8 FILLER_23_704 ();
 sg13g2_decap_8 FILLER_23_711 ();
 sg13g2_decap_8 FILLER_23_718 ();
 sg13g2_decap_8 FILLER_23_725 ();
 sg13g2_decap_8 FILLER_23_732 ();
 sg13g2_decap_8 FILLER_23_739 ();
 sg13g2_decap_8 FILLER_23_746 ();
 sg13g2_decap_8 FILLER_23_753 ();
 sg13g2_decap_8 FILLER_23_760 ();
 sg13g2_decap_8 FILLER_23_767 ();
 sg13g2_decap_8 FILLER_23_774 ();
 sg13g2_decap_8 FILLER_23_781 ();
 sg13g2_decap_8 FILLER_23_788 ();
 sg13g2_decap_8 FILLER_23_795 ();
 sg13g2_decap_8 FILLER_23_802 ();
 sg13g2_decap_8 FILLER_23_809 ();
 sg13g2_decap_8 FILLER_23_816 ();
 sg13g2_decap_8 FILLER_23_823 ();
 sg13g2_decap_8 FILLER_23_830 ();
 sg13g2_decap_8 FILLER_23_837 ();
 sg13g2_decap_8 FILLER_23_844 ();
 sg13g2_decap_8 FILLER_23_851 ();
 sg13g2_decap_8 FILLER_23_858 ();
 sg13g2_decap_8 FILLER_23_865 ();
 sg13g2_decap_8 FILLER_23_872 ();
 sg13g2_decap_8 FILLER_23_879 ();
 sg13g2_decap_8 FILLER_23_886 ();
 sg13g2_decap_8 FILLER_23_893 ();
 sg13g2_decap_8 FILLER_23_900 ();
 sg13g2_decap_8 FILLER_23_907 ();
 sg13g2_decap_8 FILLER_23_914 ();
 sg13g2_decap_8 FILLER_23_921 ();
 sg13g2_decap_8 FILLER_23_928 ();
 sg13g2_decap_8 FILLER_23_935 ();
 sg13g2_decap_8 FILLER_23_942 ();
 sg13g2_decap_8 FILLER_23_949 ();
 sg13g2_decap_8 FILLER_23_956 ();
 sg13g2_decap_8 FILLER_23_963 ();
 sg13g2_decap_8 FILLER_23_970 ();
 sg13g2_decap_8 FILLER_23_977 ();
 sg13g2_decap_8 FILLER_23_984 ();
 sg13g2_decap_8 FILLER_23_991 ();
 sg13g2_decap_8 FILLER_23_998 ();
 sg13g2_decap_8 FILLER_23_1005 ();
 sg13g2_decap_8 FILLER_23_1012 ();
 sg13g2_decap_8 FILLER_23_1019 ();
 sg13g2_fill_2 FILLER_23_1026 ();
 sg13g2_fill_1 FILLER_23_1028 ();
 sg13g2_decap_8 FILLER_24_4 ();
 sg13g2_decap_8 FILLER_24_11 ();
 sg13g2_decap_8 FILLER_24_18 ();
 sg13g2_decap_8 FILLER_24_25 ();
 sg13g2_decap_8 FILLER_24_32 ();
 sg13g2_decap_8 FILLER_24_39 ();
 sg13g2_decap_8 FILLER_24_46 ();
 sg13g2_decap_8 FILLER_24_53 ();
 sg13g2_decap_8 FILLER_24_60 ();
 sg13g2_decap_8 FILLER_24_67 ();
 sg13g2_decap_8 FILLER_24_74 ();
 sg13g2_decap_8 FILLER_24_81 ();
 sg13g2_decap_8 FILLER_24_88 ();
 sg13g2_decap_8 FILLER_24_95 ();
 sg13g2_decap_8 FILLER_24_102 ();
 sg13g2_decap_8 FILLER_24_109 ();
 sg13g2_decap_8 FILLER_24_116 ();
 sg13g2_decap_8 FILLER_24_123 ();
 sg13g2_decap_8 FILLER_24_130 ();
 sg13g2_decap_8 FILLER_24_137 ();
 sg13g2_decap_8 FILLER_24_144 ();
 sg13g2_decap_8 FILLER_24_151 ();
 sg13g2_decap_8 FILLER_24_158 ();
 sg13g2_decap_8 FILLER_24_165 ();
 sg13g2_decap_8 FILLER_24_172 ();
 sg13g2_decap_8 FILLER_24_179 ();
 sg13g2_decap_8 FILLER_24_186 ();
 sg13g2_decap_8 FILLER_24_193 ();
 sg13g2_decap_8 FILLER_24_200 ();
 sg13g2_decap_8 FILLER_24_207 ();
 sg13g2_decap_8 FILLER_24_214 ();
 sg13g2_decap_8 FILLER_24_221 ();
 sg13g2_decap_8 FILLER_24_228 ();
 sg13g2_decap_8 FILLER_24_235 ();
 sg13g2_decap_8 FILLER_24_242 ();
 sg13g2_decap_8 FILLER_24_249 ();
 sg13g2_decap_8 FILLER_24_256 ();
 sg13g2_decap_8 FILLER_24_263 ();
 sg13g2_decap_8 FILLER_24_270 ();
 sg13g2_decap_8 FILLER_24_277 ();
 sg13g2_decap_8 FILLER_24_284 ();
 sg13g2_decap_8 FILLER_24_291 ();
 sg13g2_decap_8 FILLER_24_298 ();
 sg13g2_decap_8 FILLER_24_305 ();
 sg13g2_decap_8 FILLER_24_312 ();
 sg13g2_decap_8 FILLER_24_319 ();
 sg13g2_decap_8 FILLER_24_326 ();
 sg13g2_decap_8 FILLER_24_333 ();
 sg13g2_decap_8 FILLER_24_340 ();
 sg13g2_decap_8 FILLER_24_347 ();
 sg13g2_decap_8 FILLER_24_354 ();
 sg13g2_decap_8 FILLER_24_361 ();
 sg13g2_decap_8 FILLER_24_368 ();
 sg13g2_decap_8 FILLER_24_375 ();
 sg13g2_decap_8 FILLER_24_382 ();
 sg13g2_decap_8 FILLER_24_389 ();
 sg13g2_decap_8 FILLER_24_396 ();
 sg13g2_decap_8 FILLER_24_403 ();
 sg13g2_decap_8 FILLER_24_410 ();
 sg13g2_decap_8 FILLER_24_417 ();
 sg13g2_decap_8 FILLER_24_424 ();
 sg13g2_decap_8 FILLER_24_431 ();
 sg13g2_decap_8 FILLER_24_438 ();
 sg13g2_decap_8 FILLER_24_445 ();
 sg13g2_decap_8 FILLER_24_452 ();
 sg13g2_decap_8 FILLER_24_459 ();
 sg13g2_decap_8 FILLER_24_466 ();
 sg13g2_decap_8 FILLER_24_473 ();
 sg13g2_decap_8 FILLER_24_480 ();
 sg13g2_decap_8 FILLER_24_487 ();
 sg13g2_decap_8 FILLER_24_494 ();
 sg13g2_decap_8 FILLER_24_501 ();
 sg13g2_decap_8 FILLER_24_508 ();
 sg13g2_decap_8 FILLER_24_515 ();
 sg13g2_decap_8 FILLER_24_522 ();
 sg13g2_decap_8 FILLER_24_529 ();
 sg13g2_decap_8 FILLER_24_536 ();
 sg13g2_decap_8 FILLER_24_543 ();
 sg13g2_decap_8 FILLER_24_550 ();
 sg13g2_decap_8 FILLER_24_557 ();
 sg13g2_decap_8 FILLER_24_564 ();
 sg13g2_decap_8 FILLER_24_571 ();
 sg13g2_decap_8 FILLER_24_578 ();
 sg13g2_decap_8 FILLER_24_585 ();
 sg13g2_decap_8 FILLER_24_592 ();
 sg13g2_decap_8 FILLER_24_599 ();
 sg13g2_decap_8 FILLER_24_606 ();
 sg13g2_decap_8 FILLER_24_613 ();
 sg13g2_decap_8 FILLER_24_620 ();
 sg13g2_decap_8 FILLER_24_627 ();
 sg13g2_decap_8 FILLER_24_634 ();
 sg13g2_decap_8 FILLER_24_641 ();
 sg13g2_decap_8 FILLER_24_648 ();
 sg13g2_decap_8 FILLER_24_655 ();
 sg13g2_decap_8 FILLER_24_662 ();
 sg13g2_decap_8 FILLER_24_669 ();
 sg13g2_decap_8 FILLER_24_676 ();
 sg13g2_decap_8 FILLER_24_683 ();
 sg13g2_decap_8 FILLER_24_690 ();
 sg13g2_decap_8 FILLER_24_697 ();
 sg13g2_decap_8 FILLER_24_704 ();
 sg13g2_decap_8 FILLER_24_711 ();
 sg13g2_decap_8 FILLER_24_718 ();
 sg13g2_decap_8 FILLER_24_725 ();
 sg13g2_decap_8 FILLER_24_732 ();
 sg13g2_decap_8 FILLER_24_739 ();
 sg13g2_decap_8 FILLER_24_746 ();
 sg13g2_decap_8 FILLER_24_753 ();
 sg13g2_decap_8 FILLER_24_760 ();
 sg13g2_decap_8 FILLER_24_767 ();
 sg13g2_decap_8 FILLER_24_774 ();
 sg13g2_decap_8 FILLER_24_781 ();
 sg13g2_decap_8 FILLER_24_788 ();
 sg13g2_decap_8 FILLER_24_795 ();
 sg13g2_decap_8 FILLER_24_802 ();
 sg13g2_decap_8 FILLER_24_809 ();
 sg13g2_decap_8 FILLER_24_816 ();
 sg13g2_decap_8 FILLER_24_823 ();
 sg13g2_decap_8 FILLER_24_830 ();
 sg13g2_decap_8 FILLER_24_837 ();
 sg13g2_decap_8 FILLER_24_844 ();
 sg13g2_decap_8 FILLER_24_851 ();
 sg13g2_decap_8 FILLER_24_858 ();
 sg13g2_decap_8 FILLER_24_865 ();
 sg13g2_decap_8 FILLER_24_872 ();
 sg13g2_decap_8 FILLER_24_879 ();
 sg13g2_decap_8 FILLER_24_886 ();
 sg13g2_decap_8 FILLER_24_893 ();
 sg13g2_decap_8 FILLER_24_900 ();
 sg13g2_decap_8 FILLER_24_907 ();
 sg13g2_decap_8 FILLER_24_914 ();
 sg13g2_decap_8 FILLER_24_921 ();
 sg13g2_decap_8 FILLER_24_928 ();
 sg13g2_decap_8 FILLER_24_935 ();
 sg13g2_decap_8 FILLER_24_942 ();
 sg13g2_decap_8 FILLER_24_949 ();
 sg13g2_decap_8 FILLER_24_956 ();
 sg13g2_decap_8 FILLER_24_963 ();
 sg13g2_decap_8 FILLER_24_970 ();
 sg13g2_decap_8 FILLER_24_977 ();
 sg13g2_decap_8 FILLER_24_984 ();
 sg13g2_decap_8 FILLER_24_991 ();
 sg13g2_decap_8 FILLER_24_998 ();
 sg13g2_decap_8 FILLER_24_1005 ();
 sg13g2_decap_8 FILLER_24_1012 ();
 sg13g2_decap_8 FILLER_24_1019 ();
 sg13g2_fill_2 FILLER_24_1026 ();
 sg13g2_fill_1 FILLER_24_1028 ();
 sg13g2_decap_8 FILLER_25_4 ();
 sg13g2_decap_8 FILLER_25_11 ();
 sg13g2_decap_8 FILLER_25_18 ();
 sg13g2_decap_8 FILLER_25_25 ();
 sg13g2_decap_8 FILLER_25_32 ();
 sg13g2_decap_8 FILLER_25_39 ();
 sg13g2_decap_8 FILLER_25_46 ();
 sg13g2_decap_8 FILLER_25_53 ();
 sg13g2_decap_8 FILLER_25_60 ();
 sg13g2_decap_8 FILLER_25_67 ();
 sg13g2_decap_8 FILLER_25_74 ();
 sg13g2_decap_8 FILLER_25_81 ();
 sg13g2_decap_8 FILLER_25_88 ();
 sg13g2_decap_8 FILLER_25_95 ();
 sg13g2_decap_8 FILLER_25_102 ();
 sg13g2_decap_8 FILLER_25_109 ();
 sg13g2_decap_8 FILLER_25_116 ();
 sg13g2_decap_8 FILLER_25_123 ();
 sg13g2_decap_8 FILLER_25_130 ();
 sg13g2_decap_8 FILLER_25_137 ();
 sg13g2_decap_8 FILLER_25_144 ();
 sg13g2_decap_8 FILLER_25_151 ();
 sg13g2_decap_8 FILLER_25_158 ();
 sg13g2_decap_8 FILLER_25_165 ();
 sg13g2_decap_8 FILLER_25_172 ();
 sg13g2_decap_8 FILLER_25_179 ();
 sg13g2_decap_8 FILLER_25_186 ();
 sg13g2_decap_8 FILLER_25_193 ();
 sg13g2_decap_8 FILLER_25_200 ();
 sg13g2_decap_8 FILLER_25_207 ();
 sg13g2_decap_8 FILLER_25_214 ();
 sg13g2_decap_8 FILLER_25_221 ();
 sg13g2_decap_8 FILLER_25_228 ();
 sg13g2_decap_8 FILLER_25_235 ();
 sg13g2_decap_8 FILLER_25_242 ();
 sg13g2_decap_8 FILLER_25_249 ();
 sg13g2_decap_8 FILLER_25_256 ();
 sg13g2_decap_8 FILLER_25_263 ();
 sg13g2_decap_8 FILLER_25_270 ();
 sg13g2_decap_8 FILLER_25_277 ();
 sg13g2_decap_8 FILLER_25_284 ();
 sg13g2_decap_8 FILLER_25_291 ();
 sg13g2_decap_8 FILLER_25_298 ();
 sg13g2_decap_8 FILLER_25_305 ();
 sg13g2_decap_8 FILLER_25_312 ();
 sg13g2_decap_8 FILLER_25_319 ();
 sg13g2_decap_8 FILLER_25_326 ();
 sg13g2_decap_8 FILLER_25_333 ();
 sg13g2_decap_8 FILLER_25_340 ();
 sg13g2_decap_8 FILLER_25_347 ();
 sg13g2_decap_8 FILLER_25_354 ();
 sg13g2_decap_8 FILLER_25_361 ();
 sg13g2_decap_8 FILLER_25_368 ();
 sg13g2_decap_8 FILLER_25_375 ();
 sg13g2_decap_8 FILLER_25_382 ();
 sg13g2_decap_8 FILLER_25_389 ();
 sg13g2_decap_8 FILLER_25_396 ();
 sg13g2_decap_8 FILLER_25_403 ();
 sg13g2_decap_8 FILLER_25_410 ();
 sg13g2_decap_8 FILLER_25_417 ();
 sg13g2_decap_8 FILLER_25_424 ();
 sg13g2_decap_8 FILLER_25_431 ();
 sg13g2_decap_8 FILLER_25_438 ();
 sg13g2_decap_8 FILLER_25_445 ();
 sg13g2_decap_8 FILLER_25_452 ();
 sg13g2_decap_8 FILLER_25_459 ();
 sg13g2_decap_8 FILLER_25_466 ();
 sg13g2_decap_8 FILLER_25_473 ();
 sg13g2_decap_8 FILLER_25_480 ();
 sg13g2_decap_8 FILLER_25_487 ();
 sg13g2_decap_8 FILLER_25_494 ();
 sg13g2_decap_8 FILLER_25_501 ();
 sg13g2_decap_8 FILLER_25_508 ();
 sg13g2_decap_8 FILLER_25_515 ();
 sg13g2_decap_8 FILLER_25_522 ();
 sg13g2_decap_8 FILLER_25_529 ();
 sg13g2_decap_8 FILLER_25_536 ();
 sg13g2_decap_8 FILLER_25_543 ();
 sg13g2_decap_8 FILLER_25_550 ();
 sg13g2_decap_8 FILLER_25_557 ();
 sg13g2_decap_8 FILLER_25_564 ();
 sg13g2_decap_8 FILLER_25_571 ();
 sg13g2_decap_8 FILLER_25_578 ();
 sg13g2_decap_8 FILLER_25_585 ();
 sg13g2_decap_8 FILLER_25_592 ();
 sg13g2_decap_8 FILLER_25_599 ();
 sg13g2_decap_8 FILLER_25_606 ();
 sg13g2_decap_8 FILLER_25_613 ();
 sg13g2_decap_8 FILLER_25_620 ();
 sg13g2_decap_8 FILLER_25_627 ();
 sg13g2_decap_8 FILLER_25_634 ();
 sg13g2_decap_8 FILLER_25_641 ();
 sg13g2_decap_8 FILLER_25_648 ();
 sg13g2_decap_8 FILLER_25_655 ();
 sg13g2_decap_8 FILLER_25_662 ();
 sg13g2_decap_8 FILLER_25_669 ();
 sg13g2_decap_8 FILLER_25_676 ();
 sg13g2_decap_8 FILLER_25_683 ();
 sg13g2_decap_8 FILLER_25_690 ();
 sg13g2_decap_8 FILLER_25_697 ();
 sg13g2_decap_8 FILLER_25_704 ();
 sg13g2_decap_8 FILLER_25_711 ();
 sg13g2_decap_8 FILLER_25_718 ();
 sg13g2_decap_8 FILLER_25_725 ();
 sg13g2_decap_8 FILLER_25_732 ();
 sg13g2_decap_8 FILLER_25_739 ();
 sg13g2_decap_8 FILLER_25_746 ();
 sg13g2_decap_8 FILLER_25_753 ();
 sg13g2_decap_8 FILLER_25_760 ();
 sg13g2_decap_8 FILLER_25_767 ();
 sg13g2_decap_8 FILLER_25_774 ();
 sg13g2_decap_8 FILLER_25_781 ();
 sg13g2_decap_8 FILLER_25_788 ();
 sg13g2_decap_8 FILLER_25_795 ();
 sg13g2_decap_8 FILLER_25_802 ();
 sg13g2_decap_8 FILLER_25_809 ();
 sg13g2_decap_8 FILLER_25_816 ();
 sg13g2_decap_8 FILLER_25_823 ();
 sg13g2_decap_8 FILLER_25_830 ();
 sg13g2_decap_8 FILLER_25_837 ();
 sg13g2_decap_8 FILLER_25_844 ();
 sg13g2_decap_8 FILLER_25_851 ();
 sg13g2_decap_8 FILLER_25_858 ();
 sg13g2_decap_8 FILLER_25_865 ();
 sg13g2_decap_8 FILLER_25_872 ();
 sg13g2_decap_8 FILLER_25_879 ();
 sg13g2_decap_8 FILLER_25_886 ();
 sg13g2_decap_8 FILLER_25_893 ();
 sg13g2_decap_8 FILLER_25_900 ();
 sg13g2_decap_8 FILLER_25_907 ();
 sg13g2_decap_8 FILLER_25_914 ();
 sg13g2_decap_8 FILLER_25_921 ();
 sg13g2_decap_8 FILLER_25_928 ();
 sg13g2_decap_8 FILLER_25_935 ();
 sg13g2_decap_8 FILLER_25_942 ();
 sg13g2_decap_8 FILLER_25_949 ();
 sg13g2_decap_8 FILLER_25_956 ();
 sg13g2_decap_8 FILLER_25_963 ();
 sg13g2_decap_8 FILLER_25_970 ();
 sg13g2_decap_8 FILLER_25_977 ();
 sg13g2_decap_8 FILLER_25_984 ();
 sg13g2_decap_8 FILLER_25_991 ();
 sg13g2_decap_8 FILLER_25_998 ();
 sg13g2_decap_8 FILLER_25_1005 ();
 sg13g2_decap_8 FILLER_25_1012 ();
 sg13g2_decap_8 FILLER_25_1019 ();
 sg13g2_fill_2 FILLER_25_1026 ();
 sg13g2_fill_1 FILLER_25_1028 ();
 sg13g2_decap_8 FILLER_26_4 ();
 sg13g2_decap_8 FILLER_26_11 ();
 sg13g2_decap_8 FILLER_26_18 ();
 sg13g2_decap_8 FILLER_26_25 ();
 sg13g2_decap_8 FILLER_26_32 ();
 sg13g2_decap_8 FILLER_26_39 ();
 sg13g2_decap_8 FILLER_26_46 ();
 sg13g2_fill_1 FILLER_26_53 ();
 sg13g2_decap_8 FILLER_26_62 ();
 sg13g2_decap_8 FILLER_26_69 ();
 sg13g2_decap_8 FILLER_26_76 ();
 sg13g2_decap_8 FILLER_26_83 ();
 sg13g2_decap_8 FILLER_26_90 ();
 sg13g2_decap_8 FILLER_26_97 ();
 sg13g2_decap_8 FILLER_26_104 ();
 sg13g2_decap_8 FILLER_26_111 ();
 sg13g2_decap_8 FILLER_26_118 ();
 sg13g2_decap_8 FILLER_26_125 ();
 sg13g2_decap_8 FILLER_26_132 ();
 sg13g2_decap_8 FILLER_26_139 ();
 sg13g2_decap_8 FILLER_26_146 ();
 sg13g2_decap_8 FILLER_26_153 ();
 sg13g2_decap_8 FILLER_26_160 ();
 sg13g2_decap_8 FILLER_26_167 ();
 sg13g2_decap_8 FILLER_26_174 ();
 sg13g2_decap_8 FILLER_26_181 ();
 sg13g2_decap_8 FILLER_26_188 ();
 sg13g2_decap_8 FILLER_26_195 ();
 sg13g2_decap_8 FILLER_26_202 ();
 sg13g2_decap_8 FILLER_26_209 ();
 sg13g2_decap_8 FILLER_26_216 ();
 sg13g2_decap_8 FILLER_26_223 ();
 sg13g2_decap_8 FILLER_26_230 ();
 sg13g2_decap_8 FILLER_26_237 ();
 sg13g2_decap_8 FILLER_26_244 ();
 sg13g2_decap_8 FILLER_26_251 ();
 sg13g2_decap_8 FILLER_26_258 ();
 sg13g2_decap_8 FILLER_26_265 ();
 sg13g2_decap_8 FILLER_26_272 ();
 sg13g2_decap_8 FILLER_26_279 ();
 sg13g2_decap_8 FILLER_26_286 ();
 sg13g2_decap_8 FILLER_26_293 ();
 sg13g2_decap_8 FILLER_26_300 ();
 sg13g2_decap_8 FILLER_26_307 ();
 sg13g2_decap_8 FILLER_26_314 ();
 sg13g2_decap_8 FILLER_26_321 ();
 sg13g2_decap_8 FILLER_26_328 ();
 sg13g2_decap_8 FILLER_26_335 ();
 sg13g2_decap_8 FILLER_26_342 ();
 sg13g2_decap_8 FILLER_26_349 ();
 sg13g2_decap_8 FILLER_26_356 ();
 sg13g2_decap_8 FILLER_26_363 ();
 sg13g2_decap_8 FILLER_26_370 ();
 sg13g2_decap_8 FILLER_26_377 ();
 sg13g2_decap_8 FILLER_26_384 ();
 sg13g2_decap_8 FILLER_26_391 ();
 sg13g2_decap_8 FILLER_26_398 ();
 sg13g2_decap_8 FILLER_26_405 ();
 sg13g2_decap_8 FILLER_26_412 ();
 sg13g2_decap_8 FILLER_26_419 ();
 sg13g2_decap_8 FILLER_26_426 ();
 sg13g2_decap_8 FILLER_26_433 ();
 sg13g2_decap_8 FILLER_26_440 ();
 sg13g2_decap_8 FILLER_26_447 ();
 sg13g2_decap_8 FILLER_26_454 ();
 sg13g2_decap_8 FILLER_26_461 ();
 sg13g2_decap_8 FILLER_26_468 ();
 sg13g2_decap_8 FILLER_26_475 ();
 sg13g2_decap_8 FILLER_26_482 ();
 sg13g2_decap_8 FILLER_26_489 ();
 sg13g2_decap_8 FILLER_26_496 ();
 sg13g2_decap_8 FILLER_26_503 ();
 sg13g2_decap_8 FILLER_26_510 ();
 sg13g2_decap_8 FILLER_26_517 ();
 sg13g2_decap_8 FILLER_26_524 ();
 sg13g2_decap_8 FILLER_26_531 ();
 sg13g2_decap_8 FILLER_26_538 ();
 sg13g2_decap_8 FILLER_26_545 ();
 sg13g2_decap_8 FILLER_26_552 ();
 sg13g2_decap_8 FILLER_26_559 ();
 sg13g2_decap_8 FILLER_26_566 ();
 sg13g2_decap_8 FILLER_26_573 ();
 sg13g2_decap_8 FILLER_26_580 ();
 sg13g2_decap_8 FILLER_26_587 ();
 sg13g2_decap_8 FILLER_26_594 ();
 sg13g2_decap_8 FILLER_26_601 ();
 sg13g2_decap_8 FILLER_26_608 ();
 sg13g2_decap_8 FILLER_26_615 ();
 sg13g2_decap_8 FILLER_26_622 ();
 sg13g2_decap_8 FILLER_26_629 ();
 sg13g2_decap_8 FILLER_26_636 ();
 sg13g2_decap_8 FILLER_26_643 ();
 sg13g2_decap_8 FILLER_26_650 ();
 sg13g2_decap_8 FILLER_26_657 ();
 sg13g2_decap_8 FILLER_26_664 ();
 sg13g2_decap_8 FILLER_26_671 ();
 sg13g2_decap_8 FILLER_26_678 ();
 sg13g2_decap_8 FILLER_26_685 ();
 sg13g2_decap_8 FILLER_26_692 ();
 sg13g2_decap_8 FILLER_26_699 ();
 sg13g2_decap_8 FILLER_26_706 ();
 sg13g2_decap_8 FILLER_26_713 ();
 sg13g2_decap_8 FILLER_26_720 ();
 sg13g2_decap_8 FILLER_26_727 ();
 sg13g2_decap_8 FILLER_26_734 ();
 sg13g2_decap_8 FILLER_26_741 ();
 sg13g2_decap_8 FILLER_26_748 ();
 sg13g2_decap_8 FILLER_26_755 ();
 sg13g2_decap_8 FILLER_26_762 ();
 sg13g2_decap_8 FILLER_26_769 ();
 sg13g2_decap_8 FILLER_26_776 ();
 sg13g2_decap_8 FILLER_26_783 ();
 sg13g2_decap_8 FILLER_26_790 ();
 sg13g2_decap_8 FILLER_26_797 ();
 sg13g2_decap_8 FILLER_26_804 ();
 sg13g2_decap_8 FILLER_26_811 ();
 sg13g2_decap_8 FILLER_26_818 ();
 sg13g2_decap_8 FILLER_26_825 ();
 sg13g2_decap_8 FILLER_26_832 ();
 sg13g2_decap_8 FILLER_26_839 ();
 sg13g2_decap_8 FILLER_26_846 ();
 sg13g2_decap_8 FILLER_26_853 ();
 sg13g2_decap_8 FILLER_26_860 ();
 sg13g2_decap_8 FILLER_26_867 ();
 sg13g2_decap_8 FILLER_26_874 ();
 sg13g2_decap_8 FILLER_26_881 ();
 sg13g2_decap_8 FILLER_26_888 ();
 sg13g2_decap_8 FILLER_26_895 ();
 sg13g2_decap_8 FILLER_26_902 ();
 sg13g2_decap_8 FILLER_26_909 ();
 sg13g2_decap_8 FILLER_26_916 ();
 sg13g2_decap_8 FILLER_26_923 ();
 sg13g2_decap_8 FILLER_26_930 ();
 sg13g2_decap_8 FILLER_26_937 ();
 sg13g2_decap_8 FILLER_26_944 ();
 sg13g2_decap_8 FILLER_26_951 ();
 sg13g2_decap_8 FILLER_26_958 ();
 sg13g2_decap_8 FILLER_26_965 ();
 sg13g2_decap_8 FILLER_26_972 ();
 sg13g2_decap_8 FILLER_26_979 ();
 sg13g2_decap_8 FILLER_26_986 ();
 sg13g2_decap_8 FILLER_26_993 ();
 sg13g2_decap_8 FILLER_26_1000 ();
 sg13g2_decap_8 FILLER_26_1007 ();
 sg13g2_decap_8 FILLER_26_1014 ();
 sg13g2_decap_8 FILLER_26_1021 ();
 sg13g2_fill_1 FILLER_26_1028 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_4 FILLER_27_14 ();
 sg13g2_fill_1 FILLER_27_18 ();
 sg13g2_decap_8 FILLER_27_32 ();
 sg13g2_decap_8 FILLER_27_39 ();
 sg13g2_decap_4 FILLER_27_46 ();
 sg13g2_fill_1 FILLER_27_50 ();
 sg13g2_decap_8 FILLER_27_67 ();
 sg13g2_decap_8 FILLER_27_74 ();
 sg13g2_decap_8 FILLER_27_81 ();
 sg13g2_decap_8 FILLER_27_88 ();
 sg13g2_decap_8 FILLER_27_95 ();
 sg13g2_decap_8 FILLER_27_102 ();
 sg13g2_decap_4 FILLER_27_109 ();
 sg13g2_decap_8 FILLER_27_121 ();
 sg13g2_decap_8 FILLER_27_128 ();
 sg13g2_decap_8 FILLER_27_135 ();
 sg13g2_decap_8 FILLER_27_142 ();
 sg13g2_decap_8 FILLER_27_149 ();
 sg13g2_decap_8 FILLER_27_156 ();
 sg13g2_decap_8 FILLER_27_163 ();
 sg13g2_decap_8 FILLER_27_170 ();
 sg13g2_decap_8 FILLER_27_177 ();
 sg13g2_decap_8 FILLER_27_184 ();
 sg13g2_decap_8 FILLER_27_191 ();
 sg13g2_decap_8 FILLER_27_198 ();
 sg13g2_decap_8 FILLER_27_205 ();
 sg13g2_decap_8 FILLER_27_212 ();
 sg13g2_decap_8 FILLER_27_219 ();
 sg13g2_decap_8 FILLER_27_226 ();
 sg13g2_decap_8 FILLER_27_233 ();
 sg13g2_decap_8 FILLER_27_240 ();
 sg13g2_decap_8 FILLER_27_247 ();
 sg13g2_decap_8 FILLER_27_254 ();
 sg13g2_decap_8 FILLER_27_261 ();
 sg13g2_decap_8 FILLER_27_268 ();
 sg13g2_decap_8 FILLER_27_275 ();
 sg13g2_decap_8 FILLER_27_282 ();
 sg13g2_decap_8 FILLER_27_289 ();
 sg13g2_decap_8 FILLER_27_296 ();
 sg13g2_decap_8 FILLER_27_303 ();
 sg13g2_decap_8 FILLER_27_310 ();
 sg13g2_decap_8 FILLER_27_317 ();
 sg13g2_decap_8 FILLER_27_324 ();
 sg13g2_decap_8 FILLER_27_331 ();
 sg13g2_decap_8 FILLER_27_338 ();
 sg13g2_decap_8 FILLER_27_345 ();
 sg13g2_decap_8 FILLER_27_352 ();
 sg13g2_decap_8 FILLER_27_359 ();
 sg13g2_decap_8 FILLER_27_366 ();
 sg13g2_decap_8 FILLER_27_373 ();
 sg13g2_decap_8 FILLER_27_380 ();
 sg13g2_decap_8 FILLER_27_387 ();
 sg13g2_decap_8 FILLER_27_394 ();
 sg13g2_decap_8 FILLER_27_401 ();
 sg13g2_decap_8 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_27_415 ();
 sg13g2_decap_8 FILLER_27_422 ();
 sg13g2_decap_8 FILLER_27_429 ();
 sg13g2_decap_8 FILLER_27_436 ();
 sg13g2_decap_8 FILLER_27_443 ();
 sg13g2_decap_8 FILLER_27_450 ();
 sg13g2_decap_8 FILLER_27_457 ();
 sg13g2_decap_8 FILLER_27_464 ();
 sg13g2_decap_8 FILLER_27_471 ();
 sg13g2_decap_8 FILLER_27_478 ();
 sg13g2_decap_8 FILLER_27_485 ();
 sg13g2_decap_8 FILLER_27_492 ();
 sg13g2_decap_8 FILLER_27_499 ();
 sg13g2_decap_8 FILLER_27_506 ();
 sg13g2_decap_8 FILLER_27_513 ();
 sg13g2_decap_8 FILLER_27_520 ();
 sg13g2_decap_8 FILLER_27_527 ();
 sg13g2_decap_8 FILLER_27_534 ();
 sg13g2_decap_8 FILLER_27_541 ();
 sg13g2_decap_8 FILLER_27_548 ();
 sg13g2_decap_8 FILLER_27_555 ();
 sg13g2_decap_8 FILLER_27_562 ();
 sg13g2_decap_8 FILLER_27_569 ();
 sg13g2_decap_8 FILLER_27_576 ();
 sg13g2_decap_8 FILLER_27_583 ();
 sg13g2_decap_8 FILLER_27_590 ();
 sg13g2_decap_8 FILLER_27_597 ();
 sg13g2_decap_8 FILLER_27_604 ();
 sg13g2_decap_8 FILLER_27_611 ();
 sg13g2_decap_8 FILLER_27_618 ();
 sg13g2_decap_8 FILLER_27_625 ();
 sg13g2_decap_8 FILLER_27_632 ();
 sg13g2_decap_8 FILLER_27_639 ();
 sg13g2_decap_8 FILLER_27_646 ();
 sg13g2_decap_8 FILLER_27_653 ();
 sg13g2_decap_8 FILLER_27_660 ();
 sg13g2_decap_8 FILLER_27_667 ();
 sg13g2_decap_8 FILLER_27_674 ();
 sg13g2_decap_8 FILLER_27_681 ();
 sg13g2_decap_8 FILLER_27_688 ();
 sg13g2_decap_8 FILLER_27_695 ();
 sg13g2_decap_8 FILLER_27_702 ();
 sg13g2_decap_8 FILLER_27_709 ();
 sg13g2_decap_8 FILLER_27_716 ();
 sg13g2_decap_8 FILLER_27_723 ();
 sg13g2_decap_8 FILLER_27_730 ();
 sg13g2_decap_8 FILLER_27_737 ();
 sg13g2_decap_8 FILLER_27_744 ();
 sg13g2_decap_8 FILLER_27_751 ();
 sg13g2_decap_8 FILLER_27_758 ();
 sg13g2_decap_8 FILLER_27_765 ();
 sg13g2_decap_8 FILLER_27_772 ();
 sg13g2_decap_8 FILLER_27_779 ();
 sg13g2_decap_8 FILLER_27_786 ();
 sg13g2_decap_8 FILLER_27_793 ();
 sg13g2_decap_8 FILLER_27_800 ();
 sg13g2_decap_8 FILLER_27_807 ();
 sg13g2_decap_8 FILLER_27_814 ();
 sg13g2_decap_8 FILLER_27_821 ();
 sg13g2_decap_8 FILLER_27_828 ();
 sg13g2_decap_8 FILLER_27_835 ();
 sg13g2_decap_8 FILLER_27_842 ();
 sg13g2_decap_8 FILLER_27_849 ();
 sg13g2_decap_8 FILLER_27_856 ();
 sg13g2_decap_8 FILLER_27_863 ();
 sg13g2_decap_8 FILLER_27_870 ();
 sg13g2_decap_8 FILLER_27_877 ();
 sg13g2_decap_8 FILLER_27_884 ();
 sg13g2_decap_8 FILLER_27_891 ();
 sg13g2_decap_8 FILLER_27_898 ();
 sg13g2_decap_8 FILLER_27_905 ();
 sg13g2_decap_8 FILLER_27_912 ();
 sg13g2_decap_8 FILLER_27_919 ();
 sg13g2_decap_8 FILLER_27_926 ();
 sg13g2_decap_8 FILLER_27_933 ();
 sg13g2_decap_8 FILLER_27_940 ();
 sg13g2_decap_8 FILLER_27_947 ();
 sg13g2_decap_8 FILLER_27_954 ();
 sg13g2_decap_8 FILLER_27_961 ();
 sg13g2_decap_8 FILLER_27_968 ();
 sg13g2_decap_8 FILLER_27_975 ();
 sg13g2_decap_8 FILLER_27_982 ();
 sg13g2_decap_8 FILLER_27_989 ();
 sg13g2_decap_8 FILLER_27_996 ();
 sg13g2_decap_8 FILLER_27_1003 ();
 sg13g2_decap_8 FILLER_27_1010 ();
 sg13g2_decap_8 FILLER_27_1017 ();
 sg13g2_decap_4 FILLER_27_1024 ();
 sg13g2_fill_1 FILLER_27_1028 ();
 sg13g2_decap_8 FILLER_28_4 ();
 sg13g2_decap_8 FILLER_28_11 ();
 sg13g2_decap_8 FILLER_28_18 ();
 sg13g2_decap_8 FILLER_28_25 ();
 sg13g2_decap_8 FILLER_28_32 ();
 sg13g2_decap_8 FILLER_28_39 ();
 sg13g2_decap_8 FILLER_28_46 ();
 sg13g2_fill_2 FILLER_28_53 ();
 sg13g2_fill_1 FILLER_28_55 ();
 sg13g2_decap_8 FILLER_28_61 ();
 sg13g2_decap_8 FILLER_28_68 ();
 sg13g2_decap_8 FILLER_28_75 ();
 sg13g2_decap_8 FILLER_28_82 ();
 sg13g2_decap_8 FILLER_28_89 ();
 sg13g2_fill_2 FILLER_28_96 ();
 sg13g2_decap_8 FILLER_28_106 ();
 sg13g2_fill_2 FILLER_28_117 ();
 sg13g2_decap_4 FILLER_28_124 ();
 sg13g2_decap_4 FILLER_28_132 ();
 sg13g2_fill_2 FILLER_28_136 ();
 sg13g2_decap_8 FILLER_28_146 ();
 sg13g2_decap_8 FILLER_28_153 ();
 sg13g2_decap_8 FILLER_28_160 ();
 sg13g2_decap_8 FILLER_28_167 ();
 sg13g2_decap_8 FILLER_28_174 ();
 sg13g2_decap_8 FILLER_28_181 ();
 sg13g2_decap_8 FILLER_28_188 ();
 sg13g2_decap_8 FILLER_28_195 ();
 sg13g2_decap_8 FILLER_28_202 ();
 sg13g2_decap_8 FILLER_28_209 ();
 sg13g2_decap_8 FILLER_28_216 ();
 sg13g2_decap_8 FILLER_28_223 ();
 sg13g2_decap_8 FILLER_28_230 ();
 sg13g2_decap_8 FILLER_28_237 ();
 sg13g2_decap_8 FILLER_28_244 ();
 sg13g2_decap_8 FILLER_28_251 ();
 sg13g2_decap_8 FILLER_28_258 ();
 sg13g2_decap_8 FILLER_28_265 ();
 sg13g2_decap_8 FILLER_28_272 ();
 sg13g2_decap_8 FILLER_28_279 ();
 sg13g2_decap_8 FILLER_28_286 ();
 sg13g2_decap_8 FILLER_28_293 ();
 sg13g2_decap_8 FILLER_28_300 ();
 sg13g2_decap_8 FILLER_28_307 ();
 sg13g2_decap_8 FILLER_28_314 ();
 sg13g2_decap_8 FILLER_28_321 ();
 sg13g2_decap_8 FILLER_28_328 ();
 sg13g2_decap_8 FILLER_28_335 ();
 sg13g2_decap_8 FILLER_28_342 ();
 sg13g2_decap_8 FILLER_28_349 ();
 sg13g2_decap_8 FILLER_28_356 ();
 sg13g2_decap_8 FILLER_28_363 ();
 sg13g2_decap_8 FILLER_28_370 ();
 sg13g2_decap_8 FILLER_28_377 ();
 sg13g2_decap_8 FILLER_28_384 ();
 sg13g2_decap_8 FILLER_28_391 ();
 sg13g2_decap_8 FILLER_28_398 ();
 sg13g2_decap_8 FILLER_28_405 ();
 sg13g2_decap_8 FILLER_28_412 ();
 sg13g2_decap_8 FILLER_28_419 ();
 sg13g2_decap_8 FILLER_28_426 ();
 sg13g2_decap_8 FILLER_28_433 ();
 sg13g2_decap_8 FILLER_28_440 ();
 sg13g2_decap_8 FILLER_28_447 ();
 sg13g2_decap_8 FILLER_28_454 ();
 sg13g2_decap_8 FILLER_28_461 ();
 sg13g2_decap_8 FILLER_28_468 ();
 sg13g2_decap_8 FILLER_28_475 ();
 sg13g2_decap_8 FILLER_28_482 ();
 sg13g2_decap_8 FILLER_28_489 ();
 sg13g2_decap_8 FILLER_28_496 ();
 sg13g2_decap_8 FILLER_28_503 ();
 sg13g2_decap_8 FILLER_28_510 ();
 sg13g2_decap_8 FILLER_28_517 ();
 sg13g2_decap_8 FILLER_28_524 ();
 sg13g2_decap_8 FILLER_28_531 ();
 sg13g2_decap_8 FILLER_28_538 ();
 sg13g2_decap_8 FILLER_28_545 ();
 sg13g2_decap_8 FILLER_28_552 ();
 sg13g2_decap_8 FILLER_28_559 ();
 sg13g2_decap_8 FILLER_28_566 ();
 sg13g2_decap_8 FILLER_28_573 ();
 sg13g2_decap_8 FILLER_28_580 ();
 sg13g2_decap_8 FILLER_28_587 ();
 sg13g2_decap_8 FILLER_28_594 ();
 sg13g2_decap_8 FILLER_28_601 ();
 sg13g2_decap_8 FILLER_28_608 ();
 sg13g2_decap_8 FILLER_28_615 ();
 sg13g2_decap_8 FILLER_28_622 ();
 sg13g2_decap_8 FILLER_28_629 ();
 sg13g2_decap_8 FILLER_28_636 ();
 sg13g2_decap_8 FILLER_28_643 ();
 sg13g2_decap_8 FILLER_28_650 ();
 sg13g2_decap_8 FILLER_28_657 ();
 sg13g2_decap_8 FILLER_28_664 ();
 sg13g2_decap_8 FILLER_28_671 ();
 sg13g2_decap_8 FILLER_28_678 ();
 sg13g2_decap_8 FILLER_28_685 ();
 sg13g2_decap_8 FILLER_28_692 ();
 sg13g2_decap_8 FILLER_28_699 ();
 sg13g2_decap_8 FILLER_28_706 ();
 sg13g2_decap_8 FILLER_28_713 ();
 sg13g2_decap_8 FILLER_28_720 ();
 sg13g2_decap_8 FILLER_28_727 ();
 sg13g2_decap_8 FILLER_28_734 ();
 sg13g2_decap_8 FILLER_28_741 ();
 sg13g2_decap_8 FILLER_28_748 ();
 sg13g2_decap_8 FILLER_28_755 ();
 sg13g2_decap_8 FILLER_28_762 ();
 sg13g2_decap_8 FILLER_28_769 ();
 sg13g2_decap_8 FILLER_28_776 ();
 sg13g2_decap_8 FILLER_28_783 ();
 sg13g2_decap_8 FILLER_28_790 ();
 sg13g2_decap_8 FILLER_28_797 ();
 sg13g2_decap_8 FILLER_28_804 ();
 sg13g2_decap_8 FILLER_28_811 ();
 sg13g2_decap_8 FILLER_28_818 ();
 sg13g2_decap_8 FILLER_28_825 ();
 sg13g2_decap_8 FILLER_28_832 ();
 sg13g2_decap_8 FILLER_28_839 ();
 sg13g2_decap_8 FILLER_28_846 ();
 sg13g2_decap_8 FILLER_28_853 ();
 sg13g2_decap_8 FILLER_28_860 ();
 sg13g2_decap_8 FILLER_28_867 ();
 sg13g2_decap_8 FILLER_28_874 ();
 sg13g2_decap_8 FILLER_28_881 ();
 sg13g2_decap_8 FILLER_28_888 ();
 sg13g2_decap_8 FILLER_28_895 ();
 sg13g2_decap_8 FILLER_28_902 ();
 sg13g2_decap_8 FILLER_28_909 ();
 sg13g2_decap_8 FILLER_28_916 ();
 sg13g2_decap_8 FILLER_28_923 ();
 sg13g2_decap_8 FILLER_28_930 ();
 sg13g2_decap_8 FILLER_28_937 ();
 sg13g2_decap_8 FILLER_28_944 ();
 sg13g2_decap_8 FILLER_28_951 ();
 sg13g2_decap_8 FILLER_28_958 ();
 sg13g2_decap_8 FILLER_28_965 ();
 sg13g2_decap_8 FILLER_28_972 ();
 sg13g2_decap_8 FILLER_28_979 ();
 sg13g2_decap_8 FILLER_28_986 ();
 sg13g2_decap_8 FILLER_28_993 ();
 sg13g2_decap_8 FILLER_28_1000 ();
 sg13g2_decap_8 FILLER_28_1007 ();
 sg13g2_decap_8 FILLER_28_1014 ();
 sg13g2_decap_8 FILLER_28_1021 ();
 sg13g2_fill_1 FILLER_28_1028 ();
 sg13g2_decap_8 FILLER_29_4 ();
 sg13g2_decap_8 FILLER_29_11 ();
 sg13g2_decap_8 FILLER_29_18 ();
 sg13g2_decap_8 FILLER_29_25 ();
 sg13g2_decap_8 FILLER_29_32 ();
 sg13g2_decap_8 FILLER_29_39 ();
 sg13g2_decap_8 FILLER_29_46 ();
 sg13g2_decap_8 FILLER_29_53 ();
 sg13g2_decap_8 FILLER_29_60 ();
 sg13g2_decap_8 FILLER_29_67 ();
 sg13g2_decap_8 FILLER_29_74 ();
 sg13g2_decap_8 FILLER_29_81 ();
 sg13g2_decap_8 FILLER_29_88 ();
 sg13g2_decap_8 FILLER_29_95 ();
 sg13g2_decap_8 FILLER_29_102 ();
 sg13g2_decap_8 FILLER_29_109 ();
 sg13g2_decap_8 FILLER_29_116 ();
 sg13g2_decap_8 FILLER_29_123 ();
 sg13g2_decap_8 FILLER_29_130 ();
 sg13g2_decap_8 FILLER_29_137 ();
 sg13g2_decap_8 FILLER_29_144 ();
 sg13g2_decap_8 FILLER_29_151 ();
 sg13g2_decap_8 FILLER_29_158 ();
 sg13g2_decap_8 FILLER_29_165 ();
 sg13g2_decap_8 FILLER_29_172 ();
 sg13g2_decap_8 FILLER_29_179 ();
 sg13g2_decap_8 FILLER_29_186 ();
 sg13g2_decap_8 FILLER_29_193 ();
 sg13g2_decap_8 FILLER_29_200 ();
 sg13g2_decap_8 FILLER_29_207 ();
 sg13g2_decap_8 FILLER_29_214 ();
 sg13g2_decap_8 FILLER_29_221 ();
 sg13g2_decap_8 FILLER_29_228 ();
 sg13g2_decap_8 FILLER_29_235 ();
 sg13g2_decap_8 FILLER_29_242 ();
 sg13g2_decap_8 FILLER_29_249 ();
 sg13g2_decap_8 FILLER_29_256 ();
 sg13g2_decap_8 FILLER_29_263 ();
 sg13g2_decap_8 FILLER_29_270 ();
 sg13g2_decap_8 FILLER_29_277 ();
 sg13g2_decap_8 FILLER_29_284 ();
 sg13g2_decap_8 FILLER_29_291 ();
 sg13g2_decap_8 FILLER_29_298 ();
 sg13g2_decap_8 FILLER_29_305 ();
 sg13g2_decap_8 FILLER_29_312 ();
 sg13g2_decap_8 FILLER_29_319 ();
 sg13g2_decap_8 FILLER_29_326 ();
 sg13g2_decap_8 FILLER_29_333 ();
 sg13g2_decap_8 FILLER_29_340 ();
 sg13g2_decap_8 FILLER_29_347 ();
 sg13g2_decap_8 FILLER_29_354 ();
 sg13g2_decap_8 FILLER_29_361 ();
 sg13g2_decap_8 FILLER_29_368 ();
 sg13g2_decap_8 FILLER_29_375 ();
 sg13g2_decap_8 FILLER_29_382 ();
 sg13g2_decap_8 FILLER_29_389 ();
 sg13g2_decap_8 FILLER_29_396 ();
 sg13g2_decap_8 FILLER_29_403 ();
 sg13g2_decap_8 FILLER_29_410 ();
 sg13g2_decap_8 FILLER_29_417 ();
 sg13g2_decap_8 FILLER_29_424 ();
 sg13g2_decap_8 FILLER_29_431 ();
 sg13g2_decap_8 FILLER_29_438 ();
 sg13g2_decap_8 FILLER_29_445 ();
 sg13g2_decap_8 FILLER_29_452 ();
 sg13g2_decap_8 FILLER_29_459 ();
 sg13g2_decap_8 FILLER_29_466 ();
 sg13g2_decap_8 FILLER_29_473 ();
 sg13g2_decap_8 FILLER_29_480 ();
 sg13g2_decap_8 FILLER_29_487 ();
 sg13g2_decap_8 FILLER_29_494 ();
 sg13g2_decap_8 FILLER_29_501 ();
 sg13g2_decap_8 FILLER_29_508 ();
 sg13g2_decap_8 FILLER_29_515 ();
 sg13g2_decap_8 FILLER_29_522 ();
 sg13g2_decap_8 FILLER_29_529 ();
 sg13g2_decap_8 FILLER_29_536 ();
 sg13g2_decap_8 FILLER_29_543 ();
 sg13g2_decap_8 FILLER_29_550 ();
 sg13g2_decap_8 FILLER_29_557 ();
 sg13g2_decap_8 FILLER_29_564 ();
 sg13g2_decap_8 FILLER_29_571 ();
 sg13g2_decap_8 FILLER_29_578 ();
 sg13g2_decap_8 FILLER_29_585 ();
 sg13g2_decap_8 FILLER_29_592 ();
 sg13g2_decap_8 FILLER_29_599 ();
 sg13g2_decap_8 FILLER_29_606 ();
 sg13g2_decap_8 FILLER_29_613 ();
 sg13g2_decap_8 FILLER_29_620 ();
 sg13g2_decap_8 FILLER_29_627 ();
 sg13g2_decap_8 FILLER_29_634 ();
 sg13g2_decap_8 FILLER_29_641 ();
 sg13g2_decap_8 FILLER_29_648 ();
 sg13g2_decap_8 FILLER_29_655 ();
 sg13g2_decap_8 FILLER_29_662 ();
 sg13g2_decap_8 FILLER_29_669 ();
 sg13g2_decap_8 FILLER_29_676 ();
 sg13g2_decap_8 FILLER_29_683 ();
 sg13g2_decap_8 FILLER_29_690 ();
 sg13g2_decap_8 FILLER_29_697 ();
 sg13g2_decap_8 FILLER_29_704 ();
 sg13g2_decap_8 FILLER_29_711 ();
 sg13g2_decap_8 FILLER_29_718 ();
 sg13g2_decap_8 FILLER_29_725 ();
 sg13g2_decap_8 FILLER_29_732 ();
 sg13g2_decap_8 FILLER_29_739 ();
 sg13g2_decap_8 FILLER_29_746 ();
 sg13g2_decap_8 FILLER_29_753 ();
 sg13g2_decap_8 FILLER_29_760 ();
 sg13g2_decap_8 FILLER_29_767 ();
 sg13g2_decap_8 FILLER_29_774 ();
 sg13g2_decap_8 FILLER_29_781 ();
 sg13g2_decap_8 FILLER_29_788 ();
 sg13g2_decap_8 FILLER_29_795 ();
 sg13g2_decap_8 FILLER_29_802 ();
 sg13g2_decap_8 FILLER_29_809 ();
 sg13g2_decap_8 FILLER_29_816 ();
 sg13g2_decap_8 FILLER_29_823 ();
 sg13g2_decap_8 FILLER_29_830 ();
 sg13g2_decap_8 FILLER_29_837 ();
 sg13g2_decap_8 FILLER_29_844 ();
 sg13g2_decap_8 FILLER_29_851 ();
 sg13g2_decap_8 FILLER_29_858 ();
 sg13g2_decap_8 FILLER_29_865 ();
 sg13g2_decap_8 FILLER_29_872 ();
 sg13g2_decap_8 FILLER_29_879 ();
 sg13g2_decap_8 FILLER_29_886 ();
 sg13g2_decap_8 FILLER_29_893 ();
 sg13g2_decap_8 FILLER_29_900 ();
 sg13g2_decap_8 FILLER_29_907 ();
 sg13g2_decap_8 FILLER_29_914 ();
 sg13g2_decap_8 FILLER_29_921 ();
 sg13g2_decap_8 FILLER_29_928 ();
 sg13g2_decap_8 FILLER_29_935 ();
 sg13g2_decap_8 FILLER_29_942 ();
 sg13g2_decap_8 FILLER_29_949 ();
 sg13g2_decap_8 FILLER_29_956 ();
 sg13g2_decap_8 FILLER_29_963 ();
 sg13g2_decap_8 FILLER_29_970 ();
 sg13g2_decap_8 FILLER_29_977 ();
 sg13g2_decap_8 FILLER_29_984 ();
 sg13g2_decap_8 FILLER_29_991 ();
 sg13g2_decap_8 FILLER_29_998 ();
 sg13g2_decap_8 FILLER_29_1005 ();
 sg13g2_decap_8 FILLER_29_1012 ();
 sg13g2_decap_8 FILLER_29_1019 ();
 sg13g2_fill_2 FILLER_29_1026 ();
 sg13g2_fill_1 FILLER_29_1028 ();
 sg13g2_decap_8 FILLER_30_4 ();
 sg13g2_decap_8 FILLER_30_11 ();
 sg13g2_decap_8 FILLER_30_18 ();
 sg13g2_decap_8 FILLER_30_25 ();
 sg13g2_decap_8 FILLER_30_32 ();
 sg13g2_decap_8 FILLER_30_39 ();
 sg13g2_decap_8 FILLER_30_46 ();
 sg13g2_decap_8 FILLER_30_53 ();
 sg13g2_decap_8 FILLER_30_60 ();
 sg13g2_decap_8 FILLER_30_67 ();
 sg13g2_decap_8 FILLER_30_74 ();
 sg13g2_decap_8 FILLER_30_81 ();
 sg13g2_decap_8 FILLER_30_88 ();
 sg13g2_decap_8 FILLER_30_95 ();
 sg13g2_decap_8 FILLER_30_102 ();
 sg13g2_decap_8 FILLER_30_109 ();
 sg13g2_fill_2 FILLER_30_116 ();
 sg13g2_decap_8 FILLER_30_123 ();
 sg13g2_decap_8 FILLER_30_130 ();
 sg13g2_decap_8 FILLER_30_137 ();
 sg13g2_decap_8 FILLER_30_144 ();
 sg13g2_decap_8 FILLER_30_151 ();
 sg13g2_decap_8 FILLER_30_158 ();
 sg13g2_decap_8 FILLER_30_165 ();
 sg13g2_decap_8 FILLER_30_172 ();
 sg13g2_decap_8 FILLER_30_179 ();
 sg13g2_decap_8 FILLER_30_186 ();
 sg13g2_decap_8 FILLER_30_193 ();
 sg13g2_decap_8 FILLER_30_200 ();
 sg13g2_decap_8 FILLER_30_207 ();
 sg13g2_decap_8 FILLER_30_214 ();
 sg13g2_decap_8 FILLER_30_221 ();
 sg13g2_decap_8 FILLER_30_228 ();
 sg13g2_decap_8 FILLER_30_235 ();
 sg13g2_decap_8 FILLER_30_242 ();
 sg13g2_decap_8 FILLER_30_249 ();
 sg13g2_decap_8 FILLER_30_256 ();
 sg13g2_decap_8 FILLER_30_263 ();
 sg13g2_decap_8 FILLER_30_270 ();
 sg13g2_decap_8 FILLER_30_277 ();
 sg13g2_decap_8 FILLER_30_284 ();
 sg13g2_decap_8 FILLER_30_291 ();
 sg13g2_decap_8 FILLER_30_298 ();
 sg13g2_decap_8 FILLER_30_305 ();
 sg13g2_decap_8 FILLER_30_312 ();
 sg13g2_decap_8 FILLER_30_319 ();
 sg13g2_decap_8 FILLER_30_326 ();
 sg13g2_decap_8 FILLER_30_333 ();
 sg13g2_decap_8 FILLER_30_340 ();
 sg13g2_decap_8 FILLER_30_347 ();
 sg13g2_decap_8 FILLER_30_354 ();
 sg13g2_decap_8 FILLER_30_361 ();
 sg13g2_decap_8 FILLER_30_368 ();
 sg13g2_decap_8 FILLER_30_375 ();
 sg13g2_decap_8 FILLER_30_382 ();
 sg13g2_decap_8 FILLER_30_389 ();
 sg13g2_decap_8 FILLER_30_396 ();
 sg13g2_decap_8 FILLER_30_403 ();
 sg13g2_decap_8 FILLER_30_410 ();
 sg13g2_decap_8 FILLER_30_417 ();
 sg13g2_decap_8 FILLER_30_424 ();
 sg13g2_decap_8 FILLER_30_431 ();
 sg13g2_decap_8 FILLER_30_438 ();
 sg13g2_decap_8 FILLER_30_445 ();
 sg13g2_decap_8 FILLER_30_452 ();
 sg13g2_decap_8 FILLER_30_459 ();
 sg13g2_decap_8 FILLER_30_466 ();
 sg13g2_decap_8 FILLER_30_473 ();
 sg13g2_decap_8 FILLER_30_480 ();
 sg13g2_decap_8 FILLER_30_487 ();
 sg13g2_decap_8 FILLER_30_494 ();
 sg13g2_decap_8 FILLER_30_501 ();
 sg13g2_decap_8 FILLER_30_508 ();
 sg13g2_decap_8 FILLER_30_515 ();
 sg13g2_decap_8 FILLER_30_522 ();
 sg13g2_decap_8 FILLER_30_529 ();
 sg13g2_decap_8 FILLER_30_536 ();
 sg13g2_decap_8 FILLER_30_543 ();
 sg13g2_decap_8 FILLER_30_550 ();
 sg13g2_decap_8 FILLER_30_557 ();
 sg13g2_decap_8 FILLER_30_564 ();
 sg13g2_decap_8 FILLER_30_571 ();
 sg13g2_decap_8 FILLER_30_578 ();
 sg13g2_decap_8 FILLER_30_585 ();
 sg13g2_decap_8 FILLER_30_592 ();
 sg13g2_decap_8 FILLER_30_599 ();
 sg13g2_decap_8 FILLER_30_606 ();
 sg13g2_decap_8 FILLER_30_613 ();
 sg13g2_decap_8 FILLER_30_620 ();
 sg13g2_decap_8 FILLER_30_627 ();
 sg13g2_decap_8 FILLER_30_634 ();
 sg13g2_decap_8 FILLER_30_641 ();
 sg13g2_decap_8 FILLER_30_648 ();
 sg13g2_decap_8 FILLER_30_655 ();
 sg13g2_decap_8 FILLER_30_662 ();
 sg13g2_decap_8 FILLER_30_669 ();
 sg13g2_decap_8 FILLER_30_676 ();
 sg13g2_decap_8 FILLER_30_683 ();
 sg13g2_decap_8 FILLER_30_690 ();
 sg13g2_decap_8 FILLER_30_697 ();
 sg13g2_decap_8 FILLER_30_704 ();
 sg13g2_decap_8 FILLER_30_711 ();
 sg13g2_decap_8 FILLER_30_718 ();
 sg13g2_decap_8 FILLER_30_725 ();
 sg13g2_decap_8 FILLER_30_732 ();
 sg13g2_decap_8 FILLER_30_739 ();
 sg13g2_decap_8 FILLER_30_746 ();
 sg13g2_decap_8 FILLER_30_753 ();
 sg13g2_decap_8 FILLER_30_760 ();
 sg13g2_decap_8 FILLER_30_767 ();
 sg13g2_decap_8 FILLER_30_774 ();
 sg13g2_decap_8 FILLER_30_781 ();
 sg13g2_decap_8 FILLER_30_788 ();
 sg13g2_decap_8 FILLER_30_795 ();
 sg13g2_decap_8 FILLER_30_802 ();
 sg13g2_decap_8 FILLER_30_809 ();
 sg13g2_decap_8 FILLER_30_816 ();
 sg13g2_decap_8 FILLER_30_823 ();
 sg13g2_decap_8 FILLER_30_830 ();
 sg13g2_decap_8 FILLER_30_837 ();
 sg13g2_decap_8 FILLER_30_844 ();
 sg13g2_decap_8 FILLER_30_851 ();
 sg13g2_decap_8 FILLER_30_858 ();
 sg13g2_decap_8 FILLER_30_865 ();
 sg13g2_decap_8 FILLER_30_872 ();
 sg13g2_decap_8 FILLER_30_879 ();
 sg13g2_decap_8 FILLER_30_886 ();
 sg13g2_decap_8 FILLER_30_893 ();
 sg13g2_decap_8 FILLER_30_900 ();
 sg13g2_decap_8 FILLER_30_907 ();
 sg13g2_decap_8 FILLER_30_914 ();
 sg13g2_decap_8 FILLER_30_921 ();
 sg13g2_decap_8 FILLER_30_928 ();
 sg13g2_decap_8 FILLER_30_935 ();
 sg13g2_decap_8 FILLER_30_942 ();
 sg13g2_decap_8 FILLER_30_949 ();
 sg13g2_decap_8 FILLER_30_956 ();
 sg13g2_decap_8 FILLER_30_963 ();
 sg13g2_decap_8 FILLER_30_970 ();
 sg13g2_decap_8 FILLER_30_977 ();
 sg13g2_decap_8 FILLER_30_984 ();
 sg13g2_decap_8 FILLER_30_991 ();
 sg13g2_decap_8 FILLER_30_998 ();
 sg13g2_decap_8 FILLER_30_1005 ();
 sg13g2_decap_8 FILLER_30_1012 ();
 sg13g2_decap_8 FILLER_30_1019 ();
 sg13g2_fill_2 FILLER_30_1026 ();
 sg13g2_fill_1 FILLER_30_1028 ();
 sg13g2_decap_8 FILLER_31_4 ();
 sg13g2_decap_8 FILLER_31_11 ();
 sg13g2_decap_8 FILLER_31_18 ();
 sg13g2_decap_8 FILLER_31_25 ();
 sg13g2_decap_8 FILLER_31_32 ();
 sg13g2_decap_8 FILLER_31_39 ();
 sg13g2_decap_8 FILLER_31_46 ();
 sg13g2_decap_8 FILLER_31_53 ();
 sg13g2_decap_8 FILLER_31_60 ();
 sg13g2_decap_8 FILLER_31_67 ();
 sg13g2_decap_8 FILLER_31_74 ();
 sg13g2_decap_8 FILLER_31_81 ();
 sg13g2_decap_8 FILLER_31_88 ();
 sg13g2_decap_8 FILLER_31_95 ();
 sg13g2_decap_8 FILLER_31_102 ();
 sg13g2_decap_8 FILLER_31_114 ();
 sg13g2_decap_8 FILLER_31_121 ();
 sg13g2_fill_1 FILLER_31_128 ();
 sg13g2_fill_1 FILLER_31_134 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_decap_8 FILLER_31_182 ();
 sg13g2_decap_8 FILLER_31_189 ();
 sg13g2_decap_8 FILLER_31_196 ();
 sg13g2_decap_8 FILLER_31_203 ();
 sg13g2_decap_8 FILLER_31_210 ();
 sg13g2_decap_8 FILLER_31_217 ();
 sg13g2_decap_8 FILLER_31_224 ();
 sg13g2_decap_8 FILLER_31_231 ();
 sg13g2_decap_8 FILLER_31_238 ();
 sg13g2_decap_8 FILLER_31_245 ();
 sg13g2_decap_8 FILLER_31_252 ();
 sg13g2_decap_8 FILLER_31_259 ();
 sg13g2_decap_8 FILLER_31_266 ();
 sg13g2_decap_8 FILLER_31_273 ();
 sg13g2_decap_8 FILLER_31_280 ();
 sg13g2_decap_8 FILLER_31_287 ();
 sg13g2_decap_8 FILLER_31_294 ();
 sg13g2_decap_8 FILLER_31_301 ();
 sg13g2_decap_8 FILLER_31_308 ();
 sg13g2_decap_8 FILLER_31_315 ();
 sg13g2_decap_8 FILLER_31_322 ();
 sg13g2_decap_8 FILLER_31_329 ();
 sg13g2_decap_8 FILLER_31_336 ();
 sg13g2_decap_8 FILLER_31_343 ();
 sg13g2_decap_8 FILLER_31_350 ();
 sg13g2_decap_8 FILLER_31_357 ();
 sg13g2_decap_8 FILLER_31_364 ();
 sg13g2_decap_8 FILLER_31_371 ();
 sg13g2_decap_8 FILLER_31_378 ();
 sg13g2_decap_8 FILLER_31_385 ();
 sg13g2_decap_8 FILLER_31_392 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_decap_8 FILLER_31_406 ();
 sg13g2_decap_8 FILLER_31_413 ();
 sg13g2_decap_8 FILLER_31_420 ();
 sg13g2_decap_8 FILLER_31_427 ();
 sg13g2_decap_8 FILLER_31_434 ();
 sg13g2_decap_8 FILLER_31_441 ();
 sg13g2_decap_8 FILLER_31_448 ();
 sg13g2_decap_8 FILLER_31_455 ();
 sg13g2_decap_8 FILLER_31_462 ();
 sg13g2_decap_8 FILLER_31_469 ();
 sg13g2_decap_8 FILLER_31_476 ();
 sg13g2_decap_8 FILLER_31_483 ();
 sg13g2_decap_8 FILLER_31_490 ();
 sg13g2_decap_8 FILLER_31_497 ();
 sg13g2_decap_8 FILLER_31_504 ();
 sg13g2_decap_8 FILLER_31_511 ();
 sg13g2_decap_8 FILLER_31_518 ();
 sg13g2_decap_8 FILLER_31_525 ();
 sg13g2_decap_8 FILLER_31_532 ();
 sg13g2_decap_8 FILLER_31_539 ();
 sg13g2_decap_8 FILLER_31_546 ();
 sg13g2_decap_8 FILLER_31_553 ();
 sg13g2_decap_8 FILLER_31_560 ();
 sg13g2_decap_8 FILLER_31_567 ();
 sg13g2_decap_8 FILLER_31_574 ();
 sg13g2_decap_8 FILLER_31_581 ();
 sg13g2_decap_8 FILLER_31_588 ();
 sg13g2_decap_8 FILLER_31_595 ();
 sg13g2_decap_8 FILLER_31_602 ();
 sg13g2_decap_8 FILLER_31_609 ();
 sg13g2_decap_8 FILLER_31_616 ();
 sg13g2_decap_8 FILLER_31_623 ();
 sg13g2_decap_8 FILLER_31_630 ();
 sg13g2_decap_8 FILLER_31_637 ();
 sg13g2_decap_8 FILLER_31_644 ();
 sg13g2_decap_8 FILLER_31_651 ();
 sg13g2_decap_8 FILLER_31_658 ();
 sg13g2_decap_8 FILLER_31_665 ();
 sg13g2_decap_8 FILLER_31_672 ();
 sg13g2_decap_8 FILLER_31_679 ();
 sg13g2_decap_8 FILLER_31_686 ();
 sg13g2_decap_8 FILLER_31_693 ();
 sg13g2_decap_8 FILLER_31_700 ();
 sg13g2_decap_8 FILLER_31_707 ();
 sg13g2_decap_8 FILLER_31_714 ();
 sg13g2_decap_8 FILLER_31_721 ();
 sg13g2_decap_8 FILLER_31_728 ();
 sg13g2_decap_8 FILLER_31_735 ();
 sg13g2_decap_8 FILLER_31_742 ();
 sg13g2_decap_8 FILLER_31_749 ();
 sg13g2_decap_8 FILLER_31_756 ();
 sg13g2_decap_8 FILLER_31_763 ();
 sg13g2_decap_8 FILLER_31_770 ();
 sg13g2_decap_8 FILLER_31_777 ();
 sg13g2_decap_8 FILLER_31_784 ();
 sg13g2_decap_8 FILLER_31_791 ();
 sg13g2_decap_8 FILLER_31_798 ();
 sg13g2_decap_8 FILLER_31_805 ();
 sg13g2_decap_8 FILLER_31_812 ();
 sg13g2_decap_8 FILLER_31_819 ();
 sg13g2_decap_8 FILLER_31_826 ();
 sg13g2_decap_8 FILLER_31_833 ();
 sg13g2_decap_8 FILLER_31_840 ();
 sg13g2_decap_8 FILLER_31_847 ();
 sg13g2_decap_8 FILLER_31_854 ();
 sg13g2_decap_8 FILLER_31_861 ();
 sg13g2_decap_8 FILLER_31_868 ();
 sg13g2_decap_8 FILLER_31_875 ();
 sg13g2_decap_8 FILLER_31_882 ();
 sg13g2_decap_8 FILLER_31_889 ();
 sg13g2_decap_8 FILLER_31_896 ();
 sg13g2_decap_8 FILLER_31_903 ();
 sg13g2_decap_8 FILLER_31_910 ();
 sg13g2_decap_8 FILLER_31_917 ();
 sg13g2_decap_8 FILLER_31_924 ();
 sg13g2_decap_8 FILLER_31_931 ();
 sg13g2_decap_8 FILLER_31_938 ();
 sg13g2_decap_8 FILLER_31_945 ();
 sg13g2_decap_8 FILLER_31_952 ();
 sg13g2_decap_8 FILLER_31_959 ();
 sg13g2_decap_8 FILLER_31_966 ();
 sg13g2_decap_8 FILLER_31_973 ();
 sg13g2_decap_8 FILLER_31_980 ();
 sg13g2_decap_8 FILLER_31_987 ();
 sg13g2_decap_8 FILLER_31_994 ();
 sg13g2_decap_8 FILLER_31_1001 ();
 sg13g2_decap_8 FILLER_31_1008 ();
 sg13g2_decap_8 FILLER_31_1015 ();
 sg13g2_decap_8 FILLER_31_1022 ();
 sg13g2_decap_8 FILLER_32_4 ();
 sg13g2_decap_8 FILLER_32_11 ();
 sg13g2_decap_8 FILLER_32_18 ();
 sg13g2_decap_8 FILLER_32_25 ();
 sg13g2_decap_4 FILLER_32_32 ();
 sg13g2_fill_1 FILLER_32_36 ();
 sg13g2_decap_8 FILLER_32_45 ();
 sg13g2_decap_8 FILLER_32_52 ();
 sg13g2_decap_8 FILLER_32_59 ();
 sg13g2_decap_8 FILLER_32_66 ();
 sg13g2_decap_8 FILLER_32_73 ();
 sg13g2_decap_8 FILLER_32_80 ();
 sg13g2_decap_8 FILLER_32_87 ();
 sg13g2_decap_8 FILLER_32_94 ();
 sg13g2_decap_8 FILLER_32_101 ();
 sg13g2_decap_8 FILLER_32_108 ();
 sg13g2_decap_8 FILLER_32_115 ();
 sg13g2_decap_8 FILLER_32_122 ();
 sg13g2_fill_2 FILLER_32_129 ();
 sg13g2_decap_8 FILLER_32_144 ();
 sg13g2_decap_8 FILLER_32_151 ();
 sg13g2_decap_8 FILLER_32_158 ();
 sg13g2_decap_8 FILLER_32_165 ();
 sg13g2_decap_8 FILLER_32_172 ();
 sg13g2_decap_8 FILLER_32_179 ();
 sg13g2_decap_8 FILLER_32_186 ();
 sg13g2_decap_8 FILLER_32_193 ();
 sg13g2_decap_8 FILLER_32_200 ();
 sg13g2_decap_8 FILLER_32_207 ();
 sg13g2_decap_8 FILLER_32_214 ();
 sg13g2_decap_8 FILLER_32_221 ();
 sg13g2_decap_8 FILLER_32_228 ();
 sg13g2_decap_8 FILLER_32_235 ();
 sg13g2_decap_8 FILLER_32_242 ();
 sg13g2_decap_8 FILLER_32_249 ();
 sg13g2_decap_8 FILLER_32_256 ();
 sg13g2_decap_8 FILLER_32_263 ();
 sg13g2_decap_8 FILLER_32_270 ();
 sg13g2_decap_8 FILLER_32_277 ();
 sg13g2_decap_8 FILLER_32_284 ();
 sg13g2_decap_8 FILLER_32_291 ();
 sg13g2_decap_8 FILLER_32_298 ();
 sg13g2_decap_8 FILLER_32_305 ();
 sg13g2_decap_8 FILLER_32_312 ();
 sg13g2_decap_8 FILLER_32_319 ();
 sg13g2_decap_8 FILLER_32_326 ();
 sg13g2_decap_8 FILLER_32_333 ();
 sg13g2_decap_8 FILLER_32_340 ();
 sg13g2_decap_8 FILLER_32_347 ();
 sg13g2_decap_8 FILLER_32_354 ();
 sg13g2_decap_8 FILLER_32_361 ();
 sg13g2_decap_8 FILLER_32_368 ();
 sg13g2_decap_8 FILLER_32_375 ();
 sg13g2_decap_8 FILLER_32_382 ();
 sg13g2_decap_8 FILLER_32_389 ();
 sg13g2_decap_8 FILLER_32_396 ();
 sg13g2_decap_8 FILLER_32_403 ();
 sg13g2_decap_8 FILLER_32_410 ();
 sg13g2_decap_8 FILLER_32_417 ();
 sg13g2_decap_8 FILLER_32_424 ();
 sg13g2_decap_8 FILLER_32_431 ();
 sg13g2_decap_8 FILLER_32_438 ();
 sg13g2_decap_8 FILLER_32_445 ();
 sg13g2_decap_8 FILLER_32_452 ();
 sg13g2_decap_8 FILLER_32_459 ();
 sg13g2_decap_8 FILLER_32_466 ();
 sg13g2_decap_8 FILLER_32_473 ();
 sg13g2_decap_8 FILLER_32_480 ();
 sg13g2_decap_8 FILLER_32_487 ();
 sg13g2_decap_8 FILLER_32_494 ();
 sg13g2_decap_8 FILLER_32_501 ();
 sg13g2_decap_8 FILLER_32_508 ();
 sg13g2_decap_8 FILLER_32_515 ();
 sg13g2_decap_8 FILLER_32_522 ();
 sg13g2_decap_8 FILLER_32_529 ();
 sg13g2_decap_8 FILLER_32_536 ();
 sg13g2_decap_8 FILLER_32_543 ();
 sg13g2_decap_8 FILLER_32_550 ();
 sg13g2_decap_8 FILLER_32_557 ();
 sg13g2_decap_8 FILLER_32_564 ();
 sg13g2_decap_8 FILLER_32_571 ();
 sg13g2_decap_8 FILLER_32_578 ();
 sg13g2_decap_8 FILLER_32_585 ();
 sg13g2_decap_8 FILLER_32_592 ();
 sg13g2_decap_8 FILLER_32_599 ();
 sg13g2_decap_8 FILLER_32_606 ();
 sg13g2_decap_8 FILLER_32_613 ();
 sg13g2_decap_8 FILLER_32_620 ();
 sg13g2_decap_8 FILLER_32_627 ();
 sg13g2_decap_8 FILLER_32_634 ();
 sg13g2_decap_8 FILLER_32_641 ();
 sg13g2_decap_8 FILLER_32_648 ();
 sg13g2_decap_8 FILLER_32_655 ();
 sg13g2_decap_8 FILLER_32_662 ();
 sg13g2_decap_8 FILLER_32_669 ();
 sg13g2_decap_8 FILLER_32_676 ();
 sg13g2_decap_8 FILLER_32_683 ();
 sg13g2_decap_8 FILLER_32_690 ();
 sg13g2_decap_8 FILLER_32_697 ();
 sg13g2_decap_8 FILLER_32_704 ();
 sg13g2_decap_8 FILLER_32_711 ();
 sg13g2_decap_8 FILLER_32_718 ();
 sg13g2_decap_8 FILLER_32_725 ();
 sg13g2_decap_8 FILLER_32_732 ();
 sg13g2_decap_8 FILLER_32_739 ();
 sg13g2_decap_8 FILLER_32_746 ();
 sg13g2_decap_8 FILLER_32_753 ();
 sg13g2_decap_8 FILLER_32_760 ();
 sg13g2_decap_8 FILLER_32_767 ();
 sg13g2_decap_8 FILLER_32_774 ();
 sg13g2_decap_8 FILLER_32_781 ();
 sg13g2_decap_8 FILLER_32_788 ();
 sg13g2_decap_8 FILLER_32_795 ();
 sg13g2_decap_8 FILLER_32_802 ();
 sg13g2_decap_8 FILLER_32_809 ();
 sg13g2_decap_8 FILLER_32_816 ();
 sg13g2_decap_8 FILLER_32_823 ();
 sg13g2_decap_8 FILLER_32_830 ();
 sg13g2_decap_8 FILLER_32_837 ();
 sg13g2_decap_8 FILLER_32_844 ();
 sg13g2_decap_8 FILLER_32_851 ();
 sg13g2_decap_8 FILLER_32_858 ();
 sg13g2_decap_8 FILLER_32_865 ();
 sg13g2_decap_8 FILLER_32_872 ();
 sg13g2_decap_8 FILLER_32_879 ();
 sg13g2_decap_8 FILLER_32_886 ();
 sg13g2_decap_8 FILLER_32_893 ();
 sg13g2_decap_8 FILLER_32_900 ();
 sg13g2_decap_8 FILLER_32_907 ();
 sg13g2_decap_8 FILLER_32_914 ();
 sg13g2_decap_8 FILLER_32_921 ();
 sg13g2_decap_8 FILLER_32_928 ();
 sg13g2_decap_8 FILLER_32_935 ();
 sg13g2_decap_8 FILLER_32_942 ();
 sg13g2_decap_8 FILLER_32_949 ();
 sg13g2_decap_8 FILLER_32_956 ();
 sg13g2_decap_8 FILLER_32_963 ();
 sg13g2_decap_8 FILLER_32_970 ();
 sg13g2_decap_8 FILLER_32_977 ();
 sg13g2_decap_8 FILLER_32_984 ();
 sg13g2_decap_8 FILLER_32_991 ();
 sg13g2_decap_8 FILLER_32_998 ();
 sg13g2_decap_8 FILLER_32_1005 ();
 sg13g2_decap_8 FILLER_32_1012 ();
 sg13g2_decap_8 FILLER_32_1019 ();
 sg13g2_fill_2 FILLER_32_1026 ();
 sg13g2_fill_1 FILLER_32_1028 ();
 sg13g2_decap_8 FILLER_33_4 ();
 sg13g2_decap_8 FILLER_33_11 ();
 sg13g2_fill_2 FILLER_33_18 ();
 sg13g2_fill_2 FILLER_33_32 ();
 sg13g2_decap_8 FILLER_33_41 ();
 sg13g2_decap_8 FILLER_33_48 ();
 sg13g2_decap_8 FILLER_33_55 ();
 sg13g2_decap_8 FILLER_33_62 ();
 sg13g2_decap_4 FILLER_33_69 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_210 ();
 sg13g2_decap_8 FILLER_33_217 ();
 sg13g2_decap_8 FILLER_33_224 ();
 sg13g2_decap_8 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_238 ();
 sg13g2_decap_8 FILLER_33_245 ();
 sg13g2_decap_8 FILLER_33_252 ();
 sg13g2_decap_8 FILLER_33_259 ();
 sg13g2_decap_8 FILLER_33_266 ();
 sg13g2_decap_8 FILLER_33_273 ();
 sg13g2_decap_8 FILLER_33_280 ();
 sg13g2_decap_8 FILLER_33_287 ();
 sg13g2_decap_8 FILLER_33_294 ();
 sg13g2_decap_8 FILLER_33_301 ();
 sg13g2_decap_8 FILLER_33_308 ();
 sg13g2_decap_8 FILLER_33_315 ();
 sg13g2_decap_8 FILLER_33_322 ();
 sg13g2_decap_8 FILLER_33_329 ();
 sg13g2_decap_8 FILLER_33_336 ();
 sg13g2_decap_8 FILLER_33_343 ();
 sg13g2_decap_8 FILLER_33_350 ();
 sg13g2_decap_8 FILLER_33_357 ();
 sg13g2_decap_8 FILLER_33_364 ();
 sg13g2_decap_8 FILLER_33_371 ();
 sg13g2_decap_8 FILLER_33_378 ();
 sg13g2_decap_8 FILLER_33_385 ();
 sg13g2_decap_8 FILLER_33_392 ();
 sg13g2_decap_8 FILLER_33_399 ();
 sg13g2_decap_8 FILLER_33_406 ();
 sg13g2_decap_8 FILLER_33_413 ();
 sg13g2_decap_8 FILLER_33_420 ();
 sg13g2_decap_8 FILLER_33_427 ();
 sg13g2_decap_8 FILLER_33_434 ();
 sg13g2_decap_8 FILLER_33_441 ();
 sg13g2_decap_8 FILLER_33_448 ();
 sg13g2_decap_8 FILLER_33_455 ();
 sg13g2_decap_8 FILLER_33_462 ();
 sg13g2_decap_8 FILLER_33_469 ();
 sg13g2_decap_8 FILLER_33_476 ();
 sg13g2_decap_8 FILLER_33_483 ();
 sg13g2_decap_8 FILLER_33_490 ();
 sg13g2_decap_8 FILLER_33_497 ();
 sg13g2_decap_8 FILLER_33_504 ();
 sg13g2_decap_8 FILLER_33_511 ();
 sg13g2_decap_8 FILLER_33_518 ();
 sg13g2_decap_8 FILLER_33_525 ();
 sg13g2_decap_8 FILLER_33_532 ();
 sg13g2_decap_8 FILLER_33_539 ();
 sg13g2_decap_8 FILLER_33_546 ();
 sg13g2_decap_8 FILLER_33_553 ();
 sg13g2_decap_8 FILLER_33_560 ();
 sg13g2_decap_8 FILLER_33_567 ();
 sg13g2_decap_8 FILLER_33_574 ();
 sg13g2_decap_8 FILLER_33_581 ();
 sg13g2_decap_8 FILLER_33_588 ();
 sg13g2_decap_8 FILLER_33_595 ();
 sg13g2_decap_8 FILLER_33_602 ();
 sg13g2_decap_8 FILLER_33_609 ();
 sg13g2_decap_8 FILLER_33_616 ();
 sg13g2_decap_8 FILLER_33_623 ();
 sg13g2_decap_8 FILLER_33_630 ();
 sg13g2_decap_8 FILLER_33_637 ();
 sg13g2_decap_8 FILLER_33_644 ();
 sg13g2_decap_8 FILLER_33_651 ();
 sg13g2_decap_8 FILLER_33_658 ();
 sg13g2_decap_8 FILLER_33_665 ();
 sg13g2_decap_8 FILLER_33_672 ();
 sg13g2_decap_8 FILLER_33_679 ();
 sg13g2_decap_8 FILLER_33_686 ();
 sg13g2_decap_8 FILLER_33_693 ();
 sg13g2_decap_8 FILLER_33_700 ();
 sg13g2_decap_8 FILLER_33_707 ();
 sg13g2_decap_8 FILLER_33_714 ();
 sg13g2_decap_8 FILLER_33_721 ();
 sg13g2_decap_8 FILLER_33_728 ();
 sg13g2_decap_8 FILLER_33_735 ();
 sg13g2_decap_8 FILLER_33_742 ();
 sg13g2_decap_8 FILLER_33_749 ();
 sg13g2_decap_8 FILLER_33_756 ();
 sg13g2_decap_8 FILLER_33_763 ();
 sg13g2_decap_8 FILLER_33_770 ();
 sg13g2_decap_8 FILLER_33_777 ();
 sg13g2_decap_8 FILLER_33_784 ();
 sg13g2_decap_8 FILLER_33_791 ();
 sg13g2_decap_8 FILLER_33_798 ();
 sg13g2_decap_8 FILLER_33_805 ();
 sg13g2_decap_8 FILLER_33_812 ();
 sg13g2_decap_8 FILLER_33_819 ();
 sg13g2_decap_8 FILLER_33_826 ();
 sg13g2_decap_8 FILLER_33_833 ();
 sg13g2_decap_8 FILLER_33_840 ();
 sg13g2_decap_8 FILLER_33_847 ();
 sg13g2_decap_8 FILLER_33_854 ();
 sg13g2_decap_8 FILLER_33_861 ();
 sg13g2_decap_8 FILLER_33_868 ();
 sg13g2_decap_8 FILLER_33_875 ();
 sg13g2_decap_8 FILLER_33_882 ();
 sg13g2_decap_8 FILLER_33_889 ();
 sg13g2_decap_8 FILLER_33_896 ();
 sg13g2_decap_8 FILLER_33_903 ();
 sg13g2_decap_8 FILLER_33_910 ();
 sg13g2_decap_8 FILLER_33_917 ();
 sg13g2_decap_8 FILLER_33_924 ();
 sg13g2_decap_8 FILLER_33_931 ();
 sg13g2_decap_8 FILLER_33_938 ();
 sg13g2_decap_8 FILLER_33_945 ();
 sg13g2_decap_8 FILLER_33_952 ();
 sg13g2_decap_8 FILLER_33_959 ();
 sg13g2_decap_8 FILLER_33_966 ();
 sg13g2_decap_8 FILLER_33_973 ();
 sg13g2_decap_8 FILLER_33_980 ();
 sg13g2_decap_8 FILLER_33_987 ();
 sg13g2_decap_8 FILLER_33_994 ();
 sg13g2_decap_8 FILLER_33_1001 ();
 sg13g2_decap_8 FILLER_33_1008 ();
 sg13g2_decap_8 FILLER_33_1015 ();
 sg13g2_decap_8 FILLER_33_1022 ();
 sg13g2_decap_8 FILLER_34_4 ();
 sg13g2_decap_8 FILLER_34_11 ();
 sg13g2_decap_8 FILLER_34_18 ();
 sg13g2_decap_4 FILLER_34_25 ();
 sg13g2_fill_1 FILLER_34_29 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_4 FILLER_34_56 ();
 sg13g2_decap_4 FILLER_34_64 ();
 sg13g2_fill_1 FILLER_34_68 ();
 sg13g2_decap_8 FILLER_34_89 ();
 sg13g2_decap_8 FILLER_34_96 ();
 sg13g2_decap_8 FILLER_34_103 ();
 sg13g2_decap_8 FILLER_34_110 ();
 sg13g2_decap_8 FILLER_34_117 ();
 sg13g2_decap_8 FILLER_34_124 ();
 sg13g2_decap_8 FILLER_34_131 ();
 sg13g2_decap_8 FILLER_34_138 ();
 sg13g2_decap_8 FILLER_34_145 ();
 sg13g2_decap_8 FILLER_34_152 ();
 sg13g2_decap_8 FILLER_34_159 ();
 sg13g2_decap_8 FILLER_34_166 ();
 sg13g2_decap_8 FILLER_34_173 ();
 sg13g2_decap_8 FILLER_34_180 ();
 sg13g2_decap_8 FILLER_34_187 ();
 sg13g2_decap_8 FILLER_34_194 ();
 sg13g2_decap_8 FILLER_34_201 ();
 sg13g2_decap_8 FILLER_34_208 ();
 sg13g2_decap_8 FILLER_34_215 ();
 sg13g2_decap_8 FILLER_34_222 ();
 sg13g2_decap_8 FILLER_34_229 ();
 sg13g2_decap_8 FILLER_34_236 ();
 sg13g2_decap_8 FILLER_34_243 ();
 sg13g2_decap_8 FILLER_34_250 ();
 sg13g2_decap_8 FILLER_34_257 ();
 sg13g2_decap_8 FILLER_34_264 ();
 sg13g2_decap_8 FILLER_34_271 ();
 sg13g2_decap_8 FILLER_34_278 ();
 sg13g2_decap_8 FILLER_34_285 ();
 sg13g2_decap_8 FILLER_34_292 ();
 sg13g2_decap_8 FILLER_34_299 ();
 sg13g2_decap_8 FILLER_34_306 ();
 sg13g2_decap_8 FILLER_34_313 ();
 sg13g2_decap_8 FILLER_34_320 ();
 sg13g2_decap_8 FILLER_34_327 ();
 sg13g2_decap_8 FILLER_34_334 ();
 sg13g2_decap_8 FILLER_34_341 ();
 sg13g2_decap_8 FILLER_34_348 ();
 sg13g2_decap_8 FILLER_34_355 ();
 sg13g2_decap_8 FILLER_34_362 ();
 sg13g2_decap_8 FILLER_34_369 ();
 sg13g2_decap_8 FILLER_34_376 ();
 sg13g2_decap_8 FILLER_34_383 ();
 sg13g2_decap_8 FILLER_34_390 ();
 sg13g2_decap_8 FILLER_34_397 ();
 sg13g2_decap_8 FILLER_34_404 ();
 sg13g2_decap_8 FILLER_34_411 ();
 sg13g2_decap_8 FILLER_34_418 ();
 sg13g2_decap_8 FILLER_34_425 ();
 sg13g2_decap_8 FILLER_34_432 ();
 sg13g2_decap_8 FILLER_34_439 ();
 sg13g2_decap_8 FILLER_34_446 ();
 sg13g2_decap_8 FILLER_34_453 ();
 sg13g2_decap_8 FILLER_34_460 ();
 sg13g2_decap_8 FILLER_34_467 ();
 sg13g2_decap_8 FILLER_34_474 ();
 sg13g2_decap_8 FILLER_34_481 ();
 sg13g2_decap_8 FILLER_34_488 ();
 sg13g2_decap_8 FILLER_34_495 ();
 sg13g2_decap_8 FILLER_34_502 ();
 sg13g2_decap_8 FILLER_34_509 ();
 sg13g2_decap_8 FILLER_34_516 ();
 sg13g2_decap_8 FILLER_34_523 ();
 sg13g2_decap_8 FILLER_34_530 ();
 sg13g2_decap_8 FILLER_34_537 ();
 sg13g2_decap_8 FILLER_34_544 ();
 sg13g2_decap_8 FILLER_34_551 ();
 sg13g2_decap_8 FILLER_34_558 ();
 sg13g2_decap_8 FILLER_34_565 ();
 sg13g2_decap_8 FILLER_34_572 ();
 sg13g2_decap_8 FILLER_34_579 ();
 sg13g2_decap_8 FILLER_34_586 ();
 sg13g2_decap_8 FILLER_34_593 ();
 sg13g2_decap_8 FILLER_34_600 ();
 sg13g2_decap_8 FILLER_34_607 ();
 sg13g2_decap_8 FILLER_34_614 ();
 sg13g2_decap_8 FILLER_34_621 ();
 sg13g2_decap_8 FILLER_34_628 ();
 sg13g2_decap_8 FILLER_34_635 ();
 sg13g2_decap_8 FILLER_34_642 ();
 sg13g2_decap_8 FILLER_34_649 ();
 sg13g2_decap_8 FILLER_34_656 ();
 sg13g2_decap_8 FILLER_34_663 ();
 sg13g2_decap_8 FILLER_34_670 ();
 sg13g2_decap_8 FILLER_34_677 ();
 sg13g2_decap_8 FILLER_34_684 ();
 sg13g2_decap_8 FILLER_34_691 ();
 sg13g2_decap_8 FILLER_34_698 ();
 sg13g2_decap_8 FILLER_34_705 ();
 sg13g2_decap_8 FILLER_34_712 ();
 sg13g2_decap_8 FILLER_34_719 ();
 sg13g2_decap_8 FILLER_34_726 ();
 sg13g2_decap_8 FILLER_34_733 ();
 sg13g2_decap_8 FILLER_34_740 ();
 sg13g2_decap_8 FILLER_34_747 ();
 sg13g2_decap_8 FILLER_34_754 ();
 sg13g2_decap_8 FILLER_34_761 ();
 sg13g2_decap_8 FILLER_34_768 ();
 sg13g2_decap_8 FILLER_34_775 ();
 sg13g2_decap_8 FILLER_34_782 ();
 sg13g2_decap_8 FILLER_34_789 ();
 sg13g2_decap_8 FILLER_34_796 ();
 sg13g2_decap_8 FILLER_34_803 ();
 sg13g2_decap_8 FILLER_34_810 ();
 sg13g2_decap_8 FILLER_34_817 ();
 sg13g2_decap_8 FILLER_34_824 ();
 sg13g2_decap_8 FILLER_34_831 ();
 sg13g2_decap_8 FILLER_34_838 ();
 sg13g2_decap_8 FILLER_34_845 ();
 sg13g2_decap_8 FILLER_34_852 ();
 sg13g2_decap_8 FILLER_34_859 ();
 sg13g2_decap_8 FILLER_34_866 ();
 sg13g2_decap_8 FILLER_34_873 ();
 sg13g2_decap_8 FILLER_34_880 ();
 sg13g2_decap_8 FILLER_34_887 ();
 sg13g2_decap_8 FILLER_34_894 ();
 sg13g2_decap_8 FILLER_34_901 ();
 sg13g2_decap_8 FILLER_34_908 ();
 sg13g2_decap_8 FILLER_34_915 ();
 sg13g2_decap_8 FILLER_34_922 ();
 sg13g2_decap_8 FILLER_34_929 ();
 sg13g2_decap_8 FILLER_34_936 ();
 sg13g2_decap_8 FILLER_34_943 ();
 sg13g2_decap_8 FILLER_34_950 ();
 sg13g2_decap_8 FILLER_34_957 ();
 sg13g2_decap_8 FILLER_34_964 ();
 sg13g2_decap_8 FILLER_34_971 ();
 sg13g2_decap_8 FILLER_34_978 ();
 sg13g2_decap_8 FILLER_34_985 ();
 sg13g2_decap_8 FILLER_34_992 ();
 sg13g2_decap_8 FILLER_34_999 ();
 sg13g2_decap_8 FILLER_34_1006 ();
 sg13g2_decap_8 FILLER_34_1013 ();
 sg13g2_decap_8 FILLER_34_1020 ();
 sg13g2_fill_2 FILLER_34_1027 ();
 sg13g2_decap_8 FILLER_35_4 ();
 sg13g2_decap_8 FILLER_35_11 ();
 sg13g2_decap_8 FILLER_35_18 ();
 sg13g2_decap_8 FILLER_35_25 ();
 sg13g2_decap_8 FILLER_35_32 ();
 sg13g2_decap_8 FILLER_35_39 ();
 sg13g2_decap_8 FILLER_35_46 ();
 sg13g2_decap_8 FILLER_35_53 ();
 sg13g2_decap_8 FILLER_35_60 ();
 sg13g2_decap_8 FILLER_35_67 ();
 sg13g2_decap_8 FILLER_35_74 ();
 sg13g2_decap_8 FILLER_35_81 ();
 sg13g2_decap_8 FILLER_35_88 ();
 sg13g2_decap_8 FILLER_35_95 ();
 sg13g2_decap_8 FILLER_35_102 ();
 sg13g2_decap_8 FILLER_35_109 ();
 sg13g2_decap_8 FILLER_35_116 ();
 sg13g2_decap_8 FILLER_35_123 ();
 sg13g2_decap_8 FILLER_35_130 ();
 sg13g2_decap_8 FILLER_35_137 ();
 sg13g2_decap_8 FILLER_35_144 ();
 sg13g2_decap_8 FILLER_35_151 ();
 sg13g2_decap_8 FILLER_35_158 ();
 sg13g2_decap_8 FILLER_35_165 ();
 sg13g2_decap_8 FILLER_35_172 ();
 sg13g2_decap_8 FILLER_35_179 ();
 sg13g2_decap_8 FILLER_35_186 ();
 sg13g2_decap_8 FILLER_35_193 ();
 sg13g2_decap_8 FILLER_35_200 ();
 sg13g2_decap_8 FILLER_35_207 ();
 sg13g2_decap_8 FILLER_35_214 ();
 sg13g2_decap_8 FILLER_35_221 ();
 sg13g2_decap_8 FILLER_35_228 ();
 sg13g2_decap_8 FILLER_35_235 ();
 sg13g2_decap_8 FILLER_35_242 ();
 sg13g2_decap_8 FILLER_35_249 ();
 sg13g2_decap_8 FILLER_35_256 ();
 sg13g2_decap_8 FILLER_35_263 ();
 sg13g2_decap_8 FILLER_35_270 ();
 sg13g2_decap_8 FILLER_35_277 ();
 sg13g2_decap_8 FILLER_35_284 ();
 sg13g2_decap_8 FILLER_35_291 ();
 sg13g2_decap_8 FILLER_35_298 ();
 sg13g2_decap_8 FILLER_35_305 ();
 sg13g2_decap_8 FILLER_35_312 ();
 sg13g2_decap_8 FILLER_35_319 ();
 sg13g2_decap_8 FILLER_35_326 ();
 sg13g2_decap_8 FILLER_35_333 ();
 sg13g2_decap_8 FILLER_35_340 ();
 sg13g2_decap_8 FILLER_35_347 ();
 sg13g2_decap_8 FILLER_35_354 ();
 sg13g2_decap_8 FILLER_35_361 ();
 sg13g2_decap_8 FILLER_35_368 ();
 sg13g2_decap_8 FILLER_35_375 ();
 sg13g2_decap_8 FILLER_35_382 ();
 sg13g2_decap_8 FILLER_35_389 ();
 sg13g2_decap_8 FILLER_35_396 ();
 sg13g2_decap_8 FILLER_35_403 ();
 sg13g2_decap_8 FILLER_35_410 ();
 sg13g2_decap_8 FILLER_35_417 ();
 sg13g2_decap_8 FILLER_35_424 ();
 sg13g2_decap_8 FILLER_35_431 ();
 sg13g2_decap_8 FILLER_35_438 ();
 sg13g2_decap_8 FILLER_35_445 ();
 sg13g2_decap_8 FILLER_35_452 ();
 sg13g2_decap_8 FILLER_35_459 ();
 sg13g2_decap_8 FILLER_35_466 ();
 sg13g2_decap_8 FILLER_35_473 ();
 sg13g2_decap_8 FILLER_35_480 ();
 sg13g2_decap_8 FILLER_35_487 ();
 sg13g2_decap_8 FILLER_35_494 ();
 sg13g2_decap_8 FILLER_35_501 ();
 sg13g2_decap_8 FILLER_35_508 ();
 sg13g2_decap_8 FILLER_35_515 ();
 sg13g2_decap_8 FILLER_35_522 ();
 sg13g2_decap_8 FILLER_35_529 ();
 sg13g2_decap_8 FILLER_35_536 ();
 sg13g2_decap_8 FILLER_35_543 ();
 sg13g2_decap_8 FILLER_35_550 ();
 sg13g2_decap_8 FILLER_35_557 ();
 sg13g2_decap_8 FILLER_35_564 ();
 sg13g2_decap_8 FILLER_35_571 ();
 sg13g2_decap_8 FILLER_35_578 ();
 sg13g2_decap_8 FILLER_35_585 ();
 sg13g2_decap_8 FILLER_35_592 ();
 sg13g2_decap_8 FILLER_35_599 ();
 sg13g2_decap_8 FILLER_35_606 ();
 sg13g2_decap_8 FILLER_35_613 ();
 sg13g2_decap_8 FILLER_35_620 ();
 sg13g2_decap_8 FILLER_35_627 ();
 sg13g2_decap_8 FILLER_35_634 ();
 sg13g2_decap_8 FILLER_35_641 ();
 sg13g2_decap_8 FILLER_35_648 ();
 sg13g2_decap_8 FILLER_35_655 ();
 sg13g2_decap_8 FILLER_35_662 ();
 sg13g2_decap_8 FILLER_35_669 ();
 sg13g2_decap_8 FILLER_35_676 ();
 sg13g2_decap_8 FILLER_35_683 ();
 sg13g2_decap_8 FILLER_35_690 ();
 sg13g2_decap_8 FILLER_35_697 ();
 sg13g2_decap_8 FILLER_35_704 ();
 sg13g2_decap_8 FILLER_35_711 ();
 sg13g2_decap_8 FILLER_35_718 ();
 sg13g2_decap_8 FILLER_35_725 ();
 sg13g2_decap_8 FILLER_35_732 ();
 sg13g2_decap_8 FILLER_35_739 ();
 sg13g2_decap_8 FILLER_35_746 ();
 sg13g2_decap_8 FILLER_35_753 ();
 sg13g2_decap_8 FILLER_35_760 ();
 sg13g2_decap_8 FILLER_35_767 ();
 sg13g2_decap_8 FILLER_35_774 ();
 sg13g2_decap_8 FILLER_35_781 ();
 sg13g2_decap_8 FILLER_35_788 ();
 sg13g2_decap_8 FILLER_35_795 ();
 sg13g2_decap_8 FILLER_35_802 ();
 sg13g2_decap_8 FILLER_35_809 ();
 sg13g2_decap_8 FILLER_35_816 ();
 sg13g2_decap_8 FILLER_35_823 ();
 sg13g2_decap_8 FILLER_35_830 ();
 sg13g2_decap_8 FILLER_35_837 ();
 sg13g2_decap_8 FILLER_35_844 ();
 sg13g2_decap_8 FILLER_35_851 ();
 sg13g2_decap_8 FILLER_35_858 ();
 sg13g2_decap_8 FILLER_35_865 ();
 sg13g2_decap_8 FILLER_35_872 ();
 sg13g2_decap_8 FILLER_35_879 ();
 sg13g2_decap_8 FILLER_35_886 ();
 sg13g2_decap_8 FILLER_35_893 ();
 sg13g2_decap_8 FILLER_35_900 ();
 sg13g2_decap_8 FILLER_35_907 ();
 sg13g2_decap_8 FILLER_35_914 ();
 sg13g2_decap_8 FILLER_35_921 ();
 sg13g2_decap_8 FILLER_35_928 ();
 sg13g2_decap_8 FILLER_35_935 ();
 sg13g2_decap_8 FILLER_35_942 ();
 sg13g2_decap_8 FILLER_35_949 ();
 sg13g2_decap_8 FILLER_35_956 ();
 sg13g2_decap_8 FILLER_35_963 ();
 sg13g2_decap_8 FILLER_35_970 ();
 sg13g2_decap_8 FILLER_35_977 ();
 sg13g2_decap_8 FILLER_35_984 ();
 sg13g2_decap_8 FILLER_35_991 ();
 sg13g2_decap_8 FILLER_35_998 ();
 sg13g2_decap_8 FILLER_35_1005 ();
 sg13g2_decap_8 FILLER_35_1012 ();
 sg13g2_decap_8 FILLER_35_1019 ();
 sg13g2_fill_2 FILLER_35_1026 ();
 sg13g2_fill_1 FILLER_35_1028 ();
 sg13g2_decap_8 FILLER_36_4 ();
 sg13g2_decap_8 FILLER_36_11 ();
 sg13g2_decap_8 FILLER_36_18 ();
 sg13g2_decap_8 FILLER_36_25 ();
 sg13g2_decap_8 FILLER_36_32 ();
 sg13g2_decap_8 FILLER_36_39 ();
 sg13g2_decap_8 FILLER_36_46 ();
 sg13g2_decap_8 FILLER_36_53 ();
 sg13g2_decap_8 FILLER_36_60 ();
 sg13g2_decap_8 FILLER_36_67 ();
 sg13g2_decap_8 FILLER_36_74 ();
 sg13g2_decap_8 FILLER_36_81 ();
 sg13g2_decap_8 FILLER_36_88 ();
 sg13g2_decap_8 FILLER_36_95 ();
 sg13g2_decap_8 FILLER_36_102 ();
 sg13g2_decap_8 FILLER_36_109 ();
 sg13g2_decap_8 FILLER_36_116 ();
 sg13g2_decap_8 FILLER_36_123 ();
 sg13g2_decap_8 FILLER_36_130 ();
 sg13g2_decap_8 FILLER_36_137 ();
 sg13g2_decap_8 FILLER_36_144 ();
 sg13g2_decap_8 FILLER_36_151 ();
 sg13g2_decap_8 FILLER_36_158 ();
 sg13g2_decap_8 FILLER_36_165 ();
 sg13g2_decap_8 FILLER_36_172 ();
 sg13g2_decap_8 FILLER_36_179 ();
 sg13g2_decap_8 FILLER_36_186 ();
 sg13g2_decap_8 FILLER_36_193 ();
 sg13g2_decap_8 FILLER_36_200 ();
 sg13g2_decap_8 FILLER_36_207 ();
 sg13g2_decap_8 FILLER_36_214 ();
 sg13g2_decap_8 FILLER_36_221 ();
 sg13g2_decap_8 FILLER_36_228 ();
 sg13g2_decap_8 FILLER_36_235 ();
 sg13g2_decap_8 FILLER_36_242 ();
 sg13g2_decap_8 FILLER_36_249 ();
 sg13g2_decap_8 FILLER_36_256 ();
 sg13g2_decap_8 FILLER_36_263 ();
 sg13g2_decap_8 FILLER_36_270 ();
 sg13g2_decap_8 FILLER_36_277 ();
 sg13g2_decap_8 FILLER_36_284 ();
 sg13g2_decap_8 FILLER_36_291 ();
 sg13g2_decap_8 FILLER_36_298 ();
 sg13g2_decap_8 FILLER_36_305 ();
 sg13g2_decap_8 FILLER_36_312 ();
 sg13g2_decap_8 FILLER_36_319 ();
 sg13g2_decap_8 FILLER_36_326 ();
 sg13g2_decap_8 FILLER_36_333 ();
 sg13g2_decap_8 FILLER_36_340 ();
 sg13g2_decap_8 FILLER_36_347 ();
 sg13g2_decap_8 FILLER_36_354 ();
 sg13g2_decap_8 FILLER_36_361 ();
 sg13g2_decap_8 FILLER_36_368 ();
 sg13g2_decap_8 FILLER_36_375 ();
 sg13g2_decap_8 FILLER_36_382 ();
 sg13g2_decap_8 FILLER_36_389 ();
 sg13g2_decap_8 FILLER_36_396 ();
 sg13g2_decap_8 FILLER_36_403 ();
 sg13g2_decap_8 FILLER_36_410 ();
 sg13g2_decap_8 FILLER_36_417 ();
 sg13g2_decap_8 FILLER_36_424 ();
 sg13g2_decap_8 FILLER_36_431 ();
 sg13g2_decap_8 FILLER_36_438 ();
 sg13g2_decap_8 FILLER_36_445 ();
 sg13g2_decap_8 FILLER_36_452 ();
 sg13g2_decap_8 FILLER_36_459 ();
 sg13g2_decap_8 FILLER_36_466 ();
 sg13g2_decap_8 FILLER_36_473 ();
 sg13g2_decap_8 FILLER_36_480 ();
 sg13g2_decap_8 FILLER_36_487 ();
 sg13g2_decap_8 FILLER_36_494 ();
 sg13g2_decap_8 FILLER_36_501 ();
 sg13g2_decap_8 FILLER_36_508 ();
 sg13g2_decap_8 FILLER_36_515 ();
 sg13g2_decap_8 FILLER_36_522 ();
 sg13g2_decap_8 FILLER_36_529 ();
 sg13g2_decap_8 FILLER_36_536 ();
 sg13g2_decap_8 FILLER_36_543 ();
 sg13g2_decap_8 FILLER_36_550 ();
 sg13g2_decap_8 FILLER_36_557 ();
 sg13g2_decap_8 FILLER_36_564 ();
 sg13g2_decap_8 FILLER_36_571 ();
 sg13g2_decap_8 FILLER_36_578 ();
 sg13g2_decap_8 FILLER_36_585 ();
 sg13g2_decap_8 FILLER_36_592 ();
 sg13g2_decap_8 FILLER_36_599 ();
 sg13g2_decap_8 FILLER_36_606 ();
 sg13g2_decap_8 FILLER_36_613 ();
 sg13g2_decap_8 FILLER_36_620 ();
 sg13g2_decap_8 FILLER_36_627 ();
 sg13g2_decap_8 FILLER_36_634 ();
 sg13g2_decap_8 FILLER_36_641 ();
 sg13g2_decap_8 FILLER_36_648 ();
 sg13g2_decap_8 FILLER_36_655 ();
 sg13g2_decap_8 FILLER_36_662 ();
 sg13g2_decap_8 FILLER_36_669 ();
 sg13g2_decap_8 FILLER_36_676 ();
 sg13g2_decap_8 FILLER_36_683 ();
 sg13g2_decap_8 FILLER_36_690 ();
 sg13g2_decap_8 FILLER_36_697 ();
 sg13g2_decap_8 FILLER_36_704 ();
 sg13g2_decap_8 FILLER_36_711 ();
 sg13g2_decap_8 FILLER_36_718 ();
 sg13g2_decap_8 FILLER_36_725 ();
 sg13g2_decap_8 FILLER_36_732 ();
 sg13g2_decap_8 FILLER_36_739 ();
 sg13g2_decap_8 FILLER_36_746 ();
 sg13g2_decap_8 FILLER_36_753 ();
 sg13g2_decap_8 FILLER_36_760 ();
 sg13g2_decap_8 FILLER_36_767 ();
 sg13g2_decap_8 FILLER_36_774 ();
 sg13g2_decap_8 FILLER_36_781 ();
 sg13g2_decap_8 FILLER_36_788 ();
 sg13g2_decap_8 FILLER_36_795 ();
 sg13g2_decap_8 FILLER_36_802 ();
 sg13g2_decap_8 FILLER_36_809 ();
 sg13g2_decap_8 FILLER_36_816 ();
 sg13g2_decap_8 FILLER_36_823 ();
 sg13g2_decap_8 FILLER_36_830 ();
 sg13g2_decap_8 FILLER_36_837 ();
 sg13g2_decap_8 FILLER_36_844 ();
 sg13g2_decap_8 FILLER_36_851 ();
 sg13g2_decap_8 FILLER_36_858 ();
 sg13g2_decap_8 FILLER_36_865 ();
 sg13g2_decap_8 FILLER_36_872 ();
 sg13g2_decap_8 FILLER_36_879 ();
 sg13g2_decap_8 FILLER_36_886 ();
 sg13g2_decap_8 FILLER_36_893 ();
 sg13g2_decap_8 FILLER_36_900 ();
 sg13g2_decap_8 FILLER_36_907 ();
 sg13g2_decap_8 FILLER_36_914 ();
 sg13g2_decap_8 FILLER_36_921 ();
 sg13g2_decap_8 FILLER_36_928 ();
 sg13g2_decap_8 FILLER_36_935 ();
 sg13g2_decap_8 FILLER_36_942 ();
 sg13g2_decap_8 FILLER_36_949 ();
 sg13g2_decap_8 FILLER_36_956 ();
 sg13g2_decap_8 FILLER_36_963 ();
 sg13g2_decap_8 FILLER_36_970 ();
 sg13g2_decap_8 FILLER_36_977 ();
 sg13g2_decap_8 FILLER_36_984 ();
 sg13g2_decap_8 FILLER_36_991 ();
 sg13g2_decap_8 FILLER_36_998 ();
 sg13g2_decap_8 FILLER_36_1005 ();
 sg13g2_decap_8 FILLER_36_1012 ();
 sg13g2_decap_8 FILLER_36_1019 ();
 sg13g2_fill_2 FILLER_36_1026 ();
 sg13g2_fill_1 FILLER_36_1028 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_8 FILLER_37_231 ();
 sg13g2_decap_8 FILLER_37_238 ();
 sg13g2_decap_8 FILLER_37_245 ();
 sg13g2_decap_8 FILLER_37_252 ();
 sg13g2_decap_8 FILLER_37_259 ();
 sg13g2_decap_8 FILLER_37_266 ();
 sg13g2_decap_8 FILLER_37_273 ();
 sg13g2_decap_8 FILLER_37_280 ();
 sg13g2_decap_8 FILLER_37_287 ();
 sg13g2_decap_8 FILLER_37_294 ();
 sg13g2_decap_8 FILLER_37_301 ();
 sg13g2_decap_8 FILLER_37_308 ();
 sg13g2_decap_8 FILLER_37_315 ();
 sg13g2_decap_8 FILLER_37_322 ();
 sg13g2_decap_8 FILLER_37_329 ();
 sg13g2_decap_8 FILLER_37_336 ();
 sg13g2_decap_8 FILLER_37_343 ();
 sg13g2_decap_8 FILLER_37_350 ();
 sg13g2_decap_8 FILLER_37_357 ();
 sg13g2_decap_8 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_371 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_decap_8 FILLER_37_406 ();
 sg13g2_decap_8 FILLER_37_413 ();
 sg13g2_decap_8 FILLER_37_420 ();
 sg13g2_decap_8 FILLER_37_427 ();
 sg13g2_decap_8 FILLER_37_434 ();
 sg13g2_decap_8 FILLER_37_441 ();
 sg13g2_decap_8 FILLER_37_448 ();
 sg13g2_decap_8 FILLER_37_455 ();
 sg13g2_decap_8 FILLER_37_462 ();
 sg13g2_decap_8 FILLER_37_469 ();
 sg13g2_decap_8 FILLER_37_476 ();
 sg13g2_decap_8 FILLER_37_483 ();
 sg13g2_decap_8 FILLER_37_490 ();
 sg13g2_decap_8 FILLER_37_497 ();
 sg13g2_decap_8 FILLER_37_504 ();
 sg13g2_decap_8 FILLER_37_511 ();
 sg13g2_decap_8 FILLER_37_518 ();
 sg13g2_decap_8 FILLER_37_525 ();
 sg13g2_decap_8 FILLER_37_532 ();
 sg13g2_decap_8 FILLER_37_539 ();
 sg13g2_decap_8 FILLER_37_546 ();
 sg13g2_decap_8 FILLER_37_553 ();
 sg13g2_decap_8 FILLER_37_560 ();
 sg13g2_decap_8 FILLER_37_567 ();
 sg13g2_decap_8 FILLER_37_574 ();
 sg13g2_decap_8 FILLER_37_581 ();
 sg13g2_decap_8 FILLER_37_588 ();
 sg13g2_decap_8 FILLER_37_595 ();
 sg13g2_decap_8 FILLER_37_602 ();
 sg13g2_decap_8 FILLER_37_609 ();
 sg13g2_decap_8 FILLER_37_616 ();
 sg13g2_decap_8 FILLER_37_623 ();
 sg13g2_decap_8 FILLER_37_630 ();
 sg13g2_decap_8 FILLER_37_637 ();
 sg13g2_decap_8 FILLER_37_644 ();
 sg13g2_decap_8 FILLER_37_651 ();
 sg13g2_decap_8 FILLER_37_658 ();
 sg13g2_decap_8 FILLER_37_665 ();
 sg13g2_decap_8 FILLER_37_672 ();
 sg13g2_decap_8 FILLER_37_679 ();
 sg13g2_decap_8 FILLER_37_686 ();
 sg13g2_decap_8 FILLER_37_693 ();
 sg13g2_decap_8 FILLER_37_700 ();
 sg13g2_decap_8 FILLER_37_707 ();
 sg13g2_decap_8 FILLER_37_714 ();
 sg13g2_decap_8 FILLER_37_721 ();
 sg13g2_decap_8 FILLER_37_728 ();
 sg13g2_decap_8 FILLER_37_735 ();
 sg13g2_decap_8 FILLER_37_742 ();
 sg13g2_decap_8 FILLER_37_749 ();
 sg13g2_decap_8 FILLER_37_756 ();
 sg13g2_decap_8 FILLER_37_763 ();
 sg13g2_decap_8 FILLER_37_770 ();
 sg13g2_decap_8 FILLER_37_777 ();
 sg13g2_decap_8 FILLER_37_784 ();
 sg13g2_decap_8 FILLER_37_791 ();
 sg13g2_decap_8 FILLER_37_798 ();
 sg13g2_decap_8 FILLER_37_805 ();
 sg13g2_decap_8 FILLER_37_812 ();
 sg13g2_decap_8 FILLER_37_819 ();
 sg13g2_decap_8 FILLER_37_826 ();
 sg13g2_decap_8 FILLER_37_833 ();
 sg13g2_decap_8 FILLER_37_840 ();
 sg13g2_decap_8 FILLER_37_847 ();
 sg13g2_decap_8 FILLER_37_854 ();
 sg13g2_decap_8 FILLER_37_861 ();
 sg13g2_decap_8 FILLER_37_868 ();
 sg13g2_decap_8 FILLER_37_875 ();
 sg13g2_decap_8 FILLER_37_882 ();
 sg13g2_decap_8 FILLER_37_889 ();
 sg13g2_decap_8 FILLER_37_896 ();
 sg13g2_decap_8 FILLER_37_903 ();
 sg13g2_decap_8 FILLER_37_910 ();
 sg13g2_decap_8 FILLER_37_917 ();
 sg13g2_decap_8 FILLER_37_924 ();
 sg13g2_decap_8 FILLER_37_931 ();
 sg13g2_decap_8 FILLER_37_938 ();
 sg13g2_decap_8 FILLER_37_945 ();
 sg13g2_decap_8 FILLER_37_952 ();
 sg13g2_decap_8 FILLER_37_959 ();
 sg13g2_decap_8 FILLER_37_966 ();
 sg13g2_decap_8 FILLER_37_973 ();
 sg13g2_decap_8 FILLER_37_980 ();
 sg13g2_decap_8 FILLER_37_987 ();
 sg13g2_decap_8 FILLER_37_994 ();
 sg13g2_decap_8 FILLER_37_1001 ();
 sg13g2_decap_8 FILLER_37_1008 ();
 sg13g2_decap_8 FILLER_37_1015 ();
 sg13g2_decap_8 FILLER_37_1022 ();
 sg13g2_decap_8 FILLER_38_4 ();
 sg13g2_decap_8 FILLER_38_11 ();
 sg13g2_decap_8 FILLER_38_18 ();
 sg13g2_decap_8 FILLER_38_25 ();
 sg13g2_decap_8 FILLER_38_32 ();
 sg13g2_decap_8 FILLER_38_39 ();
 sg13g2_decap_8 FILLER_38_46 ();
 sg13g2_decap_8 FILLER_38_53 ();
 sg13g2_decap_8 FILLER_38_60 ();
 sg13g2_decap_8 FILLER_38_67 ();
 sg13g2_decap_8 FILLER_38_74 ();
 sg13g2_decap_8 FILLER_38_81 ();
 sg13g2_decap_8 FILLER_38_88 ();
 sg13g2_decap_8 FILLER_38_95 ();
 sg13g2_decap_8 FILLER_38_102 ();
 sg13g2_decap_8 FILLER_38_109 ();
 sg13g2_decap_8 FILLER_38_116 ();
 sg13g2_decap_8 FILLER_38_123 ();
 sg13g2_decap_8 FILLER_38_130 ();
 sg13g2_decap_8 FILLER_38_137 ();
 sg13g2_decap_8 FILLER_38_144 ();
 sg13g2_decap_8 FILLER_38_151 ();
 sg13g2_decap_8 FILLER_38_158 ();
 sg13g2_decap_8 FILLER_38_165 ();
 sg13g2_decap_8 FILLER_38_172 ();
 sg13g2_decap_8 FILLER_38_179 ();
 sg13g2_decap_8 FILLER_38_186 ();
 sg13g2_decap_8 FILLER_38_193 ();
 sg13g2_decap_8 FILLER_38_200 ();
 sg13g2_decap_8 FILLER_38_207 ();
 sg13g2_decap_8 FILLER_38_214 ();
 sg13g2_decap_8 FILLER_38_221 ();
 sg13g2_decap_8 FILLER_38_228 ();
 sg13g2_decap_8 FILLER_38_235 ();
 sg13g2_decap_8 FILLER_38_242 ();
 sg13g2_decap_8 FILLER_38_249 ();
 sg13g2_decap_8 FILLER_38_256 ();
 sg13g2_decap_8 FILLER_38_263 ();
 sg13g2_decap_8 FILLER_38_270 ();
 sg13g2_decap_8 FILLER_38_277 ();
 sg13g2_decap_8 FILLER_38_284 ();
 sg13g2_decap_8 FILLER_38_291 ();
 sg13g2_decap_8 FILLER_38_298 ();
 sg13g2_decap_8 FILLER_38_305 ();
 sg13g2_decap_8 FILLER_38_312 ();
 sg13g2_decap_8 FILLER_38_319 ();
 sg13g2_decap_8 FILLER_38_326 ();
 sg13g2_decap_8 FILLER_38_333 ();
 sg13g2_decap_8 FILLER_38_340 ();
 sg13g2_decap_8 FILLER_38_347 ();
 sg13g2_decap_8 FILLER_38_354 ();
 sg13g2_decap_8 FILLER_38_361 ();
 sg13g2_decap_8 FILLER_38_368 ();
 sg13g2_decap_8 FILLER_38_375 ();
 sg13g2_decap_8 FILLER_38_382 ();
 sg13g2_decap_8 FILLER_38_389 ();
 sg13g2_decap_8 FILLER_38_396 ();
 sg13g2_decap_8 FILLER_38_403 ();
 sg13g2_decap_8 FILLER_38_410 ();
 sg13g2_decap_8 FILLER_38_417 ();
 sg13g2_decap_8 FILLER_38_424 ();
 sg13g2_decap_8 FILLER_38_431 ();
 sg13g2_decap_8 FILLER_38_438 ();
 sg13g2_decap_8 FILLER_38_445 ();
 sg13g2_decap_8 FILLER_38_452 ();
 sg13g2_decap_8 FILLER_38_459 ();
 sg13g2_decap_8 FILLER_38_466 ();
 sg13g2_decap_8 FILLER_38_473 ();
 sg13g2_decap_8 FILLER_38_480 ();
 sg13g2_decap_8 FILLER_38_487 ();
 sg13g2_decap_8 FILLER_38_494 ();
 sg13g2_decap_8 FILLER_38_501 ();
 sg13g2_decap_8 FILLER_38_508 ();
 sg13g2_decap_8 FILLER_38_515 ();
 sg13g2_decap_8 FILLER_38_522 ();
 sg13g2_decap_8 FILLER_38_529 ();
 sg13g2_decap_8 FILLER_38_536 ();
 sg13g2_decap_8 FILLER_38_543 ();
 sg13g2_decap_8 FILLER_38_550 ();
 sg13g2_decap_8 FILLER_38_557 ();
 sg13g2_decap_8 FILLER_38_564 ();
 sg13g2_decap_8 FILLER_38_571 ();
 sg13g2_decap_8 FILLER_38_578 ();
 sg13g2_decap_8 FILLER_38_585 ();
 sg13g2_decap_8 FILLER_38_592 ();
 sg13g2_decap_8 FILLER_38_599 ();
 sg13g2_decap_8 FILLER_38_606 ();
 sg13g2_decap_8 FILLER_38_613 ();
 sg13g2_decap_8 FILLER_38_620 ();
 sg13g2_decap_8 FILLER_38_627 ();
 sg13g2_decap_8 FILLER_38_634 ();
 sg13g2_decap_8 FILLER_38_641 ();
 sg13g2_decap_8 FILLER_38_648 ();
 sg13g2_decap_8 FILLER_38_655 ();
 sg13g2_decap_8 FILLER_38_662 ();
 sg13g2_decap_8 FILLER_38_669 ();
 sg13g2_decap_8 FILLER_38_676 ();
 sg13g2_decap_8 FILLER_38_683 ();
 sg13g2_decap_8 FILLER_38_690 ();
 sg13g2_decap_8 FILLER_38_697 ();
 sg13g2_decap_8 FILLER_38_704 ();
 sg13g2_decap_8 FILLER_38_711 ();
 sg13g2_decap_8 FILLER_38_718 ();
 sg13g2_decap_8 FILLER_38_725 ();
 sg13g2_decap_8 FILLER_38_732 ();
 sg13g2_decap_8 FILLER_38_739 ();
 sg13g2_decap_8 FILLER_38_746 ();
 sg13g2_decap_8 FILLER_38_753 ();
 sg13g2_decap_8 FILLER_38_760 ();
 sg13g2_decap_8 FILLER_38_767 ();
 sg13g2_decap_8 FILLER_38_774 ();
 sg13g2_decap_8 FILLER_38_781 ();
 sg13g2_decap_8 FILLER_38_788 ();
 sg13g2_decap_8 FILLER_38_795 ();
 sg13g2_decap_8 FILLER_38_802 ();
 sg13g2_decap_8 FILLER_38_809 ();
 sg13g2_decap_8 FILLER_38_816 ();
 sg13g2_decap_8 FILLER_38_823 ();
 sg13g2_decap_8 FILLER_38_830 ();
 sg13g2_decap_8 FILLER_38_837 ();
 sg13g2_decap_8 FILLER_38_844 ();
 sg13g2_decap_8 FILLER_38_851 ();
 sg13g2_decap_8 FILLER_38_858 ();
 sg13g2_decap_8 FILLER_38_865 ();
 sg13g2_decap_8 FILLER_38_872 ();
 sg13g2_decap_8 FILLER_38_879 ();
 sg13g2_decap_8 FILLER_38_886 ();
 sg13g2_decap_8 FILLER_38_893 ();
 sg13g2_decap_8 FILLER_38_900 ();
 sg13g2_decap_8 FILLER_38_907 ();
 sg13g2_decap_8 FILLER_38_914 ();
 sg13g2_decap_8 FILLER_38_921 ();
 sg13g2_decap_8 FILLER_38_928 ();
 sg13g2_decap_8 FILLER_38_935 ();
 sg13g2_decap_8 FILLER_38_942 ();
 sg13g2_decap_8 FILLER_38_949 ();
 sg13g2_decap_8 FILLER_38_956 ();
 sg13g2_decap_8 FILLER_38_963 ();
 sg13g2_decap_8 FILLER_38_970 ();
 sg13g2_decap_8 FILLER_38_977 ();
 sg13g2_decap_8 FILLER_38_984 ();
 sg13g2_decap_8 FILLER_38_991 ();
 sg13g2_decap_8 FILLER_38_998 ();
 sg13g2_decap_8 FILLER_38_1005 ();
 sg13g2_decap_8 FILLER_38_1012 ();
 sg13g2_decap_8 FILLER_38_1019 ();
 sg13g2_fill_2 FILLER_38_1026 ();
 sg13g2_fill_1 FILLER_38_1028 ();
 sg13g2_decap_8 FILLER_39_4 ();
 sg13g2_decap_8 FILLER_39_11 ();
 sg13g2_decap_8 FILLER_39_18 ();
 sg13g2_decap_8 FILLER_39_25 ();
 sg13g2_decap_8 FILLER_39_32 ();
 sg13g2_decap_8 FILLER_39_39 ();
 sg13g2_decap_8 FILLER_39_46 ();
 sg13g2_decap_8 FILLER_39_53 ();
 sg13g2_decap_8 FILLER_39_60 ();
 sg13g2_fill_2 FILLER_39_67 ();
 sg13g2_fill_1 FILLER_39_69 ();
 sg13g2_decap_8 FILLER_39_78 ();
 sg13g2_decap_8 FILLER_39_85 ();
 sg13g2_decap_8 FILLER_39_92 ();
 sg13g2_decap_8 FILLER_39_99 ();
 sg13g2_decap_8 FILLER_39_106 ();
 sg13g2_decap_8 FILLER_39_113 ();
 sg13g2_decap_8 FILLER_39_120 ();
 sg13g2_decap_8 FILLER_39_127 ();
 sg13g2_decap_8 FILLER_39_134 ();
 sg13g2_decap_8 FILLER_39_141 ();
 sg13g2_decap_8 FILLER_39_148 ();
 sg13g2_decap_8 FILLER_39_155 ();
 sg13g2_decap_8 FILLER_39_162 ();
 sg13g2_decap_8 FILLER_39_169 ();
 sg13g2_decap_8 FILLER_39_176 ();
 sg13g2_decap_8 FILLER_39_183 ();
 sg13g2_decap_8 FILLER_39_190 ();
 sg13g2_decap_8 FILLER_39_197 ();
 sg13g2_decap_8 FILLER_39_204 ();
 sg13g2_decap_8 FILLER_39_211 ();
 sg13g2_decap_8 FILLER_39_218 ();
 sg13g2_decap_8 FILLER_39_225 ();
 sg13g2_decap_8 FILLER_39_232 ();
 sg13g2_decap_8 FILLER_39_239 ();
 sg13g2_decap_8 FILLER_39_246 ();
 sg13g2_decap_8 FILLER_39_253 ();
 sg13g2_decap_8 FILLER_39_260 ();
 sg13g2_decap_8 FILLER_39_267 ();
 sg13g2_decap_8 FILLER_39_274 ();
 sg13g2_decap_8 FILLER_39_281 ();
 sg13g2_decap_8 FILLER_39_288 ();
 sg13g2_decap_8 FILLER_39_295 ();
 sg13g2_decap_8 FILLER_39_302 ();
 sg13g2_decap_8 FILLER_39_309 ();
 sg13g2_decap_8 FILLER_39_316 ();
 sg13g2_decap_8 FILLER_39_323 ();
 sg13g2_decap_8 FILLER_39_330 ();
 sg13g2_decap_8 FILLER_39_337 ();
 sg13g2_decap_8 FILLER_39_344 ();
 sg13g2_decap_8 FILLER_39_351 ();
 sg13g2_decap_8 FILLER_39_358 ();
 sg13g2_decap_8 FILLER_39_365 ();
 sg13g2_decap_8 FILLER_39_372 ();
 sg13g2_decap_8 FILLER_39_379 ();
 sg13g2_decap_8 FILLER_39_386 ();
 sg13g2_decap_8 FILLER_39_393 ();
 sg13g2_decap_8 FILLER_39_400 ();
 sg13g2_decap_8 FILLER_39_407 ();
 sg13g2_decap_8 FILLER_39_414 ();
 sg13g2_decap_8 FILLER_39_421 ();
 sg13g2_decap_8 FILLER_39_428 ();
 sg13g2_decap_8 FILLER_39_435 ();
 sg13g2_decap_8 FILLER_39_442 ();
 sg13g2_decap_8 FILLER_39_449 ();
 sg13g2_decap_8 FILLER_39_456 ();
 sg13g2_decap_8 FILLER_39_463 ();
 sg13g2_decap_8 FILLER_39_470 ();
 sg13g2_decap_8 FILLER_39_477 ();
 sg13g2_decap_8 FILLER_39_484 ();
 sg13g2_decap_8 FILLER_39_491 ();
 sg13g2_decap_8 FILLER_39_498 ();
 sg13g2_decap_8 FILLER_39_505 ();
 sg13g2_decap_8 FILLER_39_512 ();
 sg13g2_decap_8 FILLER_39_519 ();
 sg13g2_decap_8 FILLER_39_526 ();
 sg13g2_decap_8 FILLER_39_533 ();
 sg13g2_decap_8 FILLER_39_540 ();
 sg13g2_decap_8 FILLER_39_547 ();
 sg13g2_decap_8 FILLER_39_554 ();
 sg13g2_decap_8 FILLER_39_561 ();
 sg13g2_decap_8 FILLER_39_568 ();
 sg13g2_decap_8 FILLER_39_575 ();
 sg13g2_decap_8 FILLER_39_582 ();
 sg13g2_decap_8 FILLER_39_589 ();
 sg13g2_decap_8 FILLER_39_596 ();
 sg13g2_decap_8 FILLER_39_603 ();
 sg13g2_decap_8 FILLER_39_610 ();
 sg13g2_decap_8 FILLER_39_617 ();
 sg13g2_decap_8 FILLER_39_624 ();
 sg13g2_decap_8 FILLER_39_631 ();
 sg13g2_decap_8 FILLER_39_638 ();
 sg13g2_decap_8 FILLER_39_645 ();
 sg13g2_decap_8 FILLER_39_652 ();
 sg13g2_decap_8 FILLER_39_659 ();
 sg13g2_decap_8 FILLER_39_666 ();
 sg13g2_decap_8 FILLER_39_673 ();
 sg13g2_decap_8 FILLER_39_680 ();
 sg13g2_decap_8 FILLER_39_687 ();
 sg13g2_decap_8 FILLER_39_694 ();
 sg13g2_decap_8 FILLER_39_701 ();
 sg13g2_decap_8 FILLER_39_708 ();
 sg13g2_decap_8 FILLER_39_715 ();
 sg13g2_decap_8 FILLER_39_722 ();
 sg13g2_decap_8 FILLER_39_729 ();
 sg13g2_decap_8 FILLER_39_736 ();
 sg13g2_decap_8 FILLER_39_743 ();
 sg13g2_decap_8 FILLER_39_750 ();
 sg13g2_decap_8 FILLER_39_757 ();
 sg13g2_decap_8 FILLER_39_764 ();
 sg13g2_decap_8 FILLER_39_771 ();
 sg13g2_decap_8 FILLER_39_778 ();
 sg13g2_decap_8 FILLER_39_785 ();
 sg13g2_decap_8 FILLER_39_792 ();
 sg13g2_decap_8 FILLER_39_799 ();
 sg13g2_decap_8 FILLER_39_806 ();
 sg13g2_decap_8 FILLER_39_813 ();
 sg13g2_decap_8 FILLER_39_820 ();
 sg13g2_decap_8 FILLER_39_827 ();
 sg13g2_decap_8 FILLER_39_834 ();
 sg13g2_decap_8 FILLER_39_841 ();
 sg13g2_decap_8 FILLER_39_848 ();
 sg13g2_decap_8 FILLER_39_855 ();
 sg13g2_decap_8 FILLER_39_862 ();
 sg13g2_decap_8 FILLER_39_869 ();
 sg13g2_decap_8 FILLER_39_876 ();
 sg13g2_decap_8 FILLER_39_883 ();
 sg13g2_decap_8 FILLER_39_890 ();
 sg13g2_decap_8 FILLER_39_897 ();
 sg13g2_decap_8 FILLER_39_904 ();
 sg13g2_decap_8 FILLER_39_911 ();
 sg13g2_decap_8 FILLER_39_918 ();
 sg13g2_decap_8 FILLER_39_925 ();
 sg13g2_decap_8 FILLER_39_932 ();
 sg13g2_decap_8 FILLER_39_939 ();
 sg13g2_decap_8 FILLER_39_946 ();
 sg13g2_decap_8 FILLER_39_953 ();
 sg13g2_decap_8 FILLER_39_960 ();
 sg13g2_decap_8 FILLER_39_967 ();
 sg13g2_decap_8 FILLER_39_974 ();
 sg13g2_decap_8 FILLER_39_981 ();
 sg13g2_decap_8 FILLER_39_988 ();
 sg13g2_decap_8 FILLER_39_995 ();
 sg13g2_decap_8 FILLER_39_1002 ();
 sg13g2_decap_8 FILLER_39_1009 ();
 sg13g2_decap_8 FILLER_39_1016 ();
 sg13g2_decap_4 FILLER_39_1023 ();
 sg13g2_fill_2 FILLER_39_1027 ();
 sg13g2_decap_8 FILLER_40_4 ();
 sg13g2_decap_8 FILLER_40_11 ();
 sg13g2_decap_8 FILLER_40_18 ();
 sg13g2_decap_8 FILLER_40_25 ();
 sg13g2_decap_8 FILLER_40_32 ();
 sg13g2_decap_8 FILLER_40_39 ();
 sg13g2_decap_8 FILLER_40_46 ();
 sg13g2_decap_8 FILLER_40_53 ();
 sg13g2_decap_4 FILLER_40_60 ();
 sg13g2_fill_1 FILLER_40_76 ();
 sg13g2_fill_2 FILLER_40_82 ();
 sg13g2_decap_8 FILLER_40_100 ();
 sg13g2_decap_8 FILLER_40_107 ();
 sg13g2_decap_8 FILLER_40_114 ();
 sg13g2_decap_8 FILLER_40_121 ();
 sg13g2_decap_8 FILLER_40_128 ();
 sg13g2_decap_8 FILLER_40_135 ();
 sg13g2_decap_8 FILLER_40_142 ();
 sg13g2_decap_8 FILLER_40_149 ();
 sg13g2_decap_8 FILLER_40_156 ();
 sg13g2_decap_8 FILLER_40_163 ();
 sg13g2_decap_8 FILLER_40_170 ();
 sg13g2_decap_8 FILLER_40_177 ();
 sg13g2_decap_8 FILLER_40_184 ();
 sg13g2_decap_8 FILLER_40_191 ();
 sg13g2_decap_8 FILLER_40_198 ();
 sg13g2_decap_8 FILLER_40_205 ();
 sg13g2_decap_8 FILLER_40_212 ();
 sg13g2_decap_8 FILLER_40_219 ();
 sg13g2_decap_8 FILLER_40_226 ();
 sg13g2_decap_8 FILLER_40_233 ();
 sg13g2_decap_8 FILLER_40_240 ();
 sg13g2_decap_8 FILLER_40_247 ();
 sg13g2_decap_8 FILLER_40_254 ();
 sg13g2_decap_8 FILLER_40_261 ();
 sg13g2_decap_8 FILLER_40_268 ();
 sg13g2_decap_8 FILLER_40_275 ();
 sg13g2_decap_8 FILLER_40_282 ();
 sg13g2_decap_8 FILLER_40_289 ();
 sg13g2_decap_8 FILLER_40_296 ();
 sg13g2_decap_8 FILLER_40_303 ();
 sg13g2_decap_8 FILLER_40_310 ();
 sg13g2_decap_8 FILLER_40_317 ();
 sg13g2_decap_8 FILLER_40_324 ();
 sg13g2_decap_8 FILLER_40_331 ();
 sg13g2_decap_8 FILLER_40_338 ();
 sg13g2_decap_8 FILLER_40_345 ();
 sg13g2_decap_8 FILLER_40_352 ();
 sg13g2_decap_8 FILLER_40_359 ();
 sg13g2_decap_8 FILLER_40_366 ();
 sg13g2_decap_8 FILLER_40_373 ();
 sg13g2_decap_8 FILLER_40_380 ();
 sg13g2_decap_8 FILLER_40_387 ();
 sg13g2_decap_8 FILLER_40_394 ();
 sg13g2_decap_8 FILLER_40_401 ();
 sg13g2_decap_8 FILLER_40_408 ();
 sg13g2_decap_8 FILLER_40_415 ();
 sg13g2_decap_8 FILLER_40_422 ();
 sg13g2_decap_8 FILLER_40_429 ();
 sg13g2_decap_8 FILLER_40_436 ();
 sg13g2_decap_8 FILLER_40_443 ();
 sg13g2_decap_8 FILLER_40_450 ();
 sg13g2_decap_8 FILLER_40_457 ();
 sg13g2_decap_8 FILLER_40_464 ();
 sg13g2_decap_8 FILLER_40_471 ();
 sg13g2_decap_8 FILLER_40_478 ();
 sg13g2_decap_8 FILLER_40_485 ();
 sg13g2_decap_8 FILLER_40_492 ();
 sg13g2_decap_8 FILLER_40_499 ();
 sg13g2_decap_8 FILLER_40_506 ();
 sg13g2_decap_8 FILLER_40_513 ();
 sg13g2_decap_8 FILLER_40_520 ();
 sg13g2_decap_8 FILLER_40_527 ();
 sg13g2_decap_8 FILLER_40_534 ();
 sg13g2_decap_8 FILLER_40_541 ();
 sg13g2_decap_8 FILLER_40_548 ();
 sg13g2_decap_8 FILLER_40_555 ();
 sg13g2_decap_8 FILLER_40_562 ();
 sg13g2_decap_8 FILLER_40_569 ();
 sg13g2_decap_8 FILLER_40_576 ();
 sg13g2_decap_8 FILLER_40_583 ();
 sg13g2_decap_8 FILLER_40_590 ();
 sg13g2_decap_8 FILLER_40_597 ();
 sg13g2_decap_8 FILLER_40_604 ();
 sg13g2_decap_8 FILLER_40_611 ();
 sg13g2_decap_8 FILLER_40_618 ();
 sg13g2_decap_8 FILLER_40_625 ();
 sg13g2_decap_8 FILLER_40_632 ();
 sg13g2_decap_8 FILLER_40_639 ();
 sg13g2_decap_8 FILLER_40_646 ();
 sg13g2_decap_8 FILLER_40_653 ();
 sg13g2_decap_8 FILLER_40_660 ();
 sg13g2_decap_8 FILLER_40_667 ();
 sg13g2_decap_8 FILLER_40_674 ();
 sg13g2_decap_8 FILLER_40_681 ();
 sg13g2_decap_8 FILLER_40_688 ();
 sg13g2_decap_8 FILLER_40_695 ();
 sg13g2_decap_8 FILLER_40_702 ();
 sg13g2_decap_8 FILLER_40_709 ();
 sg13g2_decap_8 FILLER_40_716 ();
 sg13g2_decap_8 FILLER_40_723 ();
 sg13g2_decap_8 FILLER_40_730 ();
 sg13g2_decap_8 FILLER_40_737 ();
 sg13g2_decap_8 FILLER_40_744 ();
 sg13g2_decap_8 FILLER_40_751 ();
 sg13g2_decap_8 FILLER_40_758 ();
 sg13g2_decap_8 FILLER_40_765 ();
 sg13g2_decap_8 FILLER_40_772 ();
 sg13g2_decap_8 FILLER_40_779 ();
 sg13g2_decap_8 FILLER_40_786 ();
 sg13g2_decap_8 FILLER_40_793 ();
 sg13g2_decap_8 FILLER_40_800 ();
 sg13g2_decap_8 FILLER_40_807 ();
 sg13g2_decap_8 FILLER_40_814 ();
 sg13g2_decap_8 FILLER_40_821 ();
 sg13g2_decap_8 FILLER_40_828 ();
 sg13g2_decap_8 FILLER_40_835 ();
 sg13g2_decap_8 FILLER_40_842 ();
 sg13g2_decap_8 FILLER_40_849 ();
 sg13g2_decap_8 FILLER_40_856 ();
 sg13g2_decap_8 FILLER_40_863 ();
 sg13g2_decap_8 FILLER_40_870 ();
 sg13g2_decap_8 FILLER_40_877 ();
 sg13g2_decap_8 FILLER_40_884 ();
 sg13g2_decap_8 FILLER_40_891 ();
 sg13g2_decap_8 FILLER_40_898 ();
 sg13g2_decap_8 FILLER_40_905 ();
 sg13g2_decap_8 FILLER_40_912 ();
 sg13g2_decap_8 FILLER_40_919 ();
 sg13g2_decap_8 FILLER_40_926 ();
 sg13g2_decap_8 FILLER_40_933 ();
 sg13g2_decap_8 FILLER_40_940 ();
 sg13g2_decap_8 FILLER_40_947 ();
 sg13g2_decap_8 FILLER_40_954 ();
 sg13g2_decap_8 FILLER_40_961 ();
 sg13g2_decap_8 FILLER_40_968 ();
 sg13g2_decap_8 FILLER_40_975 ();
 sg13g2_decap_8 FILLER_40_982 ();
 sg13g2_decap_8 FILLER_40_989 ();
 sg13g2_decap_8 FILLER_40_996 ();
 sg13g2_decap_8 FILLER_40_1003 ();
 sg13g2_decap_8 FILLER_40_1010 ();
 sg13g2_decap_8 FILLER_40_1017 ();
 sg13g2_decap_4 FILLER_40_1024 ();
 sg13g2_fill_1 FILLER_40_1028 ();
 sg13g2_decap_8 FILLER_41_4 ();
 sg13g2_decap_8 FILLER_41_11 ();
 sg13g2_decap_8 FILLER_41_18 ();
 sg13g2_decap_8 FILLER_41_25 ();
 sg13g2_decap_8 FILLER_41_32 ();
 sg13g2_decap_8 FILLER_41_39 ();
 sg13g2_decap_8 FILLER_41_46 ();
 sg13g2_decap_8 FILLER_41_53 ();
 sg13g2_decap_8 FILLER_41_60 ();
 sg13g2_decap_4 FILLER_41_67 ();
 sg13g2_fill_2 FILLER_41_71 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_decap_8 FILLER_41_133 ();
 sg13g2_decap_8 FILLER_41_140 ();
 sg13g2_decap_8 FILLER_41_147 ();
 sg13g2_decap_8 FILLER_41_154 ();
 sg13g2_decap_8 FILLER_41_161 ();
 sg13g2_decap_8 FILLER_41_168 ();
 sg13g2_decap_8 FILLER_41_175 ();
 sg13g2_decap_8 FILLER_41_182 ();
 sg13g2_decap_8 FILLER_41_189 ();
 sg13g2_decap_8 FILLER_41_196 ();
 sg13g2_decap_8 FILLER_41_203 ();
 sg13g2_decap_8 FILLER_41_210 ();
 sg13g2_decap_8 FILLER_41_217 ();
 sg13g2_decap_8 FILLER_41_224 ();
 sg13g2_decap_8 FILLER_41_231 ();
 sg13g2_decap_8 FILLER_41_238 ();
 sg13g2_decap_8 FILLER_41_245 ();
 sg13g2_decap_8 FILLER_41_252 ();
 sg13g2_decap_8 FILLER_41_259 ();
 sg13g2_decap_8 FILLER_41_266 ();
 sg13g2_decap_8 FILLER_41_273 ();
 sg13g2_decap_8 FILLER_41_280 ();
 sg13g2_decap_8 FILLER_41_287 ();
 sg13g2_decap_8 FILLER_41_294 ();
 sg13g2_decap_8 FILLER_41_301 ();
 sg13g2_decap_8 FILLER_41_308 ();
 sg13g2_decap_8 FILLER_41_315 ();
 sg13g2_decap_8 FILLER_41_322 ();
 sg13g2_decap_8 FILLER_41_329 ();
 sg13g2_decap_8 FILLER_41_336 ();
 sg13g2_decap_8 FILLER_41_343 ();
 sg13g2_decap_8 FILLER_41_350 ();
 sg13g2_decap_8 FILLER_41_357 ();
 sg13g2_decap_8 FILLER_41_364 ();
 sg13g2_decap_8 FILLER_41_371 ();
 sg13g2_decap_8 FILLER_41_378 ();
 sg13g2_decap_8 FILLER_41_385 ();
 sg13g2_decap_8 FILLER_41_392 ();
 sg13g2_decap_8 FILLER_41_399 ();
 sg13g2_decap_8 FILLER_41_406 ();
 sg13g2_decap_8 FILLER_41_413 ();
 sg13g2_decap_8 FILLER_41_420 ();
 sg13g2_decap_8 FILLER_41_427 ();
 sg13g2_decap_8 FILLER_41_434 ();
 sg13g2_decap_8 FILLER_41_441 ();
 sg13g2_decap_8 FILLER_41_448 ();
 sg13g2_decap_8 FILLER_41_455 ();
 sg13g2_decap_8 FILLER_41_462 ();
 sg13g2_decap_8 FILLER_41_469 ();
 sg13g2_decap_8 FILLER_41_476 ();
 sg13g2_decap_8 FILLER_41_483 ();
 sg13g2_decap_8 FILLER_41_490 ();
 sg13g2_decap_8 FILLER_41_497 ();
 sg13g2_decap_8 FILLER_41_504 ();
 sg13g2_decap_8 FILLER_41_511 ();
 sg13g2_decap_8 FILLER_41_518 ();
 sg13g2_decap_8 FILLER_41_525 ();
 sg13g2_decap_8 FILLER_41_532 ();
 sg13g2_decap_8 FILLER_41_539 ();
 sg13g2_decap_8 FILLER_41_546 ();
 sg13g2_decap_8 FILLER_41_553 ();
 sg13g2_decap_8 FILLER_41_560 ();
 sg13g2_decap_8 FILLER_41_567 ();
 sg13g2_decap_8 FILLER_41_574 ();
 sg13g2_decap_8 FILLER_41_581 ();
 sg13g2_decap_8 FILLER_41_588 ();
 sg13g2_decap_8 FILLER_41_595 ();
 sg13g2_decap_8 FILLER_41_602 ();
 sg13g2_decap_8 FILLER_41_609 ();
 sg13g2_decap_8 FILLER_41_616 ();
 sg13g2_decap_8 FILLER_41_623 ();
 sg13g2_decap_8 FILLER_41_630 ();
 sg13g2_decap_8 FILLER_41_637 ();
 sg13g2_decap_8 FILLER_41_644 ();
 sg13g2_decap_8 FILLER_41_651 ();
 sg13g2_decap_8 FILLER_41_658 ();
 sg13g2_decap_8 FILLER_41_665 ();
 sg13g2_decap_8 FILLER_41_672 ();
 sg13g2_decap_8 FILLER_41_679 ();
 sg13g2_decap_8 FILLER_41_686 ();
 sg13g2_decap_8 FILLER_41_693 ();
 sg13g2_decap_8 FILLER_41_700 ();
 sg13g2_decap_8 FILLER_41_707 ();
 sg13g2_decap_8 FILLER_41_714 ();
 sg13g2_decap_8 FILLER_41_721 ();
 sg13g2_decap_8 FILLER_41_728 ();
 sg13g2_decap_8 FILLER_41_735 ();
 sg13g2_decap_8 FILLER_41_742 ();
 sg13g2_decap_8 FILLER_41_749 ();
 sg13g2_decap_8 FILLER_41_756 ();
 sg13g2_decap_8 FILLER_41_763 ();
 sg13g2_decap_8 FILLER_41_770 ();
 sg13g2_decap_8 FILLER_41_777 ();
 sg13g2_decap_8 FILLER_41_784 ();
 sg13g2_decap_8 FILLER_41_791 ();
 sg13g2_decap_8 FILLER_41_798 ();
 sg13g2_decap_8 FILLER_41_805 ();
 sg13g2_decap_8 FILLER_41_812 ();
 sg13g2_decap_8 FILLER_41_819 ();
 sg13g2_decap_8 FILLER_41_826 ();
 sg13g2_decap_8 FILLER_41_833 ();
 sg13g2_decap_8 FILLER_41_840 ();
 sg13g2_decap_8 FILLER_41_847 ();
 sg13g2_decap_8 FILLER_41_854 ();
 sg13g2_decap_8 FILLER_41_861 ();
 sg13g2_decap_8 FILLER_41_868 ();
 sg13g2_decap_8 FILLER_41_875 ();
 sg13g2_decap_8 FILLER_41_882 ();
 sg13g2_decap_8 FILLER_41_889 ();
 sg13g2_decap_8 FILLER_41_896 ();
 sg13g2_decap_8 FILLER_41_903 ();
 sg13g2_decap_8 FILLER_41_910 ();
 sg13g2_decap_8 FILLER_41_917 ();
 sg13g2_decap_8 FILLER_41_924 ();
 sg13g2_decap_8 FILLER_41_931 ();
 sg13g2_decap_8 FILLER_41_938 ();
 sg13g2_decap_8 FILLER_41_945 ();
 sg13g2_decap_8 FILLER_41_952 ();
 sg13g2_decap_8 FILLER_41_959 ();
 sg13g2_decap_8 FILLER_41_966 ();
 sg13g2_decap_8 FILLER_41_973 ();
 sg13g2_decap_8 FILLER_41_980 ();
 sg13g2_decap_8 FILLER_41_987 ();
 sg13g2_decap_8 FILLER_41_994 ();
 sg13g2_decap_8 FILLER_41_1001 ();
 sg13g2_decap_8 FILLER_41_1008 ();
 sg13g2_decap_8 FILLER_41_1015 ();
 sg13g2_decap_8 FILLER_41_1022 ();
 sg13g2_decap_8 FILLER_42_4 ();
 sg13g2_decap_8 FILLER_42_11 ();
 sg13g2_decap_8 FILLER_42_18 ();
 sg13g2_decap_8 FILLER_42_25 ();
 sg13g2_decap_8 FILLER_42_32 ();
 sg13g2_decap_8 FILLER_42_39 ();
 sg13g2_decap_8 FILLER_42_46 ();
 sg13g2_decap_8 FILLER_42_53 ();
 sg13g2_decap_8 FILLER_42_60 ();
 sg13g2_decap_8 FILLER_42_67 ();
 sg13g2_decap_8 FILLER_42_74 ();
 sg13g2_decap_8 FILLER_42_81 ();
 sg13g2_decap_8 FILLER_42_88 ();
 sg13g2_decap_8 FILLER_42_95 ();
 sg13g2_decap_8 FILLER_42_102 ();
 sg13g2_decap_8 FILLER_42_109 ();
 sg13g2_decap_8 FILLER_42_116 ();
 sg13g2_decap_8 FILLER_42_123 ();
 sg13g2_decap_8 FILLER_42_130 ();
 sg13g2_decap_8 FILLER_42_137 ();
 sg13g2_decap_8 FILLER_42_144 ();
 sg13g2_decap_8 FILLER_42_151 ();
 sg13g2_decap_8 FILLER_42_158 ();
 sg13g2_decap_8 FILLER_42_165 ();
 sg13g2_decap_8 FILLER_42_172 ();
 sg13g2_decap_8 FILLER_42_179 ();
 sg13g2_decap_8 FILLER_42_186 ();
 sg13g2_decap_8 FILLER_42_193 ();
 sg13g2_decap_8 FILLER_42_200 ();
 sg13g2_decap_8 FILLER_42_207 ();
 sg13g2_decap_8 FILLER_42_214 ();
 sg13g2_decap_8 FILLER_42_221 ();
 sg13g2_decap_8 FILLER_42_228 ();
 sg13g2_decap_8 FILLER_42_235 ();
 sg13g2_decap_8 FILLER_42_242 ();
 sg13g2_decap_8 FILLER_42_249 ();
 sg13g2_decap_8 FILLER_42_256 ();
 sg13g2_decap_8 FILLER_42_263 ();
 sg13g2_decap_8 FILLER_42_270 ();
 sg13g2_decap_8 FILLER_42_277 ();
 sg13g2_decap_8 FILLER_42_284 ();
 sg13g2_decap_8 FILLER_42_291 ();
 sg13g2_decap_8 FILLER_42_298 ();
 sg13g2_decap_8 FILLER_42_305 ();
 sg13g2_decap_8 FILLER_42_312 ();
 sg13g2_decap_8 FILLER_42_319 ();
 sg13g2_decap_8 FILLER_42_326 ();
 sg13g2_decap_8 FILLER_42_333 ();
 sg13g2_decap_8 FILLER_42_340 ();
 sg13g2_decap_8 FILLER_42_347 ();
 sg13g2_decap_8 FILLER_42_354 ();
 sg13g2_decap_8 FILLER_42_361 ();
 sg13g2_decap_8 FILLER_42_368 ();
 sg13g2_decap_8 FILLER_42_375 ();
 sg13g2_decap_8 FILLER_42_382 ();
 sg13g2_decap_8 FILLER_42_389 ();
 sg13g2_decap_8 FILLER_42_396 ();
 sg13g2_decap_8 FILLER_42_403 ();
 sg13g2_decap_8 FILLER_42_410 ();
 sg13g2_decap_8 FILLER_42_417 ();
 sg13g2_decap_8 FILLER_42_424 ();
 sg13g2_decap_8 FILLER_42_431 ();
 sg13g2_decap_8 FILLER_42_438 ();
 sg13g2_decap_8 FILLER_42_445 ();
 sg13g2_decap_8 FILLER_42_452 ();
 sg13g2_decap_8 FILLER_42_459 ();
 sg13g2_decap_8 FILLER_42_466 ();
 sg13g2_decap_8 FILLER_42_473 ();
 sg13g2_decap_8 FILLER_42_480 ();
 sg13g2_decap_8 FILLER_42_487 ();
 sg13g2_decap_8 FILLER_42_494 ();
 sg13g2_decap_8 FILLER_42_501 ();
 sg13g2_decap_8 FILLER_42_508 ();
 sg13g2_decap_8 FILLER_42_515 ();
 sg13g2_decap_8 FILLER_42_522 ();
 sg13g2_decap_8 FILLER_42_529 ();
 sg13g2_decap_8 FILLER_42_536 ();
 sg13g2_decap_8 FILLER_42_543 ();
 sg13g2_decap_8 FILLER_42_550 ();
 sg13g2_decap_8 FILLER_42_557 ();
 sg13g2_decap_8 FILLER_42_564 ();
 sg13g2_decap_8 FILLER_42_571 ();
 sg13g2_decap_8 FILLER_42_578 ();
 sg13g2_decap_8 FILLER_42_585 ();
 sg13g2_decap_8 FILLER_42_592 ();
 sg13g2_decap_8 FILLER_42_599 ();
 sg13g2_decap_8 FILLER_42_606 ();
 sg13g2_decap_8 FILLER_42_613 ();
 sg13g2_decap_8 FILLER_42_620 ();
 sg13g2_decap_8 FILLER_42_627 ();
 sg13g2_decap_8 FILLER_42_634 ();
 sg13g2_decap_8 FILLER_42_641 ();
 sg13g2_decap_8 FILLER_42_648 ();
 sg13g2_decap_8 FILLER_42_655 ();
 sg13g2_decap_8 FILLER_42_662 ();
 sg13g2_decap_8 FILLER_42_669 ();
 sg13g2_decap_8 FILLER_42_676 ();
 sg13g2_decap_8 FILLER_42_683 ();
 sg13g2_decap_8 FILLER_42_690 ();
 sg13g2_decap_8 FILLER_42_697 ();
 sg13g2_decap_8 FILLER_42_704 ();
 sg13g2_decap_8 FILLER_42_711 ();
 sg13g2_decap_8 FILLER_42_718 ();
 sg13g2_decap_8 FILLER_42_725 ();
 sg13g2_decap_8 FILLER_42_732 ();
 sg13g2_decap_8 FILLER_42_739 ();
 sg13g2_decap_8 FILLER_42_746 ();
 sg13g2_decap_8 FILLER_42_753 ();
 sg13g2_decap_8 FILLER_42_760 ();
 sg13g2_decap_8 FILLER_42_767 ();
 sg13g2_decap_8 FILLER_42_774 ();
 sg13g2_decap_8 FILLER_42_781 ();
 sg13g2_decap_8 FILLER_42_788 ();
 sg13g2_decap_8 FILLER_42_795 ();
 sg13g2_decap_8 FILLER_42_802 ();
 sg13g2_decap_8 FILLER_42_809 ();
 sg13g2_decap_8 FILLER_42_816 ();
 sg13g2_decap_8 FILLER_42_823 ();
 sg13g2_decap_8 FILLER_42_830 ();
 sg13g2_decap_8 FILLER_42_837 ();
 sg13g2_decap_8 FILLER_42_844 ();
 sg13g2_decap_8 FILLER_42_851 ();
 sg13g2_decap_8 FILLER_42_858 ();
 sg13g2_decap_8 FILLER_42_865 ();
 sg13g2_decap_8 FILLER_42_872 ();
 sg13g2_decap_8 FILLER_42_879 ();
 sg13g2_decap_8 FILLER_42_886 ();
 sg13g2_decap_8 FILLER_42_893 ();
 sg13g2_decap_8 FILLER_42_900 ();
 sg13g2_decap_8 FILLER_42_907 ();
 sg13g2_decap_8 FILLER_42_914 ();
 sg13g2_decap_8 FILLER_42_921 ();
 sg13g2_decap_8 FILLER_42_928 ();
 sg13g2_decap_8 FILLER_42_935 ();
 sg13g2_decap_8 FILLER_42_942 ();
 sg13g2_decap_8 FILLER_42_949 ();
 sg13g2_decap_8 FILLER_42_956 ();
 sg13g2_decap_8 FILLER_42_963 ();
 sg13g2_decap_8 FILLER_42_970 ();
 sg13g2_decap_8 FILLER_42_977 ();
 sg13g2_decap_8 FILLER_42_984 ();
 sg13g2_decap_8 FILLER_42_991 ();
 sg13g2_decap_8 FILLER_42_998 ();
 sg13g2_decap_8 FILLER_42_1005 ();
 sg13g2_decap_8 FILLER_42_1012 ();
 sg13g2_decap_8 FILLER_42_1019 ();
 sg13g2_fill_2 FILLER_42_1026 ();
 sg13g2_fill_1 FILLER_42_1028 ();
 sg13g2_decap_8 FILLER_43_4 ();
 sg13g2_decap_8 FILLER_43_11 ();
 sg13g2_decap_8 FILLER_43_18 ();
 sg13g2_decap_8 FILLER_43_25 ();
 sg13g2_decap_8 FILLER_43_32 ();
 sg13g2_decap_8 FILLER_43_39 ();
 sg13g2_decap_8 FILLER_43_46 ();
 sg13g2_decap_8 FILLER_43_53 ();
 sg13g2_decap_8 FILLER_43_60 ();
 sg13g2_decap_8 FILLER_43_67 ();
 sg13g2_decap_8 FILLER_43_74 ();
 sg13g2_decap_8 FILLER_43_81 ();
 sg13g2_decap_8 FILLER_43_88 ();
 sg13g2_decap_8 FILLER_43_95 ();
 sg13g2_decap_8 FILLER_43_102 ();
 sg13g2_decap_8 FILLER_43_109 ();
 sg13g2_decap_8 FILLER_43_116 ();
 sg13g2_decap_8 FILLER_43_123 ();
 sg13g2_decap_8 FILLER_43_130 ();
 sg13g2_decap_8 FILLER_43_137 ();
 sg13g2_decap_8 FILLER_43_144 ();
 sg13g2_decap_8 FILLER_43_151 ();
 sg13g2_decap_8 FILLER_43_158 ();
 sg13g2_decap_8 FILLER_43_165 ();
 sg13g2_decap_8 FILLER_43_172 ();
 sg13g2_decap_8 FILLER_43_179 ();
 sg13g2_decap_8 FILLER_43_186 ();
 sg13g2_decap_8 FILLER_43_193 ();
 sg13g2_decap_8 FILLER_43_200 ();
 sg13g2_decap_8 FILLER_43_207 ();
 sg13g2_decap_8 FILLER_43_214 ();
 sg13g2_decap_8 FILLER_43_221 ();
 sg13g2_decap_8 FILLER_43_228 ();
 sg13g2_decap_8 FILLER_43_235 ();
 sg13g2_decap_8 FILLER_43_242 ();
 sg13g2_decap_8 FILLER_43_249 ();
 sg13g2_decap_8 FILLER_43_256 ();
 sg13g2_decap_8 FILLER_43_263 ();
 sg13g2_decap_8 FILLER_43_270 ();
 sg13g2_decap_8 FILLER_43_277 ();
 sg13g2_decap_8 FILLER_43_284 ();
 sg13g2_decap_8 FILLER_43_291 ();
 sg13g2_decap_8 FILLER_43_298 ();
 sg13g2_decap_8 FILLER_43_305 ();
 sg13g2_decap_8 FILLER_43_312 ();
 sg13g2_decap_8 FILLER_43_319 ();
 sg13g2_decap_8 FILLER_43_326 ();
 sg13g2_decap_8 FILLER_43_333 ();
 sg13g2_decap_8 FILLER_43_340 ();
 sg13g2_decap_8 FILLER_43_347 ();
 sg13g2_decap_8 FILLER_43_354 ();
 sg13g2_decap_8 FILLER_43_361 ();
 sg13g2_decap_8 FILLER_43_368 ();
 sg13g2_decap_8 FILLER_43_375 ();
 sg13g2_decap_8 FILLER_43_382 ();
 sg13g2_decap_8 FILLER_43_389 ();
 sg13g2_decap_8 FILLER_43_396 ();
 sg13g2_decap_8 FILLER_43_403 ();
 sg13g2_decap_8 FILLER_43_410 ();
 sg13g2_decap_8 FILLER_43_417 ();
 sg13g2_decap_8 FILLER_43_424 ();
 sg13g2_decap_8 FILLER_43_431 ();
 sg13g2_decap_8 FILLER_43_438 ();
 sg13g2_decap_8 FILLER_43_445 ();
 sg13g2_decap_8 FILLER_43_452 ();
 sg13g2_decap_8 FILLER_43_459 ();
 sg13g2_decap_8 FILLER_43_466 ();
 sg13g2_decap_8 FILLER_43_473 ();
 sg13g2_decap_8 FILLER_43_480 ();
 sg13g2_decap_8 FILLER_43_487 ();
 sg13g2_decap_8 FILLER_43_494 ();
 sg13g2_decap_8 FILLER_43_501 ();
 sg13g2_decap_8 FILLER_43_508 ();
 sg13g2_decap_8 FILLER_43_515 ();
 sg13g2_decap_8 FILLER_43_522 ();
 sg13g2_decap_8 FILLER_43_529 ();
 sg13g2_decap_8 FILLER_43_536 ();
 sg13g2_decap_8 FILLER_43_543 ();
 sg13g2_decap_8 FILLER_43_550 ();
 sg13g2_decap_8 FILLER_43_557 ();
 sg13g2_decap_8 FILLER_43_564 ();
 sg13g2_decap_8 FILLER_43_571 ();
 sg13g2_decap_8 FILLER_43_578 ();
 sg13g2_decap_8 FILLER_43_585 ();
 sg13g2_decap_8 FILLER_43_592 ();
 sg13g2_decap_8 FILLER_43_599 ();
 sg13g2_decap_8 FILLER_43_606 ();
 sg13g2_decap_8 FILLER_43_613 ();
 sg13g2_decap_8 FILLER_43_620 ();
 sg13g2_decap_8 FILLER_43_627 ();
 sg13g2_decap_8 FILLER_43_634 ();
 sg13g2_decap_8 FILLER_43_641 ();
 sg13g2_decap_8 FILLER_43_648 ();
 sg13g2_decap_8 FILLER_43_655 ();
 sg13g2_decap_8 FILLER_43_662 ();
 sg13g2_decap_8 FILLER_43_669 ();
 sg13g2_decap_8 FILLER_43_676 ();
 sg13g2_decap_8 FILLER_43_683 ();
 sg13g2_decap_8 FILLER_43_690 ();
 sg13g2_decap_8 FILLER_43_697 ();
 sg13g2_decap_8 FILLER_43_704 ();
 sg13g2_decap_8 FILLER_43_711 ();
 sg13g2_decap_8 FILLER_43_718 ();
 sg13g2_decap_8 FILLER_43_725 ();
 sg13g2_decap_8 FILLER_43_732 ();
 sg13g2_decap_8 FILLER_43_739 ();
 sg13g2_decap_8 FILLER_43_746 ();
 sg13g2_decap_8 FILLER_43_753 ();
 sg13g2_decap_8 FILLER_43_760 ();
 sg13g2_decap_8 FILLER_43_767 ();
 sg13g2_decap_8 FILLER_43_774 ();
 sg13g2_decap_8 FILLER_43_781 ();
 sg13g2_decap_8 FILLER_43_788 ();
 sg13g2_decap_8 FILLER_43_795 ();
 sg13g2_decap_8 FILLER_43_802 ();
 sg13g2_decap_8 FILLER_43_809 ();
 sg13g2_decap_8 FILLER_43_816 ();
 sg13g2_decap_8 FILLER_43_823 ();
 sg13g2_decap_8 FILLER_43_830 ();
 sg13g2_decap_8 FILLER_43_837 ();
 sg13g2_decap_8 FILLER_43_844 ();
 sg13g2_decap_8 FILLER_43_851 ();
 sg13g2_decap_8 FILLER_43_858 ();
 sg13g2_decap_8 FILLER_43_865 ();
 sg13g2_decap_8 FILLER_43_872 ();
 sg13g2_decap_8 FILLER_43_879 ();
 sg13g2_decap_8 FILLER_43_886 ();
 sg13g2_decap_8 FILLER_43_893 ();
 sg13g2_decap_8 FILLER_43_900 ();
 sg13g2_decap_8 FILLER_43_907 ();
 sg13g2_decap_8 FILLER_43_914 ();
 sg13g2_decap_8 FILLER_43_921 ();
 sg13g2_decap_8 FILLER_43_928 ();
 sg13g2_decap_8 FILLER_43_935 ();
 sg13g2_decap_8 FILLER_43_942 ();
 sg13g2_decap_8 FILLER_43_949 ();
 sg13g2_decap_8 FILLER_43_956 ();
 sg13g2_decap_8 FILLER_43_963 ();
 sg13g2_decap_8 FILLER_43_970 ();
 sg13g2_decap_8 FILLER_43_977 ();
 sg13g2_decap_8 FILLER_43_984 ();
 sg13g2_decap_8 FILLER_43_991 ();
 sg13g2_decap_8 FILLER_43_998 ();
 sg13g2_decap_8 FILLER_43_1005 ();
 sg13g2_decap_8 FILLER_43_1012 ();
 sg13g2_decap_8 FILLER_43_1019 ();
 sg13g2_fill_2 FILLER_43_1026 ();
 sg13g2_fill_1 FILLER_43_1028 ();
 sg13g2_decap_8 FILLER_44_4 ();
 sg13g2_decap_8 FILLER_44_11 ();
 sg13g2_decap_8 FILLER_44_18 ();
 sg13g2_decap_8 FILLER_44_25 ();
 sg13g2_decap_8 FILLER_44_32 ();
 sg13g2_decap_8 FILLER_44_39 ();
 sg13g2_decap_8 FILLER_44_46 ();
 sg13g2_decap_8 FILLER_44_53 ();
 sg13g2_decap_8 FILLER_44_60 ();
 sg13g2_decap_8 FILLER_44_67 ();
 sg13g2_decap_8 FILLER_44_74 ();
 sg13g2_decap_8 FILLER_44_81 ();
 sg13g2_decap_8 FILLER_44_88 ();
 sg13g2_decap_8 FILLER_44_95 ();
 sg13g2_decap_8 FILLER_44_102 ();
 sg13g2_decap_8 FILLER_44_109 ();
 sg13g2_decap_8 FILLER_44_116 ();
 sg13g2_decap_8 FILLER_44_123 ();
 sg13g2_decap_8 FILLER_44_130 ();
 sg13g2_decap_8 FILLER_44_137 ();
 sg13g2_decap_8 FILLER_44_144 ();
 sg13g2_decap_8 FILLER_44_151 ();
 sg13g2_decap_8 FILLER_44_158 ();
 sg13g2_decap_8 FILLER_44_165 ();
 sg13g2_decap_8 FILLER_44_172 ();
 sg13g2_decap_8 FILLER_44_179 ();
 sg13g2_decap_8 FILLER_44_186 ();
 sg13g2_decap_8 FILLER_44_193 ();
 sg13g2_decap_8 FILLER_44_200 ();
 sg13g2_decap_8 FILLER_44_207 ();
 sg13g2_decap_8 FILLER_44_214 ();
 sg13g2_decap_8 FILLER_44_221 ();
 sg13g2_decap_8 FILLER_44_228 ();
 sg13g2_decap_8 FILLER_44_235 ();
 sg13g2_decap_8 FILLER_44_242 ();
 sg13g2_decap_8 FILLER_44_249 ();
 sg13g2_decap_8 FILLER_44_256 ();
 sg13g2_decap_8 FILLER_44_263 ();
 sg13g2_decap_8 FILLER_44_270 ();
 sg13g2_decap_8 FILLER_44_277 ();
 sg13g2_decap_8 FILLER_44_284 ();
 sg13g2_decap_8 FILLER_44_291 ();
 sg13g2_decap_8 FILLER_44_298 ();
 sg13g2_decap_8 FILLER_44_305 ();
 sg13g2_decap_8 FILLER_44_312 ();
 sg13g2_decap_8 FILLER_44_319 ();
 sg13g2_decap_8 FILLER_44_326 ();
 sg13g2_decap_8 FILLER_44_333 ();
 sg13g2_decap_8 FILLER_44_340 ();
 sg13g2_decap_8 FILLER_44_347 ();
 sg13g2_decap_8 FILLER_44_354 ();
 sg13g2_decap_8 FILLER_44_361 ();
 sg13g2_decap_8 FILLER_44_368 ();
 sg13g2_decap_8 FILLER_44_375 ();
 sg13g2_decap_8 FILLER_44_382 ();
 sg13g2_decap_8 FILLER_44_389 ();
 sg13g2_decap_8 FILLER_44_396 ();
 sg13g2_decap_8 FILLER_44_403 ();
 sg13g2_decap_8 FILLER_44_410 ();
 sg13g2_decap_8 FILLER_44_417 ();
 sg13g2_decap_8 FILLER_44_424 ();
 sg13g2_decap_8 FILLER_44_431 ();
 sg13g2_decap_8 FILLER_44_438 ();
 sg13g2_decap_8 FILLER_44_445 ();
 sg13g2_decap_8 FILLER_44_452 ();
 sg13g2_decap_8 FILLER_44_459 ();
 sg13g2_decap_8 FILLER_44_466 ();
 sg13g2_decap_8 FILLER_44_473 ();
 sg13g2_decap_8 FILLER_44_480 ();
 sg13g2_decap_8 FILLER_44_487 ();
 sg13g2_decap_8 FILLER_44_494 ();
 sg13g2_decap_8 FILLER_44_501 ();
 sg13g2_decap_8 FILLER_44_508 ();
 sg13g2_decap_8 FILLER_44_515 ();
 sg13g2_decap_8 FILLER_44_522 ();
 sg13g2_decap_8 FILLER_44_529 ();
 sg13g2_decap_8 FILLER_44_536 ();
 sg13g2_decap_8 FILLER_44_543 ();
 sg13g2_decap_8 FILLER_44_550 ();
 sg13g2_decap_8 FILLER_44_557 ();
 sg13g2_decap_8 FILLER_44_564 ();
 sg13g2_decap_8 FILLER_44_571 ();
 sg13g2_decap_8 FILLER_44_578 ();
 sg13g2_decap_8 FILLER_44_585 ();
 sg13g2_decap_8 FILLER_44_592 ();
 sg13g2_decap_8 FILLER_44_599 ();
 sg13g2_decap_8 FILLER_44_606 ();
 sg13g2_decap_8 FILLER_44_613 ();
 sg13g2_decap_8 FILLER_44_620 ();
 sg13g2_decap_8 FILLER_44_627 ();
 sg13g2_decap_8 FILLER_44_634 ();
 sg13g2_decap_8 FILLER_44_641 ();
 sg13g2_decap_8 FILLER_44_648 ();
 sg13g2_decap_8 FILLER_44_655 ();
 sg13g2_decap_8 FILLER_44_662 ();
 sg13g2_decap_8 FILLER_44_669 ();
 sg13g2_decap_8 FILLER_44_676 ();
 sg13g2_decap_8 FILLER_44_683 ();
 sg13g2_decap_8 FILLER_44_690 ();
 sg13g2_decap_8 FILLER_44_697 ();
 sg13g2_decap_8 FILLER_44_704 ();
 sg13g2_decap_8 FILLER_44_711 ();
 sg13g2_decap_8 FILLER_44_718 ();
 sg13g2_decap_8 FILLER_44_725 ();
 sg13g2_decap_8 FILLER_44_732 ();
 sg13g2_decap_8 FILLER_44_739 ();
 sg13g2_decap_8 FILLER_44_746 ();
 sg13g2_decap_8 FILLER_44_753 ();
 sg13g2_decap_8 FILLER_44_760 ();
 sg13g2_decap_8 FILLER_44_767 ();
 sg13g2_decap_8 FILLER_44_774 ();
 sg13g2_decap_8 FILLER_44_781 ();
 sg13g2_decap_8 FILLER_44_788 ();
 sg13g2_decap_8 FILLER_44_795 ();
 sg13g2_decap_8 FILLER_44_802 ();
 sg13g2_decap_8 FILLER_44_809 ();
 sg13g2_decap_8 FILLER_44_816 ();
 sg13g2_decap_8 FILLER_44_823 ();
 sg13g2_decap_8 FILLER_44_830 ();
 sg13g2_decap_8 FILLER_44_837 ();
 sg13g2_decap_8 FILLER_44_844 ();
 sg13g2_decap_8 FILLER_44_851 ();
 sg13g2_decap_8 FILLER_44_858 ();
 sg13g2_decap_8 FILLER_44_865 ();
 sg13g2_decap_8 FILLER_44_872 ();
 sg13g2_decap_8 FILLER_44_879 ();
 sg13g2_decap_8 FILLER_44_886 ();
 sg13g2_decap_8 FILLER_44_893 ();
 sg13g2_decap_8 FILLER_44_900 ();
 sg13g2_decap_8 FILLER_44_907 ();
 sg13g2_decap_8 FILLER_44_914 ();
 sg13g2_decap_8 FILLER_44_921 ();
 sg13g2_decap_8 FILLER_44_928 ();
 sg13g2_decap_8 FILLER_44_935 ();
 sg13g2_decap_8 FILLER_44_942 ();
 sg13g2_decap_8 FILLER_44_949 ();
 sg13g2_decap_8 FILLER_44_956 ();
 sg13g2_decap_8 FILLER_44_963 ();
 sg13g2_decap_8 FILLER_44_970 ();
 sg13g2_decap_8 FILLER_44_977 ();
 sg13g2_decap_8 FILLER_44_984 ();
 sg13g2_decap_8 FILLER_44_991 ();
 sg13g2_decap_8 FILLER_44_998 ();
 sg13g2_decap_8 FILLER_44_1005 ();
 sg13g2_decap_8 FILLER_44_1012 ();
 sg13g2_decap_8 FILLER_44_1019 ();
 sg13g2_fill_2 FILLER_44_1026 ();
 sg13g2_fill_1 FILLER_44_1028 ();
 sg13g2_decap_8 FILLER_45_4 ();
 sg13g2_decap_8 FILLER_45_11 ();
 sg13g2_decap_8 FILLER_45_18 ();
 sg13g2_decap_8 FILLER_45_25 ();
 sg13g2_decap_8 FILLER_45_32 ();
 sg13g2_decap_8 FILLER_45_39 ();
 sg13g2_decap_8 FILLER_45_46 ();
 sg13g2_decap_8 FILLER_45_53 ();
 sg13g2_decap_8 FILLER_45_60 ();
 sg13g2_decap_8 FILLER_45_67 ();
 sg13g2_decap_8 FILLER_45_74 ();
 sg13g2_decap_8 FILLER_45_81 ();
 sg13g2_decap_8 FILLER_45_88 ();
 sg13g2_decap_8 FILLER_45_95 ();
 sg13g2_decap_8 FILLER_45_102 ();
 sg13g2_decap_8 FILLER_45_109 ();
 sg13g2_decap_8 FILLER_45_116 ();
 sg13g2_decap_8 FILLER_45_123 ();
 sg13g2_decap_8 FILLER_45_130 ();
 sg13g2_decap_8 FILLER_45_137 ();
 sg13g2_decap_8 FILLER_45_144 ();
 sg13g2_decap_8 FILLER_45_151 ();
 sg13g2_decap_8 FILLER_45_158 ();
 sg13g2_decap_8 FILLER_45_165 ();
 sg13g2_decap_8 FILLER_45_172 ();
 sg13g2_decap_8 FILLER_45_179 ();
 sg13g2_decap_8 FILLER_45_186 ();
 sg13g2_decap_8 FILLER_45_193 ();
 sg13g2_decap_8 FILLER_45_200 ();
 sg13g2_decap_8 FILLER_45_207 ();
 sg13g2_decap_8 FILLER_45_214 ();
 sg13g2_decap_8 FILLER_45_221 ();
 sg13g2_decap_8 FILLER_45_228 ();
 sg13g2_decap_8 FILLER_45_235 ();
 sg13g2_decap_8 FILLER_45_242 ();
 sg13g2_decap_8 FILLER_45_249 ();
 sg13g2_decap_8 FILLER_45_256 ();
 sg13g2_decap_8 FILLER_45_263 ();
 sg13g2_decap_8 FILLER_45_270 ();
 sg13g2_decap_8 FILLER_45_277 ();
 sg13g2_decap_8 FILLER_45_284 ();
 sg13g2_decap_8 FILLER_45_291 ();
 sg13g2_decap_8 FILLER_45_298 ();
 sg13g2_decap_8 FILLER_45_305 ();
 sg13g2_decap_8 FILLER_45_312 ();
 sg13g2_decap_8 FILLER_45_319 ();
 sg13g2_decap_8 FILLER_45_326 ();
 sg13g2_decap_8 FILLER_45_333 ();
 sg13g2_decap_8 FILLER_45_340 ();
 sg13g2_decap_8 FILLER_45_347 ();
 sg13g2_decap_8 FILLER_45_354 ();
 sg13g2_decap_8 FILLER_45_361 ();
 sg13g2_decap_8 FILLER_45_368 ();
 sg13g2_decap_8 FILLER_45_375 ();
 sg13g2_decap_8 FILLER_45_382 ();
 sg13g2_decap_8 FILLER_45_389 ();
 sg13g2_decap_8 FILLER_45_396 ();
 sg13g2_decap_8 FILLER_45_403 ();
 sg13g2_decap_8 FILLER_45_410 ();
 sg13g2_decap_8 FILLER_45_417 ();
 sg13g2_decap_8 FILLER_45_424 ();
 sg13g2_decap_8 FILLER_45_431 ();
 sg13g2_decap_8 FILLER_45_438 ();
 sg13g2_decap_8 FILLER_45_445 ();
 sg13g2_decap_8 FILLER_45_452 ();
 sg13g2_decap_8 FILLER_45_459 ();
 sg13g2_decap_8 FILLER_45_466 ();
 sg13g2_decap_8 FILLER_45_473 ();
 sg13g2_decap_8 FILLER_45_480 ();
 sg13g2_decap_8 FILLER_45_487 ();
 sg13g2_decap_8 FILLER_45_494 ();
 sg13g2_decap_8 FILLER_45_501 ();
 sg13g2_decap_8 FILLER_45_508 ();
 sg13g2_decap_8 FILLER_45_515 ();
 sg13g2_decap_8 FILLER_45_522 ();
 sg13g2_decap_8 FILLER_45_529 ();
 sg13g2_decap_8 FILLER_45_536 ();
 sg13g2_decap_8 FILLER_45_543 ();
 sg13g2_decap_8 FILLER_45_550 ();
 sg13g2_decap_8 FILLER_45_557 ();
 sg13g2_decap_8 FILLER_45_564 ();
 sg13g2_decap_8 FILLER_45_571 ();
 sg13g2_decap_8 FILLER_45_578 ();
 sg13g2_decap_8 FILLER_45_585 ();
 sg13g2_decap_8 FILLER_45_592 ();
 sg13g2_decap_8 FILLER_45_599 ();
 sg13g2_decap_8 FILLER_45_606 ();
 sg13g2_decap_8 FILLER_45_613 ();
 sg13g2_decap_8 FILLER_45_620 ();
 sg13g2_decap_8 FILLER_45_627 ();
 sg13g2_decap_8 FILLER_45_634 ();
 sg13g2_decap_8 FILLER_45_641 ();
 sg13g2_decap_8 FILLER_45_648 ();
 sg13g2_decap_8 FILLER_45_655 ();
 sg13g2_decap_8 FILLER_45_662 ();
 sg13g2_decap_8 FILLER_45_669 ();
 sg13g2_decap_8 FILLER_45_676 ();
 sg13g2_decap_8 FILLER_45_683 ();
 sg13g2_decap_8 FILLER_45_690 ();
 sg13g2_decap_8 FILLER_45_697 ();
 sg13g2_decap_8 FILLER_45_704 ();
 sg13g2_decap_8 FILLER_45_711 ();
 sg13g2_decap_8 FILLER_45_718 ();
 sg13g2_decap_8 FILLER_45_725 ();
 sg13g2_decap_8 FILLER_45_732 ();
 sg13g2_decap_8 FILLER_45_739 ();
 sg13g2_decap_8 FILLER_45_746 ();
 sg13g2_decap_8 FILLER_45_753 ();
 sg13g2_decap_8 FILLER_45_760 ();
 sg13g2_decap_8 FILLER_45_767 ();
 sg13g2_decap_8 FILLER_45_774 ();
 sg13g2_decap_8 FILLER_45_781 ();
 sg13g2_decap_8 FILLER_45_788 ();
 sg13g2_decap_8 FILLER_45_795 ();
 sg13g2_decap_8 FILLER_45_802 ();
 sg13g2_decap_8 FILLER_45_809 ();
 sg13g2_decap_8 FILLER_45_816 ();
 sg13g2_decap_8 FILLER_45_823 ();
 sg13g2_decap_8 FILLER_45_830 ();
 sg13g2_decap_8 FILLER_45_837 ();
 sg13g2_decap_8 FILLER_45_844 ();
 sg13g2_decap_8 FILLER_45_851 ();
 sg13g2_decap_8 FILLER_45_858 ();
 sg13g2_decap_8 FILLER_45_865 ();
 sg13g2_decap_8 FILLER_45_872 ();
 sg13g2_decap_8 FILLER_45_879 ();
 sg13g2_decap_8 FILLER_45_886 ();
 sg13g2_decap_8 FILLER_45_893 ();
 sg13g2_decap_8 FILLER_45_900 ();
 sg13g2_decap_8 FILLER_45_907 ();
 sg13g2_decap_8 FILLER_45_914 ();
 sg13g2_decap_8 FILLER_45_921 ();
 sg13g2_decap_8 FILLER_45_928 ();
 sg13g2_decap_8 FILLER_45_935 ();
 sg13g2_decap_8 FILLER_45_942 ();
 sg13g2_decap_8 FILLER_45_949 ();
 sg13g2_decap_8 FILLER_45_956 ();
 sg13g2_decap_8 FILLER_45_963 ();
 sg13g2_decap_8 FILLER_45_970 ();
 sg13g2_decap_8 FILLER_45_977 ();
 sg13g2_decap_8 FILLER_45_984 ();
 sg13g2_decap_8 FILLER_45_991 ();
 sg13g2_decap_8 FILLER_45_998 ();
 sg13g2_decap_8 FILLER_45_1005 ();
 sg13g2_decap_8 FILLER_45_1012 ();
 sg13g2_decap_8 FILLER_45_1019 ();
 sg13g2_fill_2 FILLER_45_1026 ();
 sg13g2_fill_1 FILLER_45_1028 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_decap_8 FILLER_46_119 ();
 sg13g2_decap_8 FILLER_46_126 ();
 sg13g2_decap_8 FILLER_46_133 ();
 sg13g2_decap_8 FILLER_46_140 ();
 sg13g2_decap_8 FILLER_46_147 ();
 sg13g2_decap_8 FILLER_46_154 ();
 sg13g2_decap_8 FILLER_46_161 ();
 sg13g2_decap_8 FILLER_46_168 ();
 sg13g2_decap_8 FILLER_46_175 ();
 sg13g2_decap_8 FILLER_46_182 ();
 sg13g2_decap_8 FILLER_46_189 ();
 sg13g2_decap_8 FILLER_46_196 ();
 sg13g2_decap_8 FILLER_46_203 ();
 sg13g2_decap_8 FILLER_46_210 ();
 sg13g2_decap_8 FILLER_46_217 ();
 sg13g2_decap_8 FILLER_46_224 ();
 sg13g2_decap_8 FILLER_46_231 ();
 sg13g2_decap_8 FILLER_46_238 ();
 sg13g2_decap_8 FILLER_46_245 ();
 sg13g2_decap_8 FILLER_46_252 ();
 sg13g2_decap_8 FILLER_46_259 ();
 sg13g2_decap_8 FILLER_46_266 ();
 sg13g2_decap_8 FILLER_46_273 ();
 sg13g2_decap_8 FILLER_46_280 ();
 sg13g2_decap_8 FILLER_46_287 ();
 sg13g2_decap_8 FILLER_46_294 ();
 sg13g2_decap_8 FILLER_46_301 ();
 sg13g2_decap_8 FILLER_46_308 ();
 sg13g2_decap_8 FILLER_46_315 ();
 sg13g2_decap_8 FILLER_46_322 ();
 sg13g2_decap_8 FILLER_46_329 ();
 sg13g2_decap_8 FILLER_46_336 ();
 sg13g2_decap_8 FILLER_46_343 ();
 sg13g2_decap_8 FILLER_46_350 ();
 sg13g2_decap_8 FILLER_46_357 ();
 sg13g2_decap_8 FILLER_46_364 ();
 sg13g2_decap_8 FILLER_46_371 ();
 sg13g2_decap_8 FILLER_46_378 ();
 sg13g2_decap_8 FILLER_46_385 ();
 sg13g2_decap_8 FILLER_46_392 ();
 sg13g2_decap_8 FILLER_46_399 ();
 sg13g2_decap_8 FILLER_46_406 ();
 sg13g2_decap_8 FILLER_46_413 ();
 sg13g2_decap_8 FILLER_46_420 ();
 sg13g2_decap_8 FILLER_46_427 ();
 sg13g2_decap_8 FILLER_46_434 ();
 sg13g2_decap_8 FILLER_46_441 ();
 sg13g2_decap_8 FILLER_46_448 ();
 sg13g2_decap_8 FILLER_46_455 ();
 sg13g2_decap_8 FILLER_46_462 ();
 sg13g2_decap_8 FILLER_46_469 ();
 sg13g2_decap_8 FILLER_46_476 ();
 sg13g2_decap_8 FILLER_46_483 ();
 sg13g2_decap_8 FILLER_46_490 ();
 sg13g2_decap_8 FILLER_46_497 ();
 sg13g2_decap_8 FILLER_46_504 ();
 sg13g2_decap_8 FILLER_46_511 ();
 sg13g2_decap_8 FILLER_46_518 ();
 sg13g2_decap_8 FILLER_46_525 ();
 sg13g2_decap_8 FILLER_46_532 ();
 sg13g2_decap_8 FILLER_46_539 ();
 sg13g2_decap_8 FILLER_46_546 ();
 sg13g2_decap_8 FILLER_46_553 ();
 sg13g2_decap_8 FILLER_46_560 ();
 sg13g2_decap_8 FILLER_46_567 ();
 sg13g2_decap_8 FILLER_46_574 ();
 sg13g2_decap_8 FILLER_46_581 ();
 sg13g2_decap_8 FILLER_46_588 ();
 sg13g2_decap_8 FILLER_46_595 ();
 sg13g2_decap_8 FILLER_46_602 ();
 sg13g2_decap_8 FILLER_46_609 ();
 sg13g2_decap_8 FILLER_46_616 ();
 sg13g2_decap_8 FILLER_46_623 ();
 sg13g2_decap_8 FILLER_46_630 ();
 sg13g2_decap_8 FILLER_46_637 ();
 sg13g2_decap_8 FILLER_46_644 ();
 sg13g2_decap_8 FILLER_46_651 ();
 sg13g2_decap_8 FILLER_46_658 ();
 sg13g2_decap_8 FILLER_46_665 ();
 sg13g2_decap_8 FILLER_46_672 ();
 sg13g2_decap_8 FILLER_46_679 ();
 sg13g2_decap_8 FILLER_46_686 ();
 sg13g2_decap_8 FILLER_46_693 ();
 sg13g2_decap_8 FILLER_46_700 ();
 sg13g2_decap_8 FILLER_46_707 ();
 sg13g2_decap_8 FILLER_46_714 ();
 sg13g2_decap_8 FILLER_46_721 ();
 sg13g2_decap_8 FILLER_46_728 ();
 sg13g2_decap_8 FILLER_46_735 ();
 sg13g2_decap_8 FILLER_46_742 ();
 sg13g2_decap_8 FILLER_46_749 ();
 sg13g2_decap_8 FILLER_46_756 ();
 sg13g2_decap_8 FILLER_46_763 ();
 sg13g2_decap_8 FILLER_46_770 ();
 sg13g2_decap_8 FILLER_46_777 ();
 sg13g2_decap_8 FILLER_46_784 ();
 sg13g2_decap_8 FILLER_46_791 ();
 sg13g2_decap_8 FILLER_46_798 ();
 sg13g2_decap_8 FILLER_46_805 ();
 sg13g2_decap_8 FILLER_46_812 ();
 sg13g2_decap_8 FILLER_46_819 ();
 sg13g2_decap_8 FILLER_46_826 ();
 sg13g2_decap_8 FILLER_46_833 ();
 sg13g2_decap_8 FILLER_46_840 ();
 sg13g2_decap_8 FILLER_46_847 ();
 sg13g2_decap_8 FILLER_46_854 ();
 sg13g2_decap_8 FILLER_46_861 ();
 sg13g2_decap_8 FILLER_46_868 ();
 sg13g2_decap_8 FILLER_46_875 ();
 sg13g2_decap_8 FILLER_46_882 ();
 sg13g2_decap_8 FILLER_46_889 ();
 sg13g2_decap_8 FILLER_46_896 ();
 sg13g2_decap_8 FILLER_46_903 ();
 sg13g2_decap_8 FILLER_46_910 ();
 sg13g2_decap_8 FILLER_46_917 ();
 sg13g2_decap_8 FILLER_46_924 ();
 sg13g2_decap_8 FILLER_46_931 ();
 sg13g2_decap_8 FILLER_46_938 ();
 sg13g2_decap_8 FILLER_46_945 ();
 sg13g2_decap_8 FILLER_46_952 ();
 sg13g2_decap_8 FILLER_46_959 ();
 sg13g2_decap_8 FILLER_46_966 ();
 sg13g2_decap_8 FILLER_46_973 ();
 sg13g2_decap_8 FILLER_46_980 ();
 sg13g2_decap_8 FILLER_46_987 ();
 sg13g2_decap_8 FILLER_46_994 ();
 sg13g2_decap_8 FILLER_46_1001 ();
 sg13g2_decap_8 FILLER_46_1008 ();
 sg13g2_decap_8 FILLER_46_1015 ();
 sg13g2_decap_8 FILLER_46_1022 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_decap_8 FILLER_47_119 ();
 sg13g2_decap_8 FILLER_47_126 ();
 sg13g2_decap_8 FILLER_47_133 ();
 sg13g2_decap_8 FILLER_47_140 ();
 sg13g2_decap_8 FILLER_47_147 ();
 sg13g2_decap_8 FILLER_47_154 ();
 sg13g2_decap_8 FILLER_47_161 ();
 sg13g2_decap_8 FILLER_47_168 ();
 sg13g2_decap_8 FILLER_47_175 ();
 sg13g2_decap_8 FILLER_47_182 ();
 sg13g2_decap_8 FILLER_47_189 ();
 sg13g2_decap_8 FILLER_47_196 ();
 sg13g2_decap_8 FILLER_47_203 ();
 sg13g2_decap_8 FILLER_47_210 ();
 sg13g2_decap_8 FILLER_47_217 ();
 sg13g2_decap_8 FILLER_47_224 ();
 sg13g2_decap_8 FILLER_47_231 ();
 sg13g2_decap_8 FILLER_47_238 ();
 sg13g2_decap_8 FILLER_47_245 ();
 sg13g2_decap_8 FILLER_47_252 ();
 sg13g2_decap_8 FILLER_47_259 ();
 sg13g2_decap_8 FILLER_47_266 ();
 sg13g2_decap_8 FILLER_47_273 ();
 sg13g2_decap_8 FILLER_47_280 ();
 sg13g2_decap_8 FILLER_47_287 ();
 sg13g2_decap_8 FILLER_47_294 ();
 sg13g2_decap_8 FILLER_47_301 ();
 sg13g2_decap_8 FILLER_47_308 ();
 sg13g2_decap_8 FILLER_47_315 ();
 sg13g2_decap_8 FILLER_47_322 ();
 sg13g2_decap_8 FILLER_47_329 ();
 sg13g2_decap_8 FILLER_47_336 ();
 sg13g2_decap_8 FILLER_47_343 ();
 sg13g2_decap_8 FILLER_47_350 ();
 sg13g2_decap_8 FILLER_47_357 ();
 sg13g2_decap_8 FILLER_47_364 ();
 sg13g2_decap_8 FILLER_47_371 ();
 sg13g2_decap_8 FILLER_47_378 ();
 sg13g2_decap_8 FILLER_47_385 ();
 sg13g2_decap_8 FILLER_47_392 ();
 sg13g2_decap_8 FILLER_47_399 ();
 sg13g2_decap_8 FILLER_47_406 ();
 sg13g2_decap_8 FILLER_47_413 ();
 sg13g2_decap_8 FILLER_47_420 ();
 sg13g2_decap_8 FILLER_47_427 ();
 sg13g2_decap_8 FILLER_47_434 ();
 sg13g2_decap_8 FILLER_47_441 ();
 sg13g2_decap_8 FILLER_47_448 ();
 sg13g2_decap_8 FILLER_47_455 ();
 sg13g2_decap_8 FILLER_47_462 ();
 sg13g2_decap_8 FILLER_47_469 ();
 sg13g2_decap_8 FILLER_47_476 ();
 sg13g2_decap_8 FILLER_47_483 ();
 sg13g2_decap_8 FILLER_47_490 ();
 sg13g2_decap_8 FILLER_47_497 ();
 sg13g2_decap_8 FILLER_47_504 ();
 sg13g2_decap_8 FILLER_47_511 ();
 sg13g2_decap_8 FILLER_47_518 ();
 sg13g2_decap_8 FILLER_47_525 ();
 sg13g2_decap_8 FILLER_47_532 ();
 sg13g2_decap_8 FILLER_47_539 ();
 sg13g2_decap_8 FILLER_47_546 ();
 sg13g2_decap_8 FILLER_47_553 ();
 sg13g2_decap_8 FILLER_47_560 ();
 sg13g2_decap_8 FILLER_47_567 ();
 sg13g2_decap_8 FILLER_47_574 ();
 sg13g2_decap_8 FILLER_47_581 ();
 sg13g2_decap_8 FILLER_47_588 ();
 sg13g2_decap_8 FILLER_47_595 ();
 sg13g2_decap_8 FILLER_47_602 ();
 sg13g2_decap_8 FILLER_47_609 ();
 sg13g2_decap_8 FILLER_47_616 ();
 sg13g2_decap_8 FILLER_47_623 ();
 sg13g2_decap_8 FILLER_47_630 ();
 sg13g2_decap_8 FILLER_47_637 ();
 sg13g2_decap_8 FILLER_47_644 ();
 sg13g2_decap_8 FILLER_47_651 ();
 sg13g2_decap_8 FILLER_47_658 ();
 sg13g2_decap_8 FILLER_47_665 ();
 sg13g2_decap_8 FILLER_47_672 ();
 sg13g2_decap_8 FILLER_47_679 ();
 sg13g2_decap_8 FILLER_47_686 ();
 sg13g2_decap_8 FILLER_47_693 ();
 sg13g2_decap_8 FILLER_47_700 ();
 sg13g2_decap_8 FILLER_47_707 ();
 sg13g2_decap_8 FILLER_47_714 ();
 sg13g2_decap_8 FILLER_47_721 ();
 sg13g2_decap_8 FILLER_47_728 ();
 sg13g2_decap_8 FILLER_47_735 ();
 sg13g2_decap_8 FILLER_47_742 ();
 sg13g2_decap_8 FILLER_47_749 ();
 sg13g2_decap_8 FILLER_47_756 ();
 sg13g2_decap_8 FILLER_47_763 ();
 sg13g2_decap_8 FILLER_47_770 ();
 sg13g2_decap_8 FILLER_47_777 ();
 sg13g2_decap_8 FILLER_47_784 ();
 sg13g2_decap_8 FILLER_47_791 ();
 sg13g2_decap_8 FILLER_47_798 ();
 sg13g2_decap_8 FILLER_47_805 ();
 sg13g2_decap_8 FILLER_47_812 ();
 sg13g2_decap_8 FILLER_47_819 ();
 sg13g2_decap_8 FILLER_47_826 ();
 sg13g2_decap_8 FILLER_47_833 ();
 sg13g2_decap_8 FILLER_47_840 ();
 sg13g2_decap_8 FILLER_47_847 ();
 sg13g2_decap_8 FILLER_47_854 ();
 sg13g2_decap_8 FILLER_47_861 ();
 sg13g2_decap_8 FILLER_47_868 ();
 sg13g2_decap_8 FILLER_47_875 ();
 sg13g2_decap_8 FILLER_47_882 ();
 sg13g2_decap_8 FILLER_47_889 ();
 sg13g2_decap_8 FILLER_47_896 ();
 sg13g2_decap_8 FILLER_47_903 ();
 sg13g2_decap_8 FILLER_47_910 ();
 sg13g2_decap_8 FILLER_47_917 ();
 sg13g2_decap_8 FILLER_47_924 ();
 sg13g2_decap_8 FILLER_47_931 ();
 sg13g2_decap_8 FILLER_47_938 ();
 sg13g2_decap_8 FILLER_47_945 ();
 sg13g2_decap_8 FILLER_47_952 ();
 sg13g2_decap_8 FILLER_47_959 ();
 sg13g2_decap_8 FILLER_47_966 ();
 sg13g2_decap_8 FILLER_47_973 ();
 sg13g2_decap_8 FILLER_47_980 ();
 sg13g2_decap_8 FILLER_47_987 ();
 sg13g2_decap_8 FILLER_47_994 ();
 sg13g2_decap_8 FILLER_47_1001 ();
 sg13g2_decap_8 FILLER_47_1008 ();
 sg13g2_decap_8 FILLER_47_1015 ();
 sg13g2_decap_8 FILLER_47_1022 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_119 ();
 sg13g2_decap_8 FILLER_48_126 ();
 sg13g2_decap_8 FILLER_48_133 ();
 sg13g2_decap_8 FILLER_48_140 ();
 sg13g2_decap_8 FILLER_48_147 ();
 sg13g2_decap_8 FILLER_48_154 ();
 sg13g2_decap_8 FILLER_48_161 ();
 sg13g2_decap_8 FILLER_48_168 ();
 sg13g2_decap_8 FILLER_48_175 ();
 sg13g2_decap_8 FILLER_48_182 ();
 sg13g2_decap_8 FILLER_48_189 ();
 sg13g2_decap_8 FILLER_48_196 ();
 sg13g2_decap_8 FILLER_48_203 ();
 sg13g2_decap_8 FILLER_48_210 ();
 sg13g2_decap_8 FILLER_48_217 ();
 sg13g2_decap_8 FILLER_48_224 ();
 sg13g2_decap_8 FILLER_48_231 ();
 sg13g2_decap_8 FILLER_48_238 ();
 sg13g2_decap_8 FILLER_48_245 ();
 sg13g2_decap_8 FILLER_48_252 ();
 sg13g2_decap_8 FILLER_48_259 ();
 sg13g2_decap_8 FILLER_48_266 ();
 sg13g2_decap_8 FILLER_48_273 ();
 sg13g2_decap_8 FILLER_48_280 ();
 sg13g2_decap_8 FILLER_48_287 ();
 sg13g2_decap_8 FILLER_48_294 ();
 sg13g2_decap_8 FILLER_48_301 ();
 sg13g2_decap_8 FILLER_48_308 ();
 sg13g2_decap_8 FILLER_48_315 ();
 sg13g2_decap_8 FILLER_48_322 ();
 sg13g2_decap_8 FILLER_48_329 ();
 sg13g2_decap_8 FILLER_48_336 ();
 sg13g2_decap_8 FILLER_48_343 ();
 sg13g2_decap_8 FILLER_48_350 ();
 sg13g2_decap_8 FILLER_48_357 ();
 sg13g2_decap_8 FILLER_48_364 ();
 sg13g2_decap_8 FILLER_48_371 ();
 sg13g2_decap_8 FILLER_48_378 ();
 sg13g2_decap_8 FILLER_48_385 ();
 sg13g2_decap_8 FILLER_48_392 ();
 sg13g2_decap_8 FILLER_48_399 ();
 sg13g2_decap_8 FILLER_48_406 ();
 sg13g2_decap_8 FILLER_48_413 ();
 sg13g2_decap_8 FILLER_48_420 ();
 sg13g2_decap_8 FILLER_48_427 ();
 sg13g2_decap_8 FILLER_48_434 ();
 sg13g2_decap_8 FILLER_48_441 ();
 sg13g2_decap_8 FILLER_48_448 ();
 sg13g2_decap_8 FILLER_48_455 ();
 sg13g2_decap_8 FILLER_48_462 ();
 sg13g2_decap_8 FILLER_48_469 ();
 sg13g2_decap_8 FILLER_48_476 ();
 sg13g2_decap_8 FILLER_48_483 ();
 sg13g2_decap_8 FILLER_48_490 ();
 sg13g2_decap_8 FILLER_48_497 ();
 sg13g2_decap_8 FILLER_48_504 ();
 sg13g2_decap_8 FILLER_48_511 ();
 sg13g2_decap_8 FILLER_48_518 ();
 sg13g2_decap_8 FILLER_48_525 ();
 sg13g2_decap_8 FILLER_48_532 ();
 sg13g2_decap_8 FILLER_48_539 ();
 sg13g2_decap_8 FILLER_48_546 ();
 sg13g2_decap_8 FILLER_48_553 ();
 sg13g2_decap_8 FILLER_48_560 ();
 sg13g2_decap_8 FILLER_48_567 ();
 sg13g2_decap_8 FILLER_48_574 ();
 sg13g2_decap_8 FILLER_48_581 ();
 sg13g2_decap_8 FILLER_48_588 ();
 sg13g2_decap_8 FILLER_48_595 ();
 sg13g2_decap_8 FILLER_48_602 ();
 sg13g2_decap_8 FILLER_48_609 ();
 sg13g2_decap_8 FILLER_48_616 ();
 sg13g2_decap_8 FILLER_48_623 ();
 sg13g2_decap_8 FILLER_48_630 ();
 sg13g2_decap_8 FILLER_48_637 ();
 sg13g2_decap_8 FILLER_48_644 ();
 sg13g2_decap_8 FILLER_48_651 ();
 sg13g2_decap_8 FILLER_48_658 ();
 sg13g2_decap_8 FILLER_48_665 ();
 sg13g2_decap_8 FILLER_48_672 ();
 sg13g2_decap_8 FILLER_48_679 ();
 sg13g2_decap_8 FILLER_48_686 ();
 sg13g2_decap_8 FILLER_48_693 ();
 sg13g2_decap_8 FILLER_48_700 ();
 sg13g2_decap_8 FILLER_48_707 ();
 sg13g2_decap_8 FILLER_48_714 ();
 sg13g2_decap_8 FILLER_48_721 ();
 sg13g2_decap_8 FILLER_48_728 ();
 sg13g2_decap_8 FILLER_48_735 ();
 sg13g2_decap_8 FILLER_48_742 ();
 sg13g2_decap_8 FILLER_48_749 ();
 sg13g2_decap_8 FILLER_48_756 ();
 sg13g2_decap_8 FILLER_48_763 ();
 sg13g2_decap_8 FILLER_48_770 ();
 sg13g2_decap_8 FILLER_48_777 ();
 sg13g2_decap_8 FILLER_48_784 ();
 sg13g2_decap_8 FILLER_48_791 ();
 sg13g2_decap_8 FILLER_48_798 ();
 sg13g2_decap_8 FILLER_48_805 ();
 sg13g2_decap_8 FILLER_48_812 ();
 sg13g2_decap_8 FILLER_48_819 ();
 sg13g2_decap_8 FILLER_48_826 ();
 sg13g2_decap_8 FILLER_48_833 ();
 sg13g2_decap_8 FILLER_48_840 ();
 sg13g2_decap_8 FILLER_48_847 ();
 sg13g2_decap_8 FILLER_48_854 ();
 sg13g2_decap_8 FILLER_48_861 ();
 sg13g2_decap_8 FILLER_48_868 ();
 sg13g2_decap_8 FILLER_48_875 ();
 sg13g2_decap_8 FILLER_48_882 ();
 sg13g2_decap_8 FILLER_48_889 ();
 sg13g2_decap_8 FILLER_48_896 ();
 sg13g2_decap_8 FILLER_48_903 ();
 sg13g2_decap_8 FILLER_48_910 ();
 sg13g2_decap_8 FILLER_48_917 ();
 sg13g2_decap_8 FILLER_48_924 ();
 sg13g2_decap_8 FILLER_48_931 ();
 sg13g2_decap_8 FILLER_48_938 ();
 sg13g2_decap_8 FILLER_48_945 ();
 sg13g2_decap_8 FILLER_48_952 ();
 sg13g2_decap_8 FILLER_48_959 ();
 sg13g2_decap_8 FILLER_48_966 ();
 sg13g2_decap_8 FILLER_48_973 ();
 sg13g2_decap_8 FILLER_48_980 ();
 sg13g2_decap_8 FILLER_48_987 ();
 sg13g2_decap_8 FILLER_48_994 ();
 sg13g2_decap_8 FILLER_48_1001 ();
 sg13g2_decap_8 FILLER_48_1008 ();
 sg13g2_decap_8 FILLER_48_1015 ();
 sg13g2_decap_8 FILLER_48_1022 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_decap_8 FILLER_49_112 ();
 sg13g2_decap_8 FILLER_49_119 ();
 sg13g2_decap_8 FILLER_49_126 ();
 sg13g2_decap_8 FILLER_49_133 ();
 sg13g2_decap_8 FILLER_49_140 ();
 sg13g2_decap_8 FILLER_49_147 ();
 sg13g2_decap_8 FILLER_49_154 ();
 sg13g2_decap_8 FILLER_49_161 ();
 sg13g2_decap_8 FILLER_49_168 ();
 sg13g2_decap_8 FILLER_49_175 ();
 sg13g2_decap_8 FILLER_49_182 ();
 sg13g2_decap_8 FILLER_49_189 ();
 sg13g2_decap_8 FILLER_49_196 ();
 sg13g2_decap_8 FILLER_49_203 ();
 sg13g2_decap_8 FILLER_49_210 ();
 sg13g2_decap_8 FILLER_49_217 ();
 sg13g2_decap_8 FILLER_49_224 ();
 sg13g2_decap_8 FILLER_49_231 ();
 sg13g2_decap_8 FILLER_49_238 ();
 sg13g2_decap_8 FILLER_49_245 ();
 sg13g2_decap_8 FILLER_49_252 ();
 sg13g2_decap_8 FILLER_49_259 ();
 sg13g2_decap_8 FILLER_49_266 ();
 sg13g2_decap_8 FILLER_49_273 ();
 sg13g2_decap_8 FILLER_49_280 ();
 sg13g2_decap_8 FILLER_49_287 ();
 sg13g2_decap_8 FILLER_49_294 ();
 sg13g2_decap_8 FILLER_49_301 ();
 sg13g2_decap_8 FILLER_49_308 ();
 sg13g2_decap_8 FILLER_49_315 ();
 sg13g2_decap_8 FILLER_49_322 ();
 sg13g2_decap_8 FILLER_49_329 ();
 sg13g2_decap_8 FILLER_49_336 ();
 sg13g2_decap_8 FILLER_49_343 ();
 sg13g2_decap_8 FILLER_49_350 ();
 sg13g2_decap_8 FILLER_49_357 ();
 sg13g2_decap_8 FILLER_49_364 ();
 sg13g2_decap_8 FILLER_49_371 ();
 sg13g2_decap_8 FILLER_49_378 ();
 sg13g2_decap_8 FILLER_49_385 ();
 sg13g2_decap_8 FILLER_49_392 ();
 sg13g2_decap_8 FILLER_49_399 ();
 sg13g2_decap_8 FILLER_49_406 ();
 sg13g2_decap_8 FILLER_49_413 ();
 sg13g2_decap_8 FILLER_49_420 ();
 sg13g2_decap_8 FILLER_49_427 ();
 sg13g2_decap_8 FILLER_49_434 ();
 sg13g2_decap_8 FILLER_49_441 ();
 sg13g2_decap_8 FILLER_49_448 ();
 sg13g2_decap_8 FILLER_49_455 ();
 sg13g2_decap_8 FILLER_49_462 ();
 sg13g2_decap_8 FILLER_49_469 ();
 sg13g2_decap_8 FILLER_49_476 ();
 sg13g2_decap_8 FILLER_49_483 ();
 sg13g2_decap_8 FILLER_49_490 ();
 sg13g2_decap_8 FILLER_49_497 ();
 sg13g2_decap_8 FILLER_49_504 ();
 sg13g2_decap_8 FILLER_49_511 ();
 sg13g2_decap_8 FILLER_49_518 ();
 sg13g2_decap_8 FILLER_49_525 ();
 sg13g2_decap_8 FILLER_49_532 ();
 sg13g2_decap_8 FILLER_49_539 ();
 sg13g2_decap_8 FILLER_49_546 ();
 sg13g2_decap_8 FILLER_49_553 ();
 sg13g2_decap_8 FILLER_49_560 ();
 sg13g2_decap_8 FILLER_49_567 ();
 sg13g2_decap_8 FILLER_49_574 ();
 sg13g2_decap_8 FILLER_49_581 ();
 sg13g2_decap_8 FILLER_49_588 ();
 sg13g2_decap_8 FILLER_49_595 ();
 sg13g2_decap_8 FILLER_49_602 ();
 sg13g2_decap_8 FILLER_49_609 ();
 sg13g2_decap_8 FILLER_49_616 ();
 sg13g2_decap_8 FILLER_49_623 ();
 sg13g2_decap_8 FILLER_49_630 ();
 sg13g2_decap_8 FILLER_49_637 ();
 sg13g2_decap_8 FILLER_49_644 ();
 sg13g2_decap_8 FILLER_49_651 ();
 sg13g2_decap_8 FILLER_49_658 ();
 sg13g2_decap_8 FILLER_49_665 ();
 sg13g2_decap_8 FILLER_49_672 ();
 sg13g2_decap_8 FILLER_49_679 ();
 sg13g2_decap_8 FILLER_49_686 ();
 sg13g2_decap_8 FILLER_49_693 ();
 sg13g2_decap_8 FILLER_49_700 ();
 sg13g2_decap_8 FILLER_49_707 ();
 sg13g2_decap_8 FILLER_49_714 ();
 sg13g2_decap_8 FILLER_49_721 ();
 sg13g2_decap_8 FILLER_49_728 ();
 sg13g2_decap_8 FILLER_49_735 ();
 sg13g2_decap_8 FILLER_49_742 ();
 sg13g2_decap_8 FILLER_49_749 ();
 sg13g2_decap_8 FILLER_49_756 ();
 sg13g2_decap_8 FILLER_49_763 ();
 sg13g2_decap_8 FILLER_49_770 ();
 sg13g2_decap_8 FILLER_49_777 ();
 sg13g2_decap_8 FILLER_49_784 ();
 sg13g2_decap_8 FILLER_49_791 ();
 sg13g2_decap_8 FILLER_49_798 ();
 sg13g2_decap_8 FILLER_49_805 ();
 sg13g2_decap_8 FILLER_49_812 ();
 sg13g2_decap_8 FILLER_49_819 ();
 sg13g2_decap_8 FILLER_49_826 ();
 sg13g2_decap_8 FILLER_49_833 ();
 sg13g2_decap_8 FILLER_49_840 ();
 sg13g2_decap_8 FILLER_49_847 ();
 sg13g2_decap_8 FILLER_49_854 ();
 sg13g2_decap_8 FILLER_49_861 ();
 sg13g2_decap_8 FILLER_49_868 ();
 sg13g2_decap_8 FILLER_49_875 ();
 sg13g2_decap_8 FILLER_49_882 ();
 sg13g2_decap_8 FILLER_49_889 ();
 sg13g2_decap_8 FILLER_49_896 ();
 sg13g2_decap_8 FILLER_49_903 ();
 sg13g2_decap_8 FILLER_49_910 ();
 sg13g2_decap_8 FILLER_49_917 ();
 sg13g2_decap_8 FILLER_49_924 ();
 sg13g2_decap_8 FILLER_49_931 ();
 sg13g2_decap_8 FILLER_49_938 ();
 sg13g2_decap_8 FILLER_49_945 ();
 sg13g2_decap_8 FILLER_49_952 ();
 sg13g2_decap_8 FILLER_49_959 ();
 sg13g2_decap_8 FILLER_49_966 ();
 sg13g2_decap_8 FILLER_49_973 ();
 sg13g2_decap_8 FILLER_49_980 ();
 sg13g2_decap_8 FILLER_49_987 ();
 sg13g2_decap_8 FILLER_49_994 ();
 sg13g2_decap_8 FILLER_49_1001 ();
 sg13g2_decap_8 FILLER_49_1008 ();
 sg13g2_decap_8 FILLER_49_1015 ();
 sg13g2_decap_8 FILLER_49_1022 ();
 assign uio_oe[0] = net25;
 assign uio_oe[1] = net26;
 assign uio_oe[2] = net27;
 assign uio_oe[3] = net28;
 assign uio_oe[4] = net29;
 assign uio_oe[5] = net30;
 assign uio_oe[6] = net31;
 assign uio_oe[7] = net32;
 assign uio_out[0] = net33;
 assign uio_out[1] = net34;
 assign uio_out[2] = net35;
 assign uio_out[3] = net36;
 assign uio_out[4] = net37;
 assign uio_out[5] = net38;
 assign uio_out[6] = net39;
 assign uio_out[7] = net40;
endmodule
