module N_IO (A_I_top,
    A_O_top,
    A_T_top,
    A_config_C_bit0,
    A_config_C_bit1,
    A_config_C_bit2,
    A_config_C_bit3,
    B_I_top,
    B_O_top,
    B_T_top,
    B_config_C_bit0,
    B_config_C_bit1,
    B_config_C_bit2,
    B_config_C_bit3,
    Ci,
    UserCLK,
    UserCLKo,
    VPWR,
    VGND,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1END,
    N2END,
    N2MID,
    N4END,
    NN4END,
    S1BEG,
    S2BEG,
    S2BEGb,
    S4BEG,
    SS4BEG);
 output A_I_top;
 input A_O_top;
 output A_T_top;
 output A_config_C_bit0;
 output A_config_C_bit1;
 output A_config_C_bit2;
 output A_config_C_bit3;
 output B_I_top;
 input B_O_top;
 output B_T_top;
 output B_config_C_bit0;
 output B_config_C_bit1;
 output B_config_C_bit2;
 output B_config_C_bit3;
 input Ci;
 input UserCLK;
 output UserCLKo;
 inout VPWR;
 inout VGND;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 input [3:0] N1END;
 input [7:0] N2END;
 input [7:0] N2MID;
 input [15:0] N4END;
 input [15:0] NN4END;
 output [3:0] S1BEG;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 output [15:0] S4BEG;
 output [15:0] SS4BEG;

 wire \Inst_A_IO_1_bidirectional_frame_config_pass.Q ;
 wire \Inst_B_IO_1_bidirectional_frame_config_pass.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Inst_N_IO_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Inst_N_IO_switch_matrix.S1BEG0 ;
 wire \Inst_N_IO_switch_matrix.S1BEG1 ;
 wire \Inst_N_IO_switch_matrix.S1BEG2 ;
 wire \Inst_N_IO_switch_matrix.S1BEG3 ;
 wire \Inst_N_IO_switch_matrix.S2BEG0 ;
 wire \Inst_N_IO_switch_matrix.S2BEG1 ;
 wire \Inst_N_IO_switch_matrix.S2BEG2 ;
 wire \Inst_N_IO_switch_matrix.S2BEG3 ;
 wire \Inst_N_IO_switch_matrix.S2BEG4 ;
 wire \Inst_N_IO_switch_matrix.S2BEG5 ;
 wire \Inst_N_IO_switch_matrix.S2BEG6 ;
 wire \Inst_N_IO_switch_matrix.S2BEG7 ;
 wire \Inst_N_IO_switch_matrix.S2BEGb0 ;
 wire \Inst_N_IO_switch_matrix.S2BEGb1 ;
 wire \Inst_N_IO_switch_matrix.S2BEGb2 ;
 wire \Inst_N_IO_switch_matrix.S2BEGb3 ;
 wire \Inst_N_IO_switch_matrix.S2BEGb4 ;
 wire \Inst_N_IO_switch_matrix.S2BEGb5 ;
 wire \Inst_N_IO_switch_matrix.S2BEGb6 ;
 wire \Inst_N_IO_switch_matrix.S2BEGb7 ;
 wire \Inst_N_IO_switch_matrix.S4BEG0 ;
 wire \Inst_N_IO_switch_matrix.S4BEG1 ;
 wire \Inst_N_IO_switch_matrix.S4BEG10 ;
 wire \Inst_N_IO_switch_matrix.S4BEG11 ;
 wire \Inst_N_IO_switch_matrix.S4BEG12 ;
 wire \Inst_N_IO_switch_matrix.S4BEG13 ;
 wire \Inst_N_IO_switch_matrix.S4BEG14 ;
 wire \Inst_N_IO_switch_matrix.S4BEG15 ;
 wire \Inst_N_IO_switch_matrix.S4BEG2 ;
 wire \Inst_N_IO_switch_matrix.S4BEG3 ;
 wire \Inst_N_IO_switch_matrix.S4BEG4 ;
 wire \Inst_N_IO_switch_matrix.S4BEG5 ;
 wire \Inst_N_IO_switch_matrix.S4BEG6 ;
 wire \Inst_N_IO_switch_matrix.S4BEG7 ;
 wire \Inst_N_IO_switch_matrix.S4BEG8 ;
 wire \Inst_N_IO_switch_matrix.S4BEG9 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG0 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG1 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG10 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG11 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG12 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG13 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG14 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG15 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG2 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG3 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG4 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG5 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG6 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG7 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG8 ;
 wire \Inst_N_IO_switch_matrix.SS4BEG9 ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire UserCLK_regs;
 wire clknet_0_UserCLK;
 wire clknet_1_0__leaf_UserCLK;
 wire clknet_0_UserCLK_regs;
 wire clknet_1_0__leaf_UserCLK_regs;
 wire clknet_1_1__leaf_UserCLK_regs;
 wire [0:0] \Inst_N_IO_switch_matrix.DEBUG_select_S1BEG0 ;
 wire [0:0] \Inst_N_IO_switch_matrix.DEBUG_select_S1BEG1 ;
 wire [0:0] \Inst_N_IO_switch_matrix.DEBUG_select_S1BEG2 ;
 wire [0:0] \Inst_N_IO_switch_matrix.DEBUG_select_S1BEG3 ;

 sg13g2_mux4_1 _047_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit18.Q ),
    .A0(N1END[2]),
    .A1(N4END[15]),
    .A2(NN4END[15]),
    .A3(A_O_top),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit19.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _048_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit16.Q ),
    .A0(N2END[0]),
    .A1(N4END[0]),
    .A2(NN4END[0]),
    .A3(NN4END[8]),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit17.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEGb7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _049_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit14.Q ),
    .A0(N2END[1]),
    .A1(N4END[1]),
    .A2(NN4END[1]),
    .A3(NN4END[9]),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit15.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEGb6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _050_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit12.Q ),
    .A0(N2END[2]),
    .A1(N4END[2]),
    .A2(NN4END[2]),
    .A3(NN4END[10]),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit13.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEGb5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _051_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit10.Q ),
    .A0(N2END[3]),
    .A1(N4END[3]),
    .A2(NN4END[3]),
    .A3(NN4END[11]),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit11.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEGb4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _052_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit8.Q ),
    .A0(N2END[4]),
    .A1(N4END[4]),
    .A2(NN4END[4]),
    .A3(NN4END[12]),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit9.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEGb3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _053_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit6.Q ),
    .A0(N2END[5]),
    .A1(N4END[5]),
    .A2(NN4END[5]),
    .A3(NN4END[13]),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit7.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEGb2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _054_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit4.Q ),
    .A0(N2END[6]),
    .A1(N4END[6]),
    .A2(NN4END[6]),
    .A3(NN4END[14]),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit5.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEGb1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _055_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit2.Q ),
    .A0(N2END[7]),
    .A1(N4END[7]),
    .A2(NN4END[7]),
    .A3(NN4END[15]),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit3.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEGb0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _056_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit0.Q ),
    .A0(N2MID[0]),
    .A1(N4END[0]),
    .A2(NN4END[0]),
    .A3(NN4END[8]),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit1.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEG7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _057_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame3_bit30.Q ),
    .A0(N2MID[1]),
    .A1(N4END[1]),
    .A2(NN4END[1]),
    .A3(NN4END[9]),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame3_bit31.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEG6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _058_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame3_bit28.Q ),
    .A0(N2MID[2]),
    .A1(N4END[2]),
    .A2(NN4END[2]),
    .A3(NN4END[10]),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame3_bit29.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEG5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _059_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame3_bit26.Q ),
    .A0(N2MID[3]),
    .A1(N4END[3]),
    .A2(NN4END[3]),
    .A3(NN4END[11]),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame3_bit27.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEG4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _060_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame3_bit24.Q ),
    .A0(N2MID[4]),
    .A1(N4END[4]),
    .A2(NN4END[4]),
    .A3(NN4END[12]),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame3_bit25.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _061_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame3_bit22.Q ),
    .A0(N2MID[5]),
    .A1(N4END[5]),
    .A2(NN4END[5]),
    .A3(NN4END[13]),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame3_bit23.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _062_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame3_bit20.Q ),
    .A0(N2MID[6]),
    .A1(N4END[6]),
    .A2(NN4END[6]),
    .A3(NN4END[14]),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame3_bit21.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _063_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame3_bit18.Q ),
    .A0(N2MID[7]),
    .A1(N4END[7]),
    .A2(NN4END[7]),
    .A3(NN4END[15]),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame3_bit19.Q ),
    .X(\Inst_N_IO_switch_matrix.S2BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _064_ (.A0(N1END[0]),
    .A1(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S(\Inst_N_IO_switch_matrix.DEBUG_select_S1BEG3 [0]),
    .X(\Inst_N_IO_switch_matrix.S1BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _065_ (.A0(N1END[1]),
    .A1(B_O_top),
    .S(\Inst_N_IO_switch_matrix.DEBUG_select_S1BEG2 [0]),
    .X(\Inst_N_IO_switch_matrix.S1BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _066_ (.A0(N1END[2]),
    .A1(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S(\Inst_N_IO_switch_matrix.DEBUG_select_S1BEG1 [0]),
    .X(\Inst_N_IO_switch_matrix.S1BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _067_ (.A0(N1END[3]),
    .A1(A_O_top),
    .S(\Inst_N_IO_switch_matrix.DEBUG_select_S1BEG0 [0]),
    .X(\Inst_N_IO_switch_matrix.S1BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _068_ (.Y(_032_),
    .B(\Inst_N_IO_ConfigMem.Inst_frame0_bit24.Q ),
    .A_N(N2END[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _069_ (.B1(_032_),
    .VDD(VPWR),
    .Y(_033_),
    .VSS(VGND),
    .A1(N2MID[7]),
    .A2(\Inst_N_IO_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_nand3_1 _070_ (.B(\Inst_N_IO_ConfigMem.Inst_frame0_bit23.Q ),
    .C(_001_),
    .A(N2END[1]),
    .Y(_034_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _071_ (.B1(_034_),
    .VDD(VPWR),
    .Y(_035_),
    .VSS(VGND),
    .A1(\Inst_N_IO_ConfigMem.Inst_frame0_bit23.Q ),
    .A2(_033_));
 sg13g2_nand3b_1 _072_ (.B(_001_),
    .C(N2END[0]),
    .Y(_036_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\Inst_N_IO_ConfigMem.Inst_frame0_bit23.Q ));
 sg13g2_o21ai_1 _073_ (.B1(\Inst_N_IO_ConfigMem.Inst_frame0_bit23.Q ),
    .VDD(VPWR),
    .Y(_037_),
    .VSS(VGND),
    .A1(N2END[2]),
    .A2(\Inst_N_IO_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_nand2_1 _074_ (.Y(_038_),
    .A(N2END[4]),
    .B(\Inst_N_IO_ConfigMem.Inst_frame0_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _075_ (.B(_036_),
    .C(_037_),
    .A(\Inst_N_IO_ConfigMem.Inst_frame0_bit22.Q ),
    .Y(_039_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_038_));
 sg13g2_o21ai_1 _076_ (.B1(_039_),
    .VDD(VPWR),
    .Y(A_T_top),
    .VSS(VGND),
    .A1(\Inst_N_IO_ConfigMem.Inst_frame0_bit22.Q ),
    .A2(_035_));
 sg13g2_nand2b_1 _077_ (.Y(_040_),
    .B(N2END[5]),
    .A_N(\Inst_N_IO_ConfigMem.Inst_frame0_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _078_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame0_bit29.Q ),
    .A0(N2MID[6]),
    .A1(N2MID[7]),
    .A2(N2END[0]),
    .A3(N2END[4]),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame0_bit30.Q ),
    .X(_041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _079_ (.B1(\Inst_N_IO_ConfigMem.Inst_frame0_bit29.Q ),
    .VDD(VPWR),
    .Y(_042_),
    .VSS(VGND),
    .A1(N2END[6]),
    .A2(\Inst_N_IO_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_o21ai_1 _080_ (.B1(\Inst_N_IO_ConfigMem.Inst_frame0_bit31.Q ),
    .VDD(VPWR),
    .Y(_043_),
    .VSS(VGND),
    .A1(\Inst_N_IO_ConfigMem.Inst_frame0_bit29.Q ),
    .A2(_040_));
 sg13g2_nand2b_1 _081_ (.Y(_044_),
    .B(_042_),
    .A_N(_043_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _082_ (.B1(_044_),
    .VDD(VPWR),
    .Y(B_T_top),
    .VSS(VGND),
    .A1(\Inst_N_IO_ConfigMem.Inst_frame0_bit31.Q ),
    .A2(_041_));
 sg13g2_inv_1 _083_ (.VDD(VPWR),
    .Y(_000_),
    .A(N2END[1]),
    .VSS(VGND));
 sg13g2_inv_1 _084_ (.VDD(VPWR),
    .Y(_001_),
    .A(\Inst_N_IO_ConfigMem.Inst_frame0_bit24.Q ),
    .VSS(VGND));
 sg13g2_mux2_1 _085_ (.A0(N2END[2]),
    .A1(N2END[3]),
    .S(\Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .X(_002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _086_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_003_),
    .B(N2END[0]),
    .A(\Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q ));
 sg13g2_a21oi_1 _087_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .A2(_000_),
    .Y(_004_),
    .B1(\Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_a221oi_1 _088_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_004_),
    .C1(\Inst_N_IO_ConfigMem.Inst_frame0_bit27.Q ),
    .B1(_003_),
    .A1(\Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .Y(_005_),
    .A2(_002_));
 sg13g2_nand2_1 _089_ (.Y(_006_),
    .A(\Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .B(N2END[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _090_ (.Y(_007_),
    .B(N2END[4]),
    .A_N(\Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _091_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_006_),
    .A2(_007_),
    .Y(_008_),
    .B1(\Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_nor2b_1 _092_ (.A(N2END[7]),
    .B_N(\Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .Y(_009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _093_ (.B1(\Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .VDD(VPWR),
    .Y(_010_),
    .VSS(VGND),
    .A1(\Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .A2(N2END[6]));
 sg13g2_o21ai_1 _094_ (.B1(\Inst_N_IO_ConfigMem.Inst_frame0_bit27.Q ),
    .VDD(VPWR),
    .Y(_011_),
    .VSS(VGND),
    .A1(_009_),
    .A2(_010_));
 sg13g2_o21ai_1 _095_ (.B1(\Inst_N_IO_ConfigMem.Inst_frame0_bit28.Q ),
    .VDD(VPWR),
    .Y(_012_),
    .VSS(VGND),
    .A1(_008_),
    .A2(_011_));
 sg13g2_mux4_1 _096_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .A0(N2MID[4]),
    .A1(N2MID[5]),
    .A2(N2MID[6]),
    .A3(N2MID[7]),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _097_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .A0(N2MID[0]),
    .A1(N2MID[1]),
    .A2(N2MID[2]),
    .A3(N2MID[3]),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .X(_014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _098_ (.A0(_014_),
    .A1(_013_),
    .S(\Inst_N_IO_ConfigMem.Inst_frame0_bit27.Q ),
    .X(_015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _099_ (.Y(_016_),
    .B(_015_),
    .A_N(\Inst_N_IO_ConfigMem.Inst_frame0_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _100_ (.B1(_016_),
    .VDD(VPWR),
    .Y(B_I_top),
    .VSS(VGND),
    .A1(_005_),
    .A2(_012_));
 sg13g2_mux2_1 _101_ (.A0(N2END[2]),
    .A1(N2END[3]),
    .S(\Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .X(_017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _102_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_018_),
    .B(\Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .A(N2END[0]));
 sg13g2_a21oi_1 _103_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_000_),
    .A2(\Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .Y(_019_),
    .B1(\Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q ));
 sg13g2_a221oi_1 _104_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_019_),
    .C1(\Inst_N_IO_ConfigMem.Inst_frame0_bit20.Q ),
    .B1(_018_),
    .A1(\Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .Y(_020_),
    .A2(_017_));
 sg13g2_nand2_1 _105_ (.Y(_021_),
    .A(N2END[5]),
    .B(\Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _106_ (.Y(_022_),
    .B(N2END[4]),
    .A_N(\Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _107_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_021_),
    .A2(_022_),
    .Y(_023_),
    .B1(\Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q ));
 sg13g2_nor2b_1 _108_ (.A(N2END[7]),
    .B_N(\Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .Y(_024_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _109_ (.B1(\Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .VDD(VPWR),
    .Y(_025_),
    .VSS(VGND),
    .A1(N2END[6]),
    .A2(\Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q ));
 sg13g2_o21ai_1 _110_ (.B1(\Inst_N_IO_ConfigMem.Inst_frame0_bit20.Q ),
    .VDD(VPWR),
    .Y(_026_),
    .VSS(VGND),
    .A1(_024_),
    .A2(_025_));
 sg13g2_o21ai_1 _111_ (.B1(\Inst_N_IO_ConfigMem.Inst_frame0_bit21.Q ),
    .VDD(VPWR),
    .Y(_027_),
    .VSS(VGND),
    .A1(_023_),
    .A2(_026_));
 sg13g2_mux4_1 _112_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .A0(N2MID[0]),
    .A1(N2MID[1]),
    .A2(N2MID[2]),
    .A3(N2MID[3]),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .X(_028_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _113_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .A0(N2MID[4]),
    .A1(N2MID[5]),
    .A2(N2MID[6]),
    .A3(N2MID[7]),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .X(_029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _114_ (.A0(_028_),
    .A1(_029_),
    .S(\Inst_N_IO_ConfigMem.Inst_frame0_bit20.Q ),
    .X(_030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _115_ (.Y(_031_),
    .B(_030_),
    .A_N(\Inst_N_IO_ConfigMem.Inst_frame0_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _116_ (.B1(_031_),
    .VDD(VPWR),
    .Y(A_I_top),
    .VSS(VGND),
    .A1(_020_),
    .A2(_027_));
 sg13g2_mux4_1 _117_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame0_bit17.Q ),
    .A0(N2MID[1]),
    .A1(N2MID[5]),
    .A2(N2MID[3]),
    .A3(N2MID[7]),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame0_bit16.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG15 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _118_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame0_bit15.Q ),
    .A0(N2MID[0]),
    .A1(N2MID[4]),
    .A2(N2MID[2]),
    .A3(N2MID[6]),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame0_bit14.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG14 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _119_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame0_bit12.Q ),
    .A0(N4END[7]),
    .A1(N4END[9]),
    .A2(N4END[11]),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame0_bit13.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG13 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _120_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame0_bit10.Q ),
    .A0(N4END[1]),
    .A1(N4END[3]),
    .A2(N4END[5]),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame0_bit11.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG12 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _121_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame0_bit8.Q ),
    .A0(N4END[6]),
    .A1(N4END[8]),
    .A2(N4END[10]),
    .A3(B_O_top),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame0_bit9.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG11 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _122_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame0_bit6.Q ),
    .A0(N4END[0]),
    .A1(N4END[2]),
    .A2(N4END[4]),
    .A3(A_O_top),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame0_bit7.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG10 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _123_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame0_bit4.Q ),
    .A0(N4END[1]),
    .A1(N4END[3]),
    .A2(N4END[5]),
    .A3(N4END[7]),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame0_bit5.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG9 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _124_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame0_bit3.Q ),
    .A0(N4END[4]),
    .A1(N4END[8]),
    .A2(N4END[6]),
    .A3(N4END[10]),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame0_bit2.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG8 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _125_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame0_bit1.Q ),
    .A0(N2MID[1]),
    .A1(N2MID[5]),
    .A2(N2MID[3]),
    .A3(N2MID[7]),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame0_bit0.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _126_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit31.Q ),
    .A0(N2MID[0]),
    .A1(N2MID[4]),
    .A2(N2MID[2]),
    .A3(N2MID[6]),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit30.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _127_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit28.Q ),
    .A0(N2END[1]),
    .A1(N2END[3]),
    .A2(N2END[5]),
    .A3(N2END[7]),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit29.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _128_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit26.Q ),
    .A0(N2END[0]),
    .A1(N2END[2]),
    .A2(N2END[4]),
    .A3(N2END[6]),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit27.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _129_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit24.Q ),
    .A0(N4END[7]),
    .A1(N4END[9]),
    .A2(N4END[11]),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit25.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _130_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit22.Q ),
    .A0(N4END[1]),
    .A1(N4END[3]),
    .A2(N4END[5]),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit23.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _131_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit20.Q ),
    .A0(N4END[6]),
    .A1(N4END[8]),
    .A2(N4END[10]),
    .A3(B_O_top),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit21.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _132_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit18.Q ),
    .A0(N4END[0]),
    .A1(N4END[2]),
    .A2(N4END[4]),
    .A3(A_O_top),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit19.Q ),
    .X(\Inst_N_IO_switch_matrix.SS4BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _133_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit16.Q ),
    .A0(N4END[0]),
    .A1(NN4END[0]),
    .A2(NN4END[12]),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit17.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG15 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _134_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit14.Q ),
    .A0(N4END[1]),
    .A1(NN4END[1]),
    .A2(NN4END[13]),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit15.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG14 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _135_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit13.Q ),
    .A0(N1END[0]),
    .A1(NN4END[4]),
    .A2(N4END[4]),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit12.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG13 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _136_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit11.Q ),
    .A0(N1END[1]),
    .A1(NN4END[5]),
    .A2(N4END[5]),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit10.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG12 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _137_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit9.Q ),
    .A0(N4END[8]),
    .A1(NN4END[12]),
    .A2(NN4END[8]),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit8.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG11 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _138_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit7.Q ),
    .A0(N4END[9]),
    .A1(NN4END[13]),
    .A2(NN4END[9]),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit6.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG10 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _139_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit4.Q ),
    .A0(N1END[0]),
    .A1(N4END[12]),
    .A2(NN4END[12]),
    .A3(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit5.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG9 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _140_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit2.Q ),
    .A0(N1END[1]),
    .A1(N4END[13]),
    .A2(NN4END[13]),
    .A3(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit3.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG8 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _141_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame1_bit0.Q ),
    .A0(N4END[2]),
    .A1(NN4END[2]),
    .A2(NN4END[14]),
    .A3(B_O_top),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame1_bit1.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _142_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit30.Q ),
    .A0(N4END[3]),
    .A1(NN4END[3]),
    .A2(NN4END[15]),
    .A3(A_O_top),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit31.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _143_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit29.Q ),
    .A0(N1END[3]),
    .A1(NN4END[6]),
    .A2(N4END[6]),
    .A3(B_O_top),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit28.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _144_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit27.Q ),
    .A0(N1END[2]),
    .A1(NN4END[7]),
    .A2(N4END[7]),
    .A3(A_O_top),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit26.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _145_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit25.Q ),
    .A0(N4END[10]),
    .A1(NN4END[14]),
    .A2(NN4END[10]),
    .A3(B_O_top),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit24.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _146_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit23.Q ),
    .A0(N4END[11]),
    .A1(NN4END[15]),
    .A2(NN4END[11]),
    .A3(A_O_top),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit22.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _147_ (.S0(\Inst_N_IO_ConfigMem.Inst_frame2_bit20.Q ),
    .A0(N1END[3]),
    .A1(N4END[14]),
    .A2(NN4END[14]),
    .A3(B_O_top),
    .S1(\Inst_N_IO_ConfigMem.Inst_frame2_bit21.Q ),
    .X(\Inst_N_IO_switch_matrix.S4BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _148_ (.D(FrameData[6]),
    .GATE(FrameStrobe[3]),
    .Q(A_config_C_bit0),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _149_ (.D(FrameData[7]),
    .GATE(FrameStrobe[3]),
    .Q(A_config_C_bit1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _150_ (.D(FrameData[8]),
    .GATE(FrameStrobe[3]),
    .Q(A_config_C_bit2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _151_ (.D(FrameData[9]),
    .GATE(FrameStrobe[3]),
    .Q(A_config_C_bit3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _152_ (.D(FrameData[10]),
    .GATE(FrameStrobe[3]),
    .Q(B_config_C_bit0),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _153_ (.D(FrameData[11]),
    .GATE(FrameStrobe[3]),
    .Q(B_config_C_bit1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _154_ (.D(FrameData[12]),
    .GATE(FrameStrobe[3]),
    .Q(B_config_C_bit2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _155_ (.D(FrameData[13]),
    .GATE(FrameStrobe[3]),
    .Q(B_config_C_bit3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _156_ (.D(FrameData[14]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO_switch_matrix.DEBUG_select_S1BEG0 [0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _157_ (.D(FrameData[15]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO_switch_matrix.DEBUG_select_S1BEG1 [0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _158_ (.D(FrameData[16]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO_switch_matrix.DEBUG_select_S1BEG2 [0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _159_ (.D(FrameData[17]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO_switch_matrix.DEBUG_select_S1BEG3 [0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _160_ (.D(FrameData[18]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _161_ (.D(FrameData[19]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _162_ (.D(FrameData[20]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _163_ (.D(FrameData[21]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _164_ (.D(FrameData[22]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _165_ (.D(FrameData[23]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _166_ (.D(FrameData[24]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _167_ (.D(FrameData[25]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _168_ (.D(FrameData[26]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _169_ (.D(FrameData[27]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _170_ (.D(FrameData[28]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _171_ (.D(FrameData[29]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _172_ (.D(FrameData[30]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _173_ (.D(FrameData[31]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame3_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _174_ (.D(FrameData[0]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _175_ (.D(FrameData[1]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _176_ (.D(FrameData[2]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _177_ (.D(FrameData[3]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _178_ (.D(FrameData[4]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _179_ (.D(FrameData[5]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _180_ (.D(FrameData[6]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _181_ (.D(FrameData[7]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _182_ (.D(FrameData[8]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _183_ (.D(FrameData[9]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _184_ (.D(FrameData[10]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _185_ (.D(FrameData[11]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _186_ (.D(FrameData[12]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _187_ (.D(FrameData[13]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _188_ (.D(FrameData[14]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _189_ (.D(FrameData[15]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _190_ (.D(FrameData[16]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _191_ (.D(FrameData[17]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _192_ (.D(FrameData[18]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _193_ (.D(FrameData[19]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _194_ (.D(FrameData[20]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _195_ (.D(FrameData[21]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _196_ (.D(FrameData[22]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _197_ (.D(FrameData[23]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _198_ (.D(FrameData[24]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _199_ (.D(FrameData[25]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _200_ (.D(FrameData[26]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _201_ (.D(FrameData[27]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _202_ (.D(FrameData[28]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _203_ (.D(FrameData[29]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _204_ (.D(FrameData[30]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _205_ (.D(FrameData[31]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame2_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _206_ (.D(FrameData[0]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _207_ (.D(FrameData[1]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _208_ (.D(FrameData[2]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _209_ (.D(FrameData[3]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _210_ (.D(FrameData[4]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _211_ (.D(FrameData[5]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _212_ (.D(FrameData[6]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _213_ (.D(FrameData[7]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _214_ (.D(FrameData[8]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _215_ (.D(FrameData[9]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _216_ (.D(FrameData[10]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _217_ (.D(FrameData[11]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _218_ (.D(FrameData[12]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _219_ (.D(FrameData[13]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _220_ (.D(FrameData[14]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _221_ (.D(FrameData[15]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _222_ (.D(FrameData[16]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _223_ (.D(FrameData[17]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _224_ (.D(FrameData[18]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _225_ (.D(FrameData[19]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _226_ (.D(FrameData[20]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _227_ (.D(FrameData[21]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _228_ (.D(FrameData[22]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _229_ (.D(FrameData[23]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _230_ (.D(FrameData[24]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _231_ (.D(FrameData[25]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _232_ (.D(FrameData[26]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _233_ (.D(FrameData[27]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _234_ (.D(FrameData[28]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _235_ (.D(FrameData[29]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _236_ (.D(FrameData[30]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _237_ (.D(FrameData[31]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame1_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _238_ (.D(FrameData[0]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _239_ (.D(FrameData[1]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _240_ (.D(FrameData[2]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _241_ (.D(FrameData[3]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _242_ (.D(FrameData[4]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _243_ (.D(FrameData[5]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _244_ (.D(FrameData[6]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _245_ (.D(FrameData[7]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _246_ (.D(FrameData[8]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _247_ (.D(FrameData[9]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _248_ (.D(FrameData[10]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _249_ (.D(FrameData[11]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _250_ (.D(FrameData[12]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _251_ (.D(FrameData[13]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _252_ (.D(FrameData[14]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _253_ (.D(FrameData[15]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _254_ (.D(FrameData[16]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _255_ (.D(FrameData[17]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _256_ (.D(FrameData[18]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _257_ (.D(FrameData[19]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _258_ (.D(FrameData[20]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _259_ (.D(FrameData[21]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _260_ (.D(FrameData[22]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _261_ (.D(FrameData[23]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _262_ (.D(FrameData[24]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _263_ (.D(FrameData[25]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _264_ (.D(FrameData[26]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _265_ (.D(FrameData[27]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _266_ (.D(FrameData[28]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _267_ (.D(FrameData[29]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _268_ (.D(FrameData[30]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _269_ (.D(FrameData[31]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_N_IO_ConfigMem.Inst_frame0_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dfrbpq_1 _270_ (.RESET_B(_045_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(A_O_top),
    .Q(\Inst_A_IO_1_bidirectional_frame_config_pass.Q ),
    .CLK(clknet_1_1__leaf_UserCLK_regs));
 sg13g2_dfrbpq_1 _271_ (.RESET_B(_046_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(B_O_top),
    .Q(\Inst_B_IO_1_bidirectional_frame_config_pass.Q ),
    .CLK(clknet_1_0__leaf_UserCLK_regs));
 sg13g2_tiehi _272_ (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(_045_));
 sg13g2_tiehi _273_ (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(_046_));
 sg13g2_buf_1 _274_ (.A(FrameData[0]),
    .X(FrameData_O[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _275_ (.A(FrameData[1]),
    .X(FrameData_O[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _276_ (.A(FrameData[2]),
    .X(FrameData_O[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _277_ (.A(FrameData[3]),
    .X(FrameData_O[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _278_ (.A(FrameData[4]),
    .X(FrameData_O[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _279_ (.A(FrameData[5]),
    .X(FrameData_O[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _280_ (.A(FrameData[6]),
    .X(FrameData_O[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _281_ (.A(FrameData[7]),
    .X(FrameData_O[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _282_ (.A(FrameData[8]),
    .X(FrameData_O[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _283_ (.A(FrameData[9]),
    .X(FrameData_O[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _284_ (.A(FrameData[10]),
    .X(FrameData_O[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _285_ (.A(FrameData[11]),
    .X(FrameData_O[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _286_ (.A(FrameData[12]),
    .X(FrameData_O[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _287_ (.A(FrameData[13]),
    .X(FrameData_O[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _288_ (.A(FrameData[14]),
    .X(FrameData_O[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _289_ (.A(FrameData[15]),
    .X(FrameData_O[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _290_ (.A(FrameData[16]),
    .X(FrameData_O[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _291_ (.A(FrameData[17]),
    .X(FrameData_O[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _292_ (.A(FrameData[18]),
    .X(FrameData_O[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _293_ (.A(FrameData[19]),
    .X(FrameData_O[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _294_ (.A(FrameData[20]),
    .X(FrameData_O[20]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _295_ (.A(FrameData[21]),
    .X(FrameData_O[21]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _296_ (.A(FrameData[22]),
    .X(FrameData_O[22]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _297_ (.A(FrameData[23]),
    .X(FrameData_O[23]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _298_ (.A(FrameData[24]),
    .X(FrameData_O[24]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _299_ (.A(FrameData[25]),
    .X(FrameData_O[25]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _300_ (.A(FrameData[26]),
    .X(FrameData_O[26]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _301_ (.A(FrameData[27]),
    .X(FrameData_O[27]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _302_ (.A(FrameData[28]),
    .X(FrameData_O[28]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _303_ (.A(FrameData[29]),
    .X(FrameData_O[29]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _304_ (.A(FrameData[30]),
    .X(FrameData_O[30]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _305_ (.A(FrameData[31]),
    .X(FrameData_O[31]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _306_ (.A(FrameStrobe[0]),
    .X(FrameStrobe_O[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _307_ (.A(FrameStrobe[1]),
    .X(FrameStrobe_O[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _308_ (.A(FrameStrobe[2]),
    .X(FrameStrobe_O[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _309_ (.A(FrameStrobe[3]),
    .X(FrameStrobe_O[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _310_ (.A(FrameStrobe[4]),
    .X(FrameStrobe_O[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _311_ (.A(FrameStrobe[5]),
    .X(FrameStrobe_O[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _312_ (.A(FrameStrobe[6]),
    .X(FrameStrobe_O[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _313_ (.A(FrameStrobe[7]),
    .X(FrameStrobe_O[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _314_ (.A(FrameStrobe[8]),
    .X(FrameStrobe_O[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _315_ (.A(FrameStrobe[9]),
    .X(FrameStrobe_O[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _316_ (.A(FrameStrobe[10]),
    .X(FrameStrobe_O[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _317_ (.A(FrameStrobe[11]),
    .X(FrameStrobe_O[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _318_ (.A(FrameStrobe[12]),
    .X(FrameStrobe_O[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _319_ (.A(FrameStrobe[13]),
    .X(FrameStrobe_O[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _320_ (.A(FrameStrobe[14]),
    .X(FrameStrobe_O[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _321_ (.A(FrameStrobe[15]),
    .X(FrameStrobe_O[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _322_ (.A(FrameStrobe[16]),
    .X(FrameStrobe_O[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _323_ (.A(FrameStrobe[17]),
    .X(FrameStrobe_O[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _324_ (.A(FrameStrobe[18]),
    .X(FrameStrobe_O[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _325_ (.A(FrameStrobe[19]),
    .X(FrameStrobe_O[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _326_ (.A(\Inst_N_IO_switch_matrix.S1BEG0 ),
    .X(S1BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _327_ (.A(\Inst_N_IO_switch_matrix.S1BEG1 ),
    .X(S1BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _328_ (.A(\Inst_N_IO_switch_matrix.S1BEG2 ),
    .X(S1BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _329_ (.A(\Inst_N_IO_switch_matrix.S1BEG3 ),
    .X(S1BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _330_ (.A(\Inst_N_IO_switch_matrix.S2BEG0 ),
    .X(S2BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _331_ (.A(\Inst_N_IO_switch_matrix.S2BEG1 ),
    .X(S2BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _332_ (.A(\Inst_N_IO_switch_matrix.S2BEG2 ),
    .X(S2BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _333_ (.A(\Inst_N_IO_switch_matrix.S2BEG3 ),
    .X(S2BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _334_ (.A(\Inst_N_IO_switch_matrix.S2BEG4 ),
    .X(S2BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _335_ (.A(\Inst_N_IO_switch_matrix.S2BEG5 ),
    .X(S2BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _336_ (.A(\Inst_N_IO_switch_matrix.S2BEG6 ),
    .X(S2BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _337_ (.A(\Inst_N_IO_switch_matrix.S2BEG7 ),
    .X(S2BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _338_ (.A(\Inst_N_IO_switch_matrix.S2BEGb0 ),
    .X(S2BEGb[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _339_ (.A(\Inst_N_IO_switch_matrix.S2BEGb1 ),
    .X(S2BEGb[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _340_ (.A(\Inst_N_IO_switch_matrix.S2BEGb2 ),
    .X(S2BEGb[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _341_ (.A(\Inst_N_IO_switch_matrix.S2BEGb3 ),
    .X(S2BEGb[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _342_ (.A(\Inst_N_IO_switch_matrix.S2BEGb4 ),
    .X(S2BEGb[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _343_ (.A(\Inst_N_IO_switch_matrix.S2BEGb5 ),
    .X(S2BEGb[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _344_ (.A(\Inst_N_IO_switch_matrix.S2BEGb6 ),
    .X(S2BEGb[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _345_ (.A(\Inst_N_IO_switch_matrix.S2BEGb7 ),
    .X(S2BEGb[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _346_ (.A(\Inst_N_IO_switch_matrix.S4BEG0 ),
    .X(S4BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _347_ (.A(\Inst_N_IO_switch_matrix.S4BEG1 ),
    .X(S4BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _348_ (.A(\Inst_N_IO_switch_matrix.S4BEG2 ),
    .X(S4BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _349_ (.A(\Inst_N_IO_switch_matrix.S4BEG3 ),
    .X(S4BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _350_ (.A(\Inst_N_IO_switch_matrix.S4BEG4 ),
    .X(S4BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _351_ (.A(\Inst_N_IO_switch_matrix.S4BEG5 ),
    .X(S4BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _352_ (.A(\Inst_N_IO_switch_matrix.S4BEG6 ),
    .X(S4BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _353_ (.A(\Inst_N_IO_switch_matrix.S4BEG7 ),
    .X(S4BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _354_ (.A(\Inst_N_IO_switch_matrix.S4BEG8 ),
    .X(S4BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _355_ (.A(\Inst_N_IO_switch_matrix.S4BEG9 ),
    .X(S4BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _356_ (.A(\Inst_N_IO_switch_matrix.S4BEG10 ),
    .X(S4BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _357_ (.A(\Inst_N_IO_switch_matrix.S4BEG11 ),
    .X(S4BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _358_ (.A(\Inst_N_IO_switch_matrix.S4BEG12 ),
    .X(S4BEG[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _359_ (.A(\Inst_N_IO_switch_matrix.S4BEG13 ),
    .X(S4BEG[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _360_ (.A(\Inst_N_IO_switch_matrix.S4BEG14 ),
    .X(S4BEG[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _361_ (.A(\Inst_N_IO_switch_matrix.S4BEG15 ),
    .X(S4BEG[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _362_ (.A(\Inst_N_IO_switch_matrix.SS4BEG0 ),
    .X(SS4BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _363_ (.A(\Inst_N_IO_switch_matrix.SS4BEG1 ),
    .X(SS4BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _364_ (.A(\Inst_N_IO_switch_matrix.SS4BEG2 ),
    .X(SS4BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _365_ (.A(\Inst_N_IO_switch_matrix.SS4BEG3 ),
    .X(SS4BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _366_ (.A(\Inst_N_IO_switch_matrix.SS4BEG4 ),
    .X(SS4BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _367_ (.A(\Inst_N_IO_switch_matrix.SS4BEG5 ),
    .X(SS4BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _368_ (.A(\Inst_N_IO_switch_matrix.SS4BEG6 ),
    .X(SS4BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _369_ (.A(\Inst_N_IO_switch_matrix.SS4BEG7 ),
    .X(SS4BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _370_ (.A(\Inst_N_IO_switch_matrix.SS4BEG8 ),
    .X(SS4BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _371_ (.A(\Inst_N_IO_switch_matrix.SS4BEG9 ),
    .X(SS4BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _372_ (.A(\Inst_N_IO_switch_matrix.SS4BEG10 ),
    .X(SS4BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _373_ (.A(\Inst_N_IO_switch_matrix.SS4BEG11 ),
    .X(SS4BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _374_ (.A(\Inst_N_IO_switch_matrix.SS4BEG12 ),
    .X(SS4BEG[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _375_ (.A(\Inst_N_IO_switch_matrix.SS4BEG13 ),
    .X(SS4BEG[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _376_ (.A(\Inst_N_IO_switch_matrix.SS4BEG14 ),
    .X(SS4BEG[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _377_ (.A(\Inst_N_IO_switch_matrix.SS4BEG15 ),
    .X(SS4BEG[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _378_ (.A(clknet_1_0__leaf_UserCLK),
    .X(UserCLKo),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_regs_0_UserCLK (.A(UserCLK),
    .X(UserCLK_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_0_UserCLK (.A(UserCLK),
    .X(clknet_0_UserCLK),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_1_0__f_UserCLK (.A(clknet_0_UserCLK),
    .X(clknet_1_0__leaf_UserCLK),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_0_UserCLK_regs (.A(UserCLK_regs),
    .X(clknet_0_UserCLK_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_1_0__f_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_1_0__leaf_UserCLK_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_1_1__f_UserCLK_regs (.A(clknet_0_UserCLK_regs),
    .X(clknet_1_1__leaf_UserCLK_regs),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_423 (.VDD(VPWR),
    .VSS(VGND));
endmodule
