* NGSPICE file created from S_IO.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlhq_1 abstract view
.subckt sg13g2_dlhq_1 D GATE Q VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux4_1 abstract view
.subckt sg13g2_mux4_1 S0 A0 A1 A2 A3 S1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

.subckt S_IO A_I_top A_O_top A_T_top A_config_C_bit0 A_config_C_bit1 A_config_C_bit2
+ A_config_C_bit3 B_I_top B_O_top B_T_top B_config_C_bit0 B_config_C_bit1 B_config_C_bit2
+ B_config_C_bit3 Co FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3]
+ N2BEG[0] N2BEG[1] N2BEG[2] N2BEG[3] N2BEG[4] N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0]
+ N2BEGb[1] N2BEGb[2] N2BEGb[3] N2BEGb[4] N2BEGb[5] N2BEGb[6] N2BEGb[7] N4BEG[0] N4BEG[10]
+ N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2] N4BEG[3] N4BEG[4]
+ N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9] NN4BEG[0] NN4BEG[10] NN4BEG[11] NN4BEG[12]
+ NN4BEG[13] NN4BEG[14] NN4BEG[15] NN4BEG[1] NN4BEG[2] NN4BEG[3] NN4BEG[4] NN4BEG[5]
+ NN4BEG[6] NN4BEG[7] NN4BEG[8] NN4BEG[9] S1END[0] S1END[1] S1END[2] S1END[3] S2END[0]
+ S2END[1] S2END[2] S2END[3] S2END[4] S2END[5] S2END[6] S2END[7] S2MID[0] S2MID[1]
+ S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6] S2MID[7] S4END[0] S4END[10] S4END[11]
+ S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3] S4END[4] S4END[5]
+ S4END[6] S4END[7] S4END[8] S4END[9] SS4END[0] SS4END[10] SS4END[11] SS4END[12] SS4END[13]
+ SS4END[14] SS4END[15] SS4END[1] SS4END[2] SS4END[3] SS4END[4] SS4END[5] SS4END[6]
+ SS4END[7] SS4END[8] SS4END[9] UserCLK UserCLKo VGND VPWR
XFILLER_7_7 VPWR VGND sg13g2_decap_8
X_363_ Inst_S_IO_switch_matrix.NN4BEG0 NN4BEG[0] VPWR VGND sg13g2_buf_1
XFILLER_9_159 VPWR VGND sg13g2_decap_4
XFILLER_9_137 VPWR VGND sg13g2_fill_1
XFILLER_9_115 VPWR VGND sg13g2_decap_4
X_294_ FrameData[19] FrameData_O[19] VPWR VGND sg13g2_buf_1
XFILLER_3_67 VPWR VGND sg13g2_decap_8
X_346_ Inst_S_IO_switch_matrix.N2BEGb7 N2BEGb[7] VPWR VGND sg13g2_buf_1
XFILLER_2_313 VPWR VGND sg13g2_fill_2
XFILLER_5_4 VPWR VGND sg13g2_fill_1
X_277_ FrameData[2] FrameData_O[2] VPWR VGND sg13g2_buf_1
XFILLER_5_151 VPWR VGND sg13g2_decap_8
XFILLER_5_195 VPWR VGND sg13g2_decap_8
XFILLER_11_423 VPWR VGND sg13g2_fill_1
XFILLER_11_412 VPWR VGND sg13g2_fill_1
X_200_ FrameData[26] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit26.Q VPWR VGND
+ sg13g2_dlhq_1
X_131_ Inst_S_IO_ConfigMem.Inst_frame1_bit20.Q S4END[6] S4END[8] S4END[10] B_O_top
+ Inst_S_IO_ConfigMem.Inst_frame1_bit21.Q Inst_S_IO_switch_matrix.NN4BEG1 VPWR VGND
+ sg13g2_mux4_1
X_062_ Inst_S_IO_ConfigMem.Inst_frame3_bit20.Q S2MID[6] S4END[6] SS4END[6] SS4END[14]
+ Inst_S_IO_ConfigMem.Inst_frame3_bit21.Q Inst_S_IO_switch_matrix.N2BEG1 VPWR VGND
+ sg13g2_mux4_1
X_329_ Inst_S_IO_switch_matrix.N1BEG2 N1BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_2_132 VPWR VGND sg13g2_decap_4
XFILLER_7_268 VPWR VGND sg13g2_fill_1
XFILLER_7_257 VPWR VGND sg13g2_decap_8
X_114_ _028_ _029_ Inst_S_IO_ConfigMem.Inst_frame0_bit20.Q _030_ VPWR VGND sg13g2_mux2_1
XFILLER_0_230 VPWR VGND sg13g2_decap_4
XFILLER_11_0 VPWR VGND sg13g2_decap_8
X_362_ Inst_S_IO_switch_matrix.N4BEG15 N4BEG[15] VPWR VGND sg13g2_buf_1
XFILLER_5_311 VPWR VGND sg13g2_decap_8
X_293_ FrameData[18] FrameData_O[18] VPWR VGND sg13g2_buf_1
XFILLER_2_336 VPWR VGND sg13g2_fill_2
X_345_ Inst_S_IO_switch_matrix.N2BEGb6 N2BEGb[6] VPWR VGND sg13g2_buf_1
X_276_ FrameData[1] FrameData_O[1] VPWR VGND sg13g2_buf_1
X_130_ Inst_S_IO_ConfigMem.Inst_frame1_bit22.Q S4END[1] S4END[3] S4END[5] Inst_A_IO_1_bidirectional_frame_config_pass.Q
+ Inst_S_IO_ConfigMem.Inst_frame1_bit23.Q Inst_S_IO_switch_matrix.NN4BEG2 VPWR VGND
+ sg13g2_mux4_1
X_328_ Inst_S_IO_switch_matrix.N1BEG1 N1BEG[1] VPWR VGND sg13g2_buf_1
X_061_ Inst_S_IO_ConfigMem.Inst_frame3_bit22.Q S2MID[5] S4END[5] SS4END[5] SS4END[13]
+ Inst_S_IO_ConfigMem.Inst_frame3_bit23.Q Inst_S_IO_switch_matrix.N2BEG2 VPWR VGND
+ sg13g2_mux4_1
X_259_ FrameData[21] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit21.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_11_265 VPWR VGND sg13g2_fill_2
X_113_ Inst_S_IO_ConfigMem.Inst_frame0_bit18.Q S2MID[4] S2MID[5] S2MID[6] S2MID[7]
+ Inst_S_IO_ConfigMem.Inst_frame0_bit19.Q _029_ VPWR VGND sg13g2_mux4_1
XFILLER_6_280 VPWR VGND sg13g2_fill_2
XFILLER_0_423 VPWR VGND sg13g2_fill_1
XFILLER_4_228 VPWR VGND sg13g2_fill_2
XFILLER_8_364 VPWR VGND sg13g2_fill_1
XFILLER_8_342 VPWR VGND sg13g2_decap_4
X_361_ Inst_S_IO_switch_matrix.N4BEG14 N4BEG[14] VPWR VGND sg13g2_buf_1
XFILLER_9_106 VPWR VGND sg13g2_fill_1
X_292_ FrameData[17] FrameData_O[17] VPWR VGND sg13g2_buf_1
X_275_ FrameData[0] FrameData_O[0] VPWR VGND sg13g2_buf_1
X_344_ Inst_S_IO_switch_matrix.N2BEGb5 N2BEGb[5] VPWR VGND sg13g2_buf_1
XFILLER_11_403 VPWR VGND sg13g2_decap_8
X_060_ Inst_S_IO_ConfigMem.Inst_frame3_bit24.Q S2MID[4] S4END[4] SS4END[4] SS4END[12]
+ Inst_S_IO_ConfigMem.Inst_frame3_bit25.Q Inst_S_IO_switch_matrix.N2BEG3 VPWR VGND
+ sg13g2_mux4_1
XFILLER_9_24 VPWR VGND sg13g2_fill_2
XFILLER_0_48 VPWR VGND sg13g2_decap_8
XFILLER_2_101 VPWR VGND sg13g2_fill_1
X_327_ Inst_S_IO_switch_matrix.N1BEG0 N1BEG[0] VPWR VGND sg13g2_buf_1
X_189_ FrameData[15] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit15.Q VPWR VGND
+ sg13g2_dlhq_1
X_258_ FrameData[20] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit20.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_11_211 VPWR VGND sg13g2_decap_8
X_112_ Inst_S_IO_ConfigMem.Inst_frame0_bit18.Q S2MID[0] S2MID[1] S2MID[2] S2MID[3]
+ Inst_S_IO_ConfigMem.Inst_frame0_bit19.Q _028_ VPWR VGND sg13g2_mux4_1
XFILLER_1_0 VPWR VGND sg13g2_decap_8
X_360_ Inst_S_IO_switch_matrix.N4BEG13 N4BEG[13] VPWR VGND sg13g2_buf_1
X_291_ FrameData[16] FrameData_O[16] VPWR VGND sg13g2_buf_1
X_274_ VPWR VGND Co sg13g2_tielo
X_343_ Inst_S_IO_switch_matrix.N2BEGb4 N2BEGb[4] VPWR VGND sg13g2_buf_1
X_188_ FrameData[14] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit14.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_9_69 VPWR VGND sg13g2_decap_8
X_257_ FrameData[19] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit19.Q VPWR VGND
+ sg13g2_dlhq_1
X_326_ FrameStrobe[19] FrameStrobe_O[19] VPWR VGND sg13g2_buf_1
XFILLER_11_223 VPWR VGND sg13g2_fill_1
X_309_ FrameStrobe[2] FrameStrobe_O[2] VPWR VGND sg13g2_buf_1
XFILLER_11_267 VPWR VGND sg13g2_fill_1
X_111_ Inst_S_IO_ConfigMem.Inst_frame0_bit21.Q VPWR _027_ VGND _023_ _026_ sg13g2_o21ai_1
XFILLER_3_400 VPWR VGND sg13g2_decap_8
XFILLER_8_300 VPWR VGND sg13g2_fill_2
XFILLER_9_119 VPWR VGND sg13g2_fill_1
X_290_ FrameData[15] FrameData_O[15] VPWR VGND sg13g2_buf_1
X_273_ VPWR VGND _046_ sg13g2_tiehi
X_342_ Inst_S_IO_switch_matrix.N2BEGb3 N2BEGb[3] VPWR VGND sg13g2_buf_1
XFILLER_5_144 VPWR VGND sg13g2_decap_8
XFILLER_5_177 VPWR VGND sg13g2_fill_1
XFILLER_2_125 VPWR VGND sg13g2_decap_8
XFILLER_2_136 VPWR VGND sg13g2_fill_1
X_325_ FrameStrobe[18] FrameStrobe_O[18] VPWR VGND sg13g2_buf_1
X_187_ FrameData[13] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit13.Q VPWR VGND
+ sg13g2_dlhq_1
X_256_ FrameData[18] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit18.Q VPWR VGND
+ sg13g2_dlhq_1
X_110_ Inst_S_IO_ConfigMem.Inst_frame0_bit20.Q VPWR _026_ VGND _024_ _025_ sg13g2_o21ai_1
X_308_ FrameStrobe[1] FrameStrobe_O[1] VPWR VGND sg13g2_buf_1
X_239_ FrameData[1] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit1.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_6_250 VPWR VGND sg13g2_decap_4
XFILLER_0_404 VPWR VGND sg13g2_decap_4
XFILLER_3_220 VPWR VGND sg13g2_fill_2
XFILLER_8_389 VPWR VGND sg13g2_decap_4
XFILLER_7_92 VPWR VGND sg13g2_fill_2
X_272_ VPWR VGND _045_ sg13g2_tiehi
X_341_ Inst_S_IO_switch_matrix.N2BEGb2 N2BEGb[2] VPWR VGND sg13g2_buf_1
XFILLER_1_384 VPWR VGND sg13g2_fill_1
XFILLER_5_134 VPWR VGND sg13g2_decap_4
XFILLER_4_93 VPWR VGND sg13g2_decap_8
X_324_ FrameStrobe[17] FrameStrobe_O[17] VPWR VGND sg13g2_buf_1
X_186_ FrameData[12] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit12.Q VPWR VGND
+ sg13g2_dlhq_1
X_255_ FrameData[17] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit17.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_6_410 VPWR VGND sg13g2_fill_2
XFILLER_6_421 VPWR VGND sg13g2_fill_2
XFILLER_11_258 VPWR VGND sg13g2_decap_8
X_169_ FrameData[27] FrameStrobe[3] Inst_S_IO_ConfigMem.Inst_frame3_bit27.Q VPWR VGND
+ sg13g2_dlhq_1
X_307_ FrameStrobe[0] FrameStrobe_O[0] VPWR VGND sg13g2_buf_1
X_238_ FrameData[0] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit0.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_6_273 VPWR VGND sg13g2_decap_8
XFILLER_6_28 VPWR VGND sg13g2_fill_2
XFILLER_6_39 VPWR VGND sg13g2_fill_2
XFILLER_8_346 VPWR VGND sg13g2_fill_1
XFILLER_5_338 VPWR VGND sg13g2_decap_8
X_271_ _046_ VGND VPWR B_O_top Inst_B_IO_1_bidirectional_frame_config_pass.Q clknet_1_0__leaf_UserCLK_regs
+ sg13g2_dfrbpq_1
X_340_ Inst_S_IO_switch_matrix.N2BEGb1 N2BEGb[1] VPWR VGND sg13g2_buf_1
X_323_ FrameStrobe[16] FrameStrobe_O[16] VPWR VGND sg13g2_buf_1
X_254_ FrameData[16] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit16.Q VPWR VGND
+ sg13g2_dlhq_1
X_185_ FrameData[11] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit11.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_1_193 VPWR VGND sg13g2_decap_8
XFILLER_11_204 VPWR VGND sg13g2_decap_8
X_306_ FrameData[31] FrameData_O[31] VPWR VGND sg13g2_buf_1
X_168_ FrameData[26] FrameStrobe[3] Inst_S_IO_ConfigMem.Inst_frame3_bit26.Q VPWR VGND
+ sg13g2_dlhq_1
X_237_ FrameData[31] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit31.Q VPWR VGND
+ sg13g2_dlhq_1
X_099_ _016_ _015_ Inst_S_IO_ConfigMem.Inst_frame0_bit28.Q VPWR VGND sg13g2_nand2b_1
XFILLER_10_71 VPWR VGND sg13g2_decap_4
XFILLER_3_222 VPWR VGND sg13g2_fill_1
XFILLER_0_269 VPWR VGND sg13g2_decap_4
XFILLER_7_94 VPWR VGND sg13g2_fill_1
XFILLER_8_188 VPWR VGND sg13g2_decap_4
X_270_ _045_ VGND VPWR A_O_top Inst_A_IO_1_bidirectional_frame_config_pass.Q clknet_1_1__leaf_UserCLK_regs
+ sg13g2_dfrbpq_1
XFILLER_1_320 VPWR VGND sg13g2_fill_2
XFILLER_5_158 VPWR VGND sg13g2_decap_4
X_322_ FrameStrobe[15] FrameStrobe_O[15] VPWR VGND sg13g2_buf_1
X_253_ FrameData[15] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit15.Q VPWR VGND
+ sg13g2_dlhq_1
X_184_ FrameData[10] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit10.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_6_412 VPWR VGND sg13g2_fill_1
XFILLER_6_423 VPWR VGND sg13g2_fill_1
X_167_ FrameData[25] FrameStrobe[3] Inst_S_IO_ConfigMem.Inst_frame3_bit25.Q VPWR VGND
+ sg13g2_dlhq_1
X_098_ _014_ _013_ Inst_S_IO_ConfigMem.Inst_frame0_bit27.Q _015_ VPWR VGND sg13g2_mux2_1
X_305_ FrameData[30] FrameData_O[30] VPWR VGND sg13g2_buf_1
XFILLER_10_282 VPWR VGND sg13g2_decap_8
X_236_ FrameData[30] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit30.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_6_286 VPWR VGND sg13g2_fill_1
X_219_ FrameData[13] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit13.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_8_337 VPWR VGND sg13g2_fill_1
XFILLER_7_370 VPWR VGND sg13g2_decap_8
XFILLER_8_134 VPWR VGND sg13g2_fill_2
XFILLER_5_318 VPWR VGND sg13g2_fill_2
XFILLER_9_421 VPWR VGND sg13g2_fill_2
X_252_ FrameData[14] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit14.Q VPWR VGND
+ sg13g2_dlhq_1
X_321_ FrameStrobe[14] FrameStrobe_O[14] VPWR VGND sg13g2_buf_1
X_183_ FrameData[9] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit9.Q VPWR VGND
+ sg13g2_dlhq_1
X_235_ FrameData[29] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit29.Q VPWR VGND
+ sg13g2_dlhq_1
X_304_ FrameData[29] FrameData_O[29] VPWR VGND sg13g2_buf_1
X_166_ FrameData[24] FrameStrobe[3] Inst_S_IO_ConfigMem.Inst_frame3_bit24.Q VPWR VGND
+ sg13g2_dlhq_1
X_097_ Inst_S_IO_ConfigMem.Inst_frame0_bit25.Q S2MID[0] S2MID[1] S2MID[2] S2MID[3]
+ Inst_S_IO_ConfigMem.Inst_frame0_bit26.Q _014_ VPWR VGND sg13g2_mux4_1
XFILLER_6_243 VPWR VGND sg13g2_decap_8
XFILLER_6_254 VPWR VGND sg13g2_fill_2
XFILLER_0_408 VPWR VGND sg13g2_fill_1
XFILLER_3_213 VPWR VGND sg13g2_decap_8
X_149_ FrameData[7] FrameStrobe[3] A_config_C_bit1 VPWR VGND sg13g2_dlhq_1
X_218_ FrameData[12] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit12.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_8_124 VPWR VGND sg13g2_decap_4
XFILLER_8_113 VPWR VGND sg13g2_decap_8
XFILLER_5_138 VPWR VGND sg13g2_fill_2
XFILLER_1_322 VPWR VGND sg13g2_fill_1
XFILLER_4_182 VPWR VGND sg13g2_decap_8
XFILLER_2_119 VPWR VGND sg13g2_fill_2
XFILLER_4_86 VPWR VGND sg13g2_decap_8
XFILLER_10_421 VPWR VGND sg13g2_fill_2
XFILLER_8_0 VPWR VGND sg13g2_decap_4
X_320_ FrameStrobe[13] FrameStrobe_O[13] VPWR VGND sg13g2_buf_1
X_182_ FrameData[8] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit8.Q VPWR VGND
+ sg13g2_dlhq_1
X_251_ FrameData[13] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit13.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_9_296 VPWR VGND sg13g2_fill_1
XFILLER_9_230 VPWR VGND sg13g2_decap_8
XFILLER_11_218 VPWR VGND sg13g2_fill_1
XFILLER_3_417 VPWR VGND sg13g2_decap_8
X_303_ FrameData[28] FrameData_O[28] VPWR VGND sg13g2_buf_1
X_234_ FrameData[28] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit28.Q VPWR VGND
+ sg13g2_dlhq_1
X_096_ Inst_S_IO_ConfigMem.Inst_frame0_bit25.Q S2MID[4] S2MID[5] S2MID[6] S2MID[7]
+ Inst_S_IO_ConfigMem.Inst_frame0_bit26.Q _013_ VPWR VGND sg13g2_mux4_1
X_165_ FrameData[23] FrameStrobe[3] Inst_S_IO_ConfigMem.Inst_frame3_bit23.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_10_96 VPWR VGND sg13g2_fill_2
X_148_ FrameData[6] FrameStrobe[3] A_config_C_bit0 VPWR VGND sg13g2_dlhq_1
X_217_ FrameData[11] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit11.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_2_291 VPWR VGND sg13g2_decap_4
X_079_ Inst_S_IO_ConfigMem.Inst_frame0_bit29.Q VPWR _042_ VGND S2END[6] Inst_S_IO_ConfigMem.Inst_frame0_bit30.Q
+ sg13g2_o21ai_1
XFILLER_7_383 VPWR VGND sg13g2_fill_2
XFILLER_8_136 VPWR VGND sg13g2_fill_1
XFILLER_4_375 VPWR VGND sg13g2_decap_4
XFILLER_9_423 VPWR VGND sg13g2_fill_1
XFILLER_1_389 VPWR VGND sg13g2_decap_8
XFILLER_5_106 VPWR VGND sg13g2_fill_2
XFILLER_4_21 VPWR VGND sg13g2_fill_2
XFILLER_4_54 VPWR VGND sg13g2_decap_4
XFILLER_10_400 VPWR VGND sg13g2_fill_1
X_181_ FrameData[7] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit7.Q VPWR VGND
+ sg13g2_dlhq_1
X_250_ FrameData[12] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit12.Q VPWR VGND
+ sg13g2_dlhq_1
X_379_ clknet_1_0__leaf_UserCLK UserCLKo VPWR VGND sg13g2_buf_1
XFILLER_3_407 VPWR VGND sg13g2_fill_2
X_233_ FrameData[27] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit27.Q VPWR VGND
+ sg13g2_dlhq_1
X_095_ Inst_S_IO_ConfigMem.Inst_frame0_bit28.Q VPWR _012_ VGND _008_ _011_ sg13g2_o21ai_1
X_302_ FrameData[27] FrameData_O[27] VPWR VGND sg13g2_buf_1
XFILLER_10_252 VPWR VGND sg13g2_fill_1
XFILLER_10_241 VPWR VGND sg13g2_fill_2
X_164_ FrameData[22] FrameStrobe[3] Inst_S_IO_ConfigMem.Inst_frame3_bit22.Q VPWR VGND
+ sg13g2_dlhq_1
X_216_ FrameData[10] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit10.Q VPWR VGND
+ sg13g2_dlhq_1
X_078_ Inst_S_IO_ConfigMem.Inst_frame0_bit29.Q S2MID[6] S2MID[7] S2END[0] S2END[4]
+ Inst_S_IO_ConfigMem.Inst_frame0_bit30.Q _041_ VPWR VGND sg13g2_mux4_1
X_147_ Inst_S_IO_ConfigMem.Inst_frame2_bit20.Q S1END[3] S4END[14] SS4END[14] B_O_top
+ Inst_S_IO_ConfigMem.Inst_frame2_bit21.Q Inst_S_IO_switch_matrix.N4BEG1 VPWR VGND
+ sg13g2_mux4_1
Xclkbuf_1_0__f_UserCLK_regs clknet_0_UserCLK_regs clknet_1_0__leaf_UserCLK_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_7_170 VPWR VGND sg13g2_fill_1
XFILLER_0_390 VPWR VGND sg13g2_decap_8
XFILLER_10_423 VPWR VGND sg13g2_fill_1
X_180_ FrameData[6] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit6.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_9_276 VPWR VGND sg13g2_fill_2
X_378_ Inst_S_IO_switch_matrix.NN4BEG15 NN4BEG[15] VPWR VGND sg13g2_buf_1
XFILLER_1_165 VPWR VGND sg13g2_fill_1
X_094_ Inst_S_IO_ConfigMem.Inst_frame0_bit27.Q VPWR _011_ VGND _009_ _010_ sg13g2_o21ai_1
X_301_ FrameData[26] FrameData_O[26] VPWR VGND sg13g2_buf_1
X_232_ FrameData[26] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit26.Q VPWR VGND
+ sg13g2_dlhq_1
X_163_ FrameData[21] FrameStrobe[3] Inst_S_IO_ConfigMem.Inst_frame3_bit21.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_10_98 VPWR VGND sg13g2_fill_1
XFILLER_10_43 VPWR VGND sg13g2_fill_1
X_146_ Inst_S_IO_ConfigMem.Inst_frame2_bit23.Q S4END[11] SS4END[15] SS4END[11] A_O_top
+ Inst_S_IO_ConfigMem.Inst_frame2_bit22.Q Inst_S_IO_switch_matrix.N4BEG2 VPWR VGND
+ sg13g2_mux4_1
X_215_ FrameData[9] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit9.Q VPWR VGND
+ sg13g2_dlhq_1
X_077_ _040_ S2END[5] Inst_S_IO_ConfigMem.Inst_frame0_bit30.Q VPWR VGND sg13g2_nand2b_1
XFILLER_8_319 VPWR VGND sg13g2_fill_1
XFILLER_7_363 VPWR VGND sg13g2_decap_8
XFILLER_7_352 VPWR VGND sg13g2_decap_8
XFILLER_7_33 VPWR VGND sg13g2_fill_1
X_129_ Inst_S_IO_ConfigMem.Inst_frame1_bit24.Q S4END[7] S4END[9] S4END[11] Inst_B_IO_1_bidirectional_frame_config_pass.Q
+ Inst_S_IO_ConfigMem.Inst_frame1_bit25.Q Inst_S_IO_switch_matrix.NN4BEG3 VPWR VGND
+ sg13g2_mux4_1
XFILLER_5_108 VPWR VGND sg13g2_fill_1
XFILLER_4_23 VPWR VGND sg13g2_fill_1
X_377_ Inst_S_IO_switch_matrix.NN4BEG14 NN4BEG[14] VPWR VGND sg13g2_buf_1
XFILLER_9_200 VPWR VGND sg13g2_decap_4
X_093_ Inst_S_IO_ConfigMem.Inst_frame0_bit26.Q VPWR _010_ VGND Inst_S_IO_ConfigMem.Inst_frame0_bit25.Q
+ S2END[6] sg13g2_o21ai_1
X_300_ FrameData[25] FrameData_O[25] VPWR VGND sg13g2_buf_1
X_231_ FrameData[25] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit25.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_6_0 VPWR VGND sg13g2_decap_4
X_162_ FrameData[20] FrameStrobe[3] Inst_S_IO_ConfigMem.Inst_frame3_bit20.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_1_24 VPWR VGND sg13g2_fill_2
X_214_ FrameData[8] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit8.Q VPWR VGND
+ sg13g2_dlhq_1
X_076_ _039_ VPWR A_T_top VGND Inst_S_IO_ConfigMem.Inst_frame0_bit22.Q _035_ sg13g2_o21ai_1
X_145_ Inst_S_IO_ConfigMem.Inst_frame2_bit25.Q S4END[10] SS4END[14] SS4END[10] B_O_top
+ Inst_S_IO_ConfigMem.Inst_frame2_bit24.Q Inst_S_IO_switch_matrix.N4BEG3 VPWR VGND
+ sg13g2_mux4_1
Xclkbuf_1_0__f_UserCLK clknet_0_UserCLK clknet_1_0__leaf_UserCLK VPWR VGND sg13g2_buf_8
X_059_ Inst_S_IO_ConfigMem.Inst_frame3_bit26.Q S2MID[3] S4END[3] SS4END[3] SS4END[11]
+ Inst_S_IO_ConfigMem.Inst_frame3_bit27.Q Inst_S_IO_switch_matrix.N2BEG4 VPWR VGND
+ sg13g2_mux4_1
X_128_ Inst_S_IO_ConfigMem.Inst_frame1_bit26.Q S2END[0] S2END[2] S2END[4] S2END[6]
+ Inst_S_IO_ConfigMem.Inst_frame1_bit27.Q Inst_S_IO_switch_matrix.NN4BEG4 VPWR VGND
+ sg13g2_mux4_1
XFILLER_8_128 VPWR VGND sg13g2_fill_2
XFILLER_4_323 VPWR VGND sg13g2_fill_2
XFILLER_7_161 VPWR VGND sg13g2_decap_8
XFILLER_4_79 VPWR VGND sg13g2_decap_8
XFILLER_4_175 VPWR VGND sg13g2_decap_8
XFILLER_8_4 VPWR VGND sg13g2_fill_1
X_376_ Inst_S_IO_switch_matrix.NN4BEG13 NN4BEG[13] VPWR VGND sg13g2_buf_1
XFILLER_9_278 VPWR VGND sg13g2_fill_1
X_230_ FrameData[24] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit24.Q VPWR VGND
+ sg13g2_dlhq_1
X_161_ FrameData[19] FrameStrobe[3] Inst_S_IO_ConfigMem.Inst_frame3_bit19.Q VPWR VGND
+ sg13g2_dlhq_1
X_359_ Inst_S_IO_switch_matrix.N4BEG12 N4BEG[12] VPWR VGND sg13g2_buf_1
X_092_ S2END[7] Inst_S_IO_ConfigMem.Inst_frame0_bit25.Q _009_ VPWR VGND sg13g2_nor2b_1
XFILLER_2_421 VPWR VGND sg13g2_fill_2
X_144_ Inst_S_IO_ConfigMem.Inst_frame2_bit27.Q S1END[2] SS4END[7] S4END[7] A_O_top
+ Inst_S_IO_ConfigMem.Inst_frame2_bit26.Q Inst_S_IO_switch_matrix.N4BEG4 VPWR VGND
+ sg13g2_mux4_1
X_213_ FrameData[7] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit7.Q VPWR VGND
+ sg13g2_dlhq_1
X_075_ _036_ _037_ Inst_S_IO_ConfigMem.Inst_frame0_bit22.Q _039_ VPWR VGND _038_ sg13g2_nand4_1
XFILLER_2_251 VPWR VGND sg13g2_fill_1
XFILLER_2_273 VPWR VGND sg13g2_fill_1
XFILLER_2_295 VPWR VGND sg13g2_fill_1
XFILLER_11_383 VPWR VGND sg13g2_fill_2
X_127_ Inst_S_IO_ConfigMem.Inst_frame1_bit28.Q S2END[1] S2END[3] S2END[5] S2END[7]
+ Inst_S_IO_ConfigMem.Inst_frame1_bit29.Q Inst_S_IO_switch_matrix.NN4BEG5 VPWR VGND
+ sg13g2_mux4_1
X_058_ Inst_S_IO_ConfigMem.Inst_frame3_bit28.Q S2MID[2] S4END[2] SS4END[2] SS4END[10]
+ Inst_S_IO_ConfigMem.Inst_frame3_bit29.Q Inst_S_IO_switch_matrix.N2BEG5 VPWR VGND
+ sg13g2_mux4_1
XFILLER_4_379 VPWR VGND sg13g2_fill_2
XFILLER_4_121 VPWR VGND sg13g2_fill_2
X_375_ Inst_S_IO_switch_matrix.NN4BEG12 NN4BEG[12] VPWR VGND sg13g2_buf_1
X_091_ VGND VPWR _006_ _007_ _008_ Inst_S_IO_ConfigMem.Inst_frame0_bit26.Q sg13g2_a21oi_1
X_160_ FrameData[18] FrameStrobe[3] Inst_S_IO_ConfigMem.Inst_frame3_bit18.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_1_59 VPWR VGND sg13g2_decap_4
XFILLER_1_26 VPWR VGND sg13g2_fill_1
Xclkbuf_regs_0_UserCLK UserCLK UserCLK_regs VPWR VGND sg13g2_buf_8
X_358_ Inst_S_IO_switch_matrix.N4BEG11 N4BEG[11] VPWR VGND sg13g2_buf_1
XFILLER_6_205 VPWR VGND sg13g2_decap_4
X_289_ FrameData[14] FrameData_O[14] VPWR VGND sg13g2_buf_1
XFILLER_5_260 VPWR VGND sg13g2_decap_8
X_143_ Inst_S_IO_ConfigMem.Inst_frame2_bit29.Q S1END[3] SS4END[6] S4END[6] B_O_top
+ Inst_S_IO_ConfigMem.Inst_frame2_bit28.Q Inst_S_IO_switch_matrix.N4BEG5 VPWR VGND
+ sg13g2_mux4_1
X_074_ _038_ S2END[4] Inst_S_IO_ConfigMem.Inst_frame0_bit24.Q VPWR VGND sg13g2_nand2_1
X_212_ FrameData[6] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit6.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_11_351 VPWR VGND sg13g2_fill_1
X_057_ Inst_S_IO_ConfigMem.Inst_frame3_bit30.Q S2MID[1] S4END[1] SS4END[1] SS4END[9]
+ Inst_S_IO_ConfigMem.Inst_frame3_bit31.Q Inst_S_IO_switch_matrix.N2BEG6 VPWR VGND
+ sg13g2_mux4_1
X_126_ Inst_S_IO_ConfigMem.Inst_frame1_bit31.Q S2MID[0] S2MID[4] S2MID[2] S2MID[6]
+ Inst_S_IO_ConfigMem.Inst_frame1_bit30.Q Inst_S_IO_switch_matrix.NN4BEG6 VPWR VGND
+ sg13g2_mux4_1
XFILLER_7_377 VPWR VGND sg13g2_fill_2
XFILLER_7_311 VPWR VGND sg13g2_fill_2
XFILLER_7_14 VPWR VGND sg13g2_fill_2
XFILLER_4_325 VPWR VGND sg13g2_fill_1
XFILLER_4_347 VPWR VGND sg13g2_fill_2
XFILLER_11_181 VPWR VGND sg13g2_fill_2
X_109_ Inst_S_IO_ConfigMem.Inst_frame0_bit19.Q VPWR _025_ VGND S2END[6] Inst_S_IO_ConfigMem.Inst_frame0_bit18.Q
+ sg13g2_o21ai_1
XFILLER_9_406 VPWR VGND sg13g2_fill_2
XFILLER_0_383 VPWR VGND sg13g2_decap_8
XFILLER_4_144 VPWR VGND sg13g2_fill_2
X_374_ Inst_S_IO_switch_matrix.NN4BEG11 NN4BEG[11] VPWR VGND sg13g2_buf_1
X_090_ _007_ S2END[4] Inst_S_IO_ConfigMem.Inst_frame0_bit25.Q VPWR VGND sg13g2_nand2b_1
XFILLER_10_202 VPWR VGND sg13g2_fill_1
XFILLER_2_423 VPWR VGND sg13g2_fill_1
Xclkbuf_0_UserCLK_regs UserCLK_regs clknet_0_UserCLK_regs VPWR VGND sg13g2_buf_8
X_357_ Inst_S_IO_switch_matrix.N4BEG10 N4BEG[10] VPWR VGND sg13g2_buf_1
X_288_ FrameData[13] FrameData_O[13] VPWR VGND sg13g2_buf_1
X_142_ Inst_S_IO_ConfigMem.Inst_frame2_bit30.Q S4END[3] SS4END[3] SS4END[15] A_O_top
+ Inst_S_IO_ConfigMem.Inst_frame2_bit31.Q Inst_S_IO_switch_matrix.N4BEG6 VPWR VGND
+ sg13g2_mux4_1
X_211_ FrameData[5] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit5.Q VPWR VGND
+ sg13g2_dlhq_1
X_073_ Inst_S_IO_ConfigMem.Inst_frame0_bit23.Q VPWR _037_ VGND S2END[2] Inst_S_IO_ConfigMem.Inst_frame0_bit24.Q
+ sg13g2_o21ai_1
XFILLER_4_0 VPWR VGND sg13g2_decap_4
XFILLER_2_81 VPWR VGND sg13g2_fill_1
XFILLER_11_385 VPWR VGND sg13g2_fill_1
X_125_ Inst_S_IO_ConfigMem.Inst_frame0_bit1.Q S2MID[1] S2MID[5] S2MID[3] S2MID[7]
+ Inst_S_IO_ConfigMem.Inst_frame0_bit0.Q Inst_S_IO_switch_matrix.NN4BEG7 VPWR VGND
+ sg13g2_mux4_1
X_056_ Inst_S_IO_ConfigMem.Inst_frame2_bit0.Q S2MID[0] S4END[0] SS4END[0] SS4END[8]
+ Inst_S_IO_ConfigMem.Inst_frame2_bit1.Q Inst_S_IO_switch_matrix.N2BEG7 VPWR VGND
+ sg13g2_mux4_1
XFILLER_4_304 VPWR VGND sg13g2_fill_2
XFILLER_11_160 VPWR VGND sg13g2_fill_2
X_108_ S2END[7] Inst_S_IO_ConfigMem.Inst_frame0_bit18.Q _024_ VPWR VGND sg13g2_nor2b_1
XFILLER_4_189 VPWR VGND sg13g2_decap_4
XFILLER_9_237 VPWR VGND sg13g2_fill_1
XFILLER_9_204 VPWR VGND sg13g2_fill_1
X_373_ Inst_S_IO_switch_matrix.NN4BEG10 NN4BEG[10] VPWR VGND sg13g2_buf_1
XFILLER_5_421 VPWR VGND sg13g2_fill_2
XFILLER_5_70 VPWR VGND sg13g2_decap_8
XFILLER_10_247 VPWR VGND sg13g2_fill_1
X_356_ Inst_S_IO_switch_matrix.N4BEG9 N4BEG[9] VPWR VGND sg13g2_buf_1
X_287_ FrameData[12] FrameData_O[12] VPWR VGND sg13g2_buf_1
X_210_ FrameData[4] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit4.Q VPWR VGND
+ sg13g2_dlhq_1
X_072_ _001_ S2END[0] _036_ VPWR VGND Inst_S_IO_ConfigMem.Inst_frame0_bit23.Q sg13g2_nand3b_1
X_141_ Inst_S_IO_ConfigMem.Inst_frame1_bit0.Q S4END[2] SS4END[2] SS4END[14] B_O_top
+ Inst_S_IO_ConfigMem.Inst_frame1_bit1.Q Inst_S_IO_switch_matrix.N4BEG7 VPWR VGND
+ sg13g2_mux4_1
X_339_ Inst_S_IO_switch_matrix.N2BEGb0 N2BEGb[0] VPWR VGND sg13g2_buf_1
XFILLER_7_313 VPWR VGND sg13g2_fill_1
X_124_ Inst_S_IO_ConfigMem.Inst_frame0_bit3.Q S4END[4] S4END[8] S4END[6] S4END[10]
+ Inst_S_IO_ConfigMem.Inst_frame0_bit2.Q Inst_S_IO_switch_matrix.NN4BEG8 VPWR VGND
+ sg13g2_mux4_1
X_055_ Inst_S_IO_ConfigMem.Inst_frame2_bit2.Q S2END[7] S4END[7] SS4END[7] SS4END[15]
+ Inst_S_IO_ConfigMem.Inst_frame2_bit3.Q Inst_S_IO_switch_matrix.N2BEGb0 VPWR VGND
+ sg13g2_mux4_1
XFILLER_4_349 VPWR VGND sg13g2_fill_1
XFILLER_3_393 VPWR VGND sg13g2_decap_8
X_107_ VGND VPWR _021_ _022_ _023_ Inst_S_IO_ConfigMem.Inst_frame0_bit19.Q sg13g2_a21oi_1
XFILLER_9_408 VPWR VGND sg13g2_fill_1
XFILLER_4_146 VPWR VGND sg13g2_fill_1
XFILLER_4_168 VPWR VGND sg13g2_decap_8
X_372_ Inst_S_IO_switch_matrix.NN4BEG9 NN4BEG[9] VPWR VGND sg13g2_buf_1
XFILLER_8_293 VPWR VGND sg13g2_decap_8
X_355_ Inst_S_IO_switch_matrix.N4BEG8 N4BEG[8] VPWR VGND sg13g2_buf_1
X_286_ FrameData[11] FrameData_O[11] VPWR VGND sg13g2_buf_1
XFILLER_5_230 VPWR VGND sg13g2_decap_4
XFILLER_10_49 VPWR VGND sg13g2_fill_1
X_071_ _034_ VPWR _035_ VGND Inst_S_IO_ConfigMem.Inst_frame0_bit23.Q _033_ sg13g2_o21ai_1
X_140_ Inst_S_IO_ConfigMem.Inst_frame1_bit2.Q S1END[1] S4END[13] SS4END[13] Inst_A_IO_1_bidirectional_frame_config_pass.Q
+ Inst_S_IO_ConfigMem.Inst_frame1_bit3.Q Inst_S_IO_switch_matrix.N4BEG8 VPWR VGND
+ sg13g2_mux4_1
X_269_ FrameData[31] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit31.Q VPWR VGND
+ sg13g2_dlhq_1
Xclkbuf_1_1__f_UserCLK_regs clknet_0_UserCLK_regs clknet_1_1__leaf_UserCLK_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_2_72 VPWR VGND sg13g2_decap_8
X_338_ Inst_S_IO_switch_matrix.N2BEG7 N2BEG[7] VPWR VGND sg13g2_buf_1
X_054_ Inst_S_IO_ConfigMem.Inst_frame2_bit4.Q S2END[6] S4END[6] SS4END[6] SS4END[14]
+ Inst_S_IO_ConfigMem.Inst_frame2_bit5.Q Inst_S_IO_switch_matrix.N2BEGb1 VPWR VGND
+ sg13g2_mux4_1
X_123_ Inst_S_IO_ConfigMem.Inst_frame0_bit4.Q S4END[1] S4END[3] S4END[5] S4END[7]
+ Inst_S_IO_ConfigMem.Inst_frame0_bit5.Q Inst_S_IO_switch_matrix.NN4BEG9 VPWR VGND
+ sg13g2_mux4_1
XFILLER_11_162 VPWR VGND sg13g2_fill_1
XFILLER_7_188 VPWR VGND sg13g2_fill_2
X_106_ _022_ S2END[4] Inst_S_IO_ConfigMem.Inst_frame0_bit18.Q VPWR VGND sg13g2_nand2b_1
XFILLER_0_397 VPWR VGND sg13g2_decap_8
X_371_ Inst_S_IO_switch_matrix.NN4BEG8 NN4BEG[8] VPWR VGND sg13g2_buf_1
XFILLER_5_423 VPWR VGND sg13g2_fill_1
X_285_ FrameData[10] FrameData_O[10] VPWR VGND sg13g2_buf_1
X_354_ Inst_S_IO_switch_matrix.N4BEG7 N4BEG[7] VPWR VGND sg13g2_buf_1
XFILLER_5_253 VPWR VGND sg13g2_decap_8
X_070_ Inst_S_IO_ConfigMem.Inst_frame0_bit23.Q _001_ S2END[1] _034_ VPWR VGND sg13g2_nand3_1
X_337_ Inst_S_IO_switch_matrix.N2BEG6 N2BEG[6] VPWR VGND sg13g2_buf_1
X_199_ FrameData[25] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit25.Q VPWR VGND
+ sg13g2_dlhq_1
X_268_ FrameData[30] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit30.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_11_377 VPWR VGND sg13g2_fill_2
XFILLER_2_0 VPWR VGND sg13g2_decap_4
X_122_ Inst_S_IO_ConfigMem.Inst_frame0_bit6.Q S4END[0] S4END[2] S4END[4] A_O_top Inst_S_IO_ConfigMem.Inst_frame0_bit7.Q
+ Inst_S_IO_switch_matrix.NN4BEG10 VPWR VGND sg13g2_mux4_1
X_053_ Inst_S_IO_ConfigMem.Inst_frame2_bit6.Q S2END[5] S4END[5] SS4END[5] SS4END[13]
+ Inst_S_IO_ConfigMem.Inst_frame2_bit7.Q Inst_S_IO_switch_matrix.N2BEGb2 VPWR VGND
+ sg13g2_mux4_1
XFILLER_11_174 VPWR VGND sg13g2_decap_8
X_105_ _021_ S2END[5] Inst_S_IO_ConfigMem.Inst_frame0_bit18.Q VPWR VGND sg13g2_nand2_1
XFILLER_8_421 VPWR VGND sg13g2_fill_2
XFILLER_8_410 VPWR VGND sg13g2_fill_2
XFILLER_0_140 VPWR VGND sg13g2_decap_8
X_370_ Inst_S_IO_switch_matrix.NN4BEG7 NN4BEG[7] VPWR VGND sg13g2_buf_1
XFILLER_5_84 VPWR VGND sg13g2_fill_1
X_353_ Inst_S_IO_switch_matrix.N4BEG6 N4BEG[6] VPWR VGND sg13g2_buf_1
XFILLER_2_405 VPWR VGND sg13g2_decap_4
X_284_ FrameData[9] FrameData_O[9] VPWR VGND sg13g2_buf_1
XFILLER_2_213 VPWR VGND sg13g2_decap_4
X_336_ Inst_S_IO_switch_matrix.N2BEG5 N2BEG[5] VPWR VGND sg13g2_buf_1
X_267_ FrameData[29] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit29.Q VPWR VGND
+ sg13g2_dlhq_1
X_198_ FrameData[24] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit24.Q VPWR VGND
+ sg13g2_dlhq_1
X_121_ Inst_S_IO_ConfigMem.Inst_frame0_bit8.Q S4END[6] S4END[8] S4END[10] B_O_top
+ Inst_S_IO_ConfigMem.Inst_frame0_bit9.Q Inst_S_IO_switch_matrix.NN4BEG11 VPWR VGND
+ sg13g2_mux4_1
X_052_ Inst_S_IO_ConfigMem.Inst_frame2_bit8.Q S2END[4] S4END[4] SS4END[4] SS4END[12]
+ Inst_S_IO_ConfigMem.Inst_frame2_bit9.Q Inst_S_IO_switch_matrix.N2BEGb3 VPWR VGND
+ sg13g2_mux4_1
X_319_ FrameStrobe[12] FrameStrobe_O[12] VPWR VGND sg13g2_buf_1
XFILLER_7_168 VPWR VGND sg13g2_fill_2
X_104_ VPWR VGND _019_ Inst_S_IO_ConfigMem.Inst_frame0_bit20.Q _018_ Inst_S_IO_ConfigMem.Inst_frame0_bit19.Q
+ _020_ _017_ sg13g2_a221oi_1
XFILLER_10_0 VPWR VGND sg13g2_decap_4
X_352_ Inst_S_IO_switch_matrix.N4BEG5 N4BEG[5] VPWR VGND sg13g2_buf_1
X_283_ FrameData[8] FrameData_O[8] VPWR VGND sg13g2_buf_1
X_266_ FrameData[28] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit28.Q VPWR VGND
+ sg13g2_dlhq_1
X_335_ Inst_S_IO_switch_matrix.N2BEG4 N2BEG[4] VPWR VGND sg13g2_buf_1
XFILLER_2_247 VPWR VGND sg13g2_decap_4
X_197_ FrameData[23] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit23.Q VPWR VGND
+ sg13g2_dlhq_1
X_120_ Inst_S_IO_ConfigMem.Inst_frame0_bit10.Q S4END[1] S4END[3] S4END[5] Inst_A_IO_1_bidirectional_frame_config_pass.Q
+ Inst_S_IO_ConfigMem.Inst_frame0_bit11.Q Inst_S_IO_switch_matrix.NN4BEG12 VPWR VGND
+ sg13g2_mux4_1
X_051_ Inst_S_IO_ConfigMem.Inst_frame2_bit10.Q S2END[3] S4END[3] SS4END[3] SS4END[11]
+ Inst_S_IO_ConfigMem.Inst_frame2_bit11.Q Inst_S_IO_switch_matrix.N2BEGb4 VPWR VGND
+ sg13g2_mux4_1
X_318_ FrameStrobe[11] FrameStrobe_O[11] VPWR VGND sg13g2_buf_1
X_249_ FrameData[11] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit11.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_11_132 VPWR VGND sg13g2_fill_2
XFILLER_3_320 VPWR VGND sg13g2_decap_4
XFILLER_3_375 VPWR VGND sg13g2_fill_1
X_103_ VGND VPWR _000_ Inst_S_IO_ConfigMem.Inst_frame0_bit18.Q _019_ Inst_S_IO_ConfigMem.Inst_frame0_bit19.Q
+ sg13g2_a21oi_1
XFILLER_8_423 VPWR VGND sg13g2_fill_1
XFILLER_8_412 VPWR VGND sg13g2_fill_1
XFILLER_0_356 VPWR VGND sg13g2_fill_2
X_351_ Inst_S_IO_switch_matrix.N4BEG4 N4BEG[4] VPWR VGND sg13g2_buf_1
X_282_ FrameData[7] FrameData_O[7] VPWR VGND sg13g2_buf_1
XFILLER_5_234 VPWR VGND sg13g2_fill_2
XFILLER_5_267 VPWR VGND sg13g2_fill_2
X_334_ Inst_S_IO_switch_matrix.N2BEG3 N2BEG[3] VPWR VGND sg13g2_buf_1
X_265_ FrameData[27] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit27.Q VPWR VGND
+ sg13g2_dlhq_1
X_196_ FrameData[22] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit22.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_11_369 VPWR VGND sg13g2_decap_4
XFILLER_11_347 VPWR VGND sg13g2_decap_4
X_050_ Inst_S_IO_ConfigMem.Inst_frame2_bit12.Q S2END[2] S4END[2] SS4END[2] SS4END[10]
+ Inst_S_IO_ConfigMem.Inst_frame2_bit13.Q Inst_S_IO_switch_matrix.N2BEGb5 VPWR VGND
+ sg13g2_mux4_1
X_317_ FrameStrobe[10] FrameStrobe_O[10] VPWR VGND sg13g2_buf_1
X_179_ FrameData[5] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit5.Q VPWR VGND
+ sg13g2_dlhq_1
X_248_ FrameData[10] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit10.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_3_310 VPWR VGND sg13g2_fill_2
X_102_ VGND VPWR _018_ Inst_S_IO_ConfigMem.Inst_frame0_bit18.Q S2END[0] sg13g2_or2_1
XFILLER_7_137 VPWR VGND sg13g2_fill_2
XFILLER_8_64 VPWR VGND sg13g2_decap_8
XFILLER_3_195 VPWR VGND sg13g2_fill_1
XFILLER_0_154 VPWR VGND sg13g2_fill_2
X_350_ Inst_S_IO_switch_matrix.N4BEG3 N4BEG[3] VPWR VGND sg13g2_buf_1
X_281_ FrameData[6] FrameData_O[6] VPWR VGND sg13g2_buf_1
XFILLER_5_202 VPWR VGND sg13g2_fill_2
X_264_ FrameData[26] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit26.Q VPWR VGND
+ sg13g2_dlhq_1
X_333_ Inst_S_IO_switch_matrix.N2BEG2 N2BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_2_99 VPWR VGND sg13g2_fill_2
X_195_ FrameData[21] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit21.Q VPWR VGND
+ sg13g2_dlhq_1
X_316_ FrameStrobe[9] FrameStrobe_O[9] VPWR VGND sg13g2_buf_1
X_247_ FrameData[9] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit9.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_2_4 VPWR VGND sg13g2_fill_2
X_178_ FrameData[4] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit4.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_11_167 VPWR VGND sg13g2_decap_8
XFILLER_11_134 VPWR VGND sg13g2_fill_1
X_101_ S2END[2] S2END[3] Inst_S_IO_ConfigMem.Inst_frame0_bit18.Q _017_ VPWR VGND sg13g2_mux2_1
XFILLER_5_22 VPWR VGND sg13g2_fill_2
XFILLER_5_77 VPWR VGND sg13g2_decap_8
X_280_ FrameData[5] FrameData_O[5] VPWR VGND sg13g2_buf_1
X_263_ FrameData[25] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit25.Q VPWR VGND
+ sg13g2_dlhq_1
X_332_ Inst_S_IO_switch_matrix.N2BEG1 N2BEG[1] VPWR VGND sg13g2_buf_1
X_194_ FrameData[20] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit20.Q VPWR VGND
+ sg13g2_dlhq_1
X_246_ FrameData[8] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit8.Q VPWR VGND
+ sg13g2_dlhq_1
X_177_ FrameData[3] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit3.Q VPWR VGND
+ sg13g2_dlhq_1
X_315_ FrameStrobe[8] FrameStrobe_O[8] VPWR VGND sg13g2_buf_1
XFILLER_6_386 VPWR VGND sg13g2_decap_8
X_100_ _016_ VPWR B_I_top VGND _005_ _012_ sg13g2_o21ai_1
XFILLER_7_139 VPWR VGND sg13g2_fill_1
XFILLER_8_22 VPWR VGND sg13g2_fill_2
X_229_ FrameData[23] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit23.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_0_178 VPWR VGND sg13g2_fill_1
XFILLER_0_156 VPWR VGND sg13g2_fill_1
XFILLER_8_234 VPWR VGND sg13g2_decap_8
XFILLER_1_421 VPWR VGND sg13g2_fill_2
XFILLER_5_204 VPWR VGND sg13g2_fill_1
X_193_ FrameData[19] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit19.Q VPWR VGND
+ sg13g2_dlhq_1
X_331_ Inst_S_IO_switch_matrix.N2BEG0 N2BEG[0] VPWR VGND sg13g2_buf_1
X_262_ FrameData[24] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit24.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_9_362 VPWR VGND sg13g2_fill_2
XFILLER_9_351 VPWR VGND sg13g2_decap_8
XFILLER_2_79 VPWR VGND sg13g2_fill_2
X_176_ FrameData[2] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit2.Q VPWR VGND
+ sg13g2_dlhq_1
X_314_ FrameStrobe[7] FrameStrobe_O[7] VPWR VGND sg13g2_buf_1
X_245_ FrameData[7] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit7.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_6_343 VPWR VGND sg13g2_fill_1
XFILLER_11_125 VPWR VGND sg13g2_decap_8
XFILLER_3_324 VPWR VGND sg13g2_fill_2
X_159_ FrameData[17] FrameStrobe[3] Inst_S_IO_switch_matrix.DEBUG_select_N1BEG3[0]
+ VPWR VGND sg13g2_dlhq_1
X_228_ FrameData[22] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit22.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_5_24 VPWR VGND sg13g2_fill_1
X_192_ FrameData[18] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit18.Q VPWR VGND
+ sg13g2_dlhq_1
X_261_ FrameData[23] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit23.Q VPWR VGND
+ sg13g2_dlhq_1
X_330_ Inst_S_IO_switch_matrix.N1BEG3 N1BEG[3] VPWR VGND sg13g2_buf_1
XFILLER_9_0 VPWR VGND sg13g2_decap_8
XFILLER_11_329 VPWR VGND sg13g2_fill_1
X_175_ FrameData[1] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit1.Q VPWR VGND
+ sg13g2_dlhq_1
X_244_ FrameData[6] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit6.Q VPWR VGND
+ sg13g2_dlhq_1
X_313_ FrameStrobe[6] FrameStrobe_O[6] VPWR VGND sg13g2_buf_1
XFILLER_3_347 VPWR VGND sg13g2_decap_8
X_089_ _006_ Inst_S_IO_ConfigMem.Inst_frame0_bit25.Q S2END[5] VPWR VGND sg13g2_nand2_1
XFILLER_8_57 VPWR VGND sg13g2_decap_8
XFILLER_8_24 VPWR VGND sg13g2_fill_1
XFILLER_2_391 VPWR VGND sg13g2_decap_8
X_227_ FrameData[21] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit21.Q VPWR VGND
+ sg13g2_dlhq_1
X_158_ FrameData[16] FrameStrobe[3] Inst_S_IO_switch_matrix.DEBUG_select_N1BEG2[0]
+ VPWR VGND sg13g2_dlhq_1
XFILLER_3_166 VPWR VGND sg13g2_decap_4
XFILLER_8_258 VPWR VGND sg13g2_fill_1
XFILLER_0_147 VPWR VGND sg13g2_decap_8
XFILLER_1_412 VPWR VGND sg13g2_fill_1
XFILLER_1_423 VPWR VGND sg13g2_fill_1
XFILLER_4_272 VPWR VGND sg13g2_fill_2
X_260_ FrameData[22] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit22.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_9_331 VPWR VGND sg13g2_fill_2
XFILLER_2_48 VPWR VGND sg13g2_decap_8
X_191_ FrameData[17] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit17.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_10_396 VPWR VGND sg13g2_decap_4
X_243_ FrameData[5] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit5.Q VPWR VGND
+ sg13g2_dlhq_1
X_312_ FrameStrobe[5] FrameStrobe_O[5] VPWR VGND sg13g2_buf_1
X_174_ FrameData[0] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit0.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_9_194 VPWR VGND sg13g2_fill_2
X_088_ VPWR VGND _004_ Inst_S_IO_ConfigMem.Inst_frame0_bit27.Q _003_ Inst_S_IO_ConfigMem.Inst_frame0_bit26.Q
+ _005_ _002_ sg13g2_a221oi_1
X_157_ FrameData[15] FrameStrobe[3] Inst_S_IO_switch_matrix.DEBUG_select_N1BEG1[0]
+ VPWR VGND sg13g2_dlhq_1
X_226_ FrameData[20] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit20.Q VPWR VGND
+ sg13g2_dlhq_1
X_209_ FrameData[3] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit3.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_4_421 VPWR VGND sg13g2_fill_2
X_190_ FrameData[16] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit16.Q VPWR VGND
+ sg13g2_dlhq_1
X_173_ FrameData[31] FrameStrobe[3] Inst_S_IO_ConfigMem.Inst_frame3_bit31.Q VPWR VGND
+ sg13g2_dlhq_1
X_242_ FrameData[4] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit4.Q VPWR VGND
+ sg13g2_dlhq_1
X_311_ FrameStrobe[4] FrameStrobe_O[4] VPWR VGND sg13g2_buf_1
XFILLER_11_139 VPWR VGND sg13g2_decap_4
XFILLER_3_81 VPWR VGND sg13g2_decap_8
X_156_ FrameData[14] FrameStrobe[3] Inst_S_IO_switch_matrix.DEBUG_select_N1BEG0[0]
+ VPWR VGND sg13g2_dlhq_1
XFILLER_10_161 VPWR VGND sg13g2_fill_2
X_225_ FrameData[19] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit19.Q VPWR VGND
+ sg13g2_dlhq_1
X_087_ VGND VPWR Inst_S_IO_ConfigMem.Inst_frame0_bit25.Q _000_ _004_ Inst_S_IO_ConfigMem.Inst_frame0_bit26.Q
+ sg13g2_a21oi_1
XFILLER_3_113 VPWR VGND sg13g2_fill_2
X_208_ FrameData[2] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit2.Q VPWR VGND
+ sg13g2_dlhq_1
X_139_ Inst_S_IO_ConfigMem.Inst_frame1_bit4.Q S1END[0] S4END[12] SS4END[12] Inst_B_IO_1_bidirectional_frame_config_pass.Q
+ Inst_S_IO_ConfigMem.Inst_frame1_bit5.Q Inst_S_IO_switch_matrix.N4BEG9 VPWR VGND
+ sg13g2_mux4_1
XFILLER_8_227 VPWR VGND sg13g2_decap_8
XFILLER_1_277 VPWR VGND sg13g2_fill_1
XFILLER_1_200 VPWR VGND sg13g2_decap_8
XFILLER_9_333 VPWR VGND sg13g2_fill_1
XFILLER_9_322 VPWR VGND sg13g2_fill_1
X_310_ FrameStrobe[3] FrameStrobe_O[3] VPWR VGND sg13g2_buf_1
X_172_ FrameData[30] FrameStrobe[3] Inst_S_IO_ConfigMem.Inst_frame3_bit30.Q VPWR VGND
+ sg13g2_dlhq_1
X_241_ FrameData[3] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit3.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_6_336 VPWR VGND sg13g2_decap_8
XFILLER_7_0 VPWR VGND sg13g2_decap_8
XFILLER_11_118 VPWR VGND sg13g2_decap_8
X_086_ VGND VPWR _003_ S2END[0] Inst_S_IO_ConfigMem.Inst_frame0_bit25.Q sg13g2_or2_1
X_224_ FrameData[18] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit18.Q VPWR VGND
+ sg13g2_dlhq_1
X_155_ FrameData[13] FrameStrobe[3] B_config_C_bit3 VPWR VGND sg13g2_dlhq_1
XFILLER_0_7 VPWR VGND sg13g2_decap_4
X_138_ Inst_S_IO_ConfigMem.Inst_frame1_bit7.Q S4END[9] SS4END[13] SS4END[9] Inst_A_IO_1_bidirectional_frame_config_pass.Q
+ Inst_S_IO_ConfigMem.Inst_frame1_bit6.Q Inst_S_IO_switch_matrix.N4BEG10 VPWR VGND
+ sg13g2_mux4_1
X_207_ FrameData[1] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit1.Q VPWR VGND
+ sg13g2_dlhq_1
X_069_ _032_ VPWR _033_ VGND S2MID[7] Inst_S_IO_ConfigMem.Inst_frame0_bit24.Q sg13g2_o21ai_1
XFILLER_4_423 VPWR VGND sg13g2_fill_1
X_171_ FrameData[29] FrameStrobe[3] Inst_S_IO_ConfigMem.Inst_frame3_bit29.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_10_355 VPWR VGND sg13g2_fill_2
XFILLER_10_344 VPWR VGND sg13g2_fill_1
XFILLER_10_322 VPWR VGND sg13g2_fill_1
X_240_ FrameData[2] FrameStrobe[0] Inst_S_IO_ConfigMem.Inst_frame0_bit2.Q VPWR VGND
+ sg13g2_dlhq_1
X_369_ Inst_S_IO_switch_matrix.NN4BEG6 NN4BEG[6] VPWR VGND sg13g2_buf_1
XFILLER_3_50 VPWR VGND sg13g2_decap_8
X_223_ FrameData[17] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit17.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_10_163 VPWR VGND sg13g2_fill_1
X_085_ S2END[2] S2END[3] Inst_S_IO_ConfigMem.Inst_frame0_bit25.Q _002_ VPWR VGND sg13g2_mux2_1
X_154_ FrameData[12] FrameStrobe[3] B_config_C_bit2 VPWR VGND sg13g2_dlhq_1
XFILLER_6_112 VPWR VGND sg13g2_decap_8
XFILLER_7_421 VPWR VGND sg13g2_fill_2
XFILLER_7_410 VPWR VGND sg13g2_fill_2
X_068_ _032_ Inst_S_IO_ConfigMem.Inst_frame0_bit24.Q S2END[3] VPWR VGND sg13g2_nand2b_1
X_137_ Inst_S_IO_ConfigMem.Inst_frame1_bit9.Q S4END[8] SS4END[12] SS4END[8] Inst_B_IO_1_bidirectional_frame_config_pass.Q
+ Inst_S_IO_ConfigMem.Inst_frame1_bit8.Q Inst_S_IO_switch_matrix.N4BEG11 VPWR VGND
+ sg13g2_mux4_1
X_206_ FrameData[0] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit0.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_4_402 VPWR VGND sg13g2_decap_8
XFILLER_4_221 VPWR VGND sg13g2_decap_8
X_170_ FrameData[28] FrameStrobe[3] Inst_S_IO_ConfigMem.Inst_frame3_bit28.Q VPWR VGND
+ sg13g2_dlhq_1
X_368_ Inst_S_IO_switch_matrix.NN4BEG5 NN4BEG[5] VPWR VGND sg13g2_buf_1
X_299_ FrameData[24] FrameData_O[24] VPWR VGND sg13g2_buf_1
XFILLER_10_120 VPWR VGND sg13g2_fill_2
X_153_ FrameData[11] FrameStrobe[3] B_config_C_bit1 VPWR VGND sg13g2_dlhq_1
X_084_ VPWR _001_ Inst_S_IO_ConfigMem.Inst_frame0_bit24.Q VGND sg13g2_inv_1
X_222_ FrameData[16] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit16.Q VPWR VGND
+ sg13g2_dlhq_1
X_205_ FrameData[31] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit31.Q VPWR VGND
+ sg13g2_dlhq_1
X_136_ Inst_S_IO_ConfigMem.Inst_frame1_bit11.Q S1END[1] SS4END[5] S4END[5] Inst_A_IO_1_bidirectional_frame_config_pass.Q
+ Inst_S_IO_ConfigMem.Inst_frame1_bit10.Q Inst_S_IO_switch_matrix.N4BEG12 VPWR VGND
+ sg13g2_mux4_1
X_067_ S1END[3] A_O_top Inst_S_IO_switch_matrix.DEBUG_select_N1BEG0[0] Inst_S_IO_switch_matrix.N1BEG0
+ VPWR VGND sg13g2_mux2_1
XFILLER_9_83 VPWR VGND sg13g2_fill_2
XFILLER_0_41 VPWR VGND sg13g2_decap_8
XFILLER_0_30 VPWR VGND sg13g2_fill_1
XFILLER_11_292 VPWR VGND sg13g2_decap_4
X_119_ Inst_S_IO_ConfigMem.Inst_frame0_bit12.Q S4END[7] S4END[9] S4END[11] Inst_B_IO_1_bidirectional_frame_config_pass.Q
+ Inst_S_IO_ConfigMem.Inst_frame0_bit13.Q Inst_S_IO_switch_matrix.NN4BEG13 VPWR VGND
+ sg13g2_mux4_1
XFILLER_9_358 VPWR VGND sg13g2_decap_4
XFILLER_10_357 VPWR VGND sg13g2_fill_1
X_298_ FrameData[23] FrameData_O[23] VPWR VGND sg13g2_buf_1
X_367_ Inst_S_IO_switch_matrix.NN4BEG4 NN4BEG[4] VPWR VGND sg13g2_buf_1
XFILLER_3_74 VPWR VGND sg13g2_decap_8
X_221_ FrameData[15] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit15.Q VPWR VGND
+ sg13g2_dlhq_1
X_152_ FrameData[10] FrameStrobe[3] B_config_C_bit0 VPWR VGND sg13g2_dlhq_1
XFILLER_5_0 VPWR VGND sg13g2_decap_4
X_083_ VPWR _000_ S2END[1] VGND sg13g2_inv_1
X_204_ FrameData[30] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit30.Q VPWR VGND
+ sg13g2_dlhq_1
X_066_ S1END[2] Inst_A_IO_1_bidirectional_frame_config_pass.Q Inst_S_IO_switch_matrix.DEBUG_select_N1BEG1[0]
+ Inst_S_IO_switch_matrix.N1BEG1 VPWR VGND sg13g2_mux2_1
XFILLER_7_423 VPWR VGND sg13g2_fill_1
XFILLER_7_412 VPWR VGND sg13g2_fill_1
X_135_ Inst_S_IO_ConfigMem.Inst_frame1_bit13.Q S1END[0] SS4END[4] S4END[4] Inst_B_IO_1_bidirectional_frame_config_pass.Q
+ Inst_S_IO_ConfigMem.Inst_frame1_bit12.Q Inst_S_IO_switch_matrix.N4BEG13 VPWR VGND
+ sg13g2_mux4_1
XFILLER_8_209 VPWR VGND sg13g2_fill_1
X_049_ Inst_S_IO_ConfigMem.Inst_frame2_bit14.Q S2END[1] S4END[1] SS4END[1] SS4END[9]
+ Inst_S_IO_ConfigMem.Inst_frame2_bit15.Q Inst_S_IO_switch_matrix.N2BEGb6 VPWR VGND
+ sg13g2_mux4_1
X_118_ Inst_S_IO_ConfigMem.Inst_frame0_bit15.Q S2MID[0] S2MID[4] S2MID[2] S2MID[6]
+ Inst_S_IO_ConfigMem.Inst_frame0_bit14.Q Inst_S_IO_switch_matrix.NN4BEG14 VPWR VGND
+ sg13g2_mux4_1
XFILLER_7_264 VPWR VGND sg13g2_decap_4
XFILLER_6_30 VPWR VGND sg13g2_fill_1
XFILLER_0_292 VPWR VGND sg13g2_fill_2
X_366_ Inst_S_IO_switch_matrix.NN4BEG3 NN4BEG[3] VPWR VGND sg13g2_buf_1
XFILLER_9_167 VPWR VGND sg13g2_fill_2
X_297_ FrameData[22] FrameData_O[22] VPWR VGND sg13g2_buf_1
XFILLER_5_362 VPWR VGND sg13g2_decap_8
XFILLER_5_373 VPWR VGND sg13g2_fill_2
X_220_ FrameData[14] FrameStrobe[1] Inst_S_IO_ConfigMem.Inst_frame1_bit14.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_10_122 VPWR VGND sg13g2_fill_1
X_151_ FrameData[9] FrameStrobe[3] A_config_C_bit3 VPWR VGND sg13g2_dlhq_1
XFILLER_2_332 VPWR VGND sg13g2_decap_4
XFILLER_2_398 VPWR VGND sg13g2_decap_8
X_082_ _044_ VPWR B_T_top VGND Inst_S_IO_ConfigMem.Inst_frame0_bit31.Q _041_ sg13g2_o21ai_1
X_349_ Inst_S_IO_switch_matrix.N4BEG2 N4BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_5_170 VPWR VGND sg13g2_decap_8
X_134_ Inst_S_IO_ConfigMem.Inst_frame1_bit14.Q S4END[1] SS4END[1] SS4END[13] Inst_A_IO_1_bidirectional_frame_config_pass.Q
+ Inst_S_IO_ConfigMem.Inst_frame1_bit15.Q Inst_S_IO_switch_matrix.N4BEG14 VPWR VGND
+ sg13g2_mux4_1
X_203_ FrameData[29] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit29.Q VPWR VGND
+ sg13g2_dlhq_1
X_065_ S1END[1] B_O_top Inst_S_IO_switch_matrix.DEBUG_select_N1BEG2[0] Inst_S_IO_switch_matrix.N1BEG2
+ VPWR VGND sg13g2_mux2_1
XFILLER_9_41 VPWR VGND sg13g2_fill_2
Xclkbuf_0_UserCLK UserCLK clknet_0_UserCLK VPWR VGND sg13g2_buf_8
XFILLER_7_232 VPWR VGND sg13g2_decap_4
X_117_ Inst_S_IO_ConfigMem.Inst_frame0_bit17.Q S2MID[1] S2MID[5] S2MID[3] S2MID[7]
+ Inst_S_IO_ConfigMem.Inst_frame0_bit16.Q Inst_S_IO_switch_matrix.NN4BEG15 VPWR VGND
+ sg13g2_mux4_1
X_048_ Inst_S_IO_ConfigMem.Inst_frame2_bit16.Q S2END[0] S4END[0] SS4END[0] SS4END[8]
+ Inst_S_IO_ConfigMem.Inst_frame2_bit17.Q Inst_S_IO_switch_matrix.N2BEGb7 VPWR VGND
+ sg13g2_mux4_1
XFILLER_8_382 VPWR VGND sg13g2_decap_8
X_296_ FrameData[21] FrameData_O[21] VPWR VGND sg13g2_buf_1
X_365_ Inst_S_IO_switch_matrix.NN4BEG2 NN4BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_6_308 VPWR VGND sg13g2_decap_8
XFILLER_3_21 VPWR VGND sg13g2_decap_4
XFILLER_3_43 VPWR VGND sg13g2_decap_8
X_081_ _044_ _042_ _043_ VPWR VGND sg13g2_nand2b_1
X_150_ FrameData[8] FrameStrobe[3] A_config_C_bit2 VPWR VGND sg13g2_dlhq_1
XFILLER_6_105 VPWR VGND sg13g2_decap_8
X_348_ Inst_S_IO_switch_matrix.N4BEG1 N4BEG[1] VPWR VGND sg13g2_buf_1
X_279_ FrameData[4] FrameData_O[4] VPWR VGND sg13g2_buf_1
XFILLER_2_355 VPWR VGND sg13g2_fill_2
XFILLER_11_421 VPWR VGND sg13g2_fill_2
XFILLER_11_410 VPWR VGND sg13g2_fill_2
X_202_ FrameData[28] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit28.Q VPWR VGND
+ sg13g2_dlhq_1
X_133_ Inst_S_IO_ConfigMem.Inst_frame1_bit16.Q S4END[0] SS4END[0] SS4END[12] Inst_B_IO_1_bidirectional_frame_config_pass.Q
+ Inst_S_IO_ConfigMem.Inst_frame1_bit17.Q Inst_S_IO_switch_matrix.N4BEG15 VPWR VGND
+ sg13g2_mux4_1
XFILLER_0_11 VPWR VGND sg13g2_fill_2
X_064_ S1END[0] Inst_B_IO_1_bidirectional_frame_config_pass.Q Inst_S_IO_switch_matrix.DEBUG_select_N1BEG3[0]
+ Inst_S_IO_switch_matrix.N1BEG3 VPWR VGND sg13g2_mux2_1
X_047_ Inst_S_IO_ConfigMem.Inst_frame2_bit18.Q S1END[2] S4END[15] SS4END[15] A_O_top
+ Inst_S_IO_ConfigMem.Inst_frame2_bit19.Q Inst_S_IO_switch_matrix.N4BEG0 VPWR VGND
+ sg13g2_mux4_1
X_116_ _031_ VPWR A_I_top VGND _020_ _027_ sg13g2_o21ai_1
XFILLER_4_214 VPWR VGND sg13g2_decap_8
XFILLER_6_21 VPWR VGND sg13g2_decap_8
XFILLER_3_291 VPWR VGND sg13g2_fill_2
X_295_ FrameData[20] FrameData_O[20] VPWR VGND sg13g2_buf_1
X_364_ Inst_S_IO_switch_matrix.NN4BEG1 NN4BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_5_320 VPWR VGND sg13g2_fill_1
X_080_ Inst_S_IO_ConfigMem.Inst_frame0_bit31.Q VPWR _043_ VGND Inst_S_IO_ConfigMem.Inst_frame0_bit29.Q
+ _040_ sg13g2_o21ai_1
X_347_ Inst_S_IO_switch_matrix.N4BEG0 N4BEG[0] VPWR VGND sg13g2_buf_1
X_278_ FrameData[3] FrameData_O[3] VPWR VGND sg13g2_buf_1
XFILLER_3_109 VPWR VGND sg13g2_decap_4
X_201_ FrameData[27] FrameStrobe[2] Inst_S_IO_ConfigMem.Inst_frame2_bit27.Q VPWR VGND
+ sg13g2_dlhq_1
X_132_ Inst_S_IO_ConfigMem.Inst_frame1_bit18.Q S4END[0] S4END[2] S4END[4] A_O_top
+ Inst_S_IO_ConfigMem.Inst_frame1_bit19.Q Inst_S_IO_switch_matrix.NN4BEG0 VPWR VGND
+ sg13g2_mux4_1
XFILLER_3_0 VPWR VGND sg13g2_decap_4
X_063_ Inst_S_IO_ConfigMem.Inst_frame3_bit18.Q S2MID[7] S4END[7] SS4END[7] SS4END[15]
+ Inst_S_IO_ConfigMem.Inst_frame3_bit19.Q Inst_S_IO_switch_matrix.N2BEG0 VPWR VGND
+ sg13g2_mux4_1
XFILLER_9_76 VPWR VGND sg13g2_decap_8
XFILLER_11_285 VPWR VGND sg13g2_decap_8
X_115_ _031_ _030_ Inst_S_IO_ConfigMem.Inst_frame0_bit21.Q VPWR VGND sg13g2_nand2b_1
XFILLER_0_421 VPWR VGND sg13g2_fill_2
XFILLER_9_318 VPWR VGND sg13g2_decap_4
XFILLER_1_207 VPWR VGND sg13g2_fill_2
XFILLER_0_273 VPWR VGND sg13g2_fill_2
XFILLER_0_251 VPWR VGND sg13g2_fill_1
.ends

