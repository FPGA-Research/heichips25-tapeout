VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO S_IO4
  CLASS BLOCK ;
  FOREIGN S_IO4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 215.040 BY 53.760 ;
  PIN A_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 20.440 0.000 20.840 0.400 ;
    END
  END A_I_top
  PIN A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 14.680 0.000 15.080 0.400 ;
    END
  END A_O_top
  PIN A_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 26.200 0.000 26.600 0.400 ;
    END
  END A_T_top
  PIN B_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 37.720 0.000 38.120 0.400 ;
    END
  END B_I_top
  PIN B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 31.960 0.000 32.360 0.400 ;
    END
  END B_O_top
  PIN B_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 43.480 0.000 43.880 0.400 ;
    END
  END B_T_top
  PIN C_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.615900 ;
    PORT
      LAYER Metal2 ;
        RECT 55.000 0.000 55.400 0.400 ;
    END
  END C_I_top
  PIN C_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 49.240 0.000 49.640 0.400 ;
    END
  END C_O_top
  PIN C_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 60.760 0.000 61.160 0.400 ;
    END
  END C_T_top
  PIN Co
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.299200 ;
    PORT
      LAYER Metal2 ;
        RECT 97.240 53.360 97.640 53.760 ;
    END
  END Co
  PIN D_I_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 72.280 0.000 72.680 0.400 ;
    END
  END D_I_top
  PIN D_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.601600 ;
    PORT
      LAYER Metal2 ;
        RECT 66.520 0.000 66.920 0.400 ;
    END
  END D_O_top
  PIN D_T_top
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal2 ;
        RECT 78.040 0.000 78.440 0.400 ;
    END
  END D_T_top
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.903500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 0.220 0.400 0.620 ;
    END
  END FrameData[0]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.903500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 17.020 0.400 17.420 ;
    END
  END FrameData[10]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.903500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 18.700 0.400 19.100 ;
    END
  END FrameData[11]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.903500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 20.380 0.400 20.780 ;
    END
  END FrameData[12]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.903500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 22.060 0.400 22.460 ;
    END
  END FrameData[13]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.903500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 23.740 0.400 24.140 ;
    END
  END FrameData[14]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.903500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 25.420 0.400 25.820 ;
    END
  END FrameData[15]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.903500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 27.100 0.400 27.500 ;
    END
  END FrameData[16]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.903500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 28.780 0.400 29.180 ;
    END
  END FrameData[17]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.903500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 30.460 0.400 30.860 ;
    END
  END FrameData[18]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.903500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 32.140 0.400 32.540 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.903500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1.900 0.400 2.300 ;
    END
  END FrameData[1]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.903500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 33.820 0.400 34.220 ;
    END
  END FrameData[20]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.903500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 35.500 0.400 35.900 ;
    END
  END FrameData[21]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.903500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 37.180 0.400 37.580 ;
    END
  END FrameData[22]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.903500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 38.860 0.400 39.260 ;
    END
  END FrameData[23]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.903500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 40.540 0.400 40.940 ;
    END
  END FrameData[24]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.903500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 42.220 0.400 42.620 ;
    END
  END FrameData[25]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.903500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 43.900 0.400 44.300 ;
    END
  END FrameData[26]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.903500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 45.580 0.400 45.980 ;
    END
  END FrameData[27]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.084200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 47.260 0.400 47.660 ;
    END
  END FrameData[28]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.084200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 48.940 0.400 49.340 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.903500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3.580 0.400 3.980 ;
    END
  END FrameData[2]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.084200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 50.620 0.400 51.020 ;
    END
  END FrameData[30]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.084200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 52.300 0.400 52.700 ;
    END
  END FrameData[31]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.903500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 5.260 0.400 5.660 ;
    END
  END FrameData[3]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.903500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 6.940 0.400 7.340 ;
    END
  END FrameData[4]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.903500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 8.620 0.400 9.020 ;
    END
  END FrameData[5]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.903500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 10.300 0.400 10.700 ;
    END
  END FrameData[6]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.903500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 11.980 0.400 12.380 ;
    END
  END FrameData[7]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.903500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 13.660 0.400 14.060 ;
    END
  END FrameData[8]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.903500 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 15.340 0.400 15.740 ;
    END
  END FrameData[9]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 0.220 215.040 0.620 ;
    END
  END FrameData_O[0]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 17.020 215.040 17.420 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 18.700 215.040 19.100 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 20.380 215.040 20.780 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 22.060 215.040 22.460 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 23.740 215.040 24.140 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 25.420 215.040 25.820 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 27.100 215.040 27.500 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 28.780 215.040 29.180 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 30.460 215.040 30.860 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 32.140 215.040 32.540 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 1.900 215.040 2.300 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 33.820 215.040 34.220 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 35.500 215.040 35.900 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 37.180 215.040 37.580 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 38.860 215.040 39.260 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 40.540 215.040 40.940 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 42.220 215.040 42.620 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 43.900 215.040 44.300 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 45.580 215.040 45.980 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 47.260 215.040 47.660 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 48.940 215.040 49.340 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 3.580 215.040 3.980 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 50.620 215.040 51.020 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 52.300 215.040 52.700 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 5.260 215.040 5.660 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 6.940 215.040 7.340 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 8.620 215.040 9.020 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 10.300 215.040 10.700 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 11.980 215.040 12.380 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 13.660 215.040 14.060 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 214.640 15.340 215.040 15.740 ;
    END
  END FrameData_O[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.753500 ;
    PORT
      LAYER Metal2 ;
        RECT 89.560 0.000 89.960 0.400 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 147.160 0.000 147.560 0.400 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 152.920 0.000 153.320 0.400 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 158.680 0.000 159.080 0.400 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 164.440 0.000 164.840 0.400 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 170.200 0.000 170.600 0.400 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 175.960 0.000 176.360 0.400 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 181.720 0.000 182.120 0.400 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 187.480 0.000 187.880 0.400 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 193.240 0.000 193.640 0.400 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 199.000 0.000 199.400 0.400 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.753500 ;
    PORT
      LAYER Metal2 ;
        RECT 95.320 0.000 95.720 0.400 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.753500 ;
    PORT
      LAYER Metal2 ;
        RECT 101.080 0.000 101.480 0.400 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.753500 ;
    PORT
      LAYER Metal2 ;
        RECT 106.840 0.000 107.240 0.400 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.002300 ;
    PORT
      LAYER Metal2 ;
        RECT 112.600 0.000 113.000 0.400 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 118.360 0.000 118.760 0.400 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 124.120 0.000 124.520 0.400 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 129.880 0.000 130.280 0.400 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 135.640 0.000 136.040 0.400 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 141.400 0.000 141.800 0.400 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 149.080 53.360 149.480 53.760 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 158.680 53.360 159.080 53.760 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 159.640 53.360 160.040 53.760 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 160.600 53.360 161.000 53.760 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 161.560 53.360 161.960 53.760 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 162.520 53.360 162.920 53.760 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 163.480 53.360 163.880 53.760 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 164.440 53.360 164.840 53.760 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 165.400 53.360 165.800 53.760 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 166.360 53.360 166.760 53.760 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 167.320 53.360 167.720 53.760 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 150.040 53.360 150.440 53.760 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 151.000 53.360 151.400 53.760 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 151.960 53.360 152.360 53.760 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 152.920 53.360 153.320 53.760 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 153.880 53.360 154.280 53.760 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 154.840 53.360 155.240 53.760 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 155.800 53.360 156.200 53.760 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 156.760 53.360 157.160 53.760 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 157.720 53.360 158.120 53.760 ;
    END
  END FrameStrobe_O[9]
  PIN N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 47.320 53.360 47.720 53.760 ;
    END
  END N1BEG[0]
  PIN N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 48.280 53.360 48.680 53.760 ;
    END
  END N1BEG[1]
  PIN N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 49.240 53.360 49.640 53.760 ;
    END
  END N1BEG[2]
  PIN N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 50.200 53.360 50.600 53.760 ;
    END
  END N1BEG[3]
  PIN N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 51.160 53.360 51.560 53.760 ;
    END
  END N2BEG[0]
  PIN N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 52.120 53.360 52.520 53.760 ;
    END
  END N2BEG[1]
  PIN N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 53.080 53.360 53.480 53.760 ;
    END
  END N2BEG[2]
  PIN N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 54.040 53.360 54.440 53.760 ;
    END
  END N2BEG[3]
  PIN N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 55.000 53.360 55.400 53.760 ;
    END
  END N2BEG[4]
  PIN N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 55.960 53.360 56.360 53.760 ;
    END
  END N2BEG[5]
  PIN N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 56.920 53.360 57.320 53.760 ;
    END
  END N2BEG[6]
  PIN N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 57.880 53.360 58.280 53.760 ;
    END
  END N2BEG[7]
  PIN N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 58.840 53.360 59.240 53.760 ;
    END
  END N2BEGb[0]
  PIN N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 59.800 53.360 60.200 53.760 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 60.760 53.360 61.160 53.760 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 61.720 53.360 62.120 53.760 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 62.680 53.360 63.080 53.760 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 63.640 53.360 64.040 53.760 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 64.600 53.360 65.000 53.760 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 65.560 53.360 65.960 53.760 ;
    END
  END N2BEGb[7]
  PIN N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 66.520 53.360 66.920 53.760 ;
    END
  END N4BEG[0]
  PIN N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 76.120 53.360 76.520 53.760 ;
    END
  END N4BEG[10]
  PIN N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 77.080 53.360 77.480 53.760 ;
    END
  END N4BEG[11]
  PIN N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 78.040 53.360 78.440 53.760 ;
    END
  END N4BEG[12]
  PIN N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 79.000 53.360 79.400 53.760 ;
    END
  END N4BEG[13]
  PIN N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 79.960 53.360 80.360 53.760 ;
    END
  END N4BEG[14]
  PIN N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 80.920 53.360 81.320 53.760 ;
    END
  END N4BEG[15]
  PIN N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 67.480 53.360 67.880 53.760 ;
    END
  END N4BEG[1]
  PIN N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 68.440 53.360 68.840 53.760 ;
    END
  END N4BEG[2]
  PIN N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 69.400 53.360 69.800 53.760 ;
    END
  END N4BEG[3]
  PIN N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 70.360 53.360 70.760 53.760 ;
    END
  END N4BEG[4]
  PIN N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 71.320 53.360 71.720 53.760 ;
    END
  END N4BEG[5]
  PIN N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 72.280 53.360 72.680 53.760 ;
    END
  END N4BEG[6]
  PIN N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 73.240 53.360 73.640 53.760 ;
    END
  END N4BEG[7]
  PIN N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 74.200 53.360 74.600 53.760 ;
    END
  END N4BEG[8]
  PIN N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 75.160 53.360 75.560 53.760 ;
    END
  END N4BEG[9]
  PIN NN4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 81.880 53.360 82.280 53.760 ;
    END
  END NN4BEG[0]
  PIN NN4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 91.480 53.360 91.880 53.760 ;
    END
  END NN4BEG[10]
  PIN NN4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 92.440 53.360 92.840 53.760 ;
    END
  END NN4BEG[11]
  PIN NN4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 93.400 53.360 93.800 53.760 ;
    END
  END NN4BEG[12]
  PIN NN4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 94.360 53.360 94.760 53.760 ;
    END
  END NN4BEG[13]
  PIN NN4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 95.320 53.360 95.720 53.760 ;
    END
  END NN4BEG[14]
  PIN NN4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 96.280 53.360 96.680 53.760 ;
    END
  END NN4BEG[15]
  PIN NN4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 82.840 53.360 83.240 53.760 ;
    END
  END NN4BEG[1]
  PIN NN4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 83.800 53.360 84.200 53.760 ;
    END
  END NN4BEG[2]
  PIN NN4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 84.760 53.360 85.160 53.760 ;
    END
  END NN4BEG[3]
  PIN NN4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 85.720 53.360 86.120 53.760 ;
    END
  END NN4BEG[4]
  PIN NN4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 86.680 53.360 87.080 53.760 ;
    END
  END NN4BEG[5]
  PIN NN4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 87.640 53.360 88.040 53.760 ;
    END
  END NN4BEG[6]
  PIN NN4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 88.600 53.360 89.000 53.760 ;
    END
  END NN4BEG[7]
  PIN NN4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 89.560 53.360 89.960 53.760 ;
    END
  END NN4BEG[8]
  PIN NN4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 90.520 53.360 90.920 53.760 ;
    END
  END NN4BEG[9]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal2 ;
        RECT 98.200 53.360 98.600 53.760 ;
    END
  END S1END[0]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal2 ;
        RECT 99.160 53.360 99.560 53.760 ;
    END
  END S1END[1]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal2 ;
        RECT 100.120 53.360 100.520 53.760 ;
    END
  END S1END[2]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal2 ;
        RECT 101.080 53.360 101.480 53.760 ;
    END
  END S1END[3]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.080000 ;
    PORT
      LAYER Metal2 ;
        RECT 109.720 53.360 110.120 53.760 ;
    END
  END S2END[0]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.320800 ;
    PORT
      LAYER Metal2 ;
        RECT 110.680 53.360 111.080 53.760 ;
    END
  END S2END[1]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.531400 ;
    PORT
      LAYER Metal2 ;
        RECT 111.640 53.360 112.040 53.760 ;
    END
  END S2END[2]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.560000 ;
    PORT
      LAYER Metal2 ;
        RECT 112.600 53.360 113.000 53.760 ;
    END
  END S2END[3]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.281000 ;
    PORT
      LAYER Metal2 ;
        RECT 113.560 53.360 113.960 53.760 ;
    END
  END S2END[4]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.087800 ;
    PORT
      LAYER Metal2 ;
        RECT 114.520 53.360 114.920 53.760 ;
    END
  END S2END[5]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.326600 ;
    PORT
      LAYER Metal2 ;
        RECT 115.480 53.360 115.880 53.760 ;
    END
  END S2END[6]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.378000 ;
    PORT
      LAYER Metal2 ;
        RECT 116.440 53.360 116.840 53.760 ;
    END
  END S2END[7]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.292200 ;
    PORT
      LAYER Metal2 ;
        RECT 102.040 53.360 102.440 53.760 ;
    END
  END S2MID[0]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.292200 ;
    PORT
      LAYER Metal2 ;
        RECT 103.000 53.360 103.400 53.760 ;
    END
  END S2MID[1]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.505400 ;
    PORT
      LAYER Metal2 ;
        RECT 103.960 53.360 104.360 53.760 ;
    END
  END S2MID[2]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.505400 ;
    PORT
      LAYER Metal2 ;
        RECT 104.920 53.360 105.320 53.760 ;
    END
  END S2MID[3]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.505400 ;
    PORT
      LAYER Metal2 ;
        RECT 105.880 53.360 106.280 53.760 ;
    END
  END S2MID[4]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.505400 ;
    PORT
      LAYER Metal2 ;
        RECT 106.840 53.360 107.240 53.760 ;
    END
  END S2MID[5]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.931800 ;
    PORT
      LAYER Metal2 ;
        RECT 107.800 53.360 108.200 53.760 ;
    END
  END S2MID[6]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.145000 ;
    PORT
      LAYER Metal2 ;
        RECT 108.760 53.360 109.160 53.760 ;
    END
  END S2MID[7]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal2 ;
        RECT 117.400 53.360 117.800 53.760 ;
    END
  END S4END[0]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal2 ;
        RECT 127.000 53.360 127.400 53.760 ;
    END
  END S4END[10]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.639600 ;
    PORT
      LAYER Metal2 ;
        RECT 127.960 53.360 128.360 53.760 ;
    END
  END S4END[11]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 128.920 53.360 129.320 53.760 ;
    END
  END S4END[12]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 129.880 53.360 130.280 53.760 ;
    END
  END S4END[13]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 130.840 53.360 131.240 53.760 ;
    END
  END S4END[14]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 131.800 53.360 132.200 53.760 ;
    END
  END S4END[15]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal2 ;
        RECT 118.360 53.360 118.760 53.760 ;
    END
  END S4END[1]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal2 ;
        RECT 119.320 53.360 119.720 53.760 ;
    END
  END S4END[2]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal2 ;
        RECT 120.280 53.360 120.680 53.760 ;
    END
  END S4END[3]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal2 ;
        RECT 121.240 53.360 121.640 53.760 ;
    END
  END S4END[4]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal2 ;
        RECT 122.200 53.360 122.600 53.760 ;
    END
  END S4END[5]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal2 ;
        RECT 123.160 53.360 123.560 53.760 ;
    END
  END S4END[6]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal2 ;
        RECT 124.120 53.360 124.520 53.760 ;
    END
  END S4END[7]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal2 ;
        RECT 125.080 53.360 125.480 53.760 ;
    END
  END S4END[8]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.639600 ;
    PORT
      LAYER Metal2 ;
        RECT 126.040 53.360 126.440 53.760 ;
    END
  END S4END[9]
  PIN SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.639600 ;
    PORT
      LAYER Metal2 ;
        RECT 132.760 53.360 133.160 53.760 ;
    END
  END SS4END[0]
  PIN SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.639600 ;
    PORT
      LAYER Metal2 ;
        RECT 142.360 53.360 142.760 53.760 ;
    END
  END SS4END[10]
  PIN SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.639600 ;
    PORT
      LAYER Metal2 ;
        RECT 143.320 53.360 143.720 53.760 ;
    END
  END SS4END[11]
  PIN SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.639600 ;
    PORT
      LAYER Metal2 ;
        RECT 144.280 53.360 144.680 53.760 ;
    END
  END SS4END[12]
  PIN SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.639600 ;
    PORT
      LAYER Metal2 ;
        RECT 145.240 53.360 145.640 53.760 ;
    END
  END SS4END[13]
  PIN SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.639600 ;
    PORT
      LAYER Metal2 ;
        RECT 146.200 53.360 146.600 53.760 ;
    END
  END SS4END[14]
  PIN SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.639600 ;
    PORT
      LAYER Metal2 ;
        RECT 147.160 53.360 147.560 53.760 ;
    END
  END SS4END[15]
  PIN SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.639600 ;
    PORT
      LAYER Metal2 ;
        RECT 133.720 53.360 134.120 53.760 ;
    END
  END SS4END[1]
  PIN SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.639600 ;
    PORT
      LAYER Metal2 ;
        RECT 134.680 53.360 135.080 53.760 ;
    END
  END SS4END[2]
  PIN SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.639600 ;
    PORT
      LAYER Metal2 ;
        RECT 135.640 53.360 136.040 53.760 ;
    END
  END SS4END[3]
  PIN SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.639600 ;
    PORT
      LAYER Metal2 ;
        RECT 136.600 53.360 137.000 53.760 ;
    END
  END SS4END[4]
  PIN SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.639600 ;
    PORT
      LAYER Metal2 ;
        RECT 137.560 53.360 137.960 53.760 ;
    END
  END SS4END[5]
  PIN SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.639600 ;
    PORT
      LAYER Metal2 ;
        RECT 138.520 53.360 138.920 53.760 ;
    END
  END SS4END[6]
  PIN SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.639600 ;
    PORT
      LAYER Metal2 ;
        RECT 139.480 53.360 139.880 53.760 ;
    END
  END SS4END[7]
  PIN SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.639600 ;
    PORT
      LAYER Metal2 ;
        RECT 140.440 53.360 140.840 53.760 ;
    END
  END SS4END[8]
  PIN SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.639600 ;
    PORT
      LAYER Metal2 ;
        RECT 141.400 53.360 141.800 53.760 ;
    END
  END SS4END[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.450800 ;
    PORT
      LAYER Metal2 ;
        RECT 83.800 0.000 84.200 0.400 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 148.120 53.360 148.520 53.760 ;
    END
  END UserCLKo
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER TopMetal1 ;
        RECT 24.460 0.000 26.660 53.760 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 100.060 0.000 102.260 53.760 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 175.660 0.000 177.860 53.760 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER TopMetal1 ;
        RECT 18.260 0.000 20.460 53.760 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 93.860 0.000 96.060 53.760 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 169.460 0.000 171.660 53.760 ;
    END
  END VPWR
  OBS
      LAYER GatPoly ;
        RECT 5.760 3.630 209.280 49.290 ;
      LAYER Metal1 ;
        RECT 5.760 3.560 209.280 49.360 ;
      LAYER Metal2 ;
        RECT 5.655 53.150 47.110 53.485 ;
        RECT 47.930 53.150 48.070 53.485 ;
        RECT 48.890 53.150 49.030 53.485 ;
        RECT 49.850 53.150 49.990 53.485 ;
        RECT 50.810 53.150 50.950 53.485 ;
        RECT 51.770 53.150 51.910 53.485 ;
        RECT 52.730 53.150 52.870 53.485 ;
        RECT 53.690 53.150 53.830 53.485 ;
        RECT 54.650 53.150 54.790 53.485 ;
        RECT 55.610 53.150 55.750 53.485 ;
        RECT 56.570 53.150 56.710 53.485 ;
        RECT 57.530 53.150 57.670 53.485 ;
        RECT 58.490 53.150 58.630 53.485 ;
        RECT 59.450 53.150 59.590 53.485 ;
        RECT 60.410 53.150 60.550 53.485 ;
        RECT 61.370 53.150 61.510 53.485 ;
        RECT 62.330 53.150 62.470 53.485 ;
        RECT 63.290 53.150 63.430 53.485 ;
        RECT 64.250 53.150 64.390 53.485 ;
        RECT 65.210 53.150 65.350 53.485 ;
        RECT 66.170 53.150 66.310 53.485 ;
        RECT 67.130 53.150 67.270 53.485 ;
        RECT 68.090 53.150 68.230 53.485 ;
        RECT 69.050 53.150 69.190 53.485 ;
        RECT 70.010 53.150 70.150 53.485 ;
        RECT 70.970 53.150 71.110 53.485 ;
        RECT 71.930 53.150 72.070 53.485 ;
        RECT 72.890 53.150 73.030 53.485 ;
        RECT 73.850 53.150 73.990 53.485 ;
        RECT 74.810 53.150 74.950 53.485 ;
        RECT 75.770 53.150 75.910 53.485 ;
        RECT 76.730 53.150 76.870 53.485 ;
        RECT 77.690 53.150 77.830 53.485 ;
        RECT 78.650 53.150 78.790 53.485 ;
        RECT 79.610 53.150 79.750 53.485 ;
        RECT 80.570 53.150 80.710 53.485 ;
        RECT 81.530 53.150 81.670 53.485 ;
        RECT 82.490 53.150 82.630 53.485 ;
        RECT 83.450 53.150 83.590 53.485 ;
        RECT 84.410 53.150 84.550 53.485 ;
        RECT 85.370 53.150 85.510 53.485 ;
        RECT 86.330 53.150 86.470 53.485 ;
        RECT 87.290 53.150 87.430 53.485 ;
        RECT 88.250 53.150 88.390 53.485 ;
        RECT 89.210 53.150 89.350 53.485 ;
        RECT 90.170 53.150 90.310 53.485 ;
        RECT 91.130 53.150 91.270 53.485 ;
        RECT 92.090 53.150 92.230 53.485 ;
        RECT 93.050 53.150 93.190 53.485 ;
        RECT 94.010 53.150 94.150 53.485 ;
        RECT 94.970 53.150 95.110 53.485 ;
        RECT 95.930 53.150 96.070 53.485 ;
        RECT 96.890 53.150 97.030 53.485 ;
        RECT 97.850 53.150 97.990 53.485 ;
        RECT 98.810 53.150 98.950 53.485 ;
        RECT 99.770 53.150 99.910 53.485 ;
        RECT 100.730 53.150 100.870 53.485 ;
        RECT 101.690 53.150 101.830 53.485 ;
        RECT 102.650 53.150 102.790 53.485 ;
        RECT 103.610 53.150 103.750 53.485 ;
        RECT 104.570 53.150 104.710 53.485 ;
        RECT 105.530 53.150 105.670 53.485 ;
        RECT 106.490 53.150 106.630 53.485 ;
        RECT 107.450 53.150 107.590 53.485 ;
        RECT 108.410 53.150 108.550 53.485 ;
        RECT 109.370 53.150 109.510 53.485 ;
        RECT 110.330 53.150 110.470 53.485 ;
        RECT 111.290 53.150 111.430 53.485 ;
        RECT 112.250 53.150 112.390 53.485 ;
        RECT 113.210 53.150 113.350 53.485 ;
        RECT 114.170 53.150 114.310 53.485 ;
        RECT 115.130 53.150 115.270 53.485 ;
        RECT 116.090 53.150 116.230 53.485 ;
        RECT 117.050 53.150 117.190 53.485 ;
        RECT 118.010 53.150 118.150 53.485 ;
        RECT 118.970 53.150 119.110 53.485 ;
        RECT 119.930 53.150 120.070 53.485 ;
        RECT 120.890 53.150 121.030 53.485 ;
        RECT 121.850 53.150 121.990 53.485 ;
        RECT 122.810 53.150 122.950 53.485 ;
        RECT 123.770 53.150 123.910 53.485 ;
        RECT 124.730 53.150 124.870 53.485 ;
        RECT 125.690 53.150 125.830 53.485 ;
        RECT 126.650 53.150 126.790 53.485 ;
        RECT 127.610 53.150 127.750 53.485 ;
        RECT 128.570 53.150 128.710 53.485 ;
        RECT 129.530 53.150 129.670 53.485 ;
        RECT 130.490 53.150 130.630 53.485 ;
        RECT 131.450 53.150 131.590 53.485 ;
        RECT 132.410 53.150 132.550 53.485 ;
        RECT 133.370 53.150 133.510 53.485 ;
        RECT 134.330 53.150 134.470 53.485 ;
        RECT 135.290 53.150 135.430 53.485 ;
        RECT 136.250 53.150 136.390 53.485 ;
        RECT 137.210 53.150 137.350 53.485 ;
        RECT 138.170 53.150 138.310 53.485 ;
        RECT 139.130 53.150 139.270 53.485 ;
        RECT 140.090 53.150 140.230 53.485 ;
        RECT 141.050 53.150 141.190 53.485 ;
        RECT 142.010 53.150 142.150 53.485 ;
        RECT 142.970 53.150 143.110 53.485 ;
        RECT 143.930 53.150 144.070 53.485 ;
        RECT 144.890 53.150 145.030 53.485 ;
        RECT 145.850 53.150 145.990 53.485 ;
        RECT 146.810 53.150 146.950 53.485 ;
        RECT 147.770 53.150 147.910 53.485 ;
        RECT 148.730 53.150 148.870 53.485 ;
        RECT 149.690 53.150 149.830 53.485 ;
        RECT 150.650 53.150 150.790 53.485 ;
        RECT 151.610 53.150 151.750 53.485 ;
        RECT 152.570 53.150 152.710 53.485 ;
        RECT 153.530 53.150 153.670 53.485 ;
        RECT 154.490 53.150 154.630 53.485 ;
        RECT 155.450 53.150 155.590 53.485 ;
        RECT 156.410 53.150 156.550 53.485 ;
        RECT 157.370 53.150 157.510 53.485 ;
        RECT 158.330 53.150 158.470 53.485 ;
        RECT 159.290 53.150 159.430 53.485 ;
        RECT 160.250 53.150 160.390 53.485 ;
        RECT 161.210 53.150 161.350 53.485 ;
        RECT 162.170 53.150 162.310 53.485 ;
        RECT 163.130 53.150 163.270 53.485 ;
        RECT 164.090 53.150 164.230 53.485 ;
        RECT 165.050 53.150 165.190 53.485 ;
        RECT 166.010 53.150 166.150 53.485 ;
        RECT 166.970 53.150 167.110 53.485 ;
        RECT 167.930 53.150 212.745 53.485 ;
        RECT 5.655 0.610 212.745 53.150 ;
        RECT 5.655 0.100 14.470 0.610 ;
        RECT 15.290 0.100 20.230 0.610 ;
        RECT 21.050 0.100 25.990 0.610 ;
        RECT 26.810 0.100 31.750 0.610 ;
        RECT 32.570 0.100 37.510 0.610 ;
        RECT 38.330 0.100 43.270 0.610 ;
        RECT 44.090 0.100 49.030 0.610 ;
        RECT 49.850 0.100 54.790 0.610 ;
        RECT 55.610 0.100 60.550 0.610 ;
        RECT 61.370 0.100 66.310 0.610 ;
        RECT 67.130 0.100 72.070 0.610 ;
        RECT 72.890 0.100 77.830 0.610 ;
        RECT 78.650 0.100 83.590 0.610 ;
        RECT 84.410 0.100 89.350 0.610 ;
        RECT 90.170 0.100 95.110 0.610 ;
        RECT 95.930 0.100 100.870 0.610 ;
        RECT 101.690 0.100 106.630 0.610 ;
        RECT 107.450 0.100 112.390 0.610 ;
        RECT 113.210 0.100 118.150 0.610 ;
        RECT 118.970 0.100 123.910 0.610 ;
        RECT 124.730 0.100 129.670 0.610 ;
        RECT 130.490 0.100 135.430 0.610 ;
        RECT 136.250 0.100 141.190 0.610 ;
        RECT 142.010 0.100 146.950 0.610 ;
        RECT 147.770 0.100 152.710 0.610 ;
        RECT 153.530 0.100 158.470 0.610 ;
        RECT 159.290 0.100 164.230 0.610 ;
        RECT 165.050 0.100 169.990 0.610 ;
        RECT 170.810 0.100 175.750 0.610 ;
        RECT 176.570 0.100 181.510 0.610 ;
        RECT 182.330 0.100 187.270 0.610 ;
        RECT 188.090 0.100 193.030 0.610 ;
        RECT 193.850 0.100 198.790 0.610 ;
        RECT 199.610 0.100 212.745 0.610 ;
      LAYER Metal3 ;
        RECT 0.380 52.910 214.640 53.440 ;
        RECT 0.610 52.090 214.430 52.910 ;
        RECT 0.380 51.230 214.640 52.090 ;
        RECT 0.610 50.410 214.430 51.230 ;
        RECT 0.380 49.550 214.640 50.410 ;
        RECT 0.610 48.730 214.430 49.550 ;
        RECT 0.380 47.870 214.640 48.730 ;
        RECT 0.610 47.050 214.430 47.870 ;
        RECT 0.380 46.190 214.640 47.050 ;
        RECT 0.610 45.370 214.430 46.190 ;
        RECT 0.380 44.510 214.640 45.370 ;
        RECT 0.610 43.690 214.430 44.510 ;
        RECT 0.380 42.830 214.640 43.690 ;
        RECT 0.610 42.010 214.430 42.830 ;
        RECT 0.380 41.150 214.640 42.010 ;
        RECT 0.610 40.330 214.430 41.150 ;
        RECT 0.380 39.470 214.640 40.330 ;
        RECT 0.610 38.650 214.430 39.470 ;
        RECT 0.380 37.790 214.640 38.650 ;
        RECT 0.610 36.970 214.430 37.790 ;
        RECT 0.380 36.110 214.640 36.970 ;
        RECT 0.610 35.290 214.430 36.110 ;
        RECT 0.380 34.430 214.640 35.290 ;
        RECT 0.610 33.610 214.430 34.430 ;
        RECT 0.380 32.750 214.640 33.610 ;
        RECT 0.610 31.930 214.430 32.750 ;
        RECT 0.380 31.070 214.640 31.930 ;
        RECT 0.610 30.250 214.430 31.070 ;
        RECT 0.380 29.390 214.640 30.250 ;
        RECT 0.610 28.570 214.430 29.390 ;
        RECT 0.380 27.710 214.640 28.570 ;
        RECT 0.610 26.890 214.430 27.710 ;
        RECT 0.380 26.030 214.640 26.890 ;
        RECT 0.610 25.210 214.430 26.030 ;
        RECT 0.380 24.350 214.640 25.210 ;
        RECT 0.610 23.530 214.430 24.350 ;
        RECT 0.380 22.670 214.640 23.530 ;
        RECT 0.610 21.850 214.430 22.670 ;
        RECT 0.380 20.990 214.640 21.850 ;
        RECT 0.610 20.170 214.430 20.990 ;
        RECT 0.380 19.310 214.640 20.170 ;
        RECT 0.610 18.490 214.430 19.310 ;
        RECT 0.380 17.630 214.640 18.490 ;
        RECT 0.610 16.810 214.430 17.630 ;
        RECT 0.380 15.950 214.640 16.810 ;
        RECT 0.610 15.130 214.430 15.950 ;
        RECT 0.380 14.270 214.640 15.130 ;
        RECT 0.610 13.450 214.430 14.270 ;
        RECT 0.380 12.590 214.640 13.450 ;
        RECT 0.610 11.770 214.430 12.590 ;
        RECT 0.380 10.910 214.640 11.770 ;
        RECT 0.610 10.090 214.430 10.910 ;
        RECT 0.380 9.230 214.640 10.090 ;
        RECT 0.610 8.410 214.430 9.230 ;
        RECT 0.380 7.550 214.640 8.410 ;
        RECT 0.610 6.730 214.430 7.550 ;
        RECT 0.380 5.870 214.640 6.730 ;
        RECT 0.610 5.050 214.430 5.870 ;
        RECT 0.380 4.190 214.640 5.050 ;
        RECT 0.610 3.370 214.430 4.190 ;
        RECT 0.380 2.510 214.640 3.370 ;
        RECT 0.610 1.690 214.430 2.510 ;
        RECT 0.380 0.830 214.640 1.690 ;
        RECT 0.610 0.320 214.430 0.830 ;
      LAYER Metal4 ;
        RECT 2.295 0.695 212.745 53.065 ;
      LAYER Metal5 ;
        RECT 2.255 2.420 212.785 49.450 ;
  END
END S_IO4
END LIBRARY

