* NGSPICE file created from SE_term.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

.subckt SE_term FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3]
+ N2BEG[0] N2BEG[1] N2BEG[2] N2BEG[3] N2BEG[4] N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0]
+ N2BEGb[1] N2BEGb[2] N2BEGb[3] N2BEGb[4] N2BEGb[5] N2BEGb[6] N2BEGb[7] N4BEG[0] N4BEG[10]
+ N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2] N4BEG[3] N4BEG[4]
+ N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9] S1END[0] S1END[1] S1END[2] S1END[3]
+ S2END[0] S2END[1] S2END[2] S2END[3] S2END[4] S2END[5] S2END[6] S2END[7] S2MID[0]
+ S2MID[1] S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6] S2MID[7] S4END[0] S4END[10]
+ S4END[11] S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3] S4END[4]
+ S4END[5] S4END[6] S4END[7] S4END[8] S4END[9] UserCLK UserCLKo VGND VPWR
XFILLER_7_7 VPWR VGND sg13g2_fill_1
XFILLER_9_148 VPWR VGND sg13g2_decap_8
XFILLER_3_56 VPWR VGND sg13g2_decap_8
X_83_ S4END[4] N4BEG[11] VPWR VGND sg13g2_buf_1
XFILLER_10_169 VPWR VGND sg13g2_fill_2
XFILLER_6_118 VPWR VGND sg13g2_decap_8
XFILLER_10_114 VPWR VGND sg13g2_decap_8
XFILLER_5_195 VPWR VGND sg13g2_decap_4
X_66_ S2END[5] N2BEGb[2] VPWR VGND sg13g2_buf_1
XFILLER_0_35 VPWR VGND sg13g2_decap_8
XFILLER_2_198 VPWR VGND sg13g2_fill_2
XFILLER_9_11 VPWR VGND sg13g2_fill_2
XFILLER_9_55 VPWR VGND sg13g2_decap_4
X_49_ FrameStrobe[17] FrameStrobe_O[17] VPWR VGND sg13g2_buf_1
XFILLER_6_56 VPWR VGND sg13g2_decap_8
XFILLER_11_0 VPWR VGND sg13g2_decap_8
XFILLER_3_35 VPWR VGND sg13g2_decap_8
XFILLER_8_193 VPWR VGND sg13g2_decap_8
X_82_ S4END[5] N4BEG[10] VPWR VGND sg13g2_buf_1
XFILLER_5_174 VPWR VGND sg13g2_decap_8
X_65_ S2END[6] N2BEGb[1] VPWR VGND sg13g2_buf_1
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_2_133 VPWR VGND sg13g2_decap_4
XFILLER_2_177 VPWR VGND sg13g2_decap_8
XFILLER_9_34 VPWR VGND sg13g2_decap_8
X_48_ FrameStrobe[16] FrameStrobe_O[16] VPWR VGND sg13g2_buf_1
XFILLER_6_35 VPWR VGND sg13g2_decap_8
XFILLER_9_117 VPWR VGND sg13g2_fill_2
XFILLER_3_14 VPWR VGND sg13g2_decap_8
XFILLER_8_172 VPWR VGND sg13g2_decap_8
X_81_ S4END[6] N4BEG[9] VPWR VGND sg13g2_buf_1
XFILLER_5_153 VPWR VGND sg13g2_decap_8
X_64_ S2END[7] N2BEGb[0] VPWR VGND sg13g2_buf_1
XFILLER_2_112 VPWR VGND sg13g2_decap_8
XFILLER_2_156 VPWR VGND sg13g2_decap_8
XFILLER_9_13 VPWR VGND sg13g2_fill_1
X_47_ FrameStrobe[15] FrameStrobe_O[15] VPWR VGND sg13g2_buf_1
XFILLER_9_79 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_fill_2
XFILLER_6_14 VPWR VGND sg13g2_decap_8
XFILLER_9_129 VPWR VGND sg13g2_fill_1
XFILLER_8_151 VPWR VGND sg13g2_decap_8
X_80_ S4END[7] N4BEG[8] VPWR VGND sg13g2_buf_1
XFILLER_5_7 VPWR VGND sg13g2_decap_4
XFILLER_10_128 VPWR VGND sg13g2_decap_8
XFILLER_5_132 VPWR VGND sg13g2_decap_8
X_63_ S2MID[0] N2BEG[7] VPWR VGND sg13g2_buf_1
XFILLER_0_49 VPWR VGND sg13g2_decap_8
X_46_ FrameStrobe[14] FrameStrobe_O[14] VPWR VGND sg13g2_buf_1
X_29_ FrameData[29] FrameData_O[29] VPWR VGND sg13g2_buf_1
XFILLER_3_49 VPWR VGND sg13g2_decap_8
XFILLER_9_119 VPWR VGND sg13g2_fill_1
XFILLER_8_130 VPWR VGND sg13g2_decap_8
XFILLER_5_111 VPWR VGND sg13g2_decap_8
XFILLER_5_188 VPWR VGND sg13g2_decap_8
XFILLER_5_199 VPWR VGND sg13g2_fill_1
X_62_ S2MID[1] N2BEG[6] VPWR VGND sg13g2_buf_1
XFILLER_0_28 VPWR VGND sg13g2_decap_8
XFILLER_9_26 VPWR VGND sg13g2_decap_4
XFILLER_9_48 VPWR VGND sg13g2_decap_8
XFILLER_9_59 VPWR VGND sg13g2_fill_2
X_45_ FrameStrobe[13] FrameStrobe_O[13] VPWR VGND sg13g2_buf_1
XFILLER_1_2 VPWR VGND sg13g2_fill_1
X_28_ FrameData[28] FrameData_O[28] VPWR VGND sg13g2_buf_1
XFILLER_1_93 VPWR VGND sg13g2_decap_4
XFILLER_6_49 VPWR VGND sg13g2_decap_8
XFILLER_10_91 VPWR VGND sg13g2_fill_1
XFILLER_3_28 VPWR VGND sg13g2_decap_8
XFILLER_8_186 VPWR VGND sg13g2_decap_8
XFILLER_5_167 VPWR VGND sg13g2_decap_8
X_61_ S2MID[2] N2BEG[5] VPWR VGND sg13g2_buf_1
XFILLER_4_82 VPWR VGND sg13g2_decap_8
XFILLER_4_93 VPWR VGND sg13g2_decap_8
XFILLER_2_126 VPWR VGND sg13g2_decap_8
XFILLER_2_137 VPWR VGND sg13g2_fill_1
X_44_ FrameStrobe[12] FrameStrobe_O[12] VPWR VGND sg13g2_buf_1
X_27_ FrameData[27] FrameData_O[27] VPWR VGND sg13g2_buf_1
XFILLER_1_72 VPWR VGND sg13g2_fill_2
XFILLER_6_28 VPWR VGND sg13g2_decap_8
XFILLER_7_82 VPWR VGND sg13g2_decap_8
XFILLER_8_165 VPWR VGND sg13g2_decap_8
XFILLER_5_146 VPWR VGND sg13g2_decap_8
X_60_ S2MID[3] N2BEG[4] VPWR VGND sg13g2_buf_1
XFILLER_4_61 VPWR VGND sg13g2_decap_8
XFILLER_2_105 VPWR VGND sg13g2_decap_8
XFILLER_2_149 VPWR VGND sg13g2_decap_8
XFILLER_3_7 VPWR VGND sg13g2_fill_2
X_43_ FrameStrobe[11] FrameStrobe_O[11] VPWR VGND sg13g2_buf_1
XFILLER_1_160 VPWR VGND sg13g2_decap_8
X_26_ FrameData[26] FrameData_O[26] VPWR VGND sg13g2_buf_1
XFILLER_1_40 VPWR VGND sg13g2_decap_4
XFILLER_10_82 VPWR VGND sg13g2_decap_8
X_09_ FrameData[9] FrameData_O[9] VPWR VGND sg13g2_buf_1
XFILLER_7_61 VPWR VGND sg13g2_decap_8
XFILLER_8_144 VPWR VGND sg13g2_decap_8
XFILLER_5_125 VPWR VGND sg13g2_decap_8
XFILLER_4_40 VPWR VGND sg13g2_decap_8
XFILLER_9_18 VPWR VGND sg13g2_decap_4
X_42_ FrameStrobe[10] FrameStrobe_O[10] VPWR VGND sg13g2_buf_1
XFILLER_1_85 VPWR VGND sg13g2_decap_4
X_25_ FrameData[25] FrameData_O[25] VPWR VGND sg13g2_buf_1
XFILLER_10_50 VPWR VGND sg13g2_fill_1
X_08_ FrameData[8] FrameData_O[8] VPWR VGND sg13g2_buf_1
XFILLER_11_7 VPWR VGND sg13g2_decap_8
XFILLER_7_40 VPWR VGND sg13g2_decap_8
XFILLER_8_123 VPWR VGND sg13g2_decap_8
XFILLER_5_104 VPWR VGND sg13g2_decap_8
XFILLER_3_9 VPWR VGND sg13g2_fill_1
XFILLER_1_184 VPWR VGND sg13g2_fill_2
X_41_ FrameStrobe[9] FrameStrobe_O[9] VPWR VGND sg13g2_buf_1
X_24_ FrameData[24] FrameData_O[24] VPWR VGND sg13g2_buf_1
X_07_ FrameData[7] FrameData_O[7] VPWR VGND sg13g2_buf_1
XFILLER_7_96 VPWR VGND sg13g2_decap_8
XFILLER_8_102 VPWR VGND sg13g2_decap_8
XFILLER_8_179 VPWR VGND sg13g2_decap_8
XFILLER_4_182 VPWR VGND sg13g2_decap_4
XFILLER_2_119 VPWR VGND sg13g2_decap_8
XFILLER_4_75 VPWR VGND sg13g2_decap_8
XFILLER_1_141 VPWR VGND sg13g2_decap_4
X_40_ FrameStrobe[8] FrameStrobe_O[8] VPWR VGND sg13g2_buf_1
XFILLER_8_0 VPWR VGND sg13g2_decap_8
XFILLER_1_65 VPWR VGND sg13g2_decap_8
X_23_ FrameData[23] FrameData_O[23] VPWR VGND sg13g2_buf_1
XFILLER_10_96 VPWR VGND sg13g2_fill_2
X_06_ FrameData[6] FrameData_O[6] VPWR VGND sg13g2_buf_1
XFILLER_7_75 VPWR VGND sg13g2_decap_8
XFILLER_8_158 VPWR VGND sg13g2_decap_8
XFILLER_5_139 VPWR VGND sg13g2_decap_8
XFILLER_4_54 VPWR VGND sg13g2_decap_8
XFILLER_4_161 VPWR VGND sg13g2_decap_8
XFILLER_4_194 VPWR VGND sg13g2_decap_4
XFILLER_1_44 VPWR VGND sg13g2_fill_2
X_22_ FrameData[22] FrameData_O[22] VPWR VGND sg13g2_buf_1
XFILLER_10_75 VPWR VGND sg13g2_decap_8
X_05_ FrameData[5] FrameData_O[5] VPWR VGND sg13g2_buf_1
XFILLER_7_54 VPWR VGND sg13g2_decap_8
XFILLER_8_137 VPWR VGND sg13g2_decap_8
XFILLER_5_118 VPWR VGND sg13g2_decap_8
XFILLER_4_33 VPWR VGND sg13g2_decap_8
XFILLER_4_140 VPWR VGND sg13g2_decap_8
XFILLER_1_198 VPWR VGND sg13g2_fill_2
XFILLER_1_110 VPWR VGND sg13g2_fill_1
X_21_ FrameData[21] FrameData_O[21] VPWR VGND sg13g2_buf_1
XFILLER_1_78 VPWR VGND sg13g2_decap_8
XFILLER_10_32 VPWR VGND sg13g2_fill_1
X_04_ FrameData[4] FrameData_O[4] VPWR VGND sg13g2_buf_1
XFILLER_7_33 VPWR VGND sg13g2_decap_8
XFILLER_8_116 VPWR VGND sg13g2_decap_8
XFILLER_7_193 VPWR VGND sg13g2_decap_8
XFILLER_1_177 VPWR VGND sg13g2_decap_8
XFILLER_1_155 VPWR VGND sg13g2_fill_1
XFILLER_1_122 VPWR VGND sg13g2_fill_1
XFILLER_6_0 VPWR VGND sg13g2_decap_8
X_20_ FrameData[20] FrameData_O[20] VPWR VGND sg13g2_buf_1
XFILLER_10_55 VPWR VGND sg13g2_decap_4
X_03_ FrameData[3] FrameData_O[3] VPWR VGND sg13g2_buf_1
XFILLER_7_12 VPWR VGND sg13g2_decap_8
XFILLER_7_89 VPWR VGND sg13g2_decap_8
XFILLER_7_161 VPWR VGND sg13g2_decap_8
XFILLER_7_183 VPWR VGND sg13g2_fill_2
XFILLER_4_68 VPWR VGND sg13g2_decap_8
XFILLER_4_175 VPWR VGND sg13g2_decap_8
XFILLER_1_167 VPWR VGND sg13g2_fill_2
XFILLER_1_134 VPWR VGND sg13g2_fill_2
XFILLER_1_101 VPWR VGND sg13g2_decap_8
XFILLER_1_58 VPWR VGND sg13g2_decap_8
XFILLER_1_25 VPWR VGND sg13g2_fill_2
XFILLER_10_45 VPWR VGND sg13g2_fill_1
X_79_ S4END[8] N4BEG[7] VPWR VGND sg13g2_buf_1
XFILLER_10_89 VPWR VGND sg13g2_fill_2
X_02_ FrameData[2] FrameData_O[2] VPWR VGND sg13g2_buf_1
XFILLER_7_68 VPWR VGND sg13g2_decap_8
XFILLER_11_191 VPWR VGND sg13g2_decap_8
XFILLER_4_47 VPWR VGND sg13g2_decap_8
XFILLER_4_121 VPWR VGND sg13g2_fill_1
XFILLER_4_154 VPWR VGND sg13g2_decap_8
XFILLER_4_198 VPWR VGND sg13g2_fill_2
XFILLER_5_90 VPWR VGND sg13g2_decap_8
XFILLER_1_15 VPWR VGND sg13g2_decap_4
X_78_ S4END[9] N4BEG[6] VPWR VGND sg13g2_buf_1
X_01_ FrameData[1] FrameData_O[1] VPWR VGND sg13g2_buf_1
XFILLER_2_91 VPWR VGND sg13g2_decap_8
XFILLER_7_47 VPWR VGND sg13g2_decap_8
XFILLER_7_152 VPWR VGND sg13g2_decap_4
XFILLER_4_26 VPWR VGND sg13g2_decap_8
XFILLER_4_100 VPWR VGND sg13g2_decap_8
XFILLER_4_133 VPWR VGND sg13g2_decap_8
XFILLER_1_136 VPWR VGND sg13g2_fill_1
XFILLER_1_27 VPWR VGND sg13g2_fill_1
X_77_ S4END[10] N4BEG[5] VPWR VGND sg13g2_buf_1
XFILLER_10_25 VPWR VGND sg13g2_decap_8
XFILLER_10_69 VPWR VGND sg13g2_fill_2
X_00_ FrameData[0] FrameData_O[0] VPWR VGND sg13g2_buf_1
XFILLER_4_0 VPWR VGND sg13g2_decap_8
XFILLER_2_70 VPWR VGND sg13g2_decap_8
XFILLER_7_26 VPWR VGND sg13g2_decap_8
XFILLER_8_109 VPWR VGND sg13g2_decap_8
XFILLER_11_182 VPWR VGND sg13g2_decap_4
XFILLER_7_131 VPWR VGND sg13g2_decap_8
XFILLER_1_115 VPWR VGND sg13g2_decap_8
X_76_ S4END[11] N4BEG[4] VPWR VGND sg13g2_buf_1
XFILLER_10_59 VPWR VGND sg13g2_fill_2
X_59_ S2MID[4] N2BEG[3] VPWR VGND sg13g2_buf_1
XFILLER_11_91 VPWR VGND sg13g2_decap_8
XFILLER_11_161 VPWR VGND sg13g2_decap_8
XFILLER_7_110 VPWR VGND sg13g2_decap_8
XFILLER_7_176 VPWR VGND sg13g2_decap_8
XFILLER_8_81 VPWR VGND sg13g2_decap_8
XFILLER_4_168 VPWR VGND sg13g2_decap_8
XFILLER_1_149 VPWR VGND sg13g2_fill_2
XFILLER_1_127 VPWR VGND sg13g2_decap_8
XFILLER_0_182 VPWR VGND sg13g2_decap_8
XFILLER_5_71 VPWR VGND sg13g2_decap_8
X_75_ S4END[12] N4BEG[3] VPWR VGND sg13g2_buf_1
X_58_ S2MID[5] N2BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_11_70 VPWR VGND sg13g2_decap_8
XFILLER_11_140 VPWR VGND sg13g2_decap_8
XFILLER_8_60 VPWR VGND sg13g2_decap_8
XFILLER_4_114 VPWR VGND sg13g2_decap_8
XFILLER_4_147 VPWR VGND sg13g2_decap_8
XFILLER_0_161 VPWR VGND sg13g2_decap_8
XFILLER_5_50 VPWR VGND sg13g2_decap_8
XFILLER_1_19 VPWR VGND sg13g2_fill_2
X_74_ S4END[13] N4BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_2_84 VPWR VGND sg13g2_decap_8
X_57_ S2MID[6] N2BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_2_0 VPWR VGND sg13g2_decap_8
XFILLER_7_145 VPWR VGND sg13g2_decap_8
XFILLER_7_156 VPWR VGND sg13g2_fill_1
XFILLER_4_19 VPWR VGND sg13g2_decap_8
XFILLER_4_126 VPWR VGND sg13g2_decap_8
XFILLER_0_140 VPWR VGND sg13g2_decap_8
XFILLER_6_7 VPWR VGND sg13g2_decap_8
X_73_ S4END[14] N4BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_10_18 VPWR VGND sg13g2_decap_8
XFILLER_2_63 VPWR VGND sg13g2_decap_8
X_56_ S2MID[7] N2BEG[0] VPWR VGND sg13g2_buf_1
XFILLER_7_19 VPWR VGND sg13g2_decap_8
X_39_ FrameStrobe[7] FrameStrobe_O[7] VPWR VGND sg13g2_buf_1
XFILLER_11_186 VPWR VGND sg13g2_fill_1
XFILLER_11_175 VPWR VGND sg13g2_decap_8
XFILLER_7_124 VPWR VGND sg13g2_decap_8
XFILLER_7_168 VPWR VGND sg13g2_decap_4
XFILLER_8_95 VPWR VGND sg13g2_decap_8
XFILLER_1_108 VPWR VGND sg13g2_fill_2
XFILLER_3_182 VPWR VGND sg13g2_decap_8
XFILLER_0_196 VPWR VGND sg13g2_decap_4
XFILLER_5_85 VPWR VGND sg13g2_fill_1
XFILLER_10_0 VPWR VGND sg13g2_decap_4
X_72_ S4END[15] N4BEG[0] VPWR VGND sg13g2_buf_1
XFILLER_2_42 VPWR VGND sg13g2_decap_8
X_55_ S1END[0] N1BEG[3] VPWR VGND sg13g2_buf_1
XFILLER_11_84 VPWR VGND sg13g2_decap_8
X_38_ FrameStrobe[6] FrameStrobe_O[6] VPWR VGND sg13g2_buf_1
XFILLER_11_198 VPWR VGND sg13g2_fill_2
XFILLER_11_154 VPWR VGND sg13g2_decap_8
XFILLER_7_103 VPWR VGND sg13g2_decap_8
XFILLER_8_74 VPWR VGND sg13g2_decap_8
XFILLER_3_161 VPWR VGND sg13g2_decap_8
XFILLER_0_175 VPWR VGND sg13g2_decap_8
XFILLER_5_64 VPWR VGND sg13g2_decap_8
XFILLER_5_97 VPWR VGND sg13g2_decap_8
X_71_ S2END[0] N2BEGb[7] VPWR VGND sg13g2_buf_1
XFILLER_2_21 VPWR VGND sg13g2_decap_8
XFILLER_2_98 VPWR VGND sg13g2_decap_8
X_54_ S1END[1] N1BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_11_63 VPWR VGND sg13g2_decap_8
X_37_ FrameStrobe[5] FrameStrobe_O[5] VPWR VGND sg13g2_buf_1
XFILLER_11_133 VPWR VGND sg13g2_decap_8
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_8_53 VPWR VGND sg13g2_decap_8
XFILLER_4_107 VPWR VGND sg13g2_decap_8
XFILLER_3_140 VPWR VGND sg13g2_decap_8
XFILLER_0_154 VPWR VGND sg13g2_decap_8
XFILLER_5_43 VPWR VGND sg13g2_decap_8
X_70_ S2END[1] N2BEGb[6] VPWR VGND sg13g2_buf_1
XFILLER_2_77 VPWR VGND sg13g2_decap_8
X_53_ S1END[2] N1BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_11_42 VPWR VGND sg13g2_decap_8
X_36_ FrameStrobe[4] FrameStrobe_O[4] VPWR VGND sg13g2_buf_1
XFILLER_11_112 VPWR VGND sg13g2_decap_8
XFILLER_7_138 VPWR VGND sg13g2_decap_8
XFILLER_6_160 VPWR VGND sg13g2_fill_2
XFILLER_6_193 VPWR VGND sg13g2_decap_8
XFILLER_8_32 VPWR VGND sg13g2_decap_8
X_19_ FrameData[19] FrameData_O[19] VPWR VGND sg13g2_buf_1
XFILLER_3_196 VPWR VGND sg13g2_decap_4
XFILLER_0_133 VPWR VGND sg13g2_decap_8
XFILLER_5_22 VPWR VGND sg13g2_decap_8
XFILLER_2_56 VPWR VGND sg13g2_decap_8
X_52_ S1END[3] N1BEG[0] VPWR VGND sg13g2_buf_1
XFILLER_11_98 VPWR VGND sg13g2_decap_8
XFILLER_11_21 VPWR VGND sg13g2_decap_8
X_35_ FrameStrobe[3] FrameStrobe_O[3] VPWR VGND sg13g2_buf_1
XFILLER_11_168 VPWR VGND sg13g2_decap_8
XFILLER_9_191 VPWR VGND sg13g2_decap_8
XFILLER_7_117 VPWR VGND sg13g2_decap_8
XFILLER_8_11 VPWR VGND sg13g2_decap_8
XFILLER_8_88 VPWR VGND sg13g2_decap_8
X_18_ FrameData[18] FrameData_O[18] VPWR VGND sg13g2_buf_1
XFILLER_3_175 VPWR VGND sg13g2_decap_8
XFILLER_0_189 VPWR VGND sg13g2_decap_8
XFILLER_0_112 VPWR VGND sg13g2_decap_8
XFILLER_5_78 VPWR VGND sg13g2_decap_8
XFILLER_10_4 VPWR VGND sg13g2_fill_2
XFILLER_2_35 VPWR VGND sg13g2_decap_8
X_51_ FrameStrobe[19] FrameStrobe_O[19] VPWR VGND sg13g2_buf_1
XFILLER_11_77 VPWR VGND sg13g2_decap_8
X_34_ FrameStrobe[2] FrameStrobe_O[2] VPWR VGND sg13g2_buf_1
XFILLER_11_147 VPWR VGND sg13g2_decap_8
XFILLER_8_67 VPWR VGND sg13g2_decap_8
X_17_ FrameData[17] FrameData_O[17] VPWR VGND sg13g2_buf_1
XFILLER_6_173 VPWR VGND sg13g2_decap_8
XFILLER_6_184 VPWR VGND sg13g2_decap_4
XFILLER_3_154 VPWR VGND sg13g2_decap_8
XFILLER_0_168 VPWR VGND sg13g2_decap_8
XFILLER_5_57 VPWR VGND sg13g2_decap_8
XFILLER_2_14 VPWR VGND sg13g2_decap_8
X_50_ FrameStrobe[18] FrameStrobe_O[18] VPWR VGND sg13g2_buf_1
XFILLER_9_0 VPWR VGND sg13g2_decap_8
XFILLER_11_56 VPWR VGND sg13g2_decap_8
XFILLER_2_7 VPWR VGND sg13g2_decap_8
X_33_ FrameStrobe[1] FrameStrobe_O[1] VPWR VGND sg13g2_buf_1
XFILLER_9_182 VPWR VGND sg13g2_decap_4
XFILLER_9_160 VPWR VGND sg13g2_decap_4
XFILLER_11_126 VPWR VGND sg13g2_decap_8
X_16_ FrameData[16] FrameData_O[16] VPWR VGND sg13g2_buf_1
XFILLER_8_46 VPWR VGND sg13g2_decap_8
XFILLER_3_133 VPWR VGND sg13g2_decap_8
XFILLER_0_91 VPWR VGND sg13g2_decap_8
XFILLER_0_147 VPWR VGND sg13g2_decap_8
XFILLER_5_36 VPWR VGND sg13g2_decap_8
XFILLER_11_35 VPWR VGND sg13g2_decap_8
X_32_ FrameStrobe[0] FrameStrobe_O[0] VPWR VGND sg13g2_buf_1
XFILLER_11_105 VPWR VGND sg13g2_decap_8
XFILLER_3_91 VPWR VGND sg13g2_decap_8
XFILLER_10_171 VPWR VGND sg13g2_fill_1
X_15_ FrameData[15] FrameData_O[15] VPWR VGND sg13g2_buf_1
XFILLER_6_153 VPWR VGND sg13g2_decap_8
XFILLER_8_25 VPWR VGND sg13g2_decap_8
XFILLER_3_112 VPWR VGND sg13g2_decap_8
XFILLER_3_189 VPWR VGND sg13g2_decap_8
XFILLER_0_70 VPWR VGND sg13g2_decap_8
XFILLER_0_126 VPWR VGND sg13g2_decap_8
XFILLER_5_15 VPWR VGND sg13g2_decap_8
XFILLER_6_91 VPWR VGND sg13g2_decap_8
XFILLER_2_49 VPWR VGND sg13g2_decap_8
XFILLER_11_14 VPWR VGND sg13g2_decap_8
X_31_ FrameData[31] FrameData_O[31] VPWR VGND sg13g2_buf_1
XFILLER_3_70 VPWR VGND sg13g2_decap_8
XFILLER_6_132 VPWR VGND sg13g2_decap_8
XFILLER_10_150 VPWR VGND sg13g2_decap_4
X_14_ FrameData[14] FrameData_O[14] VPWR VGND sg13g2_buf_1
XFILLER_3_168 VPWR VGND sg13g2_decap_8
XFILLER_0_105 VPWR VGND sg13g2_decap_8
XFILLER_6_70 VPWR VGND sg13g2_decap_8
XFILLER_2_28 VPWR VGND sg13g2_decap_8
X_30_ FrameData[30] FrameData_O[30] VPWR VGND sg13g2_buf_1
XFILLER_7_0 VPWR VGND sg13g2_decap_8
XFILLER_9_141 VPWR VGND sg13g2_decap_8
XFILLER_10_195 VPWR VGND sg13g2_decap_4
XFILLER_0_7 VPWR VGND sg13g2_decap_8
XFILLER_6_166 VPWR VGND sg13g2_decap_8
XFILLER_6_188 VPWR VGND sg13g2_fill_1
X_13_ FrameData[13] FrameData_O[13] VPWR VGND sg13g2_buf_1
XFILLER_3_147 VPWR VGND sg13g2_decap_8
XFILLER_2_191 VPWR VGND sg13g2_decap_8
XFILLER_11_49 VPWR VGND sg13g2_decap_8
XFILLER_11_119 VPWR VGND sg13g2_decap_8
XFILLER_9_186 VPWR VGND sg13g2_fill_1
XFILLER_9_175 VPWR VGND sg13g2_decap_8
XFILLER_8_39 VPWR VGND sg13g2_decap_8
XFILLER_10_163 VPWR VGND sg13g2_fill_2
X_12_ FrameData[12] FrameData_O[12] VPWR VGND sg13g2_buf_1
XFILLER_6_112 VPWR VGND sg13g2_fill_2
XFILLER_3_126 VPWR VGND sg13g2_decap_8
XFILLER_2_170 VPWR VGND sg13g2_decap_8
XFILLER_0_84 VPWR VGND sg13g2_decap_8
XFILLER_5_29 VPWR VGND sg13g2_decap_8
XFILLER_11_28 VPWR VGND sg13g2_decap_8
XFILLER_9_198 VPWR VGND sg13g2_fill_2
X_88_ UserCLK UserCLKo VPWR VGND sg13g2_buf_1
XFILLER_3_84 VPWR VGND sg13g2_decap_8
XFILLER_9_110 VPWR VGND sg13g2_decap_8
X_11_ FrameData[11] FrameData_O[11] VPWR VGND sg13g2_buf_1
XFILLER_6_146 VPWR VGND sg13g2_decap_8
XFILLER_8_18 VPWR VGND sg13g2_decap_8
XFILLER_3_105 VPWR VGND sg13g2_decap_8
XFILLER_0_63 VPWR VGND sg13g2_decap_8
XFILLER_0_119 VPWR VGND sg13g2_decap_8
XFILLER_6_84 VPWR VGND sg13g2_decap_8
XFILLER_9_155 VPWR VGND sg13g2_fill_1
XFILLER_3_63 VPWR VGND sg13g2_decap_8
X_87_ S4END[0] N4BEG[15] VPWR VGND sg13g2_buf_1
XFILLER_10_176 VPWR VGND sg13g2_decap_8
X_10_ FrameData[10] FrameData_O[10] VPWR VGND sg13g2_buf_1
XFILLER_5_0 VPWR VGND sg13g2_decap_8
XFILLER_6_125 VPWR VGND sg13g2_decap_8
XFILLER_10_121 VPWR VGND sg13g2_decap_8
XFILLER_10_154 VPWR VGND sg13g2_fill_1
XFILLER_0_42 VPWR VGND sg13g2_decap_8
XFILLER_9_95 VPWR VGND sg13g2_decap_8
XFILLER_6_63 VPWR VGND sg13g2_decap_8
XFILLER_9_134 VPWR VGND sg13g2_decap_8
XFILLER_3_42 VPWR VGND sg13g2_decap_8
X_86_ S4END[1] N4BEG[14] VPWR VGND sg13g2_buf_1
XFILLER_10_199 VPWR VGND sg13g2_fill_1
XFILLER_10_144 VPWR VGND sg13g2_fill_2
XFILLER_5_181 VPWR VGND sg13g2_decap_8
X_69_ S2END[2] N2BEGb[5] VPWR VGND sg13g2_buf_1
XFILLER_0_98 VPWR VGND sg13g2_decap_8
XFILLER_0_21 VPWR VGND sg13g2_decap_8
XFILLER_2_184 VPWR VGND sg13g2_decap_8
XFILLER_9_41 VPWR VGND sg13g2_decap_8
XFILLER_6_42 VPWR VGND sg13g2_decap_8
XFILLER_9_102 VPWR VGND sg13g2_decap_4
XFILLER_9_124 VPWR VGND sg13g2_fill_1
XFILLER_9_168 VPWR VGND sg13g2_decap_8
XFILLER_3_21 VPWR VGND sg13g2_decap_8
XFILLER_3_98 VPWR VGND sg13g2_decap_8
X_85_ S4END[2] N4BEG[13] VPWR VGND sg13g2_buf_1
XFILLER_6_105 VPWR VGND sg13g2_decap_8
XFILLER_5_160 VPWR VGND sg13g2_decap_8
XFILLER_3_119 VPWR VGND sg13g2_decap_8
X_68_ S2END[3] N2BEGb[4] VPWR VGND sg13g2_buf_1
XFILLER_2_163 VPWR VGND sg13g2_decap_8
XFILLER_0_77 VPWR VGND sg13g2_decap_8
XFILLER_9_86 VPWR VGND sg13g2_fill_1
XFILLER_6_21 VPWR VGND sg13g2_decap_8
XFILLER_6_98 VPWR VGND sg13g2_decap_8
XFILLER_3_77 VPWR VGND sg13g2_decap_8
X_84_ S4END[3] N4BEG[12] VPWR VGND sg13g2_buf_1
XFILLER_10_135 VPWR VGND sg13g2_fill_1
XFILLER_6_139 VPWR VGND sg13g2_decap_8
X_67_ S2END[4] N2BEGb[3] VPWR VGND sg13g2_buf_1
XFILLER_2_142 VPWR VGND sg13g2_decap_8
XFILLER_3_0 VPWR VGND sg13g2_decap_8
XFILLER_0_56 VPWR VGND sg13g2_decap_8
XFILLER_9_65 VPWR VGND sg13g2_fill_2
XFILLER_6_77 VPWR VGND sg13g2_decap_8
.ends

