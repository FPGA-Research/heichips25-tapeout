`default_nettype none

module fabric_wrapper #(
    	parameter FrameBitsPerRow = 32,
	parameter MaxFramesPerCol = 20,
	
	parameter NumColumns = 6,
	parameter NumRows = 10,
	
    parameter FABRIC_NUM_IO_NORTH = 16,
    parameter FABRIC_NUM_IO_SOUTH = 16
)(
    input clk_i,
    
    // Configuration
    input  logic [(FrameBitsPerRow*NumRows)-1:0]    FrameData_i,
    input  logic [(MaxFramesPerCol*NumColumns)-1:0] FrameStrobe_i,
    
    // Fabric is configured
    input                                 configured_i,

    // I/Os North
    input  [FABRIC_NUM_IO_NORTH-1:0]      io_north_in_i,
    output [FABRIC_NUM_IO_NORTH-1:0]      io_north_out_o,
    output [FABRIC_NUM_IO_NORTH-1:0]      io_north_oe_o,

    // I/Os South
    input  [FABRIC_NUM_IO_SOUTH-1:0]      io_south_in_i,
    output [FABRIC_NUM_IO_SOUTH-1:0]      io_south_out_o,
    output [FABRIC_NUM_IO_SOUTH-1:0]      io_south_oe_o
);
    
    // TT_PROJECT 0 (X0Y1)
    logic [7:0] tt_project_0_ui_in;
    logic [7:0] tt_project_0_uo_out;
    logic [7:0] tt_project_0_uio_in;
    logic [7:0] tt_project_0_uio_out;
    logic [7:0] tt_project_0_uio_oe;
    logic  tt_project_0_ena;
    logic  tt_project_0_clk;
    logic  tt_project_0_rst_n;

    // TT_PROJECT 1 (X0Y2)
    logic [7:0] tt_project_1_ui_in;
    logic [7:0] tt_project_1_uo_out;
    logic [7:0] tt_project_1_uio_in;
    logic [7:0] tt_project_1_uio_out;
    logic [7:0] tt_project_1_uio_oe;
    logic  tt_project_1_ena;
    logic  tt_project_1_clk;
    logic  tt_project_1_rst_n;

    // TT_PROJECT 2 (X0Y3)
    logic [7:0] tt_project_2_ui_in;
    logic [7:0] tt_project_2_uo_out;
    logic [7:0] tt_project_2_uio_in;
    logic [7:0] tt_project_2_uio_out;
    logic [7:0] tt_project_2_uio_oe;
    logic  tt_project_2_ena;
    logic  tt_project_2_clk;
    logic  tt_project_2_rst_n;

    // TT_PROJECT 3 (X0Y4)
    logic [7:0] tt_project_3_ui_in;
    logic [7:0] tt_project_3_uo_out;
    logic [7:0] tt_project_3_uio_in;
    logic [7:0] tt_project_3_uio_out;
    logic [7:0] tt_project_3_uio_oe;
    logic  tt_project_3_ena;
    logic  tt_project_3_clk;
    logic  tt_project_3_rst_n;

    // TT_PROJECT 4 (X0Y5)
    logic [7:0] tt_project_4_ui_in;
    logic [7:0] tt_project_4_uo_out;
    logic [7:0] tt_project_4_uio_in;
    logic [7:0] tt_project_4_uio_out;
    logic [7:0] tt_project_4_uio_oe;
    logic  tt_project_4_ena;
    logic  tt_project_4_clk;
    logic  tt_project_4_rst_n;

    // TT_PROJECT 5 (X0Y6)
    logic [7:0] tt_project_5_ui_in;
    logic [7:0] tt_project_5_uo_out;
    logic [7:0] tt_project_5_uio_in;
    logic [7:0] tt_project_5_uio_out;
    logic [7:0] tt_project_5_uio_oe;
    logic  tt_project_5_ena;
    logic  tt_project_5_clk;
    logic  tt_project_5_rst_n;

    // TT_PROJECT 6 (X0Y7)
    logic [7:0] tt_project_6_ui_in;
    logic [7:0] tt_project_6_uo_out;
    logic [7:0] tt_project_6_uio_in;
    logic [7:0] tt_project_6_uio_out;
    logic [7:0] tt_project_6_uio_oe;
    logic  tt_project_6_ena;
    logic  tt_project_6_clk;
    logic  tt_project_6_rst_n;

    // TT_PROJECT 7 (X0Y8)
    logic [7:0] tt_project_7_ui_in;
    logic [7:0] tt_project_7_uo_out;
    logic [7:0] tt_project_7_uio_in;
    logic [7:0] tt_project_7_uio_out;
    logic [7:0] tt_project_7_uio_oe;
    logic  tt_project_7_ena;
    logic  tt_project_7_clk;
    logic  tt_project_7_rst_n;

    // TT_PROJECT 8 (X5Y3)
    logic [7:0] tt_project_8_ui_in;
    logic [7:0] tt_project_8_uo_out;
    logic [7:0] tt_project_8_uio_in;
    logic [7:0] tt_project_8_uio_out;
    logic [7:0] tt_project_8_uio_oe;
    logic  tt_project_8_ena;
    logic  tt_project_8_clk;
    logic  tt_project_8_rst_n;

    // TT_PROJECT 9 (X5Y4)
    logic [7:0] tt_project_9_ui_in;
    logic [7:0] tt_project_9_uo_out;
    logic [7:0] tt_project_9_uio_in;
    logic [7:0] tt_project_9_uio_out;
    logic [7:0] tt_project_9_uio_oe;
    logic  tt_project_9_ena;
    logic  tt_project_9_clk;
    logic  tt_project_9_rst_n;

    // TT_PROJECT 10 (X5Y5)
    logic [7:0] tt_project_10_ui_in;
    logic [7:0] tt_project_10_uo_out;
    logic [7:0] tt_project_10_uio_in;
    logic [7:0] tt_project_10_uio_out;
    logic [7:0] tt_project_10_uio_oe;
    logic  tt_project_10_ena;
    logic  tt_project_10_clk;
    logic  tt_project_10_rst_n;

    // TT_PROJECT 11 (X5Y6)
    logic [7:0] tt_project_11_ui_in;
    logic [7:0] tt_project_11_uo_out;
    logic [7:0] tt_project_11_uio_in;
    logic [7:0] tt_project_11_uio_out;
    logic [7:0] tt_project_11_uio_oe;
    logic  tt_project_11_ena;
    logic  tt_project_11_clk;
    logic  tt_project_11_rst_n;

    // TT_PROJECT 12 (X5Y7)
    logic [7:0] tt_project_12_ui_in;
    logic [7:0] tt_project_12_uo_out;
    logic [7:0] tt_project_12_uio_in;
    logic [7:0] tt_project_12_uio_out;
    logic [7:0] tt_project_12_uio_oe;
    logic  tt_project_12_ena;
    logic  tt_project_12_clk;
    logic  tt_project_12_rst_n;

    // TT_PROJECT 13 (X5Y8)
    logic [7:0] tt_project_13_ui_in;
    logic [7:0] tt_project_13_uo_out;
    logic [7:0] tt_project_13_uio_in;
    logic [7:0] tt_project_13_uio_out;
    logic [7:0] tt_project_13_uio_oe;
    logic  tt_project_13_ena;
    logic  tt_project_13_clk;
    logic  tt_project_13_rst_n;
    
    eFPGA
    //#(
    //    .MaxFramesPerCol(MaxFramesPerCol),
    //    .FrameBitsPerRow(FrameBitsPerRow)
    //)
    eFPGA
    (
        .FrameData      (FrameData_i),
        .FrameStrobe    (FrameStrobe_i),
        .UserCLK        (clk_i),

        // North I/Os
        .Tile_X1Y0_A_O_top(io_north_in_i[0]),
        .Tile_X1Y0_A_I_top(io_north_out_o[0]),
        .Tile_X1Y0_A_T_top(io_north_oe_o[0]),

        .Tile_X1Y0_B_O_top(io_north_in_i[1]),
        .Tile_X1Y0_B_I_top(io_north_out_o[1]),
        .Tile_X1Y0_B_T_top(io_north_oe_o[1]),

        .Tile_X1Y0_C_O_top(io_north_in_i[2]),
        .Tile_X1Y0_C_I_top(io_north_out_o[2]),
        .Tile_X1Y0_C_T_top(io_north_oe_o[2]),

        .Tile_X1Y0_D_O_top(io_north_in_i[3]),
        .Tile_X1Y0_D_I_top(io_north_out_o[3]),
        .Tile_X1Y0_D_T_top(io_north_oe_o[3]),

        .Tile_X2Y0_A_O_top(io_north_in_i[4]),
        .Tile_X2Y0_A_I_top(io_north_out_o[4]),
        .Tile_X2Y0_A_T_top(io_north_oe_o[4]),

        .Tile_X2Y0_B_O_top(io_north_in_i[5]),
        .Tile_X2Y0_B_I_top(io_north_out_o[5]),
        .Tile_X2Y0_B_T_top(io_north_oe_o[5]),

        .Tile_X2Y0_C_O_top(io_north_in_i[6]),
        .Tile_X2Y0_C_I_top(io_north_out_o[6]),
        .Tile_X2Y0_C_T_top(io_north_oe_o[6]),

        .Tile_X2Y0_D_O_top(io_north_in_i[7]),
        .Tile_X2Y0_D_I_top(io_north_out_o[7]),
        .Tile_X2Y0_D_T_top(io_north_oe_o[7]),

        .Tile_X3Y0_A_O_top(io_north_in_i[8]),
        .Tile_X3Y0_A_I_top(io_north_out_o[8]),
        .Tile_X3Y0_A_T_top(io_north_oe_o[8]),

        .Tile_X3Y0_B_O_top(io_north_in_i[9]),
        .Tile_X3Y0_B_I_top(io_north_out_o[9]),
        .Tile_X3Y0_B_T_top(io_north_oe_o[9]),

        .Tile_X3Y0_C_O_top(io_north_in_i[10]),
        .Tile_X3Y0_C_I_top(io_north_out_o[10]),
        .Tile_X3Y0_C_T_top(io_north_oe_o[10]),

        .Tile_X3Y0_D_O_top(io_north_in_i[11]),
        .Tile_X3Y0_D_I_top(io_north_out_o[11]),
        .Tile_X3Y0_D_T_top(io_north_oe_o[11]),

        .Tile_X4Y0_A_O_top(io_north_in_i[12]),
        .Tile_X4Y0_A_I_top(io_north_out_o[12]),
        .Tile_X4Y0_A_T_top(io_north_oe_o[12]),

        .Tile_X4Y0_B_O_top(io_north_in_i[13]),
        .Tile_X4Y0_B_I_top(io_north_out_o[13]),
        .Tile_X4Y0_B_T_top(io_north_oe_o[13]),

        .Tile_X4Y0_C_O_top(io_north_in_i[14]),
        .Tile_X4Y0_C_I_top(io_north_out_o[14]),
        .Tile_X4Y0_C_T_top(io_north_oe_o[14]),

        .Tile_X4Y0_D_O_top(io_north_in_i[15]),
        .Tile_X4Y0_D_I_top(io_north_out_o[15]),
        .Tile_X4Y0_D_T_top(io_north_oe_o[15]),

        // South I/Os
        .Tile_X1Y9_A_O_top(io_south_in_i[0]),
        .Tile_X1Y9_A_I_top(io_south_out_o[0]),
        .Tile_X1Y9_A_T_top(io_south_oe_o[0]),

        .Tile_X1Y9_B_O_top(io_south_in_i[1]),
        .Tile_X1Y9_B_I_top(io_south_out_o[1]),
        .Tile_X1Y9_B_T_top(io_south_oe_o[1]),

        .Tile_X1Y9_C_O_top(io_south_in_i[2]),
        .Tile_X1Y9_C_I_top(io_south_out_o[2]),
        .Tile_X1Y9_C_T_top(io_south_oe_o[2]),

        .Tile_X1Y9_D_O_top(io_south_in_i[3]),
        .Tile_X1Y9_D_I_top(io_south_out_o[3]),
        .Tile_X1Y9_D_T_top(io_south_oe_o[3]),

        .Tile_X2Y9_A_O_top(io_south_in_i[4]),
        .Tile_X2Y9_A_I_top(io_south_out_o[4]),
        .Tile_X2Y9_A_T_top(io_south_oe_o[4]),

        .Tile_X2Y9_B_O_top(io_south_in_i[5]),
        .Tile_X2Y9_B_I_top(io_south_out_o[5]),
        .Tile_X2Y9_B_T_top(io_south_oe_o[5]),

        .Tile_X2Y9_C_O_top(io_south_in_i[6]),
        .Tile_X2Y9_C_I_top(io_south_out_o[6]),
        .Tile_X2Y9_C_T_top(io_south_oe_o[6]),

        .Tile_X2Y9_D_O_top(io_south_in_i[7]),
        .Tile_X2Y9_D_I_top(io_south_out_o[7]),
        .Tile_X2Y9_D_T_top(io_south_oe_o[7]),

        .Tile_X3Y9_A_O_top(io_south_in_i[8]),
        .Tile_X3Y9_A_I_top(io_south_out_o[8]),
        .Tile_X3Y9_A_T_top(io_south_oe_o[8]),

        .Tile_X3Y9_B_O_top(io_south_in_i[9]),
        .Tile_X3Y9_B_I_top(io_south_out_o[9]),
        .Tile_X3Y9_B_T_top(io_south_oe_o[9]),

        .Tile_X3Y9_C_O_top(io_south_in_i[10]),
        .Tile_X3Y9_C_I_top(io_south_out_o[10]),
        .Tile_X3Y9_C_T_top(io_south_oe_o[10]),

        .Tile_X3Y9_D_O_top(io_south_in_i[11]),
        .Tile_X3Y9_D_I_top(io_south_out_o[11]),
        .Tile_X3Y9_D_T_top(io_south_oe_o[11]),

        .Tile_X4Y9_A_O_top(io_south_in_i[12]),
        .Tile_X4Y9_A_I_top(io_south_out_o[12]),
        .Tile_X4Y9_A_T_top(io_south_oe_o[12]),

        .Tile_X4Y9_B_O_top(io_south_in_i[13]),
        .Tile_X4Y9_B_I_top(io_south_out_o[13]),
        .Tile_X4Y9_B_T_top(io_south_oe_o[13]),

        .Tile_X4Y9_C_O_top(io_south_in_i[14]),
        .Tile_X4Y9_C_I_top(io_south_out_o[14]),
        .Tile_X4Y9_C_T_top(io_south_oe_o[14]),

        .Tile_X4Y9_D_O_top(io_south_in_i[15]),
        .Tile_X4Y9_D_I_top(io_south_out_o[15]),
        .Tile_X4Y9_D_T_top(io_south_oe_o[15]),
        
        // TT_PROJECT 0 (X0Y1)
        .Tile_X0Y1_UI_IN_TT_PROJECT0(tt_project_0_ui_in[0]),
        .Tile_X0Y1_UI_IN_TT_PROJECT1(tt_project_0_ui_in[1]),
        .Tile_X0Y1_UI_IN_TT_PROJECT2(tt_project_0_ui_in[2]),
        .Tile_X0Y1_UI_IN_TT_PROJECT3(tt_project_0_ui_in[3]),
        .Tile_X0Y1_UI_IN_TT_PROJECT4(tt_project_0_ui_in[4]),
        .Tile_X0Y1_UI_IN_TT_PROJECT5(tt_project_0_ui_in[5]),
        .Tile_X0Y1_UI_IN_TT_PROJECT6(tt_project_0_ui_in[6]),
        .Tile_X0Y1_UI_IN_TT_PROJECT7(tt_project_0_ui_in[7]),
        .Tile_X0Y1_UO_OUT_TT_PROJECT0(tt_project_0_uo_out[0]),
        .Tile_X0Y1_UO_OUT_TT_PROJECT1(tt_project_0_uo_out[1]),
        .Tile_X0Y1_UO_OUT_TT_PROJECT2(tt_project_0_uo_out[2]),
        .Tile_X0Y1_UO_OUT_TT_PROJECT3(tt_project_0_uo_out[3]),
        .Tile_X0Y1_UO_OUT_TT_PROJECT4(tt_project_0_uo_out[4]),
        .Tile_X0Y1_UO_OUT_TT_PROJECT5(tt_project_0_uo_out[5]),
        .Tile_X0Y1_UO_OUT_TT_PROJECT6(tt_project_0_uo_out[6]),
        .Tile_X0Y1_UO_OUT_TT_PROJECT7(tt_project_0_uo_out[7]),
        .Tile_X0Y1_UIO_IN_TT_PROJECT0(tt_project_0_uio_in[0]),
        .Tile_X0Y1_UIO_IN_TT_PROJECT1(tt_project_0_uio_in[1]),
        .Tile_X0Y1_UIO_IN_TT_PROJECT2(tt_project_0_uio_in[2]),
        .Tile_X0Y1_UIO_IN_TT_PROJECT3(tt_project_0_uio_in[3]),
        .Tile_X0Y1_UIO_IN_TT_PROJECT4(tt_project_0_uio_in[4]),
        .Tile_X0Y1_UIO_IN_TT_PROJECT5(tt_project_0_uio_in[5]),
        .Tile_X0Y1_UIO_IN_TT_PROJECT6(tt_project_0_uio_in[6]),
        .Tile_X0Y1_UIO_IN_TT_PROJECT7(tt_project_0_uio_in[7]),
        .Tile_X0Y1_UIO_OUT_TT_PROJECT0(tt_project_0_uio_out[0]),
        .Tile_X0Y1_UIO_OUT_TT_PROJECT1(tt_project_0_uio_out[1]),
        .Tile_X0Y1_UIO_OUT_TT_PROJECT2(tt_project_0_uio_out[2]),
        .Tile_X0Y1_UIO_OUT_TT_PROJECT3(tt_project_0_uio_out[3]),
        .Tile_X0Y1_UIO_OUT_TT_PROJECT4(tt_project_0_uio_out[4]),
        .Tile_X0Y1_UIO_OUT_TT_PROJECT5(tt_project_0_uio_out[5]),
        .Tile_X0Y1_UIO_OUT_TT_PROJECT6(tt_project_0_uio_out[6]),
        .Tile_X0Y1_UIO_OUT_TT_PROJECT7(tt_project_0_uio_out[7]),
        .Tile_X0Y1_UIO_OE_TT_PROJECT0(tt_project_0_uio_oe[0]),
        .Tile_X0Y1_UIO_OE_TT_PROJECT1(tt_project_0_uio_oe[1]),
        .Tile_X0Y1_UIO_OE_TT_PROJECT2(tt_project_0_uio_oe[2]),
        .Tile_X0Y1_UIO_OE_TT_PROJECT3(tt_project_0_uio_oe[3]),
        .Tile_X0Y1_UIO_OE_TT_PROJECT4(tt_project_0_uio_oe[4]),
        .Tile_X0Y1_UIO_OE_TT_PROJECT5(tt_project_0_uio_oe[5]),
        .Tile_X0Y1_UIO_OE_TT_PROJECT6(tt_project_0_uio_oe[6]),
        .Tile_X0Y1_UIO_OE_TT_PROJECT7(tt_project_0_uio_oe[7]),
        .Tile_X0Y1_ENA_TT_PROJECT(tt_project_0_ena),
        .Tile_X0Y1_CLK_TT_PROJECT(tt_project_0_clk),
        .Tile_X0Y1_RST_N_TT_PROJECT(tt_project_0_rst_n),

        // TT_PROJECT 1 (X0Y2)
        .Tile_X0Y2_UI_IN_TT_PROJECT0(tt_project_1_ui_in[0]),
        .Tile_X0Y2_UI_IN_TT_PROJECT1(tt_project_1_ui_in[1]),
        .Tile_X0Y2_UI_IN_TT_PROJECT2(tt_project_1_ui_in[2]),
        .Tile_X0Y2_UI_IN_TT_PROJECT3(tt_project_1_ui_in[3]),
        .Tile_X0Y2_UI_IN_TT_PROJECT4(tt_project_1_ui_in[4]),
        .Tile_X0Y2_UI_IN_TT_PROJECT5(tt_project_1_ui_in[5]),
        .Tile_X0Y2_UI_IN_TT_PROJECT6(tt_project_1_ui_in[6]),
        .Tile_X0Y2_UI_IN_TT_PROJECT7(tt_project_1_ui_in[7]),
        .Tile_X0Y2_UO_OUT_TT_PROJECT0(tt_project_1_uo_out[0]),
        .Tile_X0Y2_UO_OUT_TT_PROJECT1(tt_project_1_uo_out[1]),
        .Tile_X0Y2_UO_OUT_TT_PROJECT2(tt_project_1_uo_out[2]),
        .Tile_X0Y2_UO_OUT_TT_PROJECT3(tt_project_1_uo_out[3]),
        .Tile_X0Y2_UO_OUT_TT_PROJECT4(tt_project_1_uo_out[4]),
        .Tile_X0Y2_UO_OUT_TT_PROJECT5(tt_project_1_uo_out[5]),
        .Tile_X0Y2_UO_OUT_TT_PROJECT6(tt_project_1_uo_out[6]),
        .Tile_X0Y2_UO_OUT_TT_PROJECT7(tt_project_1_uo_out[7]),
        .Tile_X0Y2_UIO_IN_TT_PROJECT0(tt_project_1_uio_in[0]),
        .Tile_X0Y2_UIO_IN_TT_PROJECT1(tt_project_1_uio_in[1]),
        .Tile_X0Y2_UIO_IN_TT_PROJECT2(tt_project_1_uio_in[2]),
        .Tile_X0Y2_UIO_IN_TT_PROJECT3(tt_project_1_uio_in[3]),
        .Tile_X0Y2_UIO_IN_TT_PROJECT4(tt_project_1_uio_in[4]),
        .Tile_X0Y2_UIO_IN_TT_PROJECT5(tt_project_1_uio_in[5]),
        .Tile_X0Y2_UIO_IN_TT_PROJECT6(tt_project_1_uio_in[6]),
        .Tile_X0Y2_UIO_IN_TT_PROJECT7(tt_project_1_uio_in[7]),
        .Tile_X0Y2_UIO_OUT_TT_PROJECT0(tt_project_1_uio_out[0]),
        .Tile_X0Y2_UIO_OUT_TT_PROJECT1(tt_project_1_uio_out[1]),
        .Tile_X0Y2_UIO_OUT_TT_PROJECT2(tt_project_1_uio_out[2]),
        .Tile_X0Y2_UIO_OUT_TT_PROJECT3(tt_project_1_uio_out[3]),
        .Tile_X0Y2_UIO_OUT_TT_PROJECT4(tt_project_1_uio_out[4]),
        .Tile_X0Y2_UIO_OUT_TT_PROJECT5(tt_project_1_uio_out[5]),
        .Tile_X0Y2_UIO_OUT_TT_PROJECT6(tt_project_1_uio_out[6]),
        .Tile_X0Y2_UIO_OUT_TT_PROJECT7(tt_project_1_uio_out[7]),
        .Tile_X0Y2_UIO_OE_TT_PROJECT0(tt_project_1_uio_oe[0]),
        .Tile_X0Y2_UIO_OE_TT_PROJECT1(tt_project_1_uio_oe[1]),
        .Tile_X0Y2_UIO_OE_TT_PROJECT2(tt_project_1_uio_oe[2]),
        .Tile_X0Y2_UIO_OE_TT_PROJECT3(tt_project_1_uio_oe[3]),
        .Tile_X0Y2_UIO_OE_TT_PROJECT4(tt_project_1_uio_oe[4]),
        .Tile_X0Y2_UIO_OE_TT_PROJECT5(tt_project_1_uio_oe[5]),
        .Tile_X0Y2_UIO_OE_TT_PROJECT6(tt_project_1_uio_oe[6]),
        .Tile_X0Y2_UIO_OE_TT_PROJECT7(tt_project_1_uio_oe[7]),
        .Tile_X0Y2_ENA_TT_PROJECT(tt_project_1_ena),
        .Tile_X0Y2_CLK_TT_PROJECT(tt_project_1_clk),
        .Tile_X0Y2_RST_N_TT_PROJECT(tt_project_1_rst_n),

        // TT_PROJECT 2 (X0Y3)
        .Tile_X0Y3_UI_IN_TT_PROJECT0(tt_project_2_ui_in[0]),
        .Tile_X0Y3_UI_IN_TT_PROJECT1(tt_project_2_ui_in[1]),
        .Tile_X0Y3_UI_IN_TT_PROJECT2(tt_project_2_ui_in[2]),
        .Tile_X0Y3_UI_IN_TT_PROJECT3(tt_project_2_ui_in[3]),
        .Tile_X0Y3_UI_IN_TT_PROJECT4(tt_project_2_ui_in[4]),
        .Tile_X0Y3_UI_IN_TT_PROJECT5(tt_project_2_ui_in[5]),
        .Tile_X0Y3_UI_IN_TT_PROJECT6(tt_project_2_ui_in[6]),
        .Tile_X0Y3_UI_IN_TT_PROJECT7(tt_project_2_ui_in[7]),
        .Tile_X0Y3_UO_OUT_TT_PROJECT0(tt_project_2_uo_out[0]),
        .Tile_X0Y3_UO_OUT_TT_PROJECT1(tt_project_2_uo_out[1]),
        .Tile_X0Y3_UO_OUT_TT_PROJECT2(tt_project_2_uo_out[2]),
        .Tile_X0Y3_UO_OUT_TT_PROJECT3(tt_project_2_uo_out[3]),
        .Tile_X0Y3_UO_OUT_TT_PROJECT4(tt_project_2_uo_out[4]),
        .Tile_X0Y3_UO_OUT_TT_PROJECT5(tt_project_2_uo_out[5]),
        .Tile_X0Y3_UO_OUT_TT_PROJECT6(tt_project_2_uo_out[6]),
        .Tile_X0Y3_UO_OUT_TT_PROJECT7(tt_project_2_uo_out[7]),
        .Tile_X0Y3_UIO_IN_TT_PROJECT0(tt_project_2_uio_in[0]),
        .Tile_X0Y3_UIO_IN_TT_PROJECT1(tt_project_2_uio_in[1]),
        .Tile_X0Y3_UIO_IN_TT_PROJECT2(tt_project_2_uio_in[2]),
        .Tile_X0Y3_UIO_IN_TT_PROJECT3(tt_project_2_uio_in[3]),
        .Tile_X0Y3_UIO_IN_TT_PROJECT4(tt_project_2_uio_in[4]),
        .Tile_X0Y3_UIO_IN_TT_PROJECT5(tt_project_2_uio_in[5]),
        .Tile_X0Y3_UIO_IN_TT_PROJECT6(tt_project_2_uio_in[6]),
        .Tile_X0Y3_UIO_IN_TT_PROJECT7(tt_project_2_uio_in[7]),
        .Tile_X0Y3_UIO_OUT_TT_PROJECT0(tt_project_2_uio_out[0]),
        .Tile_X0Y3_UIO_OUT_TT_PROJECT1(tt_project_2_uio_out[1]),
        .Tile_X0Y3_UIO_OUT_TT_PROJECT2(tt_project_2_uio_out[2]),
        .Tile_X0Y3_UIO_OUT_TT_PROJECT3(tt_project_2_uio_out[3]),
        .Tile_X0Y3_UIO_OUT_TT_PROJECT4(tt_project_2_uio_out[4]),
        .Tile_X0Y3_UIO_OUT_TT_PROJECT5(tt_project_2_uio_out[5]),
        .Tile_X0Y3_UIO_OUT_TT_PROJECT6(tt_project_2_uio_out[6]),
        .Tile_X0Y3_UIO_OUT_TT_PROJECT7(tt_project_2_uio_out[7]),
        .Tile_X0Y3_UIO_OE_TT_PROJECT0(tt_project_2_uio_oe[0]),
        .Tile_X0Y3_UIO_OE_TT_PROJECT1(tt_project_2_uio_oe[1]),
        .Tile_X0Y3_UIO_OE_TT_PROJECT2(tt_project_2_uio_oe[2]),
        .Tile_X0Y3_UIO_OE_TT_PROJECT3(tt_project_2_uio_oe[3]),
        .Tile_X0Y3_UIO_OE_TT_PROJECT4(tt_project_2_uio_oe[4]),
        .Tile_X0Y3_UIO_OE_TT_PROJECT5(tt_project_2_uio_oe[5]),
        .Tile_X0Y3_UIO_OE_TT_PROJECT6(tt_project_2_uio_oe[6]),
        .Tile_X0Y3_UIO_OE_TT_PROJECT7(tt_project_2_uio_oe[7]),
        .Tile_X0Y3_ENA_TT_PROJECT(tt_project_2_ena),
        .Tile_X0Y3_CLK_TT_PROJECT(tt_project_2_clk),
        .Tile_X0Y3_RST_N_TT_PROJECT(tt_project_2_rst_n),

        // TT_PROJECT 3 (X0Y4)
        .Tile_X0Y4_UI_IN_TT_PROJECT0(tt_project_3_ui_in[0]),
        .Tile_X0Y4_UI_IN_TT_PROJECT1(tt_project_3_ui_in[1]),
        .Tile_X0Y4_UI_IN_TT_PROJECT2(tt_project_3_ui_in[2]),
        .Tile_X0Y4_UI_IN_TT_PROJECT3(tt_project_3_ui_in[3]),
        .Tile_X0Y4_UI_IN_TT_PROJECT4(tt_project_3_ui_in[4]),
        .Tile_X0Y4_UI_IN_TT_PROJECT5(tt_project_3_ui_in[5]),
        .Tile_X0Y4_UI_IN_TT_PROJECT6(tt_project_3_ui_in[6]),
        .Tile_X0Y4_UI_IN_TT_PROJECT7(tt_project_3_ui_in[7]),
        .Tile_X0Y4_UO_OUT_TT_PROJECT0(tt_project_3_uo_out[0]),
        .Tile_X0Y4_UO_OUT_TT_PROJECT1(tt_project_3_uo_out[1]),
        .Tile_X0Y4_UO_OUT_TT_PROJECT2(tt_project_3_uo_out[2]),
        .Tile_X0Y4_UO_OUT_TT_PROJECT3(tt_project_3_uo_out[3]),
        .Tile_X0Y4_UO_OUT_TT_PROJECT4(tt_project_3_uo_out[4]),
        .Tile_X0Y4_UO_OUT_TT_PROJECT5(tt_project_3_uo_out[5]),
        .Tile_X0Y4_UO_OUT_TT_PROJECT6(tt_project_3_uo_out[6]),
        .Tile_X0Y4_UO_OUT_TT_PROJECT7(tt_project_3_uo_out[7]),
        .Tile_X0Y4_UIO_IN_TT_PROJECT0(tt_project_3_uio_in[0]),
        .Tile_X0Y4_UIO_IN_TT_PROJECT1(tt_project_3_uio_in[1]),
        .Tile_X0Y4_UIO_IN_TT_PROJECT2(tt_project_3_uio_in[2]),
        .Tile_X0Y4_UIO_IN_TT_PROJECT3(tt_project_3_uio_in[3]),
        .Tile_X0Y4_UIO_IN_TT_PROJECT4(tt_project_3_uio_in[4]),
        .Tile_X0Y4_UIO_IN_TT_PROJECT5(tt_project_3_uio_in[5]),
        .Tile_X0Y4_UIO_IN_TT_PROJECT6(tt_project_3_uio_in[6]),
        .Tile_X0Y4_UIO_IN_TT_PROJECT7(tt_project_3_uio_in[7]),
        .Tile_X0Y4_UIO_OUT_TT_PROJECT0(tt_project_3_uio_out[0]),
        .Tile_X0Y4_UIO_OUT_TT_PROJECT1(tt_project_3_uio_out[1]),
        .Tile_X0Y4_UIO_OUT_TT_PROJECT2(tt_project_3_uio_out[2]),
        .Tile_X0Y4_UIO_OUT_TT_PROJECT3(tt_project_3_uio_out[3]),
        .Tile_X0Y4_UIO_OUT_TT_PROJECT4(tt_project_3_uio_out[4]),
        .Tile_X0Y4_UIO_OUT_TT_PROJECT5(tt_project_3_uio_out[5]),
        .Tile_X0Y4_UIO_OUT_TT_PROJECT6(tt_project_3_uio_out[6]),
        .Tile_X0Y4_UIO_OUT_TT_PROJECT7(tt_project_3_uio_out[7]),
        .Tile_X0Y4_UIO_OE_TT_PROJECT0(tt_project_3_uio_oe[0]),
        .Tile_X0Y4_UIO_OE_TT_PROJECT1(tt_project_3_uio_oe[1]),
        .Tile_X0Y4_UIO_OE_TT_PROJECT2(tt_project_3_uio_oe[2]),
        .Tile_X0Y4_UIO_OE_TT_PROJECT3(tt_project_3_uio_oe[3]),
        .Tile_X0Y4_UIO_OE_TT_PROJECT4(tt_project_3_uio_oe[4]),
        .Tile_X0Y4_UIO_OE_TT_PROJECT5(tt_project_3_uio_oe[5]),
        .Tile_X0Y4_UIO_OE_TT_PROJECT6(tt_project_3_uio_oe[6]),
        .Tile_X0Y4_UIO_OE_TT_PROJECT7(tt_project_3_uio_oe[7]),
        .Tile_X0Y4_ENA_TT_PROJECT(tt_project_3_ena),
        .Tile_X0Y4_CLK_TT_PROJECT(tt_project_3_clk),
        .Tile_X0Y4_RST_N_TT_PROJECT(tt_project_3_rst_n),

        // TT_PROJECT 4 (X0Y5)
        .Tile_X0Y5_UI_IN_TT_PROJECT0(tt_project_4_ui_in[0]),
        .Tile_X0Y5_UI_IN_TT_PROJECT1(tt_project_4_ui_in[1]),
        .Tile_X0Y5_UI_IN_TT_PROJECT2(tt_project_4_ui_in[2]),
        .Tile_X0Y5_UI_IN_TT_PROJECT3(tt_project_4_ui_in[3]),
        .Tile_X0Y5_UI_IN_TT_PROJECT4(tt_project_4_ui_in[4]),
        .Tile_X0Y5_UI_IN_TT_PROJECT5(tt_project_4_ui_in[5]),
        .Tile_X0Y5_UI_IN_TT_PROJECT6(tt_project_4_ui_in[6]),
        .Tile_X0Y5_UI_IN_TT_PROJECT7(tt_project_4_ui_in[7]),
        .Tile_X0Y5_UO_OUT_TT_PROJECT0(tt_project_4_uo_out[0]),
        .Tile_X0Y5_UO_OUT_TT_PROJECT1(tt_project_4_uo_out[1]),
        .Tile_X0Y5_UO_OUT_TT_PROJECT2(tt_project_4_uo_out[2]),
        .Tile_X0Y5_UO_OUT_TT_PROJECT3(tt_project_4_uo_out[3]),
        .Tile_X0Y5_UO_OUT_TT_PROJECT4(tt_project_4_uo_out[4]),
        .Tile_X0Y5_UO_OUT_TT_PROJECT5(tt_project_4_uo_out[5]),
        .Tile_X0Y5_UO_OUT_TT_PROJECT6(tt_project_4_uo_out[6]),
        .Tile_X0Y5_UO_OUT_TT_PROJECT7(tt_project_4_uo_out[7]),
        .Tile_X0Y5_UIO_IN_TT_PROJECT0(tt_project_4_uio_in[0]),
        .Tile_X0Y5_UIO_IN_TT_PROJECT1(tt_project_4_uio_in[1]),
        .Tile_X0Y5_UIO_IN_TT_PROJECT2(tt_project_4_uio_in[2]),
        .Tile_X0Y5_UIO_IN_TT_PROJECT3(tt_project_4_uio_in[3]),
        .Tile_X0Y5_UIO_IN_TT_PROJECT4(tt_project_4_uio_in[4]),
        .Tile_X0Y5_UIO_IN_TT_PROJECT5(tt_project_4_uio_in[5]),
        .Tile_X0Y5_UIO_IN_TT_PROJECT6(tt_project_4_uio_in[6]),
        .Tile_X0Y5_UIO_IN_TT_PROJECT7(tt_project_4_uio_in[7]),
        .Tile_X0Y5_UIO_OUT_TT_PROJECT0(tt_project_4_uio_out[0]),
        .Tile_X0Y5_UIO_OUT_TT_PROJECT1(tt_project_4_uio_out[1]),
        .Tile_X0Y5_UIO_OUT_TT_PROJECT2(tt_project_4_uio_out[2]),
        .Tile_X0Y5_UIO_OUT_TT_PROJECT3(tt_project_4_uio_out[3]),
        .Tile_X0Y5_UIO_OUT_TT_PROJECT4(tt_project_4_uio_out[4]),
        .Tile_X0Y5_UIO_OUT_TT_PROJECT5(tt_project_4_uio_out[5]),
        .Tile_X0Y5_UIO_OUT_TT_PROJECT6(tt_project_4_uio_out[6]),
        .Tile_X0Y5_UIO_OUT_TT_PROJECT7(tt_project_4_uio_out[7]),
        .Tile_X0Y5_UIO_OE_TT_PROJECT0(tt_project_4_uio_oe[0]),
        .Tile_X0Y5_UIO_OE_TT_PROJECT1(tt_project_4_uio_oe[1]),
        .Tile_X0Y5_UIO_OE_TT_PROJECT2(tt_project_4_uio_oe[2]),
        .Tile_X0Y5_UIO_OE_TT_PROJECT3(tt_project_4_uio_oe[3]),
        .Tile_X0Y5_UIO_OE_TT_PROJECT4(tt_project_4_uio_oe[4]),
        .Tile_X0Y5_UIO_OE_TT_PROJECT5(tt_project_4_uio_oe[5]),
        .Tile_X0Y5_UIO_OE_TT_PROJECT6(tt_project_4_uio_oe[6]),
        .Tile_X0Y5_UIO_OE_TT_PROJECT7(tt_project_4_uio_oe[7]),
        .Tile_X0Y5_ENA_TT_PROJECT(tt_project_4_ena),
        .Tile_X0Y5_CLK_TT_PROJECT(tt_project_4_clk),
        .Tile_X0Y5_RST_N_TT_PROJECT(tt_project_4_rst_n),

        // TT_PROJECT 5 (X0Y6)
        .Tile_X0Y6_UI_IN_TT_PROJECT0(tt_project_5_ui_in[0]),
        .Tile_X0Y6_UI_IN_TT_PROJECT1(tt_project_5_ui_in[1]),
        .Tile_X0Y6_UI_IN_TT_PROJECT2(tt_project_5_ui_in[2]),
        .Tile_X0Y6_UI_IN_TT_PROJECT3(tt_project_5_ui_in[3]),
        .Tile_X0Y6_UI_IN_TT_PROJECT4(tt_project_5_ui_in[4]),
        .Tile_X0Y6_UI_IN_TT_PROJECT5(tt_project_5_ui_in[5]),
        .Tile_X0Y6_UI_IN_TT_PROJECT6(tt_project_5_ui_in[6]),
        .Tile_X0Y6_UI_IN_TT_PROJECT7(tt_project_5_ui_in[7]),
        .Tile_X0Y6_UO_OUT_TT_PROJECT0(tt_project_5_uo_out[0]),
        .Tile_X0Y6_UO_OUT_TT_PROJECT1(tt_project_5_uo_out[1]),
        .Tile_X0Y6_UO_OUT_TT_PROJECT2(tt_project_5_uo_out[2]),
        .Tile_X0Y6_UO_OUT_TT_PROJECT3(tt_project_5_uo_out[3]),
        .Tile_X0Y6_UO_OUT_TT_PROJECT4(tt_project_5_uo_out[4]),
        .Tile_X0Y6_UO_OUT_TT_PROJECT5(tt_project_5_uo_out[5]),
        .Tile_X0Y6_UO_OUT_TT_PROJECT6(tt_project_5_uo_out[6]),
        .Tile_X0Y6_UO_OUT_TT_PROJECT7(tt_project_5_uo_out[7]),
        .Tile_X0Y6_UIO_IN_TT_PROJECT0(tt_project_5_uio_in[0]),
        .Tile_X0Y6_UIO_IN_TT_PROJECT1(tt_project_5_uio_in[1]),
        .Tile_X0Y6_UIO_IN_TT_PROJECT2(tt_project_5_uio_in[2]),
        .Tile_X0Y6_UIO_IN_TT_PROJECT3(tt_project_5_uio_in[3]),
        .Tile_X0Y6_UIO_IN_TT_PROJECT4(tt_project_5_uio_in[4]),
        .Tile_X0Y6_UIO_IN_TT_PROJECT5(tt_project_5_uio_in[5]),
        .Tile_X0Y6_UIO_IN_TT_PROJECT6(tt_project_5_uio_in[6]),
        .Tile_X0Y6_UIO_IN_TT_PROJECT7(tt_project_5_uio_in[7]),
        .Tile_X0Y6_UIO_OUT_TT_PROJECT0(tt_project_5_uio_out[0]),
        .Tile_X0Y6_UIO_OUT_TT_PROJECT1(tt_project_5_uio_out[1]),
        .Tile_X0Y6_UIO_OUT_TT_PROJECT2(tt_project_5_uio_out[2]),
        .Tile_X0Y6_UIO_OUT_TT_PROJECT3(tt_project_5_uio_out[3]),
        .Tile_X0Y6_UIO_OUT_TT_PROJECT4(tt_project_5_uio_out[4]),
        .Tile_X0Y6_UIO_OUT_TT_PROJECT5(tt_project_5_uio_out[5]),
        .Tile_X0Y6_UIO_OUT_TT_PROJECT6(tt_project_5_uio_out[6]),
        .Tile_X0Y6_UIO_OUT_TT_PROJECT7(tt_project_5_uio_out[7]),
        .Tile_X0Y6_UIO_OE_TT_PROJECT0(tt_project_5_uio_oe[0]),
        .Tile_X0Y6_UIO_OE_TT_PROJECT1(tt_project_5_uio_oe[1]),
        .Tile_X0Y6_UIO_OE_TT_PROJECT2(tt_project_5_uio_oe[2]),
        .Tile_X0Y6_UIO_OE_TT_PROJECT3(tt_project_5_uio_oe[3]),
        .Tile_X0Y6_UIO_OE_TT_PROJECT4(tt_project_5_uio_oe[4]),
        .Tile_X0Y6_UIO_OE_TT_PROJECT5(tt_project_5_uio_oe[5]),
        .Tile_X0Y6_UIO_OE_TT_PROJECT6(tt_project_5_uio_oe[6]),
        .Tile_X0Y6_UIO_OE_TT_PROJECT7(tt_project_5_uio_oe[7]),
        .Tile_X0Y6_ENA_TT_PROJECT(tt_project_5_ena),
        .Tile_X0Y6_CLK_TT_PROJECT(tt_project_5_clk),
        .Tile_X0Y6_RST_N_TT_PROJECT(tt_project_5_rst_n),

        // TT_PROJECT 6 (X0Y7)
        .Tile_X0Y7_UI_IN_TT_PROJECT0(tt_project_6_ui_in[0]),
        .Tile_X0Y7_UI_IN_TT_PROJECT1(tt_project_6_ui_in[1]),
        .Tile_X0Y7_UI_IN_TT_PROJECT2(tt_project_6_ui_in[2]),
        .Tile_X0Y7_UI_IN_TT_PROJECT3(tt_project_6_ui_in[3]),
        .Tile_X0Y7_UI_IN_TT_PROJECT4(tt_project_6_ui_in[4]),
        .Tile_X0Y7_UI_IN_TT_PROJECT5(tt_project_6_ui_in[5]),
        .Tile_X0Y7_UI_IN_TT_PROJECT6(tt_project_6_ui_in[6]),
        .Tile_X0Y7_UI_IN_TT_PROJECT7(tt_project_6_ui_in[7]),
        .Tile_X0Y7_UO_OUT_TT_PROJECT0(tt_project_6_uo_out[0]),
        .Tile_X0Y7_UO_OUT_TT_PROJECT1(tt_project_6_uo_out[1]),
        .Tile_X0Y7_UO_OUT_TT_PROJECT2(tt_project_6_uo_out[2]),
        .Tile_X0Y7_UO_OUT_TT_PROJECT3(tt_project_6_uo_out[3]),
        .Tile_X0Y7_UO_OUT_TT_PROJECT4(tt_project_6_uo_out[4]),
        .Tile_X0Y7_UO_OUT_TT_PROJECT5(tt_project_6_uo_out[5]),
        .Tile_X0Y7_UO_OUT_TT_PROJECT6(tt_project_6_uo_out[6]),
        .Tile_X0Y7_UO_OUT_TT_PROJECT7(tt_project_6_uo_out[7]),
        .Tile_X0Y7_UIO_IN_TT_PROJECT0(tt_project_6_uio_in[0]),
        .Tile_X0Y7_UIO_IN_TT_PROJECT1(tt_project_6_uio_in[1]),
        .Tile_X0Y7_UIO_IN_TT_PROJECT2(tt_project_6_uio_in[2]),
        .Tile_X0Y7_UIO_IN_TT_PROJECT3(tt_project_6_uio_in[3]),
        .Tile_X0Y7_UIO_IN_TT_PROJECT4(tt_project_6_uio_in[4]),
        .Tile_X0Y7_UIO_IN_TT_PROJECT5(tt_project_6_uio_in[5]),
        .Tile_X0Y7_UIO_IN_TT_PROJECT6(tt_project_6_uio_in[6]),
        .Tile_X0Y7_UIO_IN_TT_PROJECT7(tt_project_6_uio_in[7]),
        .Tile_X0Y7_UIO_OUT_TT_PROJECT0(tt_project_6_uio_out[0]),
        .Tile_X0Y7_UIO_OUT_TT_PROJECT1(tt_project_6_uio_out[1]),
        .Tile_X0Y7_UIO_OUT_TT_PROJECT2(tt_project_6_uio_out[2]),
        .Tile_X0Y7_UIO_OUT_TT_PROJECT3(tt_project_6_uio_out[3]),
        .Tile_X0Y7_UIO_OUT_TT_PROJECT4(tt_project_6_uio_out[4]),
        .Tile_X0Y7_UIO_OUT_TT_PROJECT5(tt_project_6_uio_out[5]),
        .Tile_X0Y7_UIO_OUT_TT_PROJECT6(tt_project_6_uio_out[6]),
        .Tile_X0Y7_UIO_OUT_TT_PROJECT7(tt_project_6_uio_out[7]),
        .Tile_X0Y7_UIO_OE_TT_PROJECT0(tt_project_6_uio_oe[0]),
        .Tile_X0Y7_UIO_OE_TT_PROJECT1(tt_project_6_uio_oe[1]),
        .Tile_X0Y7_UIO_OE_TT_PROJECT2(tt_project_6_uio_oe[2]),
        .Tile_X0Y7_UIO_OE_TT_PROJECT3(tt_project_6_uio_oe[3]),
        .Tile_X0Y7_UIO_OE_TT_PROJECT4(tt_project_6_uio_oe[4]),
        .Tile_X0Y7_UIO_OE_TT_PROJECT5(tt_project_6_uio_oe[5]),
        .Tile_X0Y7_UIO_OE_TT_PROJECT6(tt_project_6_uio_oe[6]),
        .Tile_X0Y7_UIO_OE_TT_PROJECT7(tt_project_6_uio_oe[7]),
        .Tile_X0Y7_ENA_TT_PROJECT(tt_project_6_ena),
        .Tile_X0Y7_CLK_TT_PROJECT(tt_project_6_clk),
        .Tile_X0Y7_RST_N_TT_PROJECT(tt_project_6_rst_n),

        // TT_PROJECT 7 (X0Y8)
        .Tile_X0Y8_UI_IN_TT_PROJECT0(tt_project_7_ui_in[0]),
        .Tile_X0Y8_UI_IN_TT_PROJECT1(tt_project_7_ui_in[1]),
        .Tile_X0Y8_UI_IN_TT_PROJECT2(tt_project_7_ui_in[2]),
        .Tile_X0Y8_UI_IN_TT_PROJECT3(tt_project_7_ui_in[3]),
        .Tile_X0Y8_UI_IN_TT_PROJECT4(tt_project_7_ui_in[4]),
        .Tile_X0Y8_UI_IN_TT_PROJECT5(tt_project_7_ui_in[5]),
        .Tile_X0Y8_UI_IN_TT_PROJECT6(tt_project_7_ui_in[6]),
        .Tile_X0Y8_UI_IN_TT_PROJECT7(tt_project_7_ui_in[7]),
        .Tile_X0Y8_UO_OUT_TT_PROJECT0(tt_project_7_uo_out[0]),
        .Tile_X0Y8_UO_OUT_TT_PROJECT1(tt_project_7_uo_out[1]),
        .Tile_X0Y8_UO_OUT_TT_PROJECT2(tt_project_7_uo_out[2]),
        .Tile_X0Y8_UO_OUT_TT_PROJECT3(tt_project_7_uo_out[3]),
        .Tile_X0Y8_UO_OUT_TT_PROJECT4(tt_project_7_uo_out[4]),
        .Tile_X0Y8_UO_OUT_TT_PROJECT5(tt_project_7_uo_out[5]),
        .Tile_X0Y8_UO_OUT_TT_PROJECT6(tt_project_7_uo_out[6]),
        .Tile_X0Y8_UO_OUT_TT_PROJECT7(tt_project_7_uo_out[7]),
        .Tile_X0Y8_UIO_IN_TT_PROJECT0(tt_project_7_uio_in[0]),
        .Tile_X0Y8_UIO_IN_TT_PROJECT1(tt_project_7_uio_in[1]),
        .Tile_X0Y8_UIO_IN_TT_PROJECT2(tt_project_7_uio_in[2]),
        .Tile_X0Y8_UIO_IN_TT_PROJECT3(tt_project_7_uio_in[3]),
        .Tile_X0Y8_UIO_IN_TT_PROJECT4(tt_project_7_uio_in[4]),
        .Tile_X0Y8_UIO_IN_TT_PROJECT5(tt_project_7_uio_in[5]),
        .Tile_X0Y8_UIO_IN_TT_PROJECT6(tt_project_7_uio_in[6]),
        .Tile_X0Y8_UIO_IN_TT_PROJECT7(tt_project_7_uio_in[7]),
        .Tile_X0Y8_UIO_OUT_TT_PROJECT0(tt_project_7_uio_out[0]),
        .Tile_X0Y8_UIO_OUT_TT_PROJECT1(tt_project_7_uio_out[1]),
        .Tile_X0Y8_UIO_OUT_TT_PROJECT2(tt_project_7_uio_out[2]),
        .Tile_X0Y8_UIO_OUT_TT_PROJECT3(tt_project_7_uio_out[3]),
        .Tile_X0Y8_UIO_OUT_TT_PROJECT4(tt_project_7_uio_out[4]),
        .Tile_X0Y8_UIO_OUT_TT_PROJECT5(tt_project_7_uio_out[5]),
        .Tile_X0Y8_UIO_OUT_TT_PROJECT6(tt_project_7_uio_out[6]),
        .Tile_X0Y8_UIO_OUT_TT_PROJECT7(tt_project_7_uio_out[7]),
        .Tile_X0Y8_UIO_OE_TT_PROJECT0(tt_project_7_uio_oe[0]),
        .Tile_X0Y8_UIO_OE_TT_PROJECT1(tt_project_7_uio_oe[1]),
        .Tile_X0Y8_UIO_OE_TT_PROJECT2(tt_project_7_uio_oe[2]),
        .Tile_X0Y8_UIO_OE_TT_PROJECT3(tt_project_7_uio_oe[3]),
        .Tile_X0Y8_UIO_OE_TT_PROJECT4(tt_project_7_uio_oe[4]),
        .Tile_X0Y8_UIO_OE_TT_PROJECT5(tt_project_7_uio_oe[5]),
        .Tile_X0Y8_UIO_OE_TT_PROJECT6(tt_project_7_uio_oe[6]),
        .Tile_X0Y8_UIO_OE_TT_PROJECT7(tt_project_7_uio_oe[7]),
        .Tile_X0Y8_ENA_TT_PROJECT(tt_project_7_ena),
        .Tile_X0Y8_CLK_TT_PROJECT(tt_project_7_clk),
        .Tile_X0Y8_RST_N_TT_PROJECT(tt_project_7_rst_n),

        // TT_PROJECT 8 (X5Y3)
        .Tile_X5Y3_UI_IN_TT_PROJECT0(tt_project_8_ui_in[0]),
        .Tile_X5Y3_UI_IN_TT_PROJECT1(tt_project_8_ui_in[1]),
        .Tile_X5Y3_UI_IN_TT_PROJECT2(tt_project_8_ui_in[2]),
        .Tile_X5Y3_UI_IN_TT_PROJECT3(tt_project_8_ui_in[3]),
        .Tile_X5Y3_UI_IN_TT_PROJECT4(tt_project_8_ui_in[4]),
        .Tile_X5Y3_UI_IN_TT_PROJECT5(tt_project_8_ui_in[5]),
        .Tile_X5Y3_UI_IN_TT_PROJECT6(tt_project_8_ui_in[6]),
        .Tile_X5Y3_UI_IN_TT_PROJECT7(tt_project_8_ui_in[7]),
        .Tile_X5Y3_UO_OUT_TT_PROJECT0(tt_project_8_uo_out[0]),
        .Tile_X5Y3_UO_OUT_TT_PROJECT1(tt_project_8_uo_out[1]),
        .Tile_X5Y3_UO_OUT_TT_PROJECT2(tt_project_8_uo_out[2]),
        .Tile_X5Y3_UO_OUT_TT_PROJECT3(tt_project_8_uo_out[3]),
        .Tile_X5Y3_UO_OUT_TT_PROJECT4(tt_project_8_uo_out[4]),
        .Tile_X5Y3_UO_OUT_TT_PROJECT5(tt_project_8_uo_out[5]),
        .Tile_X5Y3_UO_OUT_TT_PROJECT6(tt_project_8_uo_out[6]),
        .Tile_X5Y3_UO_OUT_TT_PROJECT7(tt_project_8_uo_out[7]),
        .Tile_X5Y3_UIO_IN_TT_PROJECT0(tt_project_8_uio_in[0]),
        .Tile_X5Y3_UIO_IN_TT_PROJECT1(tt_project_8_uio_in[1]),
        .Tile_X5Y3_UIO_IN_TT_PROJECT2(tt_project_8_uio_in[2]),
        .Tile_X5Y3_UIO_IN_TT_PROJECT3(tt_project_8_uio_in[3]),
        .Tile_X5Y3_UIO_IN_TT_PROJECT4(tt_project_8_uio_in[4]),
        .Tile_X5Y3_UIO_IN_TT_PROJECT5(tt_project_8_uio_in[5]),
        .Tile_X5Y3_UIO_IN_TT_PROJECT6(tt_project_8_uio_in[6]),
        .Tile_X5Y3_UIO_IN_TT_PROJECT7(tt_project_8_uio_in[7]),
        .Tile_X5Y3_UIO_OUT_TT_PROJECT0(tt_project_8_uio_out[0]),
        .Tile_X5Y3_UIO_OUT_TT_PROJECT1(tt_project_8_uio_out[1]),
        .Tile_X5Y3_UIO_OUT_TT_PROJECT2(tt_project_8_uio_out[2]),
        .Tile_X5Y3_UIO_OUT_TT_PROJECT3(tt_project_8_uio_out[3]),
        .Tile_X5Y3_UIO_OUT_TT_PROJECT4(tt_project_8_uio_out[4]),
        .Tile_X5Y3_UIO_OUT_TT_PROJECT5(tt_project_8_uio_out[5]),
        .Tile_X5Y3_UIO_OUT_TT_PROJECT6(tt_project_8_uio_out[6]),
        .Tile_X5Y3_UIO_OUT_TT_PROJECT7(tt_project_8_uio_out[7]),
        .Tile_X5Y3_UIO_OE_TT_PROJECT0(tt_project_8_uio_oe[0]),
        .Tile_X5Y3_UIO_OE_TT_PROJECT1(tt_project_8_uio_oe[1]),
        .Tile_X5Y3_UIO_OE_TT_PROJECT2(tt_project_8_uio_oe[2]),
        .Tile_X5Y3_UIO_OE_TT_PROJECT3(tt_project_8_uio_oe[3]),
        .Tile_X5Y3_UIO_OE_TT_PROJECT4(tt_project_8_uio_oe[4]),
        .Tile_X5Y3_UIO_OE_TT_PROJECT5(tt_project_8_uio_oe[5]),
        .Tile_X5Y3_UIO_OE_TT_PROJECT6(tt_project_8_uio_oe[6]),
        .Tile_X5Y3_UIO_OE_TT_PROJECT7(tt_project_8_uio_oe[7]),
        .Tile_X5Y3_ENA_TT_PROJECT(tt_project_8_ena),
        .Tile_X5Y3_CLK_TT_PROJECT(tt_project_8_clk),
        .Tile_X5Y3_RST_N_TT_PROJECT(tt_project_8_rst_n),

        // TT_PROJECT 9 (X5Y4)
        .Tile_X5Y4_UI_IN_TT_PROJECT0(tt_project_9_ui_in[0]),
        .Tile_X5Y4_UI_IN_TT_PROJECT1(tt_project_9_ui_in[1]),
        .Tile_X5Y4_UI_IN_TT_PROJECT2(tt_project_9_ui_in[2]),
        .Tile_X5Y4_UI_IN_TT_PROJECT3(tt_project_9_ui_in[3]),
        .Tile_X5Y4_UI_IN_TT_PROJECT4(tt_project_9_ui_in[4]),
        .Tile_X5Y4_UI_IN_TT_PROJECT5(tt_project_9_ui_in[5]),
        .Tile_X5Y4_UI_IN_TT_PROJECT6(tt_project_9_ui_in[6]),
        .Tile_X5Y4_UI_IN_TT_PROJECT7(tt_project_9_ui_in[7]),
        .Tile_X5Y4_UO_OUT_TT_PROJECT0(tt_project_9_uo_out[0]),
        .Tile_X5Y4_UO_OUT_TT_PROJECT1(tt_project_9_uo_out[1]),
        .Tile_X5Y4_UO_OUT_TT_PROJECT2(tt_project_9_uo_out[2]),
        .Tile_X5Y4_UO_OUT_TT_PROJECT3(tt_project_9_uo_out[3]),
        .Tile_X5Y4_UO_OUT_TT_PROJECT4(tt_project_9_uo_out[4]),
        .Tile_X5Y4_UO_OUT_TT_PROJECT5(tt_project_9_uo_out[5]),
        .Tile_X5Y4_UO_OUT_TT_PROJECT6(tt_project_9_uo_out[6]),
        .Tile_X5Y4_UO_OUT_TT_PROJECT7(tt_project_9_uo_out[7]),
        .Tile_X5Y4_UIO_IN_TT_PROJECT0(tt_project_9_uio_in[0]),
        .Tile_X5Y4_UIO_IN_TT_PROJECT1(tt_project_9_uio_in[1]),
        .Tile_X5Y4_UIO_IN_TT_PROJECT2(tt_project_9_uio_in[2]),
        .Tile_X5Y4_UIO_IN_TT_PROJECT3(tt_project_9_uio_in[3]),
        .Tile_X5Y4_UIO_IN_TT_PROJECT4(tt_project_9_uio_in[4]),
        .Tile_X5Y4_UIO_IN_TT_PROJECT5(tt_project_9_uio_in[5]),
        .Tile_X5Y4_UIO_IN_TT_PROJECT6(tt_project_9_uio_in[6]),
        .Tile_X5Y4_UIO_IN_TT_PROJECT7(tt_project_9_uio_in[7]),
        .Tile_X5Y4_UIO_OUT_TT_PROJECT0(tt_project_9_uio_out[0]),
        .Tile_X5Y4_UIO_OUT_TT_PROJECT1(tt_project_9_uio_out[1]),
        .Tile_X5Y4_UIO_OUT_TT_PROJECT2(tt_project_9_uio_out[2]),
        .Tile_X5Y4_UIO_OUT_TT_PROJECT3(tt_project_9_uio_out[3]),
        .Tile_X5Y4_UIO_OUT_TT_PROJECT4(tt_project_9_uio_out[4]),
        .Tile_X5Y4_UIO_OUT_TT_PROJECT5(tt_project_9_uio_out[5]),
        .Tile_X5Y4_UIO_OUT_TT_PROJECT6(tt_project_9_uio_out[6]),
        .Tile_X5Y4_UIO_OUT_TT_PROJECT7(tt_project_9_uio_out[7]),
        .Tile_X5Y4_UIO_OE_TT_PROJECT0(tt_project_9_uio_oe[0]),
        .Tile_X5Y4_UIO_OE_TT_PROJECT1(tt_project_9_uio_oe[1]),
        .Tile_X5Y4_UIO_OE_TT_PROJECT2(tt_project_9_uio_oe[2]),
        .Tile_X5Y4_UIO_OE_TT_PROJECT3(tt_project_9_uio_oe[3]),
        .Tile_X5Y4_UIO_OE_TT_PROJECT4(tt_project_9_uio_oe[4]),
        .Tile_X5Y4_UIO_OE_TT_PROJECT5(tt_project_9_uio_oe[5]),
        .Tile_X5Y4_UIO_OE_TT_PROJECT6(tt_project_9_uio_oe[6]),
        .Tile_X5Y4_UIO_OE_TT_PROJECT7(tt_project_9_uio_oe[7]),
        .Tile_X5Y4_ENA_TT_PROJECT(tt_project_9_ena),
        .Tile_X5Y4_CLK_TT_PROJECT(tt_project_9_clk),
        .Tile_X5Y4_RST_N_TT_PROJECT(tt_project_9_rst_n),

        // TT_PROJECT 10 (X5Y5)
        .Tile_X5Y5_UI_IN_TT_PROJECT0(tt_project_10_ui_in[0]),
        .Tile_X5Y5_UI_IN_TT_PROJECT1(tt_project_10_ui_in[1]),
        .Tile_X5Y5_UI_IN_TT_PROJECT2(tt_project_10_ui_in[2]),
        .Tile_X5Y5_UI_IN_TT_PROJECT3(tt_project_10_ui_in[3]),
        .Tile_X5Y5_UI_IN_TT_PROJECT4(tt_project_10_ui_in[4]),
        .Tile_X5Y5_UI_IN_TT_PROJECT5(tt_project_10_ui_in[5]),
        .Tile_X5Y5_UI_IN_TT_PROJECT6(tt_project_10_ui_in[6]),
        .Tile_X5Y5_UI_IN_TT_PROJECT7(tt_project_10_ui_in[7]),
        .Tile_X5Y5_UO_OUT_TT_PROJECT0(tt_project_10_uo_out[0]),
        .Tile_X5Y5_UO_OUT_TT_PROJECT1(tt_project_10_uo_out[1]),
        .Tile_X5Y5_UO_OUT_TT_PROJECT2(tt_project_10_uo_out[2]),
        .Tile_X5Y5_UO_OUT_TT_PROJECT3(tt_project_10_uo_out[3]),
        .Tile_X5Y5_UO_OUT_TT_PROJECT4(tt_project_10_uo_out[4]),
        .Tile_X5Y5_UO_OUT_TT_PROJECT5(tt_project_10_uo_out[5]),
        .Tile_X5Y5_UO_OUT_TT_PROJECT6(tt_project_10_uo_out[6]),
        .Tile_X5Y5_UO_OUT_TT_PROJECT7(tt_project_10_uo_out[7]),
        .Tile_X5Y5_UIO_IN_TT_PROJECT0(tt_project_10_uio_in[0]),
        .Tile_X5Y5_UIO_IN_TT_PROJECT1(tt_project_10_uio_in[1]),
        .Tile_X5Y5_UIO_IN_TT_PROJECT2(tt_project_10_uio_in[2]),
        .Tile_X5Y5_UIO_IN_TT_PROJECT3(tt_project_10_uio_in[3]),
        .Tile_X5Y5_UIO_IN_TT_PROJECT4(tt_project_10_uio_in[4]),
        .Tile_X5Y5_UIO_IN_TT_PROJECT5(tt_project_10_uio_in[5]),
        .Tile_X5Y5_UIO_IN_TT_PROJECT6(tt_project_10_uio_in[6]),
        .Tile_X5Y5_UIO_IN_TT_PROJECT7(tt_project_10_uio_in[7]),
        .Tile_X5Y5_UIO_OUT_TT_PROJECT0(tt_project_10_uio_out[0]),
        .Tile_X5Y5_UIO_OUT_TT_PROJECT1(tt_project_10_uio_out[1]),
        .Tile_X5Y5_UIO_OUT_TT_PROJECT2(tt_project_10_uio_out[2]),
        .Tile_X5Y5_UIO_OUT_TT_PROJECT3(tt_project_10_uio_out[3]),
        .Tile_X5Y5_UIO_OUT_TT_PROJECT4(tt_project_10_uio_out[4]),
        .Tile_X5Y5_UIO_OUT_TT_PROJECT5(tt_project_10_uio_out[5]),
        .Tile_X5Y5_UIO_OUT_TT_PROJECT6(tt_project_10_uio_out[6]),
        .Tile_X5Y5_UIO_OUT_TT_PROJECT7(tt_project_10_uio_out[7]),
        .Tile_X5Y5_UIO_OE_TT_PROJECT0(tt_project_10_uio_oe[0]),
        .Tile_X5Y5_UIO_OE_TT_PROJECT1(tt_project_10_uio_oe[1]),
        .Tile_X5Y5_UIO_OE_TT_PROJECT2(tt_project_10_uio_oe[2]),
        .Tile_X5Y5_UIO_OE_TT_PROJECT3(tt_project_10_uio_oe[3]),
        .Tile_X5Y5_UIO_OE_TT_PROJECT4(tt_project_10_uio_oe[4]),
        .Tile_X5Y5_UIO_OE_TT_PROJECT5(tt_project_10_uio_oe[5]),
        .Tile_X5Y5_UIO_OE_TT_PROJECT6(tt_project_10_uio_oe[6]),
        .Tile_X5Y5_UIO_OE_TT_PROJECT7(tt_project_10_uio_oe[7]),
        .Tile_X5Y5_ENA_TT_PROJECT(tt_project_10_ena),
        .Tile_X5Y5_CLK_TT_PROJECT(tt_project_10_clk),
        .Tile_X5Y5_RST_N_TT_PROJECT(tt_project_10_rst_n),

        // TT_PROJECT 11 (X5Y6)
        .Tile_X5Y6_UI_IN_TT_PROJECT0(tt_project_11_ui_in[0]),
        .Tile_X5Y6_UI_IN_TT_PROJECT1(tt_project_11_ui_in[1]),
        .Tile_X5Y6_UI_IN_TT_PROJECT2(tt_project_11_ui_in[2]),
        .Tile_X5Y6_UI_IN_TT_PROJECT3(tt_project_11_ui_in[3]),
        .Tile_X5Y6_UI_IN_TT_PROJECT4(tt_project_11_ui_in[4]),
        .Tile_X5Y6_UI_IN_TT_PROJECT5(tt_project_11_ui_in[5]),
        .Tile_X5Y6_UI_IN_TT_PROJECT6(tt_project_11_ui_in[6]),
        .Tile_X5Y6_UI_IN_TT_PROJECT7(tt_project_11_ui_in[7]),
        .Tile_X5Y6_UO_OUT_TT_PROJECT0(tt_project_11_uo_out[0]),
        .Tile_X5Y6_UO_OUT_TT_PROJECT1(tt_project_11_uo_out[1]),
        .Tile_X5Y6_UO_OUT_TT_PROJECT2(tt_project_11_uo_out[2]),
        .Tile_X5Y6_UO_OUT_TT_PROJECT3(tt_project_11_uo_out[3]),
        .Tile_X5Y6_UO_OUT_TT_PROJECT4(tt_project_11_uo_out[4]),
        .Tile_X5Y6_UO_OUT_TT_PROJECT5(tt_project_11_uo_out[5]),
        .Tile_X5Y6_UO_OUT_TT_PROJECT6(tt_project_11_uo_out[6]),
        .Tile_X5Y6_UO_OUT_TT_PROJECT7(tt_project_11_uo_out[7]),
        .Tile_X5Y6_UIO_IN_TT_PROJECT0(tt_project_11_uio_in[0]),
        .Tile_X5Y6_UIO_IN_TT_PROJECT1(tt_project_11_uio_in[1]),
        .Tile_X5Y6_UIO_IN_TT_PROJECT2(tt_project_11_uio_in[2]),
        .Tile_X5Y6_UIO_IN_TT_PROJECT3(tt_project_11_uio_in[3]),
        .Tile_X5Y6_UIO_IN_TT_PROJECT4(tt_project_11_uio_in[4]),
        .Tile_X5Y6_UIO_IN_TT_PROJECT5(tt_project_11_uio_in[5]),
        .Tile_X5Y6_UIO_IN_TT_PROJECT6(tt_project_11_uio_in[6]),
        .Tile_X5Y6_UIO_IN_TT_PROJECT7(tt_project_11_uio_in[7]),
        .Tile_X5Y6_UIO_OUT_TT_PROJECT0(tt_project_11_uio_out[0]),
        .Tile_X5Y6_UIO_OUT_TT_PROJECT1(tt_project_11_uio_out[1]),
        .Tile_X5Y6_UIO_OUT_TT_PROJECT2(tt_project_11_uio_out[2]),
        .Tile_X5Y6_UIO_OUT_TT_PROJECT3(tt_project_11_uio_out[3]),
        .Tile_X5Y6_UIO_OUT_TT_PROJECT4(tt_project_11_uio_out[4]),
        .Tile_X5Y6_UIO_OUT_TT_PROJECT5(tt_project_11_uio_out[5]),
        .Tile_X5Y6_UIO_OUT_TT_PROJECT6(tt_project_11_uio_out[6]),
        .Tile_X5Y6_UIO_OUT_TT_PROJECT7(tt_project_11_uio_out[7]),
        .Tile_X5Y6_UIO_OE_TT_PROJECT0(tt_project_11_uio_oe[0]),
        .Tile_X5Y6_UIO_OE_TT_PROJECT1(tt_project_11_uio_oe[1]),
        .Tile_X5Y6_UIO_OE_TT_PROJECT2(tt_project_11_uio_oe[2]),
        .Tile_X5Y6_UIO_OE_TT_PROJECT3(tt_project_11_uio_oe[3]),
        .Tile_X5Y6_UIO_OE_TT_PROJECT4(tt_project_11_uio_oe[4]),
        .Tile_X5Y6_UIO_OE_TT_PROJECT5(tt_project_11_uio_oe[5]),
        .Tile_X5Y6_UIO_OE_TT_PROJECT6(tt_project_11_uio_oe[6]),
        .Tile_X5Y6_UIO_OE_TT_PROJECT7(tt_project_11_uio_oe[7]),
        .Tile_X5Y6_ENA_TT_PROJECT(tt_project_11_ena),
        .Tile_X5Y6_CLK_TT_PROJECT(tt_project_11_clk),
        .Tile_X5Y6_RST_N_TT_PROJECT(tt_project_11_rst_n),

        // TT_PROJECT 12 (X5Y7)
        .Tile_X5Y7_UI_IN_TT_PROJECT0(tt_project_12_ui_in[0]),
        .Tile_X5Y7_UI_IN_TT_PROJECT1(tt_project_12_ui_in[1]),
        .Tile_X5Y7_UI_IN_TT_PROJECT2(tt_project_12_ui_in[2]),
        .Tile_X5Y7_UI_IN_TT_PROJECT3(tt_project_12_ui_in[3]),
        .Tile_X5Y7_UI_IN_TT_PROJECT4(tt_project_12_ui_in[4]),
        .Tile_X5Y7_UI_IN_TT_PROJECT5(tt_project_12_ui_in[5]),
        .Tile_X5Y7_UI_IN_TT_PROJECT6(tt_project_12_ui_in[6]),
        .Tile_X5Y7_UI_IN_TT_PROJECT7(tt_project_12_ui_in[7]),
        .Tile_X5Y7_UO_OUT_TT_PROJECT0(tt_project_12_uo_out[0]),
        .Tile_X5Y7_UO_OUT_TT_PROJECT1(tt_project_12_uo_out[1]),
        .Tile_X5Y7_UO_OUT_TT_PROJECT2(tt_project_12_uo_out[2]),
        .Tile_X5Y7_UO_OUT_TT_PROJECT3(tt_project_12_uo_out[3]),
        .Tile_X5Y7_UO_OUT_TT_PROJECT4(tt_project_12_uo_out[4]),
        .Tile_X5Y7_UO_OUT_TT_PROJECT5(tt_project_12_uo_out[5]),
        .Tile_X5Y7_UO_OUT_TT_PROJECT6(tt_project_12_uo_out[6]),
        .Tile_X5Y7_UO_OUT_TT_PROJECT7(tt_project_12_uo_out[7]),
        .Tile_X5Y7_UIO_IN_TT_PROJECT0(tt_project_12_uio_in[0]),
        .Tile_X5Y7_UIO_IN_TT_PROJECT1(tt_project_12_uio_in[1]),
        .Tile_X5Y7_UIO_IN_TT_PROJECT2(tt_project_12_uio_in[2]),
        .Tile_X5Y7_UIO_IN_TT_PROJECT3(tt_project_12_uio_in[3]),
        .Tile_X5Y7_UIO_IN_TT_PROJECT4(tt_project_12_uio_in[4]),
        .Tile_X5Y7_UIO_IN_TT_PROJECT5(tt_project_12_uio_in[5]),
        .Tile_X5Y7_UIO_IN_TT_PROJECT6(tt_project_12_uio_in[6]),
        .Tile_X5Y7_UIO_IN_TT_PROJECT7(tt_project_12_uio_in[7]),
        .Tile_X5Y7_UIO_OUT_TT_PROJECT0(tt_project_12_uio_out[0]),
        .Tile_X5Y7_UIO_OUT_TT_PROJECT1(tt_project_12_uio_out[1]),
        .Tile_X5Y7_UIO_OUT_TT_PROJECT2(tt_project_12_uio_out[2]),
        .Tile_X5Y7_UIO_OUT_TT_PROJECT3(tt_project_12_uio_out[3]),
        .Tile_X5Y7_UIO_OUT_TT_PROJECT4(tt_project_12_uio_out[4]),
        .Tile_X5Y7_UIO_OUT_TT_PROJECT5(tt_project_12_uio_out[5]),
        .Tile_X5Y7_UIO_OUT_TT_PROJECT6(tt_project_12_uio_out[6]),
        .Tile_X5Y7_UIO_OUT_TT_PROJECT7(tt_project_12_uio_out[7]),
        .Tile_X5Y7_UIO_OE_TT_PROJECT0(tt_project_12_uio_oe[0]),
        .Tile_X5Y7_UIO_OE_TT_PROJECT1(tt_project_12_uio_oe[1]),
        .Tile_X5Y7_UIO_OE_TT_PROJECT2(tt_project_12_uio_oe[2]),
        .Tile_X5Y7_UIO_OE_TT_PROJECT3(tt_project_12_uio_oe[3]),
        .Tile_X5Y7_UIO_OE_TT_PROJECT4(tt_project_12_uio_oe[4]),
        .Tile_X5Y7_UIO_OE_TT_PROJECT5(tt_project_12_uio_oe[5]),
        .Tile_X5Y7_UIO_OE_TT_PROJECT6(tt_project_12_uio_oe[6]),
        .Tile_X5Y7_UIO_OE_TT_PROJECT7(tt_project_12_uio_oe[7]),
        .Tile_X5Y7_ENA_TT_PROJECT(tt_project_12_ena),
        .Tile_X5Y7_CLK_TT_PROJECT(tt_project_12_clk),
        .Tile_X5Y7_RST_N_TT_PROJECT(tt_project_12_rst_n),

        // TT_PROJECT 13 (X5Y8)
        .Tile_X5Y8_UI_IN_TT_PROJECT0(tt_project_13_ui_in[0]),
        .Tile_X5Y8_UI_IN_TT_PROJECT1(tt_project_13_ui_in[1]),
        .Tile_X5Y8_UI_IN_TT_PROJECT2(tt_project_13_ui_in[2]),
        .Tile_X5Y8_UI_IN_TT_PROJECT3(tt_project_13_ui_in[3]),
        .Tile_X5Y8_UI_IN_TT_PROJECT4(tt_project_13_ui_in[4]),
        .Tile_X5Y8_UI_IN_TT_PROJECT5(tt_project_13_ui_in[5]),
        .Tile_X5Y8_UI_IN_TT_PROJECT6(tt_project_13_ui_in[6]),
        .Tile_X5Y8_UI_IN_TT_PROJECT7(tt_project_13_ui_in[7]),
        .Tile_X5Y8_UO_OUT_TT_PROJECT0(tt_project_13_uo_out[0]),
        .Tile_X5Y8_UO_OUT_TT_PROJECT1(tt_project_13_uo_out[1]),
        .Tile_X5Y8_UO_OUT_TT_PROJECT2(tt_project_13_uo_out[2]),
        .Tile_X5Y8_UO_OUT_TT_PROJECT3(tt_project_13_uo_out[3]),
        .Tile_X5Y8_UO_OUT_TT_PROJECT4(tt_project_13_uo_out[4]),
        .Tile_X5Y8_UO_OUT_TT_PROJECT5(tt_project_13_uo_out[5]),
        .Tile_X5Y8_UO_OUT_TT_PROJECT6(tt_project_13_uo_out[6]),
        .Tile_X5Y8_UO_OUT_TT_PROJECT7(tt_project_13_uo_out[7]),
        .Tile_X5Y8_UIO_IN_TT_PROJECT0(tt_project_13_uio_in[0]),
        .Tile_X5Y8_UIO_IN_TT_PROJECT1(tt_project_13_uio_in[1]),
        .Tile_X5Y8_UIO_IN_TT_PROJECT2(tt_project_13_uio_in[2]),
        .Tile_X5Y8_UIO_IN_TT_PROJECT3(tt_project_13_uio_in[3]),
        .Tile_X5Y8_UIO_IN_TT_PROJECT4(tt_project_13_uio_in[4]),
        .Tile_X5Y8_UIO_IN_TT_PROJECT5(tt_project_13_uio_in[5]),
        .Tile_X5Y8_UIO_IN_TT_PROJECT6(tt_project_13_uio_in[6]),
        .Tile_X5Y8_UIO_IN_TT_PROJECT7(tt_project_13_uio_in[7]),
        .Tile_X5Y8_UIO_OUT_TT_PROJECT0(tt_project_13_uio_out[0]),
        .Tile_X5Y8_UIO_OUT_TT_PROJECT1(tt_project_13_uio_out[1]),
        .Tile_X5Y8_UIO_OUT_TT_PROJECT2(tt_project_13_uio_out[2]),
        .Tile_X5Y8_UIO_OUT_TT_PROJECT3(tt_project_13_uio_out[3]),
        .Tile_X5Y8_UIO_OUT_TT_PROJECT4(tt_project_13_uio_out[4]),
        .Tile_X5Y8_UIO_OUT_TT_PROJECT5(tt_project_13_uio_out[5]),
        .Tile_X5Y8_UIO_OUT_TT_PROJECT6(tt_project_13_uio_out[6]),
        .Tile_X5Y8_UIO_OUT_TT_PROJECT7(tt_project_13_uio_out[7]),
        .Tile_X5Y8_UIO_OE_TT_PROJECT0(tt_project_13_uio_oe[0]),
        .Tile_X5Y8_UIO_OE_TT_PROJECT1(tt_project_13_uio_oe[1]),
        .Tile_X5Y8_UIO_OE_TT_PROJECT2(tt_project_13_uio_oe[2]),
        .Tile_X5Y8_UIO_OE_TT_PROJECT3(tt_project_13_uio_oe[3]),
        .Tile_X5Y8_UIO_OE_TT_PROJECT4(tt_project_13_uio_oe[4]),
        .Tile_X5Y8_UIO_OE_TT_PROJECT5(tt_project_13_uio_oe[5]),
        .Tile_X5Y8_UIO_OE_TT_PROJECT6(tt_project_13_uio_oe[6]),
        .Tile_X5Y8_UIO_OE_TT_PROJECT7(tt_project_13_uio_oe[7]),
        .Tile_X5Y8_ENA_TT_PROJECT(tt_project_13_ena),
        .Tile_X5Y8_CLK_TT_PROJECT(tt_project_13_clk),
        .Tile_X5Y8_RST_N_TT_PROJECT(tt_project_13_rst_n)
    );

    // TT_PROJECT
    
    heichips25_example_small heichips25_example_small_0 (
        .clk        (tt_project_0_clk),
        .rst_n      (tt_project_0_rst_n),
        .ena        (tt_project_0_ena),
        .ui_in      (tt_project_0_ui_in),
        .uio_in     (tt_project_0_uio_in),
        .uo_out     (tt_project_0_uo_out),
        .uio_out    (tt_project_0_uio_out),
        .uio_oe     (tt_project_0_uio_oe)
    );

    heichips25_example_small heichips25_example_small_1 (
        .clk        (tt_project_1_clk),
        .rst_n      (tt_project_1_rst_n),
        .ena        (tt_project_1_ena),
        .ui_in      (tt_project_1_ui_in),
        .uio_in     (tt_project_1_uio_in),
        .uo_out     (tt_project_1_uo_out),
        .uio_out    (tt_project_1_uio_out),
        .uio_oe     (tt_project_1_uio_oe)
    );

    heichips25_example_small heichips25_example_small_2 (
        .clk        (tt_project_2_clk),
        .rst_n      (tt_project_2_rst_n),
        .ena        (tt_project_2_ena),
        .ui_in      (tt_project_2_ui_in),
        .uio_in     (tt_project_2_uio_in),
        .uo_out     (tt_project_2_uo_out),
        .uio_out    (tt_project_2_uio_out),
        .uio_oe     (tt_project_2_uio_oe)
    );

    heichips25_example_small heichips25_example_small_3 (
        .clk        (tt_project_3_clk),
        .rst_n      (tt_project_3_rst_n),
        .ena        (tt_project_3_ena),
        .ui_in      (tt_project_3_ui_in),
        .uio_in     (tt_project_3_uio_in),
        .uo_out     (tt_project_3_uo_out),
        .uio_out    (tt_project_3_uio_out),
        .uio_oe     (tt_project_3_uio_oe)
    );

    heichips25_example_small heichips25_example_small_4 (
        .clk        (tt_project_4_clk),
        .rst_n      (tt_project_4_rst_n),
        .ena        (tt_project_4_ena),
        .ui_in      (tt_project_4_ui_in),
        .uio_in     (tt_project_4_uio_in),
        .uo_out     (tt_project_4_uo_out),
        .uio_out    (tt_project_4_uio_out),
        .uio_oe     (tt_project_4_uio_oe)
    );

    heichips25_example_small heichips25_example_small_5 (
        .clk        (tt_project_5_clk),
        .rst_n      (tt_project_5_rst_n),
        .ena        (tt_project_5_ena),
        .ui_in      (tt_project_5_ui_in),
        .uio_in     (tt_project_5_uio_in),
        .uo_out     (tt_project_5_uo_out),
        .uio_out    (tt_project_5_uio_out),
        .uio_oe     (tt_project_5_uio_oe)
    );

    heichips25_example_small heichips25_example_small_6 (
        .clk        (tt_project_6_clk),
        .rst_n      (tt_project_6_rst_n),
        .ena        (tt_project_6_ena),
        .ui_in      (tt_project_6_ui_in),
        .uio_in     (tt_project_6_uio_in),
        .uo_out     (tt_project_6_uo_out),
        .uio_out    (tt_project_6_uio_out),
        .uio_oe     (tt_project_6_uio_oe)
    );

    heichips25_example_small heichips25_example_small_7 (
        .clk        (tt_project_7_clk),
        .rst_n      (tt_project_7_rst_n),
        .ena        (tt_project_7_ena),
        .ui_in      (tt_project_7_ui_in),
        .uio_in     (tt_project_7_uio_in),
        .uo_out     (tt_project_7_uo_out),
        .uio_out    (tt_project_7_uio_out),
        .uio_oe     (tt_project_7_uio_oe)
    );

    heichips25_example_small heichips25_example_small_8 (
        .clk        (tt_project_8_clk),
        .rst_n      (tt_project_8_rst_n),
        .ena        (tt_project_8_ena),
        .ui_in      (tt_project_8_ui_in),
        .uio_in     (tt_project_8_uio_in),
        .uo_out     (tt_project_8_uo_out),
        .uio_out    (tt_project_8_uio_out),
        .uio_oe     (tt_project_8_uio_oe)
    );

    heichips25_example_small heichips25_example_small_9 (
        .clk        (tt_project_9_clk),
        .rst_n      (tt_project_9_rst_n),
        .ena        (tt_project_9_ena),
        .ui_in      (tt_project_9_ui_in),
        .uio_in     (tt_project_9_uio_in),
        .uo_out     (tt_project_9_uo_out),
        .uio_out    (tt_project_9_uio_out),
        .uio_oe     (tt_project_9_uio_oe)
    );

    heichips25_example_small heichips25_example_small_10 (
        .clk        (tt_project_10_clk),
        .rst_n      (tt_project_10_rst_n),
        .ena        (tt_project_10_ena),
        .ui_in      (tt_project_10_ui_in),
        .uio_in     (tt_project_10_uio_in),
        .uo_out     (tt_project_10_uo_out),
        .uio_out    (tt_project_10_uio_out),
        .uio_oe     (tt_project_10_uio_oe)
    );

    heichips25_example_small heichips25_example_small_11 (
        .clk        (tt_project_11_clk),
        .rst_n      (tt_project_11_rst_n),
        .ena        (tt_project_11_ena),
        .ui_in      (tt_project_11_ui_in),
        .uio_in     (tt_project_11_uio_in),
        .uo_out     (tt_project_11_uo_out),
        .uio_out    (tt_project_11_uio_out),
        .uio_oe     (tt_project_11_uio_oe)
    );

    heichips25_example_small heichips25_example_small_12 (
        .clk        (tt_project_12_clk),
        .rst_n      (tt_project_12_rst_n),
        .ena        (tt_project_12_ena),
        .ui_in      (tt_project_12_ui_in),
        .uio_in     (tt_project_12_uio_in),
        .uo_out     (tt_project_12_uo_out),
        .uio_out    (tt_project_12_uio_out),
        .uio_oe     (tt_project_12_uio_oe)
    );

    heichips25_example_small heichips25_example_small_13 (
        .clk        (tt_project_13_clk),
        .rst_n      (tt_project_13_rst_n),
        .ena        (tt_project_13_ena),
        .ui_in      (tt_project_13_ui_in),
        .uio_in     (tt_project_13_uio_in),
        .uo_out     (tt_project_13_uo_out),
        .uio_out    (tt_project_13_uio_out),
        .uio_oe     (tt_project_13_uio_oe)
    );


    // SRAMs

endmodule

`default_nettype wire
