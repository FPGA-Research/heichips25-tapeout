module heichips25_example_small (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net25;

 sg13g2_and2_1 _29_ (.A(net1),
    .B(net9),
    .X(_00_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _30_ (.A(net2),
    .B(net10),
    .X(_01_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _31_ (.B(net10),
    .A(net2),
    .X(_02_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _32_ (.B(_02_),
    .A(_00_),
    .X(net18),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _33_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_01_),
    .Y(_03_),
    .A2(_02_),
    .A1(_00_));
 sg13g2_and2_1 _34_ (.A(net3),
    .B(net11),
    .X(_04_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _35_ (.Y(_05_),
    .A(net3),
    .B(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _36_ (.A(_03_),
    .B(_05_),
    .Y(_06_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _37_ (.B(_05_),
    .A(_03_),
    .X(net19),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _38_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_07_),
    .B(net12),
    .A(net4));
 sg13g2_and2_1 _39_ (.A(net4),
    .B(net12),
    .X(_08_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _40_ (.B(net12),
    .A(net4),
    .X(_09_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _41_ (.A(_04_),
    .B(_06_),
    .Y(_10_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _42_ (.Y(net20),
    .A(_09_),
    .B(_10_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _43_ (.Y(_11_),
    .B(_09_),
    .A_N(_05_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _44_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04_),
    .A2(_07_),
    .Y(_12_),
    .B1(_08_));
 sg13g2_o21ai_1 _45_ (.B1(_12_),
    .VDD(VPWR),
    .Y(_13_),
    .VSS(VGND),
    .A1(_03_),
    .A2(_11_));
 sg13g2_nand2_1 _46_ (.Y(_14_),
    .A(net5),
    .B(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _47_ (.B(net13),
    .A(net5),
    .X(_15_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _48_ (.VDD(VPWR),
    .Y(_16_),
    .A(_15_),
    .VSS(VGND));
 sg13g2_nand2_1 _49_ (.Y(_17_),
    .A(_13_),
    .B(_15_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _50_ (.Y(net21),
    .A(_13_),
    .B(_16_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _51_ (.A(net6),
    .B(net14),
    .Y(_18_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _52_ (.Y(_19_),
    .A(net6),
    .B(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _53_ (.Y(_20_),
    .A(_14_),
    .B(_17_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _54_ (.Y(net22),
    .A(_19_),
    .B(_20_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _55_ (.A(_16_),
    .B(_19_),
    .Y(_21_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _56_ (.A(_14_),
    .B(_18_),
    .Y(_22_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _57_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_21_),
    .C1(_22_),
    .B1(_13_),
    .A1(net6),
    .Y(_23_),
    .A2(net14));
 sg13g2_nand2_1 _58_ (.Y(_24_),
    .A(net7),
    .B(net15),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _59_ (.A(net7),
    .B(net15),
    .Y(_25_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _60_ (.B(net15),
    .A(net7),
    .X(_26_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _61_ (.Y(net23),
    .A(_23_),
    .B(_26_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _62_ (.B1(_24_),
    .VDD(VPWR),
    .Y(_27_),
    .VSS(VGND),
    .A1(_23_),
    .A2(_25_));
 sg13g2_xnor2_1 _63_ (.Y(_28_),
    .A(net8),
    .B(net16),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _64_ (.Y(net24),
    .A(_27_),
    .B(_28_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _65_ (.B(net9),
    .A(net1),
    .X(net17),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo heichips25_example_small_26 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net26));
 sg13g2_tielo heichips25_example_small_27 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net27));
 sg13g2_tielo heichips25_example_small_28 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net28));
 sg13g2_tielo heichips25_example_small_29 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net29));
 sg13g2_tielo heichips25_example_small_30 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net30));
 sg13g2_tielo heichips25_example_small_31 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net31));
 sg13g2_tielo heichips25_example_small_32 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net32));
 sg13g2_tielo heichips25_example_small_33 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net33));
 sg13g2_tielo heichips25_example_small_34 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net34));
 sg13g2_tielo heichips25_example_small_35 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net35));
 sg13g2_tielo heichips25_example_small_36 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net36));
 sg13g2_tielo heichips25_example_small_37 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net37));
 sg13g2_tielo heichips25_example_small_38 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net38));
 sg13g2_tielo heichips25_example_small_39 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net39));
 sg13g2_tielo heichips25_example_small_40 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net40));
 sg13g2_decap_8 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input13 (.A(uio_in[4]),
    .X(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input14 (.A(uio_in[5]),
    .X(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input15 (.A(uio_in[6]),
    .X(net15),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input16 (.A(uio_in[7]),
    .X(net16),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo heichips25_example_small_25 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net25));
 sg13g2_decap_8 FILLER_0_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1022 (.VDD(VPWR),
    .VSS(VGND));
 assign uio_oe[0] = net25;
 assign uio_oe[1] = net26;
 assign uio_oe[2] = net27;
 assign uio_oe[3] = net28;
 assign uio_oe[4] = net29;
 assign uio_oe[5] = net30;
 assign uio_oe[6] = net31;
 assign uio_oe[7] = net32;
 assign uio_out[0] = net33;
 assign uio_out[1] = net34;
 assign uio_out[2] = net35;
 assign uio_out[3] = net36;
 assign uio_out[4] = net37;
 assign uio_out[5] = net38;
 assign uio_out[6] = net39;
 assign uio_out[7] = net40;
endmodule
