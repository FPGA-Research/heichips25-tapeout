magic
tech ihp-sg13g2
magscale 1 2
timestamp 1753090738
<< metal1 >>
rect 1152 9848 41856 9872
rect 1152 9808 4928 9848
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 5296 9808 20048 9848
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20416 9808 35168 9848
rect 35208 9808 35250 9848
rect 35290 9808 35332 9848
rect 35372 9808 35414 9848
rect 35454 9808 35496 9848
rect 35536 9808 41856 9848
rect 1152 9784 41856 9808
rect 1411 9680 1469 9681
rect 1411 9640 1420 9680
rect 1460 9640 1469 9680
rect 1411 9639 1469 9640
rect 2179 9680 2237 9681
rect 2179 9640 2188 9680
rect 2228 9640 2237 9680
rect 2179 9639 2237 9640
rect 7459 9680 7517 9681
rect 7459 9640 7468 9680
rect 7508 9640 7517 9680
rect 7459 9639 7517 9640
rect 9379 9680 9437 9681
rect 9379 9640 9388 9680
rect 9428 9640 9437 9680
rect 9379 9639 9437 9640
rect 32235 9680 32277 9689
rect 32235 9640 32236 9680
rect 32276 9640 32277 9680
rect 32235 9631 32277 9640
rect 34539 9680 34581 9689
rect 34539 9640 34540 9680
rect 34580 9640 34581 9680
rect 34539 9631 34581 9640
rect 36555 9680 36597 9689
rect 36555 9640 36556 9680
rect 36596 9640 36597 9680
rect 36555 9631 36597 9640
rect 36939 9680 36981 9689
rect 36939 9640 36940 9680
rect 36980 9640 36981 9680
rect 36939 9631 36981 9640
rect 37323 9680 37365 9689
rect 37323 9640 37324 9680
rect 37364 9640 37365 9680
rect 37323 9631 37365 9640
rect 39339 9680 39381 9689
rect 39339 9640 39340 9680
rect 39380 9640 39381 9680
rect 39339 9631 39381 9640
rect 39723 9680 39765 9689
rect 39723 9640 39724 9680
rect 39764 9640 39765 9680
rect 39723 9631 39765 9640
rect 40107 9680 40149 9689
rect 40107 9640 40108 9680
rect 40148 9640 40149 9680
rect 40107 9631 40149 9640
rect 40683 9680 40725 9689
rect 40683 9640 40684 9680
rect 40724 9640 40725 9680
rect 40683 9631 40725 9640
rect 41067 9680 41109 9689
rect 41067 9640 41068 9680
rect 41108 9640 41109 9680
rect 41067 9631 41109 9640
rect 3819 9596 3861 9605
rect 3819 9556 3820 9596
rect 3860 9556 3861 9596
rect 3819 9547 3861 9556
rect 1515 9512 1557 9521
rect 1515 9472 1516 9512
rect 1556 9472 1557 9512
rect 1515 9463 1557 9472
rect 1611 9512 1653 9521
rect 1611 9472 1612 9512
rect 1652 9472 1653 9512
rect 1611 9463 1653 9472
rect 1707 9512 1749 9521
rect 1707 9472 1708 9512
rect 1748 9472 1749 9512
rect 1707 9463 1749 9472
rect 1899 9512 1941 9521
rect 1899 9472 1900 9512
rect 1940 9472 1941 9512
rect 1899 9463 1941 9472
rect 1995 9512 2037 9521
rect 1995 9472 1996 9512
rect 2036 9472 2037 9512
rect 1995 9463 2037 9472
rect 2371 9512 2429 9513
rect 2371 9472 2380 9512
rect 2420 9472 2429 9512
rect 2371 9471 2429 9472
rect 3619 9512 3677 9513
rect 3619 9472 3628 9512
rect 3668 9472 3677 9512
rect 3619 9471 3677 9472
rect 4286 9512 4344 9513
rect 4286 9472 4295 9512
rect 4335 9472 4344 9512
rect 4286 9471 4344 9472
rect 4395 9512 4437 9521
rect 4395 9472 4396 9512
rect 4436 9472 4437 9512
rect 4395 9463 4437 9472
rect 4491 9512 4533 9521
rect 4491 9472 4492 9512
rect 4532 9472 4533 9512
rect 4491 9463 4533 9472
rect 4675 9512 4733 9513
rect 4675 9472 4684 9512
rect 4724 9472 4733 9512
rect 4675 9471 4733 9472
rect 4771 9512 4829 9513
rect 4771 9472 4780 9512
rect 4820 9472 4829 9512
rect 4771 9471 4829 9472
rect 4963 9512 5021 9513
rect 4963 9472 4972 9512
rect 5012 9472 5021 9512
rect 4963 9471 5021 9472
rect 5443 9512 5501 9513
rect 5443 9472 5452 9512
rect 5492 9472 5501 9512
rect 5443 9471 5501 9472
rect 6691 9512 6749 9513
rect 6691 9472 6700 9512
rect 6740 9472 6749 9512
rect 6691 9471 6749 9472
rect 6979 9512 7037 9513
rect 6979 9472 6988 9512
rect 7028 9472 7037 9512
rect 6979 9471 7037 9472
rect 7179 9512 7221 9521
rect 7179 9472 7180 9512
rect 7220 9472 7221 9512
rect 7179 9463 7221 9472
rect 7275 9512 7317 9521
rect 7275 9472 7276 9512
rect 7316 9472 7317 9512
rect 7275 9463 7317 9472
rect 7659 9512 7701 9521
rect 7659 9472 7660 9512
rect 7700 9472 7701 9512
rect 7659 9463 7701 9472
rect 7755 9512 7797 9521
rect 7755 9472 7756 9512
rect 7796 9472 7797 9512
rect 7755 9463 7797 9472
rect 7851 9512 7893 9521
rect 7851 9472 7852 9512
rect 7892 9472 7893 9512
rect 7851 9463 7893 9472
rect 7947 9512 7989 9521
rect 7947 9472 7948 9512
rect 7988 9472 7989 9512
rect 7947 9463 7989 9472
rect 8331 9512 8373 9521
rect 8331 9472 8332 9512
rect 8372 9472 8373 9512
rect 8331 9463 8373 9472
rect 8619 9512 8661 9521
rect 8619 9472 8620 9512
rect 8660 9472 8661 9512
rect 8619 9463 8661 9472
rect 8715 9512 8757 9521
rect 8715 9472 8716 9512
rect 8756 9472 8757 9512
rect 8715 9463 8757 9472
rect 8811 9512 8853 9521
rect 8811 9472 8812 9512
rect 8852 9472 8853 9512
rect 8811 9463 8853 9472
rect 8907 9512 8949 9521
rect 8907 9472 8908 9512
rect 8948 9472 8949 9512
rect 8907 9463 8949 9472
rect 9099 9512 9141 9521
rect 9099 9472 9100 9512
rect 9140 9472 9141 9512
rect 9099 9463 9141 9472
rect 9195 9512 9237 9521
rect 9195 9472 9196 9512
rect 9236 9472 9237 9512
rect 9195 9463 9237 9472
rect 9859 9512 9917 9513
rect 9859 9472 9868 9512
rect 9908 9472 9917 9512
rect 9859 9471 9917 9472
rect 11107 9512 11165 9513
rect 11107 9472 11116 9512
rect 11156 9472 11165 9512
rect 11107 9471 11165 9472
rect 11491 9512 11549 9513
rect 11491 9472 11500 9512
rect 11540 9472 11549 9512
rect 11491 9471 11549 9472
rect 12739 9512 12797 9513
rect 12739 9472 12748 9512
rect 12788 9472 12797 9512
rect 12739 9471 12797 9472
rect 13123 9512 13181 9513
rect 13123 9472 13132 9512
rect 13172 9472 13181 9512
rect 13123 9471 13181 9472
rect 14371 9512 14429 9513
rect 14371 9472 14380 9512
rect 14420 9472 14429 9512
rect 14371 9471 14429 9472
rect 14755 9512 14813 9513
rect 14755 9472 14764 9512
rect 14804 9472 14813 9512
rect 14755 9471 14813 9472
rect 16003 9512 16061 9513
rect 16003 9472 16012 9512
rect 16052 9472 16061 9512
rect 16003 9471 16061 9472
rect 16387 9512 16445 9513
rect 16387 9472 16396 9512
rect 16436 9472 16445 9512
rect 16387 9471 16445 9472
rect 17635 9512 17693 9513
rect 17635 9472 17644 9512
rect 17684 9472 17693 9512
rect 17635 9471 17693 9472
rect 18115 9512 18173 9513
rect 18115 9472 18124 9512
rect 18164 9472 18173 9512
rect 18115 9471 18173 9472
rect 19363 9512 19421 9513
rect 19363 9472 19372 9512
rect 19412 9472 19421 9512
rect 19363 9471 19421 9472
rect 19747 9512 19805 9513
rect 19747 9472 19756 9512
rect 19796 9472 19805 9512
rect 19747 9471 19805 9472
rect 20995 9512 21053 9513
rect 20995 9472 21004 9512
rect 21044 9472 21053 9512
rect 20995 9471 21053 9472
rect 21379 9512 21437 9513
rect 21379 9472 21388 9512
rect 21428 9472 21437 9512
rect 21379 9471 21437 9472
rect 22627 9512 22685 9513
rect 22627 9472 22636 9512
rect 22676 9472 22685 9512
rect 22627 9471 22685 9472
rect 23203 9512 23261 9513
rect 23203 9472 23212 9512
rect 23252 9472 23261 9512
rect 23203 9471 23261 9472
rect 24451 9512 24509 9513
rect 24451 9472 24460 9512
rect 24500 9472 24509 9512
rect 24451 9471 24509 9472
rect 25027 9512 25085 9513
rect 25027 9472 25036 9512
rect 25076 9472 25085 9512
rect 25027 9471 25085 9472
rect 26275 9512 26333 9513
rect 26275 9472 26284 9512
rect 26324 9472 26333 9512
rect 26275 9471 26333 9472
rect 26659 9512 26717 9513
rect 26659 9472 26668 9512
rect 26708 9472 26717 9512
rect 26659 9471 26717 9472
rect 27907 9512 27965 9513
rect 27907 9472 27916 9512
rect 27956 9472 27965 9512
rect 27907 9471 27965 9472
rect 28291 9512 28349 9513
rect 28291 9472 28300 9512
rect 28340 9472 28349 9512
rect 28291 9471 28349 9472
rect 29539 9512 29597 9513
rect 29539 9472 29548 9512
rect 29588 9472 29597 9512
rect 29539 9471 29597 9472
rect 30691 9512 30749 9513
rect 30691 9472 30700 9512
rect 30740 9472 30749 9512
rect 30691 9471 30749 9472
rect 31851 9512 31893 9521
rect 31851 9472 31852 9512
rect 31892 9472 31893 9512
rect 31851 9463 31893 9472
rect 32899 9512 32957 9513
rect 32899 9472 32908 9512
rect 32948 9472 32957 9512
rect 32899 9471 32957 9472
rect 34147 9512 34205 9513
rect 34147 9472 34156 9512
rect 34196 9472 34205 9512
rect 34147 9471 34205 9472
rect 34915 9512 34973 9513
rect 34915 9472 34924 9512
rect 34964 9472 34973 9512
rect 34915 9471 34973 9472
rect 36163 9512 36221 9513
rect 36163 9472 36172 9512
rect 36212 9472 36221 9512
rect 36163 9471 36221 9472
rect 37699 9512 37757 9513
rect 37699 9472 37708 9512
rect 37748 9472 37757 9512
rect 37699 9471 37757 9472
rect 38947 9512 39005 9513
rect 38947 9472 38956 9512
rect 38996 9472 39005 9512
rect 38947 9471 39005 9472
rect 31083 9428 31125 9437
rect 31083 9388 31084 9428
rect 31124 9388 31125 9428
rect 31083 9379 31125 9388
rect 32419 9428 32477 9429
rect 32419 9388 32428 9428
rect 32468 9388 32477 9428
rect 32419 9387 32477 9388
rect 34723 9428 34781 9429
rect 34723 9388 34732 9428
rect 34772 9388 34781 9428
rect 34723 9387 34781 9388
rect 36739 9428 36797 9429
rect 36739 9388 36748 9428
rect 36788 9388 36797 9428
rect 36739 9387 36797 9388
rect 37123 9428 37181 9429
rect 37123 9388 37132 9428
rect 37172 9388 37181 9428
rect 37123 9387 37181 9388
rect 37507 9428 37565 9429
rect 37507 9388 37516 9428
rect 37556 9388 37565 9428
rect 37507 9387 37565 9388
rect 39523 9428 39581 9429
rect 39523 9388 39532 9428
rect 39572 9388 39581 9428
rect 39523 9387 39581 9388
rect 39907 9428 39965 9429
rect 39907 9388 39916 9428
rect 39956 9388 39965 9428
rect 39907 9387 39965 9388
rect 40291 9428 40349 9429
rect 40291 9388 40300 9428
rect 40340 9388 40349 9428
rect 40291 9387 40349 9388
rect 40483 9428 40541 9429
rect 40483 9388 40492 9428
rect 40532 9388 40541 9428
rect 40483 9387 40541 9388
rect 40867 9428 40925 9429
rect 40867 9388 40876 9428
rect 40916 9388 40925 9428
rect 40867 9387 40925 9388
rect 41251 9428 41309 9429
rect 41251 9388 41260 9428
rect 41300 9388 41309 9428
rect 41251 9387 41309 9388
rect 5259 9344 5301 9353
rect 5259 9304 5260 9344
rect 5300 9304 5301 9344
rect 5259 9295 5301 9304
rect 8331 9344 8373 9353
rect 8331 9304 8332 9344
rect 8372 9304 8373 9344
rect 8331 9295 8373 9304
rect 41451 9344 41493 9353
rect 41451 9304 41452 9344
rect 41492 9304 41493 9344
rect 41451 9295 41493 9304
rect 4779 9260 4821 9269
rect 4779 9220 4780 9260
rect 4820 9220 4821 9260
rect 4779 9211 4821 9220
rect 5067 9260 5109 9269
rect 5067 9220 5068 9260
rect 5108 9220 5109 9260
rect 5067 9211 5109 9220
rect 6891 9260 6933 9269
rect 6891 9220 6892 9260
rect 6932 9220 6933 9260
rect 6891 9211 6933 9220
rect 8139 9260 8181 9269
rect 8139 9220 8140 9260
rect 8180 9220 8181 9260
rect 8139 9211 8181 9220
rect 11307 9260 11349 9269
rect 11307 9220 11308 9260
rect 11348 9220 11349 9260
rect 11307 9211 11349 9220
rect 12939 9260 12981 9269
rect 12939 9220 12940 9260
rect 12980 9220 12981 9260
rect 12939 9211 12981 9220
rect 14571 9260 14613 9269
rect 14571 9220 14572 9260
rect 14612 9220 14613 9260
rect 14571 9211 14613 9220
rect 16203 9260 16245 9269
rect 16203 9220 16204 9260
rect 16244 9220 16245 9260
rect 16203 9211 16245 9220
rect 17835 9260 17877 9269
rect 17835 9220 17836 9260
rect 17876 9220 17877 9260
rect 17835 9211 17877 9220
rect 19563 9260 19605 9269
rect 19563 9220 19564 9260
rect 19604 9220 19605 9260
rect 19563 9211 19605 9220
rect 21195 9260 21237 9269
rect 21195 9220 21196 9260
rect 21236 9220 21237 9260
rect 21195 9211 21237 9220
rect 22827 9260 22869 9269
rect 22827 9220 22828 9260
rect 22868 9220 22869 9260
rect 22827 9211 22869 9220
rect 24651 9260 24693 9269
rect 24651 9220 24652 9260
rect 24692 9220 24693 9260
rect 24651 9211 24693 9220
rect 24843 9260 24885 9269
rect 24843 9220 24844 9260
rect 24884 9220 24885 9260
rect 24843 9211 24885 9220
rect 26475 9260 26517 9269
rect 26475 9220 26476 9260
rect 26516 9220 26517 9260
rect 26475 9211 26517 9220
rect 28107 9260 28149 9269
rect 28107 9220 28108 9260
rect 28148 9220 28149 9260
rect 28107 9211 28149 9220
rect 30219 9260 30261 9269
rect 30219 9220 30220 9260
rect 30260 9220 30261 9260
rect 30219 9211 30261 9220
rect 34347 9260 34389 9269
rect 34347 9220 34348 9260
rect 34388 9220 34389 9260
rect 34347 9211 34389 9220
rect 36363 9260 36405 9269
rect 36363 9220 36364 9260
rect 36404 9220 36405 9260
rect 36363 9211 36405 9220
rect 39147 9260 39189 9269
rect 39147 9220 39148 9260
rect 39188 9220 39189 9260
rect 39147 9211 39189 9220
rect 1152 9092 41856 9116
rect 1152 9052 3688 9092
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 4056 9052 18808 9092
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 19176 9052 33928 9092
rect 33968 9052 34010 9092
rect 34050 9052 34092 9092
rect 34132 9052 34174 9092
rect 34214 9052 34256 9092
rect 34296 9052 41856 9092
rect 1152 9028 41856 9052
rect 5643 8924 5685 8933
rect 5643 8884 5644 8924
rect 5684 8884 5685 8924
rect 5643 8875 5685 8884
rect 9195 8924 9237 8933
rect 9195 8884 9196 8924
rect 9236 8884 9237 8924
rect 9195 8875 9237 8884
rect 20235 8840 20277 8849
rect 20235 8800 20236 8840
rect 20276 8800 20277 8840
rect 20235 8791 20277 8800
rect 21099 8840 21141 8849
rect 21099 8800 21100 8840
rect 21140 8800 21141 8840
rect 21099 8791 21141 8800
rect 22731 8840 22773 8849
rect 22731 8800 22732 8840
rect 22772 8800 22773 8840
rect 22731 8791 22773 8800
rect 30891 8840 30933 8849
rect 30891 8800 30892 8840
rect 30932 8800 30933 8840
rect 30891 8791 30933 8800
rect 11115 8756 11157 8765
rect 11115 8716 11116 8756
rect 11156 8716 11157 8756
rect 20035 8756 20093 8757
rect 11115 8707 11157 8716
rect 19515 8714 19557 8723
rect 20035 8716 20044 8756
rect 20084 8716 20093 8756
rect 20035 8715 20093 8716
rect 20515 8756 20573 8757
rect 20515 8716 20524 8756
rect 20564 8716 20573 8756
rect 20515 8715 20573 8716
rect 20899 8756 20957 8757
rect 20899 8716 20908 8756
rect 20948 8716 20957 8756
rect 27235 8756 27293 8757
rect 20899 8715 20957 8716
rect 12075 8686 12117 8695
rect 3147 8677 3189 8686
rect 1315 8672 1373 8673
rect 1315 8632 1324 8672
rect 1364 8632 1373 8672
rect 1315 8631 1373 8632
rect 2563 8672 2621 8673
rect 2563 8632 2572 8672
rect 2612 8632 2621 8672
rect 2563 8631 2621 8632
rect 3147 8637 3148 8677
rect 3188 8637 3189 8677
rect 3147 8628 3189 8637
rect 3619 8672 3677 8673
rect 3619 8632 3628 8672
rect 3668 8632 3677 8672
rect 3619 8631 3677 8632
rect 4107 8672 4149 8681
rect 4107 8632 4108 8672
rect 4148 8632 4149 8672
rect 4107 8623 4149 8632
rect 4203 8672 4245 8681
rect 4203 8632 4204 8672
rect 4244 8632 4245 8672
rect 4203 8623 4245 8632
rect 4587 8672 4629 8681
rect 4587 8632 4588 8672
rect 4628 8632 4629 8672
rect 4587 8623 4629 8632
rect 4683 8672 4725 8681
rect 4683 8632 4684 8672
rect 4724 8632 4725 8672
rect 4683 8623 4725 8632
rect 5251 8672 5309 8673
rect 5251 8632 5260 8672
rect 5300 8632 5309 8672
rect 5251 8631 5309 8632
rect 5355 8672 5397 8681
rect 5355 8632 5356 8672
rect 5396 8632 5397 8672
rect 5355 8623 5397 8632
rect 6115 8672 6173 8673
rect 6115 8632 6124 8672
rect 6164 8632 6173 8672
rect 6115 8631 6173 8632
rect 7363 8672 7421 8673
rect 7363 8632 7372 8672
rect 7412 8632 7421 8672
rect 7363 8631 7421 8632
rect 7747 8672 7805 8673
rect 7747 8632 7756 8672
rect 7796 8632 7805 8672
rect 7747 8631 7805 8632
rect 8995 8672 9053 8673
rect 8995 8632 9004 8672
rect 9044 8632 9053 8672
rect 8995 8631 9053 8632
rect 9483 8672 9525 8681
rect 9483 8632 9484 8672
rect 9524 8632 9525 8672
rect 9483 8623 9525 8632
rect 9579 8672 9621 8681
rect 9579 8632 9580 8672
rect 9620 8632 9621 8672
rect 9579 8623 9621 8632
rect 9675 8672 9717 8681
rect 9675 8632 9676 8672
rect 9716 8632 9717 8672
rect 9675 8623 9717 8632
rect 9963 8672 10005 8681
rect 9963 8632 9964 8672
rect 10004 8632 10005 8672
rect 9963 8623 10005 8632
rect 10059 8672 10101 8681
rect 10059 8632 10060 8672
rect 10100 8632 10101 8672
rect 10059 8623 10101 8632
rect 10539 8672 10581 8681
rect 10539 8632 10540 8672
rect 10580 8632 10581 8672
rect 10539 8623 10581 8632
rect 10635 8672 10677 8681
rect 10635 8632 10636 8672
rect 10676 8632 10677 8672
rect 10635 8623 10677 8632
rect 11019 8672 11061 8681
rect 11019 8632 11020 8672
rect 11060 8632 11061 8672
rect 11019 8623 11061 8632
rect 11587 8672 11645 8673
rect 11587 8632 11596 8672
rect 11636 8632 11645 8672
rect 12075 8646 12076 8686
rect 12116 8646 12117 8686
rect 12075 8637 12117 8646
rect 12459 8672 12501 8681
rect 11587 8631 11645 8632
rect 12459 8632 12460 8672
rect 12500 8632 12501 8672
rect 12459 8623 12501 8632
rect 12555 8672 12597 8681
rect 12555 8632 12556 8672
rect 12596 8632 12597 8672
rect 12555 8623 12597 8632
rect 13131 8672 13173 8681
rect 13131 8632 13132 8672
rect 13172 8632 13173 8672
rect 13131 8623 13173 8632
rect 13227 8672 13269 8681
rect 13227 8632 13228 8672
rect 13268 8632 13269 8672
rect 13227 8623 13269 8632
rect 13515 8672 13557 8681
rect 13515 8632 13516 8672
rect 13556 8632 13557 8672
rect 13515 8623 13557 8632
rect 13611 8672 13653 8681
rect 13611 8632 13612 8672
rect 13652 8632 13653 8672
rect 13611 8623 13653 8632
rect 13995 8672 14037 8681
rect 13995 8632 13996 8672
rect 14036 8632 14037 8672
rect 13995 8623 14037 8632
rect 14091 8672 14133 8681
rect 15051 8677 15093 8686
rect 14091 8632 14092 8672
rect 14132 8632 14133 8672
rect 14091 8623 14133 8632
rect 14563 8672 14621 8673
rect 14563 8632 14572 8672
rect 14612 8632 14621 8672
rect 14563 8631 14621 8632
rect 15051 8637 15052 8677
rect 15092 8637 15093 8677
rect 15051 8628 15093 8637
rect 15435 8672 15477 8681
rect 15435 8632 15436 8672
rect 15476 8632 15477 8672
rect 15435 8623 15477 8632
rect 15531 8672 15573 8681
rect 15531 8632 15532 8672
rect 15572 8632 15573 8672
rect 15531 8623 15573 8632
rect 15627 8672 15669 8681
rect 15627 8632 15628 8672
rect 15668 8632 15669 8672
rect 15627 8623 15669 8632
rect 15723 8672 15765 8681
rect 15723 8632 15724 8672
rect 15764 8632 15765 8672
rect 15723 8623 15765 8632
rect 16195 8672 16253 8673
rect 16195 8632 16204 8672
rect 16244 8632 16253 8672
rect 16195 8631 16253 8632
rect 17443 8672 17501 8673
rect 17443 8632 17452 8672
rect 17492 8632 17501 8672
rect 17443 8631 17501 8632
rect 17931 8672 17973 8681
rect 17931 8632 17932 8672
rect 17972 8632 17973 8672
rect 17931 8623 17973 8632
rect 18027 8672 18069 8681
rect 18027 8632 18028 8672
rect 18068 8632 18069 8672
rect 18027 8623 18069 8632
rect 18411 8672 18453 8681
rect 18411 8632 18412 8672
rect 18452 8632 18453 8672
rect 18411 8623 18453 8632
rect 18507 8672 18549 8681
rect 19515 8674 19516 8714
rect 19556 8674 19557 8714
rect 24603 8714 24645 8723
rect 27235 8716 27244 8756
rect 27284 8716 27293 8756
rect 27235 8715 27293 8716
rect 38755 8756 38813 8757
rect 38755 8716 38764 8756
rect 38804 8716 38813 8756
rect 38755 8715 38813 8716
rect 40867 8756 40925 8757
rect 40867 8716 40876 8756
rect 40916 8716 40925 8756
rect 40867 8715 40925 8716
rect 41251 8756 41309 8757
rect 41251 8716 41260 8756
rect 41300 8716 41309 8756
rect 41251 8715 41309 8716
rect 18507 8632 18508 8672
rect 18548 8632 18549 8672
rect 18507 8623 18549 8632
rect 18979 8672 19037 8673
rect 18979 8632 18988 8672
rect 19028 8632 19037 8672
rect 19515 8665 19557 8674
rect 21283 8672 21341 8673
rect 18979 8631 19037 8632
rect 21283 8632 21292 8672
rect 21332 8632 21341 8672
rect 21283 8631 21341 8632
rect 22531 8672 22589 8673
rect 22531 8632 22540 8672
rect 22580 8632 22589 8672
rect 22531 8631 22589 8632
rect 23019 8672 23061 8681
rect 23019 8632 23020 8672
rect 23060 8632 23061 8672
rect 23019 8623 23061 8632
rect 23115 8672 23157 8681
rect 23115 8632 23116 8672
rect 23156 8632 23157 8672
rect 23115 8623 23157 8632
rect 23499 8672 23541 8681
rect 23499 8632 23500 8672
rect 23540 8632 23541 8672
rect 23499 8623 23541 8632
rect 23595 8672 23637 8681
rect 24603 8674 24604 8714
rect 24644 8674 24645 8714
rect 26667 8686 26709 8695
rect 23595 8632 23596 8672
rect 23636 8632 23637 8672
rect 23595 8623 23637 8632
rect 24067 8672 24125 8673
rect 24067 8632 24076 8672
rect 24116 8632 24125 8672
rect 24603 8665 24645 8674
rect 25131 8672 25173 8681
rect 24067 8631 24125 8632
rect 25131 8632 25132 8672
rect 25172 8632 25173 8672
rect 25131 8623 25173 8632
rect 25227 8672 25269 8681
rect 25227 8632 25228 8672
rect 25268 8632 25269 8672
rect 25227 8623 25269 8632
rect 25611 8672 25653 8681
rect 25611 8632 25612 8672
rect 25652 8632 25653 8672
rect 25611 8623 25653 8632
rect 25707 8672 25749 8681
rect 25707 8632 25708 8672
rect 25748 8632 25749 8672
rect 25707 8623 25749 8632
rect 26179 8672 26237 8673
rect 26179 8632 26188 8672
rect 26228 8632 26237 8672
rect 26667 8646 26668 8686
rect 26708 8646 26709 8686
rect 26667 8637 26709 8646
rect 28771 8672 28829 8673
rect 26179 8631 26237 8632
rect 28771 8632 28780 8672
rect 28820 8632 28829 8672
rect 28771 8631 28829 8632
rect 29635 8672 29693 8673
rect 29635 8632 29644 8672
rect 29684 8632 29693 8672
rect 29635 8631 29693 8632
rect 31083 8672 31125 8681
rect 31083 8632 31084 8672
rect 31124 8632 31125 8672
rect 31083 8623 31125 8632
rect 31939 8672 31997 8673
rect 31939 8632 31948 8672
rect 31988 8632 31997 8672
rect 31939 8631 31997 8632
rect 32803 8672 32861 8673
rect 32803 8632 32812 8672
rect 32852 8632 32861 8672
rect 32803 8631 32861 8632
rect 35491 8672 35549 8673
rect 35491 8632 35500 8672
rect 35540 8632 35549 8672
rect 35491 8631 35549 8632
rect 36355 8672 36413 8673
rect 36355 8632 36364 8672
rect 36404 8632 36413 8672
rect 36355 8631 36413 8632
rect 37123 8672 37181 8673
rect 37123 8632 37132 8672
rect 37172 8632 37181 8672
rect 37123 8631 37181 8632
rect 38371 8672 38429 8673
rect 38371 8632 38380 8672
rect 38420 8632 38429 8672
rect 38371 8631 38429 8632
rect 39139 8672 39197 8673
rect 39139 8632 39148 8672
rect 39188 8632 39197 8672
rect 39139 8631 39197 8632
rect 40387 8672 40445 8673
rect 40387 8632 40396 8672
rect 40436 8632 40445 8672
rect 40387 8631 40445 8632
rect 2955 8588 2997 8597
rect 2955 8548 2956 8588
rect 2996 8548 2997 8588
rect 2955 8539 2997 8548
rect 26859 8588 26901 8597
rect 26859 8548 26860 8588
rect 26900 8548 26901 8588
rect 26859 8539 26901 8548
rect 30027 8588 30069 8597
rect 30027 8548 30028 8588
rect 30068 8548 30069 8588
rect 30027 8539 30069 8548
rect 31563 8588 31605 8597
rect 31563 8548 31564 8588
rect 31604 8548 31605 8588
rect 31563 8539 31605 8548
rect 36747 8588 36789 8597
rect 36747 8548 36748 8588
rect 36788 8548 36789 8588
rect 36747 8539 36789 8548
rect 2763 8504 2805 8513
rect 2763 8464 2764 8504
rect 2804 8464 2805 8504
rect 2763 8455 2805 8464
rect 5163 8500 5205 8509
rect 5163 8460 5164 8500
rect 5204 8460 5205 8500
rect 5163 8451 5205 8460
rect 7563 8504 7605 8513
rect 7563 8464 7564 8504
rect 7604 8464 7605 8504
rect 7563 8455 7605 8464
rect 9763 8504 9821 8505
rect 9763 8464 9772 8504
rect 9812 8464 9821 8504
rect 9763 8463 9821 8464
rect 10243 8504 10301 8505
rect 10243 8464 10252 8504
rect 10292 8464 10301 8504
rect 10243 8463 10301 8464
rect 12267 8504 12309 8513
rect 12267 8464 12268 8504
rect 12308 8464 12309 8504
rect 12267 8455 12309 8464
rect 12739 8504 12797 8505
rect 12739 8464 12748 8504
rect 12788 8464 12797 8504
rect 12739 8463 12797 8464
rect 12931 8504 12989 8505
rect 12931 8464 12940 8504
rect 12980 8464 12989 8504
rect 12931 8463 12989 8464
rect 15243 8504 15285 8513
rect 15243 8464 15244 8504
rect 15284 8464 15285 8504
rect 15243 8455 15285 8464
rect 17643 8504 17685 8513
rect 17643 8464 17644 8504
rect 17684 8464 17685 8504
rect 17643 8455 17685 8464
rect 19659 8504 19701 8513
rect 19659 8464 19660 8504
rect 19700 8464 19701 8504
rect 19659 8455 19701 8464
rect 20715 8504 20757 8513
rect 20715 8464 20716 8504
rect 20756 8464 20757 8504
rect 20715 8455 20757 8464
rect 24747 8504 24789 8513
rect 24747 8464 24748 8504
rect 24788 8464 24789 8504
rect 24747 8455 24789 8464
rect 27051 8504 27093 8513
rect 27051 8464 27052 8504
rect 27092 8464 27093 8504
rect 27051 8455 27093 8464
rect 27619 8504 27677 8505
rect 27619 8464 27628 8504
rect 27668 8464 27677 8504
rect 27619 8463 27677 8464
rect 33955 8504 34013 8505
rect 33955 8464 33964 8504
rect 34004 8464 34013 8504
rect 33955 8463 34013 8464
rect 34339 8504 34397 8505
rect 34339 8464 34348 8504
rect 34388 8464 34397 8504
rect 34339 8463 34397 8464
rect 36939 8504 36981 8513
rect 36939 8464 36940 8504
rect 36980 8464 36981 8504
rect 36939 8455 36981 8464
rect 38571 8504 38613 8513
rect 38571 8464 38572 8504
rect 38612 8464 38613 8504
rect 38571 8455 38613 8464
rect 40587 8504 40629 8513
rect 40587 8464 40588 8504
rect 40628 8464 40629 8504
rect 40587 8455 40629 8464
rect 41067 8504 41109 8513
rect 41067 8464 41068 8504
rect 41108 8464 41109 8504
rect 41067 8455 41109 8464
rect 41451 8504 41493 8513
rect 41451 8464 41452 8504
rect 41492 8464 41493 8504
rect 41451 8455 41493 8464
rect 1152 8336 41856 8360
rect 1152 8296 4928 8336
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 5296 8296 20048 8336
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20416 8296 35168 8336
rect 35208 8296 35250 8336
rect 35290 8296 35332 8336
rect 35372 8296 35414 8336
rect 35454 8296 35496 8336
rect 35536 8296 41856 8336
rect 1152 8272 41856 8296
rect 2859 8168 2901 8177
rect 2859 8128 2860 8168
rect 2900 8128 2901 8168
rect 2859 8119 2901 8128
rect 3051 8168 3093 8177
rect 3051 8128 3052 8168
rect 3092 8128 3093 8168
rect 3051 8119 3093 8128
rect 8131 8168 8189 8169
rect 8131 8128 8140 8168
rect 8180 8128 8189 8168
rect 8131 8127 8189 8128
rect 9859 8168 9917 8169
rect 9859 8128 9868 8168
rect 9908 8128 9917 8168
rect 9859 8127 9917 8128
rect 10347 8168 10389 8177
rect 10347 8128 10348 8168
rect 10388 8128 10389 8168
rect 10347 8119 10389 8128
rect 13611 8168 13653 8177
rect 13611 8128 13612 8168
rect 13652 8128 13653 8168
rect 13611 8119 13653 8128
rect 15715 8168 15773 8169
rect 15715 8128 15724 8168
rect 15764 8128 15773 8168
rect 15715 8127 15773 8128
rect 18315 8168 18357 8177
rect 18315 8128 18316 8168
rect 18356 8128 18357 8168
rect 18315 8119 18357 8128
rect 22443 8168 22485 8177
rect 22443 8128 22444 8168
rect 22484 8128 22485 8168
rect 22443 8119 22485 8128
rect 38187 8168 38229 8177
rect 38187 8128 38188 8168
rect 38228 8128 38229 8168
rect 38187 8119 38229 8128
rect 40875 8168 40917 8177
rect 40875 8128 40876 8168
rect 40916 8128 40917 8168
rect 40875 8119 40917 8128
rect 26571 8084 26613 8093
rect 26571 8044 26572 8084
rect 26612 8044 26613 8084
rect 26571 8035 26613 8044
rect 28587 8084 28629 8093
rect 28587 8044 28588 8084
rect 28628 8044 28629 8084
rect 28587 8035 28629 8044
rect 40491 8084 40533 8093
rect 40491 8044 40492 8084
rect 40532 8044 40533 8084
rect 40491 8035 40533 8044
rect 1411 8000 1469 8001
rect 1411 7960 1420 8000
rect 1460 7960 1469 8000
rect 1411 7959 1469 7960
rect 2659 8000 2717 8001
rect 2659 7960 2668 8000
rect 2708 7960 2717 8000
rect 2659 7959 2717 7960
rect 3235 8000 3293 8001
rect 3235 7960 3244 8000
rect 3284 7960 3293 8000
rect 3235 7959 3293 7960
rect 4483 8000 4541 8001
rect 4483 7960 4492 8000
rect 4532 7960 4541 8000
rect 4483 7959 4541 7960
rect 4963 8000 5021 8001
rect 4963 7960 4972 8000
rect 5012 7960 5021 8000
rect 4963 7959 5021 7960
rect 5259 8000 5301 8009
rect 5259 7960 5260 8000
rect 5300 7960 5301 8000
rect 5259 7951 5301 7960
rect 5355 8000 5397 8009
rect 5355 7960 5356 8000
rect 5396 7960 5397 8000
rect 5355 7951 5397 7960
rect 5827 8000 5885 8001
rect 5827 7960 5836 8000
rect 5876 7960 5885 8000
rect 5827 7959 5885 7960
rect 7075 8000 7133 8001
rect 7075 7960 7084 8000
rect 7124 7960 7133 8000
rect 7075 7959 7133 7960
rect 7651 8000 7709 8001
rect 7651 7960 7660 8000
rect 7700 7960 7709 8000
rect 7651 7959 7709 7960
rect 7747 8000 7805 8001
rect 7747 7960 7756 8000
rect 7796 7960 7805 8000
rect 7747 7959 7805 7960
rect 7947 8000 7989 8009
rect 7947 7960 7948 8000
rect 7988 7960 7989 8000
rect 7947 7951 7989 7960
rect 8043 8000 8085 8009
rect 8043 7960 8044 8000
rect 8084 7960 8085 8000
rect 8515 8000 8573 8001
rect 8043 7951 8085 7960
rect 8200 7985 8242 7994
rect 8200 7945 8201 7985
rect 8241 7945 8242 7985
rect 8515 7960 8524 8000
rect 8564 7960 8573 8000
rect 8515 7959 8573 7960
rect 8811 8000 8853 8009
rect 8811 7960 8812 8000
rect 8852 7960 8853 8000
rect 8811 7951 8853 7960
rect 8907 8000 8949 8009
rect 8907 7960 8908 8000
rect 8948 7960 8949 8000
rect 8907 7951 8949 7960
rect 9387 8000 9429 8009
rect 9387 7960 9388 8000
rect 9428 7960 9429 8000
rect 9387 7951 9429 7960
rect 9483 8000 9525 8009
rect 9483 7960 9484 8000
rect 9524 7960 9525 8000
rect 9483 7951 9525 7960
rect 9579 8000 9621 8009
rect 9579 7960 9580 8000
rect 9620 7960 9621 8000
rect 9579 7951 9621 7960
rect 9675 8000 9717 8009
rect 9675 7960 9676 8000
rect 9716 7960 9717 8000
rect 9675 7951 9717 7960
rect 9963 8000 10005 8009
rect 9963 7960 9964 8000
rect 10004 7960 10005 8000
rect 9963 7951 10005 7960
rect 10059 8000 10101 8009
rect 10059 7960 10060 8000
rect 10100 7960 10101 8000
rect 10059 7951 10101 7960
rect 10155 8000 10197 8009
rect 10155 7960 10156 8000
rect 10196 7960 10197 8000
rect 10155 7951 10197 7960
rect 10531 8000 10589 8001
rect 10531 7960 10540 8000
rect 10580 7960 10589 8000
rect 10531 7959 10589 7960
rect 11779 8000 11837 8001
rect 11779 7960 11788 8000
rect 11828 7960 11837 8000
rect 11779 7959 11837 7960
rect 12163 8000 12221 8001
rect 12163 7960 12172 8000
rect 12212 7960 12221 8000
rect 12163 7959 12221 7960
rect 13411 8000 13469 8001
rect 13411 7960 13420 8000
rect 13460 7960 13469 8000
rect 13411 7959 13469 7960
rect 13795 8000 13853 8001
rect 13795 7960 13804 8000
rect 13844 7960 13853 8000
rect 13795 7959 13853 7960
rect 15043 8000 15101 8001
rect 15043 7960 15052 8000
rect 15092 7960 15101 8000
rect 15043 7959 15101 7960
rect 15435 8000 15477 8009
rect 15435 7960 15436 8000
rect 15476 7960 15477 8000
rect 15435 7951 15477 7960
rect 15531 8000 15573 8009
rect 15531 7960 15532 8000
rect 15572 7960 15573 8000
rect 15531 7951 15573 7960
rect 15915 8000 15957 8009
rect 15915 7960 15916 8000
rect 15956 7960 15957 8000
rect 15915 7951 15957 7960
rect 16011 8000 16053 8009
rect 16011 7960 16012 8000
rect 16052 7960 16053 8000
rect 16011 7951 16053 7960
rect 16107 8000 16149 8009
rect 16107 7960 16108 8000
rect 16148 7960 16149 8000
rect 16107 7951 16149 7960
rect 16203 8000 16245 8009
rect 16203 7960 16204 8000
rect 16244 7960 16245 8000
rect 16203 7951 16245 7960
rect 16587 8000 16629 8009
rect 16587 7960 16588 8000
rect 16628 7960 16629 8000
rect 16587 7951 16629 7960
rect 16683 8000 16725 8009
rect 16683 7960 16684 8000
rect 16724 7960 16725 8000
rect 16683 7951 16725 7960
rect 17635 8000 17693 8001
rect 17635 7960 17644 8000
rect 17684 7960 17693 8000
rect 17635 7959 17693 7960
rect 18123 7995 18165 8004
rect 18123 7955 18124 7995
rect 18164 7955 18165 7995
rect 18499 8000 18557 8001
rect 18499 7960 18508 8000
rect 18548 7960 18557 8000
rect 18499 7959 18557 7960
rect 19747 8000 19805 8001
rect 19747 7960 19756 8000
rect 19796 7960 19805 8000
rect 19747 7959 19805 7960
rect 20803 8000 20861 8001
rect 20803 7960 20812 8000
rect 20852 7960 20861 8000
rect 20803 7959 20861 7960
rect 22051 8000 22109 8001
rect 22051 7960 22060 8000
rect 22100 7960 22109 8000
rect 22051 7959 22109 7960
rect 23491 8000 23549 8001
rect 23491 7960 23500 8000
rect 23540 7960 23549 8000
rect 23491 7959 23549 7960
rect 24739 8000 24797 8001
rect 24739 7960 24748 8000
rect 24788 7960 24797 8000
rect 24739 7959 24797 7960
rect 25123 8000 25181 8001
rect 25123 7960 25132 8000
rect 25172 7960 25181 8000
rect 25123 7959 25181 7960
rect 26371 8000 26429 8001
rect 26371 7960 26380 8000
rect 26420 7960 26429 8000
rect 26371 7959 26429 7960
rect 26859 8000 26901 8009
rect 26859 7960 26860 8000
rect 26900 7960 26901 8000
rect 18123 7946 18165 7955
rect 26859 7951 26901 7960
rect 26955 8000 26997 8009
rect 26955 7960 26956 8000
rect 26996 7960 26997 8000
rect 26955 7951 26997 7960
rect 27339 8000 27381 8009
rect 27339 7960 27340 8000
rect 27380 7960 27381 8000
rect 27339 7951 27381 7960
rect 27907 8000 27965 8001
rect 27907 7960 27916 8000
rect 27956 7960 27965 8000
rect 27907 7959 27965 7960
rect 28395 7995 28437 8004
rect 28395 7955 28396 7995
rect 28436 7955 28437 7995
rect 28963 8000 29021 8001
rect 28963 7960 28972 8000
rect 29012 7960 29021 8000
rect 28963 7959 29021 7960
rect 30211 8000 30269 8001
rect 30211 7960 30220 8000
rect 30260 7960 30269 8000
rect 30211 7959 30269 7960
rect 30595 8000 30653 8001
rect 30595 7960 30604 8000
rect 30644 7960 30653 8000
rect 30595 7959 30653 7960
rect 31843 8000 31901 8001
rect 31843 7960 31852 8000
rect 31892 7960 31901 8000
rect 31843 7959 31901 7960
rect 32419 8000 32477 8001
rect 32419 7960 32428 8000
rect 32468 7960 32477 8000
rect 32419 7959 32477 7960
rect 33667 8000 33725 8001
rect 33667 7960 33676 8000
rect 33716 7960 33725 8000
rect 33667 7959 33725 7960
rect 35107 8000 35165 8001
rect 35107 7960 35116 8000
rect 35156 7960 35165 8000
rect 35107 7959 35165 7960
rect 35971 8000 36029 8001
rect 35971 7960 35980 8000
rect 36020 7960 36029 8000
rect 35971 7959 36029 7960
rect 36363 8000 36405 8009
rect 36363 7960 36364 8000
rect 36404 7960 36405 8000
rect 28395 7946 28437 7955
rect 36363 7951 36405 7960
rect 36643 8000 36701 8001
rect 36643 7960 36652 8000
rect 36692 7960 36701 8000
rect 36643 7959 36701 7960
rect 38763 8000 38805 8009
rect 38763 7960 38764 8000
rect 38804 7960 38805 8000
rect 38763 7951 38805 7960
rect 38859 8000 38901 8009
rect 38859 7960 38860 8000
rect 38900 7960 38901 8000
rect 38859 7951 38901 7960
rect 39811 8000 39869 8001
rect 39811 7960 39820 8000
rect 39860 7960 39869 8000
rect 39811 7959 39869 7960
rect 40347 7990 40389 7999
rect 40347 7950 40348 7990
rect 40388 7950 40389 7990
rect 8200 7936 8242 7945
rect 40347 7941 40389 7950
rect 17067 7916 17109 7925
rect 17067 7876 17068 7916
rect 17108 7876 17109 7916
rect 17067 7867 17109 7876
rect 17163 7916 17205 7925
rect 17163 7876 17164 7916
rect 17204 7876 17205 7916
rect 17163 7867 17205 7876
rect 20419 7916 20477 7917
rect 20419 7876 20428 7916
rect 20468 7876 20477 7916
rect 20419 7875 20477 7876
rect 22627 7916 22685 7917
rect 22627 7876 22636 7916
rect 22676 7876 22685 7916
rect 22627 7875 22685 7876
rect 27435 7916 27477 7925
rect 27435 7876 27436 7916
rect 27476 7876 27477 7916
rect 27435 7867 27477 7876
rect 38371 7916 38429 7917
rect 38371 7876 38380 7916
rect 38420 7876 38429 7916
rect 38371 7875 38429 7876
rect 39243 7916 39285 7925
rect 39243 7876 39244 7916
rect 39284 7876 39285 7916
rect 39243 7867 39285 7876
rect 39339 7916 39381 7925
rect 39339 7876 39340 7916
rect 39380 7876 39381 7916
rect 39339 7867 39381 7876
rect 40675 7916 40733 7917
rect 40675 7876 40684 7916
rect 40724 7876 40733 7916
rect 40675 7875 40733 7876
rect 41059 7916 41117 7917
rect 41059 7876 41068 7916
rect 41108 7876 41117 7916
rect 41059 7875 41117 7876
rect 41443 7916 41501 7917
rect 41443 7876 41452 7916
rect 41492 7876 41501 7916
rect 41443 7875 41501 7876
rect 9187 7832 9245 7833
rect 9187 7792 9196 7832
rect 9236 7792 9245 7832
rect 9187 7791 9245 7792
rect 37803 7832 37845 7841
rect 37803 7792 37804 7832
rect 37844 7792 37845 7832
rect 37803 7783 37845 7792
rect 41643 7832 41685 7841
rect 41643 7792 41644 7832
rect 41684 7792 41685 7832
rect 41643 7783 41685 7792
rect 5635 7748 5693 7749
rect 5635 7708 5644 7748
rect 5684 7708 5693 7748
rect 5635 7707 5693 7708
rect 7275 7748 7317 7757
rect 7275 7708 7276 7748
rect 7316 7708 7317 7748
rect 7275 7699 7317 7708
rect 15243 7748 15285 7757
rect 15243 7708 15244 7748
rect 15284 7708 15285 7748
rect 15243 7699 15285 7708
rect 19947 7748 19989 7757
rect 19947 7708 19948 7748
rect 19988 7708 19989 7748
rect 19947 7699 19989 7708
rect 20619 7748 20661 7757
rect 20619 7708 20620 7748
rect 20660 7708 20661 7748
rect 20619 7699 20661 7708
rect 22251 7748 22293 7757
rect 22251 7708 22252 7748
rect 22292 7708 22293 7748
rect 22251 7699 22293 7708
rect 24939 7748 24981 7757
rect 24939 7708 24940 7748
rect 24980 7708 24981 7748
rect 24939 7699 24981 7708
rect 30411 7748 30453 7757
rect 30411 7708 30412 7748
rect 30452 7708 30453 7748
rect 30411 7699 30453 7708
rect 32043 7748 32085 7757
rect 32043 7708 32044 7748
rect 32084 7708 32085 7748
rect 32043 7699 32085 7708
rect 32235 7748 32277 7757
rect 32235 7708 32236 7748
rect 32276 7708 32277 7748
rect 32235 7699 32277 7708
rect 33955 7748 34013 7749
rect 33955 7708 33964 7748
rect 34004 7708 34013 7748
rect 33955 7707 34013 7708
rect 36939 7748 36981 7757
rect 36939 7708 36940 7748
rect 36980 7708 36981 7748
rect 36939 7699 36981 7708
rect 41259 7748 41301 7757
rect 41259 7708 41260 7748
rect 41300 7708 41301 7748
rect 41259 7699 41301 7708
rect 1152 7580 41856 7604
rect 1152 7540 3688 7580
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 4056 7540 18808 7580
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 19176 7540 33928 7580
rect 33968 7540 34010 7580
rect 34050 7540 34092 7580
rect 34132 7540 34174 7580
rect 34214 7540 34256 7580
rect 34296 7540 41856 7580
rect 1152 7516 41856 7540
rect 3523 7412 3581 7413
rect 3523 7372 3532 7412
rect 3572 7372 3581 7412
rect 3523 7371 3581 7372
rect 9003 7412 9045 7421
rect 9003 7372 9004 7412
rect 9044 7372 9045 7412
rect 9003 7363 9045 7372
rect 9867 7412 9909 7421
rect 9867 7372 9868 7412
rect 9908 7372 9909 7412
rect 9867 7363 9909 7372
rect 32331 7412 32373 7421
rect 32331 7372 32332 7412
rect 32372 7372 32373 7412
rect 32331 7363 32373 7372
rect 37803 7412 37845 7421
rect 37803 7372 37804 7412
rect 37844 7372 37845 7412
rect 37803 7363 37845 7372
rect 2955 7328 2997 7337
rect 2955 7288 2956 7328
rect 2996 7288 2997 7328
rect 2955 7279 2997 7288
rect 29547 7328 29589 7337
rect 29547 7288 29548 7328
rect 29588 7288 29589 7328
rect 29547 7279 29589 7288
rect 3243 7244 3285 7253
rect 3243 7204 3244 7244
rect 3284 7204 3285 7244
rect 3243 7195 3285 7204
rect 5451 7244 5493 7253
rect 5451 7204 5452 7244
rect 5492 7204 5493 7244
rect 25219 7244 25277 7245
rect 5451 7195 5493 7204
rect 24699 7202 24741 7211
rect 25219 7204 25228 7244
rect 25268 7204 25277 7244
rect 25219 7203 25277 7204
rect 25603 7244 25661 7245
rect 25603 7204 25612 7244
rect 25652 7204 25661 7244
rect 25603 7203 25661 7204
rect 29347 7244 29405 7245
rect 29347 7204 29356 7244
rect 29396 7204 29405 7244
rect 32131 7244 32189 7245
rect 29347 7203 29405 7204
rect 1315 7160 1373 7161
rect 1315 7120 1324 7160
rect 1364 7120 1373 7160
rect 1315 7119 1373 7120
rect 1507 7160 1565 7161
rect 1507 7120 1516 7160
rect 1556 7120 1565 7160
rect 1507 7119 1565 7120
rect 2755 7160 2813 7161
rect 2755 7120 2764 7160
rect 2804 7120 2813 7160
rect 2755 7119 2813 7120
rect 3147 7160 3189 7169
rect 3147 7120 3148 7160
rect 3188 7120 3189 7160
rect 3147 7111 3189 7120
rect 3339 7160 3381 7169
rect 3339 7120 3340 7160
rect 3380 7120 3381 7160
rect 3339 7111 3381 7120
rect 3915 7160 3957 7169
rect 3915 7120 3916 7160
rect 3956 7120 3957 7160
rect 3915 7111 3957 7120
rect 4195 7160 4253 7161
rect 4195 7120 4204 7160
rect 4244 7120 4253 7160
rect 4195 7119 4253 7120
rect 4491 7160 4533 7169
rect 4491 7120 4492 7160
rect 4532 7120 4533 7160
rect 4491 7111 4533 7120
rect 4675 7160 4733 7161
rect 4675 7120 4684 7160
rect 4724 7120 4733 7160
rect 4675 7119 4733 7120
rect 4971 7160 5013 7169
rect 4971 7120 4972 7160
rect 5012 7120 5013 7160
rect 4971 7111 5013 7120
rect 5067 7160 5109 7169
rect 5067 7120 5068 7160
rect 5108 7120 5109 7160
rect 5067 7111 5109 7120
rect 5547 7160 5589 7169
rect 6507 7165 6549 7174
rect 5547 7120 5548 7160
rect 5588 7120 5589 7160
rect 5547 7111 5589 7120
rect 6019 7160 6077 7161
rect 6019 7120 6028 7160
rect 6068 7120 6077 7160
rect 6019 7119 6077 7120
rect 6507 7125 6508 7165
rect 6548 7125 6549 7165
rect 6507 7116 6549 7125
rect 7083 7160 7125 7169
rect 7083 7120 7084 7160
rect 7124 7120 7125 7160
rect 7083 7111 7125 7120
rect 7179 7160 7221 7169
rect 7179 7120 7180 7160
rect 7220 7120 7221 7160
rect 7179 7111 7221 7120
rect 7563 7160 7605 7169
rect 7563 7120 7564 7160
rect 7604 7120 7605 7160
rect 7563 7111 7605 7120
rect 7659 7160 7701 7169
rect 8619 7165 8661 7174
rect 7659 7120 7660 7160
rect 7700 7120 7701 7160
rect 7659 7111 7701 7120
rect 8131 7160 8189 7161
rect 8131 7120 8140 7160
rect 8180 7120 8189 7160
rect 8131 7119 8189 7120
rect 8619 7125 8620 7165
rect 8660 7125 8661 7165
rect 8619 7116 8661 7125
rect 9003 7160 9045 7169
rect 9003 7120 9004 7160
rect 9044 7120 9045 7160
rect 9003 7111 9045 7120
rect 9291 7160 9333 7169
rect 9291 7120 9292 7160
rect 9332 7120 9333 7160
rect 9291 7111 9333 7120
rect 9483 7160 9525 7169
rect 9483 7120 9484 7160
rect 9524 7120 9525 7160
rect 9483 7111 9525 7120
rect 9579 7160 9621 7169
rect 9579 7120 9580 7160
rect 9620 7120 9621 7160
rect 9579 7111 9621 7120
rect 9667 7160 9725 7161
rect 9667 7120 9676 7160
rect 9716 7120 9725 7160
rect 9667 7119 9725 7120
rect 10051 7160 10109 7161
rect 10051 7120 10060 7160
rect 10100 7120 10109 7160
rect 10051 7119 10109 7120
rect 11299 7160 11357 7161
rect 11299 7120 11308 7160
rect 11348 7120 11357 7160
rect 11299 7119 11357 7120
rect 11875 7160 11933 7161
rect 11875 7120 11884 7160
rect 11924 7120 11933 7160
rect 11875 7119 11933 7120
rect 13123 7160 13181 7161
rect 13123 7120 13132 7160
rect 13172 7120 13181 7160
rect 13123 7119 13181 7120
rect 13515 7160 13557 7169
rect 13515 7120 13516 7160
rect 13556 7120 13557 7160
rect 13515 7111 13557 7120
rect 13707 7160 13749 7169
rect 13707 7120 13708 7160
rect 13748 7120 13749 7160
rect 13707 7111 13749 7120
rect 13795 7160 13853 7161
rect 13795 7120 13804 7160
rect 13844 7120 13853 7160
rect 13795 7119 13853 7120
rect 13995 7160 14037 7169
rect 13995 7120 13996 7160
rect 14036 7120 14037 7160
rect 13995 7111 14037 7120
rect 14091 7160 14133 7169
rect 14091 7120 14092 7160
rect 14132 7120 14133 7160
rect 14091 7111 14133 7120
rect 14187 7160 14229 7169
rect 14187 7120 14188 7160
rect 14228 7120 14229 7160
rect 14187 7111 14229 7120
rect 14283 7160 14325 7169
rect 14283 7120 14284 7160
rect 14324 7120 14325 7160
rect 14283 7111 14325 7120
rect 14467 7160 14525 7161
rect 14467 7120 14476 7160
rect 14516 7120 14525 7160
rect 14467 7119 14525 7120
rect 15715 7160 15773 7161
rect 15715 7120 15724 7160
rect 15764 7120 15773 7160
rect 15715 7119 15773 7120
rect 16099 7160 16157 7161
rect 16099 7120 16108 7160
rect 16148 7120 16157 7160
rect 16099 7119 16157 7120
rect 17347 7160 17405 7161
rect 17347 7120 17356 7160
rect 17396 7120 17405 7160
rect 17347 7119 17405 7120
rect 17731 7160 17789 7161
rect 17731 7120 17740 7160
rect 17780 7120 17789 7160
rect 17731 7119 17789 7120
rect 18979 7160 19037 7161
rect 18979 7120 18988 7160
rect 19028 7120 19037 7160
rect 18979 7119 19037 7120
rect 19363 7160 19421 7161
rect 19363 7120 19372 7160
rect 19412 7120 19421 7160
rect 19363 7119 19421 7120
rect 20611 7160 20669 7161
rect 20611 7120 20620 7160
rect 20660 7120 20669 7160
rect 20611 7119 20669 7120
rect 21379 7160 21437 7161
rect 21379 7120 21388 7160
rect 21428 7120 21437 7160
rect 21379 7119 21437 7120
rect 22627 7160 22685 7161
rect 22627 7120 22636 7160
rect 22676 7120 22685 7160
rect 22627 7119 22685 7120
rect 23115 7160 23157 7169
rect 23115 7120 23116 7160
rect 23156 7120 23157 7160
rect 23115 7111 23157 7120
rect 23211 7160 23253 7169
rect 23211 7120 23212 7160
rect 23252 7120 23253 7160
rect 23211 7111 23253 7120
rect 23595 7160 23637 7169
rect 23595 7120 23596 7160
rect 23636 7120 23637 7160
rect 23595 7111 23637 7120
rect 23691 7160 23733 7169
rect 24699 7162 24700 7202
rect 24740 7162 24741 7202
rect 31611 7202 31653 7211
rect 32131 7204 32140 7244
rect 32180 7204 32189 7244
rect 32131 7203 32189 7204
rect 32515 7244 32573 7245
rect 32515 7204 32524 7244
rect 32564 7204 32573 7244
rect 32515 7203 32573 7204
rect 36459 7244 36501 7253
rect 36459 7204 36460 7244
rect 36500 7204 36501 7244
rect 23691 7120 23692 7160
rect 23732 7120 23733 7160
rect 23691 7111 23733 7120
rect 24163 7160 24221 7161
rect 24163 7120 24172 7160
rect 24212 7120 24221 7160
rect 24699 7153 24741 7162
rect 25891 7160 25949 7161
rect 24163 7119 24221 7120
rect 25891 7120 25900 7160
rect 25940 7120 25949 7160
rect 25891 7119 25949 7120
rect 27139 7160 27197 7161
rect 27139 7120 27148 7160
rect 27188 7120 27197 7160
rect 27139 7119 27197 7120
rect 27523 7160 27581 7161
rect 27523 7120 27532 7160
rect 27572 7120 27581 7160
rect 27523 7119 27581 7120
rect 28771 7160 28829 7161
rect 28771 7120 28780 7160
rect 28820 7120 28829 7160
rect 28771 7119 28829 7120
rect 30027 7160 30069 7169
rect 30027 7120 30028 7160
rect 30068 7120 30069 7160
rect 30027 7111 30069 7120
rect 30123 7160 30165 7169
rect 30123 7120 30124 7160
rect 30164 7120 30165 7160
rect 30123 7111 30165 7120
rect 30507 7160 30549 7169
rect 30507 7120 30508 7160
rect 30548 7120 30549 7160
rect 30507 7111 30549 7120
rect 30603 7160 30645 7169
rect 31611 7162 31612 7202
rect 31652 7162 31653 7202
rect 36459 7195 36501 7204
rect 37987 7244 38045 7245
rect 37987 7204 37996 7244
rect 38036 7204 38045 7244
rect 37987 7203 38045 7204
rect 39051 7244 39093 7253
rect 39051 7204 39052 7244
rect 39092 7204 39093 7244
rect 39051 7195 39093 7204
rect 40675 7244 40733 7245
rect 40675 7204 40684 7244
rect 40724 7204 40733 7244
rect 40675 7203 40733 7204
rect 40867 7244 40925 7245
rect 40867 7204 40876 7244
rect 40916 7204 40925 7244
rect 40867 7203 40925 7204
rect 41251 7244 41309 7245
rect 41251 7204 41260 7244
rect 41300 7204 41309 7244
rect 41251 7203 41309 7204
rect 37419 7174 37461 7183
rect 30603 7120 30604 7160
rect 30644 7120 30645 7160
rect 30603 7111 30645 7120
rect 31075 7160 31133 7161
rect 31075 7120 31084 7160
rect 31124 7120 31133 7160
rect 31611 7153 31653 7162
rect 32899 7160 32957 7161
rect 31075 7119 31133 7120
rect 32899 7120 32908 7160
rect 32948 7120 32957 7160
rect 32899 7119 32957 7120
rect 34147 7160 34205 7161
rect 34147 7120 34156 7160
rect 34196 7120 34205 7160
rect 34147 7119 34205 7120
rect 34531 7160 34589 7161
rect 34531 7120 34540 7160
rect 34580 7120 34589 7160
rect 34531 7119 34589 7120
rect 35491 7160 35549 7161
rect 35491 7120 35500 7160
rect 35540 7120 35549 7160
rect 35491 7119 35549 7120
rect 35883 7160 35925 7169
rect 35883 7120 35884 7160
rect 35924 7120 35925 7160
rect 35883 7111 35925 7120
rect 35979 7160 36021 7169
rect 35979 7120 35980 7160
rect 36020 7120 36021 7160
rect 35979 7111 36021 7120
rect 36363 7160 36405 7169
rect 36363 7120 36364 7160
rect 36404 7120 36405 7160
rect 36363 7111 36405 7120
rect 36931 7160 36989 7161
rect 36931 7120 36940 7160
rect 36980 7120 36989 7160
rect 37419 7134 37420 7174
rect 37460 7134 37461 7174
rect 37419 7125 37461 7134
rect 38571 7160 38613 7169
rect 36931 7119 36989 7120
rect 38571 7120 38572 7160
rect 38612 7120 38613 7160
rect 38571 7111 38613 7120
rect 38667 7160 38709 7169
rect 38667 7120 38668 7160
rect 38708 7120 38709 7160
rect 38667 7111 38709 7120
rect 39147 7160 39189 7169
rect 40107 7165 40149 7174
rect 39147 7120 39148 7160
rect 39188 7120 39189 7160
rect 39147 7111 39189 7120
rect 39619 7160 39677 7161
rect 39619 7120 39628 7160
rect 39668 7120 39677 7160
rect 39619 7119 39677 7120
rect 40107 7125 40108 7165
rect 40148 7125 40149 7165
rect 40107 7116 40149 7125
rect 3819 7076 3861 7085
rect 3819 7036 3820 7076
rect 3860 7036 3861 7076
rect 3819 7027 3861 7036
rect 4587 7076 4629 7085
rect 4587 7036 4588 7076
rect 4628 7036 4629 7076
rect 4587 7027 4629 7036
rect 6699 7076 6741 7085
rect 6699 7036 6700 7076
rect 6740 7036 6741 7076
rect 6699 7027 6741 7036
rect 8811 7076 8853 7085
rect 8811 7036 8812 7076
rect 8852 7036 8853 7076
rect 8811 7027 8853 7036
rect 13611 7076 13653 7085
rect 13611 7036 13612 7076
rect 13652 7036 13653 7076
rect 13611 7027 13653 7036
rect 22827 7076 22869 7085
rect 22827 7036 22828 7076
rect 22868 7036 22869 7076
rect 22827 7027 22869 7036
rect 24843 7076 24885 7085
rect 24843 7036 24844 7076
rect 24884 7036 24885 7076
rect 24843 7027 24885 7036
rect 31755 7076 31797 7085
rect 31755 7036 31756 7076
rect 31796 7036 31797 7076
rect 31755 7027 31797 7036
rect 1227 6992 1269 7001
rect 1227 6952 1228 6992
rect 1268 6952 1269 6992
rect 1227 6943 1269 6952
rect 13323 6992 13365 7001
rect 13323 6952 13324 6992
rect 13364 6952 13365 6992
rect 13323 6943 13365 6952
rect 15915 6992 15957 7001
rect 15915 6952 15916 6992
rect 15956 6952 15957 6992
rect 15915 6943 15957 6952
rect 17547 6992 17589 7001
rect 17547 6952 17548 6992
rect 17588 6952 17589 6992
rect 17547 6943 17589 6952
rect 19179 6992 19221 7001
rect 19179 6952 19180 6992
rect 19220 6952 19221 6992
rect 19179 6943 19221 6952
rect 20811 6992 20853 7001
rect 20811 6952 20812 6992
rect 20852 6952 20853 6992
rect 20811 6943 20853 6952
rect 25035 6992 25077 7001
rect 25035 6952 25036 6992
rect 25076 6952 25077 6992
rect 25035 6943 25077 6952
rect 25419 6992 25461 7001
rect 25419 6952 25420 6992
rect 25460 6952 25461 6992
rect 25419 6943 25461 6952
rect 27339 6992 27381 7001
rect 27339 6952 27340 6992
rect 27380 6952 27381 6992
rect 27339 6943 27381 6952
rect 28971 6992 29013 7001
rect 28971 6952 28972 6992
rect 29012 6952 29013 6992
rect 28971 6943 29013 6952
rect 29163 6992 29205 7001
rect 29163 6952 29164 6992
rect 29204 6952 29205 6992
rect 29163 6943 29205 6952
rect 31947 6992 31989 7001
rect 31947 6952 31948 6992
rect 31988 6952 31989 6992
rect 31947 6943 31989 6952
rect 34347 6992 34389 7001
rect 34347 6952 34348 6992
rect 34388 6952 34389 6992
rect 34347 6943 34389 6952
rect 35019 6992 35061 7001
rect 35019 6952 35020 6992
rect 35060 6952 35061 6992
rect 35019 6943 35061 6952
rect 37611 6992 37653 7001
rect 37611 6952 37612 6992
rect 37652 6952 37653 6992
rect 37611 6943 37653 6952
rect 40299 6992 40341 7001
rect 40299 6952 40300 6992
rect 40340 6952 40341 6992
rect 40299 6943 40341 6952
rect 40491 6992 40533 7001
rect 40491 6952 40492 6992
rect 40532 6952 40533 6992
rect 40491 6943 40533 6952
rect 41067 6992 41109 7001
rect 41067 6952 41068 6992
rect 41108 6952 41109 6992
rect 41067 6943 41109 6952
rect 41451 6992 41493 7001
rect 41451 6952 41452 6992
rect 41492 6952 41493 6992
rect 41451 6943 41493 6952
rect 1152 6824 41856 6848
rect 1152 6784 4928 6824
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 5296 6784 20048 6824
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20416 6784 35168 6824
rect 35208 6784 35250 6824
rect 35290 6784 35332 6824
rect 35372 6784 35414 6824
rect 35454 6784 35496 6824
rect 35536 6784 41856 6824
rect 1152 6760 41856 6784
rect 1219 6656 1277 6657
rect 1219 6616 1228 6656
rect 1268 6616 1277 6656
rect 1219 6615 1277 6616
rect 3147 6656 3189 6665
rect 3147 6616 3148 6656
rect 3188 6616 3189 6656
rect 3147 6607 3189 6616
rect 6691 6656 6749 6657
rect 6691 6616 6700 6656
rect 6740 6616 6749 6656
rect 6691 6615 6749 6616
rect 8811 6656 8853 6665
rect 8811 6616 8812 6656
rect 8852 6616 8853 6656
rect 8811 6607 8853 6616
rect 11683 6656 11741 6657
rect 11683 6616 11692 6656
rect 11732 6616 11741 6656
rect 11683 6615 11741 6616
rect 15915 6656 15957 6665
rect 15915 6616 15916 6656
rect 15956 6616 15957 6656
rect 15915 6607 15957 6616
rect 20043 6656 20085 6665
rect 20043 6616 20044 6656
rect 20084 6616 20085 6656
rect 20043 6607 20085 6616
rect 38763 6656 38805 6665
rect 38763 6616 38764 6656
rect 38804 6616 38805 6656
rect 38763 6607 38805 6616
rect 40587 6656 40629 6665
rect 40587 6616 40588 6656
rect 40628 6616 40629 6656
rect 40587 6607 40629 6616
rect 4971 6572 5013 6581
rect 4971 6532 4972 6572
rect 5012 6532 5013 6572
rect 4971 6523 5013 6532
rect 5739 6572 5781 6581
rect 5739 6532 5740 6572
rect 5780 6532 5781 6572
rect 5739 6523 5781 6532
rect 15339 6572 15381 6581
rect 15339 6532 15340 6572
rect 15380 6532 15381 6572
rect 15339 6523 15381 6532
rect 19851 6572 19893 6581
rect 19851 6532 19852 6572
rect 19892 6532 19893 6572
rect 19851 6523 19893 6532
rect 22923 6572 22965 6581
rect 22923 6532 22924 6572
rect 22964 6532 22965 6572
rect 22923 6523 22965 6532
rect 28779 6572 28821 6581
rect 28779 6532 28780 6572
rect 28820 6532 28821 6572
rect 28779 6523 28821 6532
rect 34155 6572 34197 6581
rect 34155 6532 34156 6572
rect 34196 6532 34197 6572
rect 34155 6523 34197 6532
rect 36171 6572 36213 6581
rect 36171 6532 36172 6572
rect 36212 6532 36213 6572
rect 36171 6523 36213 6532
rect 1419 6488 1461 6497
rect 1419 6448 1420 6488
rect 1460 6448 1461 6488
rect 1419 6439 1461 6448
rect 1515 6488 1557 6497
rect 1515 6448 1516 6488
rect 1556 6448 1557 6488
rect 1515 6439 1557 6448
rect 1699 6488 1757 6489
rect 1699 6448 1708 6488
rect 1748 6448 1757 6488
rect 1699 6447 1757 6448
rect 2947 6488 3005 6489
rect 2947 6448 2956 6488
rect 2996 6448 3005 6488
rect 2947 6447 3005 6448
rect 3819 6488 3861 6497
rect 3819 6448 3820 6488
rect 3860 6448 3861 6488
rect 3819 6439 3861 6448
rect 3915 6488 3957 6497
rect 3915 6448 3916 6488
rect 3956 6448 3957 6488
rect 3915 6439 3957 6448
rect 4195 6488 4253 6489
rect 4195 6448 4204 6488
rect 4244 6448 4253 6488
rect 4195 6447 4253 6448
rect 4579 6488 4637 6489
rect 4579 6448 4588 6488
rect 4628 6448 4637 6488
rect 4579 6447 4637 6448
rect 4875 6488 4917 6497
rect 4875 6448 4876 6488
rect 4916 6448 4917 6488
rect 4875 6439 4917 6448
rect 5835 6488 5877 6497
rect 5835 6448 5836 6488
rect 5876 6448 5877 6488
rect 5835 6439 5877 6448
rect 6115 6488 6173 6489
rect 6115 6448 6124 6488
rect 6164 6448 6173 6488
rect 6115 6447 6173 6448
rect 6499 6488 6557 6489
rect 6499 6448 6508 6488
rect 6548 6448 6557 6488
rect 6499 6447 6557 6448
rect 6603 6488 6645 6497
rect 6603 6448 6604 6488
rect 6644 6448 6645 6488
rect 6603 6439 6645 6448
rect 6795 6488 6837 6497
rect 6795 6448 6796 6488
rect 6836 6448 6837 6488
rect 6795 6439 6837 6448
rect 7083 6488 7125 6497
rect 7083 6448 7084 6488
rect 7124 6448 7125 6488
rect 7083 6439 7125 6448
rect 7179 6488 7221 6497
rect 7179 6448 7180 6488
rect 7220 6448 7221 6488
rect 7179 6439 7221 6448
rect 8131 6488 8189 6489
rect 8131 6448 8140 6488
rect 8180 6448 8189 6488
rect 9099 6488 9141 6497
rect 8131 6447 8189 6448
rect 8619 6474 8661 6483
rect 8619 6434 8620 6474
rect 8660 6434 8661 6474
rect 8619 6425 8661 6434
rect 9003 6443 9045 6452
rect 7563 6404 7605 6413
rect 7563 6364 7564 6404
rect 7604 6364 7605 6404
rect 7563 6355 7605 6364
rect 7659 6404 7701 6413
rect 7659 6364 7660 6404
rect 7700 6364 7701 6404
rect 9003 6403 9004 6443
rect 9044 6403 9045 6443
rect 9099 6448 9100 6488
rect 9140 6448 9141 6488
rect 9099 6439 9141 6448
rect 9195 6488 9237 6497
rect 9195 6448 9196 6488
rect 9236 6448 9237 6488
rect 9195 6439 9237 6448
rect 9291 6488 9333 6497
rect 9291 6448 9292 6488
rect 9332 6448 9333 6488
rect 9291 6439 9333 6448
rect 9571 6488 9629 6489
rect 9571 6448 9580 6488
rect 9620 6448 9629 6488
rect 9571 6447 9629 6448
rect 10819 6488 10877 6489
rect 10819 6448 10828 6488
rect 10868 6448 10877 6488
rect 10819 6447 10877 6448
rect 11403 6488 11445 6497
rect 11403 6448 11404 6488
rect 11444 6448 11445 6488
rect 11403 6439 11445 6448
rect 11499 6488 11541 6497
rect 11499 6448 11500 6488
rect 11540 6448 11541 6488
rect 11499 6439 11541 6448
rect 11595 6488 11637 6497
rect 11595 6448 11596 6488
rect 11636 6448 11637 6488
rect 11595 6439 11637 6448
rect 11875 6488 11933 6489
rect 11875 6448 11884 6488
rect 11924 6448 11933 6488
rect 11875 6447 11933 6448
rect 13123 6488 13181 6489
rect 13123 6448 13132 6488
rect 13172 6448 13181 6488
rect 13123 6447 13181 6448
rect 13611 6488 13653 6497
rect 13611 6448 13612 6488
rect 13652 6448 13653 6488
rect 13611 6439 13653 6448
rect 13707 6488 13749 6497
rect 13707 6448 13708 6488
rect 13748 6448 13749 6488
rect 13707 6439 13749 6448
rect 14659 6488 14717 6489
rect 14659 6448 14668 6488
rect 14708 6448 14717 6488
rect 16099 6488 16157 6489
rect 14659 6447 14717 6448
rect 15195 6478 15237 6487
rect 15195 6438 15196 6478
rect 15236 6438 15237 6478
rect 16099 6448 16108 6488
rect 16148 6448 16157 6488
rect 16099 6447 16157 6448
rect 17347 6488 17405 6489
rect 17347 6448 17356 6488
rect 17396 6448 17405 6488
rect 17347 6447 17405 6448
rect 18123 6488 18165 6497
rect 18123 6448 18124 6488
rect 18164 6448 18165 6488
rect 18123 6439 18165 6448
rect 18219 6488 18261 6497
rect 18219 6448 18220 6488
rect 18260 6448 18261 6488
rect 18219 6439 18261 6448
rect 19171 6488 19229 6489
rect 19171 6448 19180 6488
rect 19220 6448 19229 6488
rect 21195 6488 21237 6497
rect 19171 6447 19229 6448
rect 19707 6478 19749 6487
rect 15195 6429 15237 6438
rect 19707 6438 19708 6478
rect 19748 6438 19749 6478
rect 21195 6448 21196 6488
rect 21236 6448 21237 6488
rect 21195 6439 21237 6448
rect 21291 6488 21333 6497
rect 21291 6448 21292 6488
rect 21332 6448 21333 6488
rect 21291 6439 21333 6448
rect 22243 6488 22301 6489
rect 22243 6448 22252 6488
rect 22292 6448 22301 6488
rect 22243 6447 22301 6448
rect 22731 6483 22773 6492
rect 22731 6443 22732 6483
rect 22772 6443 22773 6483
rect 23107 6488 23165 6489
rect 23107 6448 23116 6488
rect 23156 6448 23165 6488
rect 23107 6447 23165 6448
rect 24355 6488 24413 6489
rect 24355 6448 24364 6488
rect 24404 6448 24413 6488
rect 24355 6447 24413 6448
rect 24931 6488 24989 6489
rect 24931 6448 24940 6488
rect 24980 6448 24989 6488
rect 24931 6447 24989 6448
rect 26179 6488 26237 6489
rect 26179 6448 26188 6488
rect 26228 6448 26237 6488
rect 26179 6447 26237 6448
rect 27051 6488 27093 6497
rect 27051 6448 27052 6488
rect 27092 6448 27093 6488
rect 19707 6429 19749 6438
rect 22731 6434 22773 6443
rect 27051 6439 27093 6448
rect 27147 6488 27189 6497
rect 27147 6448 27148 6488
rect 27188 6448 27189 6488
rect 27147 6439 27189 6448
rect 27531 6488 27573 6497
rect 27531 6448 27532 6488
rect 27572 6448 27573 6488
rect 27531 6439 27573 6448
rect 28099 6488 28157 6489
rect 28099 6448 28108 6488
rect 28148 6448 28157 6488
rect 29155 6488 29213 6489
rect 28099 6447 28157 6448
rect 28635 6478 28677 6487
rect 28635 6438 28636 6478
rect 28676 6438 28677 6478
rect 29155 6448 29164 6488
rect 29204 6448 29213 6488
rect 29155 6447 29213 6448
rect 30403 6488 30461 6489
rect 30403 6448 30412 6488
rect 30452 6448 30461 6488
rect 30403 6447 30461 6448
rect 30691 6488 30749 6489
rect 30691 6448 30700 6488
rect 30740 6448 30749 6488
rect 30691 6447 30749 6448
rect 31939 6488 31997 6489
rect 31939 6448 31948 6488
rect 31988 6448 31997 6488
rect 31939 6447 31997 6448
rect 32427 6488 32469 6497
rect 32427 6448 32428 6488
rect 32468 6448 32469 6488
rect 32427 6439 32469 6448
rect 32523 6488 32565 6497
rect 32523 6448 32524 6488
rect 32564 6448 32565 6488
rect 32523 6439 32565 6448
rect 33475 6488 33533 6489
rect 33475 6448 33484 6488
rect 33524 6448 33533 6488
rect 33475 6447 33533 6448
rect 33963 6483 34005 6492
rect 33963 6443 33964 6483
rect 34004 6443 34005 6483
rect 28635 6429 28677 6438
rect 33963 6434 34005 6443
rect 34443 6488 34485 6497
rect 34443 6448 34444 6488
rect 34484 6448 34485 6488
rect 34443 6439 34485 6448
rect 34539 6488 34581 6497
rect 34539 6448 34540 6488
rect 34580 6448 34581 6488
rect 34539 6439 34581 6448
rect 34923 6488 34965 6497
rect 34923 6448 34924 6488
rect 34964 6448 34965 6488
rect 34923 6439 34965 6448
rect 35491 6488 35549 6489
rect 35491 6448 35500 6488
rect 35540 6448 35549 6488
rect 37315 6488 37373 6489
rect 35491 6447 35549 6448
rect 36027 6478 36069 6487
rect 36027 6438 36028 6478
rect 36068 6438 36069 6478
rect 37315 6448 37324 6488
rect 37364 6448 37373 6488
rect 37315 6447 37373 6448
rect 38563 6488 38621 6489
rect 38563 6448 38572 6488
rect 38612 6448 38621 6488
rect 38563 6447 38621 6448
rect 39139 6488 39197 6489
rect 39139 6448 39148 6488
rect 39188 6448 39197 6488
rect 39139 6447 39197 6448
rect 40387 6488 40445 6489
rect 40387 6448 40396 6488
rect 40436 6448 40445 6488
rect 40387 6447 40445 6448
rect 36027 6429 36069 6438
rect 9003 6394 9045 6403
rect 14091 6404 14133 6413
rect 7659 6355 7701 6364
rect 14091 6364 14092 6404
rect 14132 6364 14133 6404
rect 14091 6355 14133 6364
rect 14187 6404 14229 6413
rect 14187 6364 14188 6404
rect 14228 6364 14229 6404
rect 14187 6355 14229 6364
rect 15715 6404 15773 6405
rect 15715 6364 15724 6404
rect 15764 6364 15773 6404
rect 15715 6363 15773 6364
rect 18603 6404 18645 6413
rect 18603 6364 18604 6404
rect 18644 6364 18645 6404
rect 18603 6355 18645 6364
rect 18699 6404 18741 6413
rect 18699 6364 18700 6404
rect 18740 6364 18741 6404
rect 18699 6355 18741 6364
rect 20227 6404 20285 6405
rect 20227 6364 20236 6404
rect 20276 6364 20285 6404
rect 20227 6363 20285 6364
rect 21675 6404 21717 6413
rect 21675 6364 21676 6404
rect 21716 6364 21717 6404
rect 21675 6355 21717 6364
rect 21771 6404 21813 6413
rect 21771 6364 21772 6404
rect 21812 6364 21813 6404
rect 21771 6355 21813 6364
rect 27627 6404 27669 6413
rect 27627 6364 27628 6404
rect 27668 6364 27669 6404
rect 27627 6355 27669 6364
rect 32907 6404 32949 6413
rect 32907 6364 32908 6404
rect 32948 6364 32949 6404
rect 32907 6355 32949 6364
rect 33003 6404 33045 6413
rect 33003 6364 33004 6404
rect 33044 6364 33045 6404
rect 33003 6355 33045 6364
rect 35019 6404 35061 6413
rect 35019 6364 35020 6404
rect 35060 6364 35061 6404
rect 35019 6355 35061 6364
rect 40867 6404 40925 6405
rect 40867 6364 40876 6404
rect 40916 6364 40925 6404
rect 40867 6363 40925 6364
rect 41251 6404 41309 6405
rect 41251 6364 41260 6404
rect 41300 6364 41309 6404
rect 41251 6363 41309 6364
rect 5251 6320 5309 6321
rect 5251 6280 5260 6320
rect 5300 6280 5309 6320
rect 5251 6279 5309 6280
rect 5443 6320 5501 6321
rect 5443 6280 5452 6320
rect 5492 6280 5501 6320
rect 5443 6279 5501 6280
rect 17547 6320 17589 6329
rect 17547 6280 17548 6320
rect 17588 6280 17589 6320
rect 17547 6271 17589 6280
rect 36363 6320 36405 6329
rect 36363 6280 36364 6320
rect 36404 6280 36405 6320
rect 36363 6271 36405 6280
rect 36747 6320 36789 6329
rect 36747 6280 36748 6320
rect 36788 6280 36789 6320
rect 36747 6271 36789 6280
rect 41067 6320 41109 6329
rect 41067 6280 41068 6320
rect 41108 6280 41109 6320
rect 41067 6271 41109 6280
rect 3523 6236 3581 6237
rect 3523 6196 3532 6236
rect 3572 6196 3581 6236
rect 3523 6195 3581 6196
rect 11019 6236 11061 6245
rect 11019 6196 11020 6236
rect 11060 6196 11061 6236
rect 11019 6187 11061 6196
rect 13323 6236 13365 6245
rect 13323 6196 13324 6236
rect 13364 6196 13365 6236
rect 13323 6187 13365 6196
rect 24555 6236 24597 6245
rect 24555 6196 24556 6236
rect 24596 6196 24597 6236
rect 24555 6187 24597 6196
rect 26379 6236 26421 6245
rect 26379 6196 26380 6236
rect 26420 6196 26421 6236
rect 26379 6187 26421 6196
rect 28971 6236 29013 6245
rect 28971 6196 28972 6236
rect 29012 6196 29013 6236
rect 28971 6187 29013 6196
rect 32139 6236 32181 6245
rect 32139 6196 32140 6236
rect 32180 6196 32181 6236
rect 32139 6187 32181 6196
rect 41451 6236 41493 6245
rect 41451 6196 41452 6236
rect 41492 6196 41493 6236
rect 41451 6187 41493 6196
rect 1152 6068 41856 6092
rect 1152 6028 3688 6068
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 4056 6028 18808 6068
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 19176 6028 33928 6068
rect 33968 6028 34010 6068
rect 34050 6028 34092 6068
rect 34132 6028 34174 6068
rect 34214 6028 34256 6068
rect 34296 6028 41856 6068
rect 1152 6004 41856 6028
rect 3147 5900 3189 5909
rect 3147 5860 3148 5900
rect 3188 5860 3189 5900
rect 3147 5851 3189 5860
rect 5827 5900 5885 5901
rect 5827 5860 5836 5900
rect 5876 5860 5885 5900
rect 5827 5859 5885 5860
rect 8131 5900 8189 5901
rect 8131 5860 8140 5900
rect 8180 5860 8189 5900
rect 8131 5859 8189 5860
rect 31659 5900 31701 5909
rect 31659 5860 31660 5900
rect 31700 5860 31701 5900
rect 31659 5851 31701 5860
rect 34251 5900 34293 5909
rect 34251 5860 34252 5900
rect 34292 5860 34293 5900
rect 34251 5851 34293 5860
rect 36171 5900 36213 5909
rect 36171 5860 36172 5900
rect 36212 5860 36213 5900
rect 36171 5851 36213 5860
rect 41451 5900 41493 5909
rect 41451 5860 41452 5900
rect 41492 5860 41493 5900
rect 41451 5851 41493 5860
rect 3715 5816 3773 5817
rect 3715 5776 3724 5816
rect 3764 5776 3773 5816
rect 3715 5775 3773 5776
rect 4683 5816 4725 5825
rect 4683 5776 4684 5816
rect 4724 5776 4725 5816
rect 4683 5767 4725 5776
rect 10059 5816 10101 5825
rect 10059 5776 10060 5816
rect 10100 5776 10101 5816
rect 10059 5767 10101 5776
rect 41067 5816 41109 5825
rect 41067 5776 41068 5816
rect 41108 5776 41109 5816
rect 41067 5767 41109 5776
rect 6603 5732 6645 5741
rect 6603 5692 6604 5732
rect 6644 5692 6645 5732
rect 6603 5683 6645 5692
rect 13227 5732 13269 5741
rect 13227 5692 13228 5732
rect 13268 5692 13269 5732
rect 13227 5683 13269 5692
rect 21099 5732 21141 5741
rect 21099 5692 21100 5732
rect 21140 5692 21141 5732
rect 21099 5683 21141 5692
rect 22819 5732 22877 5733
rect 22819 5692 22828 5732
rect 22868 5692 22877 5732
rect 22819 5691 22877 5692
rect 23203 5732 23261 5733
rect 23203 5692 23212 5732
rect 23252 5692 23261 5732
rect 23203 5691 23261 5692
rect 23875 5732 23933 5733
rect 23875 5692 23884 5732
rect 23924 5692 23933 5732
rect 26467 5732 26525 5733
rect 23875 5691 23933 5692
rect 25947 5690 25989 5699
rect 26467 5692 26476 5732
rect 26516 5692 26525 5732
rect 26467 5691 26525 5692
rect 27139 5732 27197 5733
rect 27139 5692 27148 5732
rect 27188 5692 27197 5732
rect 27139 5691 27197 5692
rect 29931 5732 29973 5741
rect 29931 5692 29932 5732
rect 29972 5692 29973 5732
rect 8523 5667 8565 5676
rect 7659 5657 7701 5666
rect 1227 5648 1269 5657
rect 1227 5608 1228 5648
rect 1268 5608 1269 5648
rect 1227 5599 1269 5608
rect 1419 5648 1461 5657
rect 1419 5608 1420 5648
rect 1460 5608 1461 5648
rect 1419 5599 1461 5608
rect 1507 5648 1565 5649
rect 1507 5608 1516 5648
rect 1556 5608 1565 5648
rect 1507 5607 1565 5608
rect 1699 5648 1757 5649
rect 1699 5608 1708 5648
rect 1748 5608 1757 5648
rect 1699 5607 1757 5608
rect 2947 5648 3005 5649
rect 2947 5608 2956 5648
rect 2996 5608 3005 5648
rect 2947 5607 3005 5608
rect 3339 5648 3381 5657
rect 3339 5608 3340 5648
rect 3380 5608 3381 5648
rect 3339 5599 3381 5608
rect 3523 5648 3581 5649
rect 3523 5608 3532 5648
rect 3572 5608 3581 5648
rect 3523 5607 3581 5608
rect 4107 5648 4149 5657
rect 4107 5608 4108 5648
rect 4148 5608 4149 5648
rect 4107 5599 4149 5608
rect 4387 5648 4445 5649
rect 4387 5608 4396 5648
rect 4436 5608 4445 5648
rect 4387 5607 4445 5608
rect 4683 5648 4725 5657
rect 4683 5608 4684 5648
rect 4724 5608 4725 5648
rect 4683 5599 4725 5608
rect 4875 5648 4917 5657
rect 4875 5608 4876 5648
rect 4916 5608 4917 5648
rect 4875 5599 4917 5608
rect 5155 5648 5213 5649
rect 5155 5608 5164 5648
rect 5204 5608 5213 5648
rect 5155 5607 5213 5608
rect 5451 5648 5493 5657
rect 5451 5608 5452 5648
rect 5492 5608 5493 5648
rect 5451 5599 5493 5608
rect 6123 5648 6165 5657
rect 6123 5608 6124 5648
rect 6164 5608 6165 5648
rect 6123 5599 6165 5608
rect 6219 5648 6261 5657
rect 6219 5608 6220 5648
rect 6260 5608 6261 5648
rect 6219 5599 6261 5608
rect 6699 5648 6741 5657
rect 6699 5608 6700 5648
rect 6740 5608 6741 5648
rect 6699 5599 6741 5608
rect 7171 5648 7229 5649
rect 7171 5608 7180 5648
rect 7220 5608 7229 5648
rect 7659 5617 7660 5657
rect 7700 5617 7701 5657
rect 8523 5627 8524 5667
rect 8564 5627 8565 5667
rect 18027 5667 18069 5676
rect 8523 5618 8565 5627
rect 8803 5648 8861 5649
rect 7659 5608 7701 5617
rect 8803 5608 8812 5648
rect 8852 5608 8861 5648
rect 7171 5607 7229 5608
rect 8803 5607 8861 5608
rect 9099 5648 9141 5657
rect 9099 5608 9100 5648
rect 9140 5608 9141 5648
rect 9099 5599 9141 5608
rect 9195 5648 9237 5657
rect 9195 5608 9196 5648
rect 9236 5608 9237 5648
rect 9195 5599 9237 5608
rect 9675 5648 9717 5657
rect 9675 5608 9676 5648
rect 9716 5608 9717 5648
rect 9675 5599 9717 5608
rect 9771 5648 9813 5657
rect 9771 5608 9772 5648
rect 9812 5608 9813 5648
rect 9771 5599 9813 5608
rect 9867 5648 9909 5657
rect 9867 5608 9868 5648
rect 9908 5608 9909 5648
rect 9867 5599 9909 5608
rect 10059 5648 10101 5657
rect 10059 5608 10060 5648
rect 10100 5608 10101 5648
rect 10059 5599 10101 5608
rect 10251 5648 10293 5657
rect 10251 5608 10252 5648
rect 10292 5608 10293 5648
rect 10251 5599 10293 5608
rect 10339 5648 10397 5649
rect 10339 5608 10348 5648
rect 10388 5608 10397 5648
rect 10339 5607 10397 5608
rect 10531 5648 10589 5649
rect 10531 5608 10540 5648
rect 10580 5608 10589 5648
rect 10531 5607 10589 5608
rect 10915 5648 10973 5649
rect 10915 5608 10924 5648
rect 10964 5608 10973 5648
rect 10915 5607 10973 5608
rect 12163 5648 12221 5649
rect 12163 5608 12172 5648
rect 12212 5608 12221 5648
rect 12163 5607 12221 5608
rect 12651 5648 12693 5657
rect 12651 5608 12652 5648
rect 12692 5608 12693 5648
rect 12651 5599 12693 5608
rect 12747 5648 12789 5657
rect 12747 5608 12748 5648
rect 12788 5608 12789 5648
rect 12747 5599 12789 5608
rect 13131 5648 13173 5657
rect 14187 5653 14229 5662
rect 13131 5608 13132 5648
rect 13172 5608 13173 5648
rect 13131 5599 13173 5608
rect 13699 5648 13757 5649
rect 13699 5608 13708 5648
rect 13748 5608 13757 5648
rect 13699 5607 13757 5608
rect 14187 5613 14188 5653
rect 14228 5613 14229 5653
rect 14187 5604 14229 5613
rect 16195 5648 16253 5649
rect 16195 5608 16204 5648
rect 16244 5608 16253 5648
rect 16195 5607 16253 5608
rect 17443 5648 17501 5649
rect 17443 5608 17452 5648
rect 17492 5608 17501 5648
rect 17443 5607 17501 5608
rect 17931 5648 17973 5657
rect 17931 5608 17932 5648
rect 17972 5608 17973 5648
rect 18027 5627 18028 5667
rect 18068 5627 18069 5667
rect 19467 5662 19509 5671
rect 18027 5618 18069 5627
rect 18411 5648 18453 5657
rect 17931 5599 17973 5608
rect 18411 5608 18412 5648
rect 18452 5608 18453 5648
rect 18411 5599 18453 5608
rect 18507 5648 18549 5657
rect 18507 5608 18508 5648
rect 18548 5608 18549 5648
rect 18507 5599 18549 5608
rect 18979 5648 19037 5649
rect 18979 5608 18988 5648
rect 19028 5608 19037 5648
rect 19467 5622 19468 5662
rect 19508 5622 19509 5662
rect 22155 5662 22197 5671
rect 19467 5613 19509 5622
rect 20619 5648 20661 5657
rect 18979 5607 19037 5608
rect 20619 5608 20620 5648
rect 20660 5608 20661 5648
rect 20619 5599 20661 5608
rect 20715 5648 20757 5657
rect 20715 5608 20716 5648
rect 20756 5608 20757 5648
rect 20715 5599 20757 5608
rect 21195 5648 21237 5657
rect 21195 5608 21196 5648
rect 21236 5608 21237 5648
rect 21195 5599 21237 5608
rect 21667 5648 21725 5649
rect 21667 5608 21676 5648
rect 21716 5608 21725 5648
rect 22155 5622 22156 5662
rect 22196 5622 22197 5662
rect 22155 5613 22197 5622
rect 24363 5648 24405 5657
rect 21667 5607 21725 5608
rect 24363 5608 24364 5648
rect 24404 5608 24405 5648
rect 24363 5599 24405 5608
rect 24459 5648 24501 5657
rect 24459 5608 24460 5648
rect 24500 5608 24501 5648
rect 24459 5599 24501 5608
rect 24843 5648 24885 5657
rect 24843 5608 24844 5648
rect 24884 5608 24885 5648
rect 24843 5599 24885 5608
rect 24939 5648 24981 5657
rect 25947 5650 25948 5690
rect 25988 5650 25989 5690
rect 29931 5683 29973 5692
rect 31459 5732 31517 5733
rect 31459 5692 31468 5732
rect 31508 5692 31517 5732
rect 31459 5691 31517 5692
rect 31843 5732 31901 5733
rect 31843 5692 31852 5732
rect 31892 5692 31901 5732
rect 31843 5691 31901 5692
rect 32811 5732 32853 5741
rect 32811 5692 32812 5732
rect 32852 5692 32853 5732
rect 32811 5683 32853 5692
rect 34435 5732 34493 5733
rect 34435 5692 34444 5732
rect 34484 5692 34493 5732
rect 34435 5691 34493 5692
rect 36547 5732 36605 5733
rect 36547 5692 36556 5732
rect 36596 5692 36605 5732
rect 36547 5691 36605 5692
rect 37219 5732 37277 5733
rect 37219 5692 37228 5732
rect 37268 5692 37277 5732
rect 37219 5691 37277 5692
rect 40099 5732 40157 5733
rect 40099 5692 40108 5732
rect 40148 5692 40157 5732
rect 40099 5691 40157 5692
rect 40483 5732 40541 5733
rect 40483 5692 40492 5732
rect 40532 5692 40541 5732
rect 40483 5691 40541 5692
rect 40867 5732 40925 5733
rect 40867 5692 40876 5732
rect 40916 5692 40925 5732
rect 40867 5691 40925 5692
rect 41251 5732 41309 5733
rect 41251 5692 41260 5732
rect 41300 5692 41309 5732
rect 41251 5691 41309 5692
rect 30939 5657 30981 5666
rect 33867 5662 33909 5671
rect 24939 5608 24940 5648
rect 24980 5608 24981 5648
rect 24939 5599 24981 5608
rect 25411 5648 25469 5649
rect 25411 5608 25420 5648
rect 25460 5608 25469 5648
rect 25947 5641 25989 5650
rect 27619 5648 27677 5649
rect 25411 5607 25469 5608
rect 27619 5608 27628 5648
rect 27668 5608 27677 5648
rect 27619 5607 27677 5608
rect 28867 5648 28925 5649
rect 28867 5608 28876 5648
rect 28916 5608 28925 5648
rect 28867 5607 28925 5608
rect 29355 5648 29397 5657
rect 29355 5608 29356 5648
rect 29396 5608 29397 5648
rect 29355 5599 29397 5608
rect 29451 5648 29493 5657
rect 29451 5608 29452 5648
rect 29492 5608 29493 5648
rect 29451 5599 29493 5608
rect 29835 5648 29877 5657
rect 29835 5608 29836 5648
rect 29876 5608 29877 5648
rect 29835 5599 29877 5608
rect 30403 5648 30461 5649
rect 30403 5608 30412 5648
rect 30452 5608 30461 5648
rect 30939 5617 30940 5657
rect 30980 5617 30981 5657
rect 30939 5608 30981 5617
rect 32331 5648 32373 5657
rect 32331 5608 32332 5648
rect 32372 5608 32373 5648
rect 30403 5607 30461 5608
rect 32331 5599 32373 5608
rect 32427 5648 32469 5657
rect 32427 5608 32428 5648
rect 32468 5608 32469 5648
rect 32427 5599 32469 5608
rect 32907 5648 32949 5657
rect 32907 5608 32908 5648
rect 32948 5608 32949 5648
rect 32907 5599 32949 5608
rect 33379 5648 33437 5649
rect 33379 5608 33388 5648
rect 33428 5608 33437 5648
rect 33867 5622 33868 5662
rect 33908 5622 33909 5662
rect 39099 5657 39141 5666
rect 33867 5613 33909 5622
rect 34723 5648 34781 5649
rect 33379 5607 33437 5608
rect 34723 5608 34732 5648
rect 34772 5608 34781 5648
rect 34723 5607 34781 5608
rect 35971 5648 36029 5649
rect 35971 5608 35980 5648
rect 36020 5608 36029 5648
rect 35971 5607 36029 5608
rect 37515 5648 37557 5657
rect 37515 5608 37516 5648
rect 37556 5608 37557 5648
rect 37515 5599 37557 5608
rect 37611 5648 37653 5657
rect 37611 5608 37612 5648
rect 37652 5608 37653 5648
rect 37611 5599 37653 5608
rect 37995 5648 38037 5657
rect 37995 5608 37996 5648
rect 38036 5608 38037 5648
rect 37995 5599 38037 5608
rect 38091 5648 38133 5657
rect 38091 5608 38092 5648
rect 38132 5608 38133 5648
rect 38091 5599 38133 5608
rect 38563 5648 38621 5649
rect 38563 5608 38572 5648
rect 38612 5608 38621 5648
rect 39099 5617 39100 5657
rect 39140 5617 39141 5657
rect 39099 5608 39141 5617
rect 38563 5607 38621 5608
rect 3435 5564 3477 5573
rect 3435 5524 3436 5564
rect 3476 5524 3477 5564
rect 3435 5515 3477 5524
rect 4011 5564 4053 5573
rect 4011 5524 4012 5564
rect 4052 5524 4053 5564
rect 4011 5515 4053 5524
rect 5547 5564 5589 5573
rect 5547 5524 5548 5564
rect 5588 5524 5589 5564
rect 5547 5515 5589 5524
rect 8427 5564 8469 5573
rect 8427 5524 8428 5564
rect 8468 5524 8469 5564
rect 8427 5515 8469 5524
rect 12363 5564 12405 5573
rect 12363 5524 12364 5564
rect 12404 5524 12405 5564
rect 12363 5515 12405 5524
rect 22347 5564 22389 5573
rect 22347 5524 22348 5564
rect 22388 5524 22389 5564
rect 22347 5515 22389 5524
rect 26091 5564 26133 5573
rect 26091 5524 26092 5564
rect 26132 5524 26133 5564
rect 26091 5515 26133 5524
rect 29067 5564 29109 5573
rect 29067 5524 29068 5564
rect 29108 5524 29109 5564
rect 29067 5515 29109 5524
rect 31083 5564 31125 5573
rect 31083 5524 31084 5564
rect 31124 5524 31125 5564
rect 31083 5515 31125 5524
rect 1315 5480 1373 5481
rect 1315 5440 1324 5480
rect 1364 5440 1373 5480
rect 1315 5439 1373 5440
rect 3147 5480 3189 5489
rect 3147 5440 3148 5480
rect 3188 5440 3189 5480
rect 3147 5431 3189 5440
rect 7851 5480 7893 5489
rect 7851 5440 7852 5480
rect 7892 5440 7893 5480
rect 7851 5431 7893 5440
rect 9379 5480 9437 5481
rect 9379 5440 9388 5480
rect 9428 5440 9437 5480
rect 9379 5439 9437 5440
rect 9571 5480 9629 5481
rect 9571 5440 9580 5480
rect 9620 5440 9629 5480
rect 9571 5439 9629 5440
rect 10635 5480 10677 5489
rect 10635 5440 10636 5480
rect 10676 5440 10677 5480
rect 10635 5431 10677 5440
rect 14379 5480 14421 5489
rect 14379 5440 14380 5480
rect 14420 5440 14421 5480
rect 14379 5431 14421 5440
rect 17643 5480 17685 5489
rect 17643 5440 17644 5480
rect 17684 5440 17685 5480
rect 17643 5431 17685 5440
rect 19659 5480 19701 5489
rect 19659 5440 19660 5480
rect 19700 5440 19701 5480
rect 19659 5431 19701 5440
rect 22635 5480 22677 5489
rect 22635 5440 22636 5480
rect 22676 5440 22677 5480
rect 22635 5431 22677 5440
rect 23019 5480 23061 5489
rect 23019 5440 23020 5480
rect 23060 5440 23061 5480
rect 23019 5431 23061 5440
rect 24075 5480 24117 5489
rect 24075 5440 24076 5480
rect 24116 5440 24117 5480
rect 24075 5431 24117 5440
rect 26283 5480 26325 5489
rect 26283 5440 26284 5480
rect 26324 5440 26325 5480
rect 26283 5431 26325 5440
rect 27339 5480 27381 5489
rect 27339 5440 27340 5480
rect 27380 5440 27381 5480
rect 27339 5431 27381 5440
rect 31275 5480 31317 5489
rect 31275 5440 31276 5480
rect 31316 5440 31317 5480
rect 31275 5431 31317 5440
rect 34059 5480 34101 5489
rect 34059 5440 34060 5480
rect 34100 5440 34101 5480
rect 34059 5431 34101 5440
rect 36363 5480 36405 5489
rect 36363 5440 36364 5480
rect 36404 5440 36405 5480
rect 36363 5431 36405 5440
rect 37035 5480 37077 5489
rect 37035 5440 37036 5480
rect 37076 5440 37077 5480
rect 37035 5431 37077 5440
rect 39243 5480 39285 5489
rect 39243 5440 39244 5480
rect 39284 5440 39285 5480
rect 39243 5431 39285 5440
rect 39915 5480 39957 5489
rect 39915 5440 39916 5480
rect 39956 5440 39957 5480
rect 39915 5431 39957 5440
rect 40683 5480 40725 5489
rect 40683 5440 40684 5480
rect 40724 5440 40725 5480
rect 40683 5431 40725 5440
rect 1152 5312 41856 5336
rect 1152 5272 4928 5312
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 5296 5272 20048 5312
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20416 5272 35168 5312
rect 35208 5272 35250 5312
rect 35290 5272 35332 5312
rect 35372 5272 35414 5312
rect 35454 5272 35496 5312
rect 35536 5272 41856 5312
rect 1152 5248 41856 5272
rect 3531 5186 3573 5195
rect 3531 5146 3532 5186
rect 3572 5146 3573 5186
rect 3531 5137 3573 5146
rect 6507 5144 6549 5153
rect 6507 5104 6508 5144
rect 6548 5104 6549 5144
rect 6507 5095 6549 5104
rect 8715 5144 8757 5153
rect 8715 5104 8716 5144
rect 8756 5104 8757 5144
rect 8715 5095 8757 5104
rect 13995 5144 14037 5153
rect 13995 5104 13996 5144
rect 14036 5104 14037 5144
rect 13995 5095 14037 5104
rect 31083 5144 31125 5153
rect 31083 5104 31084 5144
rect 31124 5104 31125 5144
rect 31083 5095 31125 5104
rect 36267 5144 36309 5153
rect 36267 5104 36268 5144
rect 36308 5104 36309 5144
rect 36267 5095 36309 5104
rect 3147 5060 3189 5069
rect 3147 5020 3148 5060
rect 3188 5020 3189 5060
rect 3147 5011 3189 5020
rect 3819 5060 3861 5069
rect 3819 5020 3820 5060
rect 3860 5020 3861 5060
rect 3819 5011 3861 5020
rect 8523 5060 8565 5069
rect 8523 5020 8524 5060
rect 8564 5020 8565 5060
rect 8523 5011 8565 5020
rect 16299 5060 16341 5069
rect 16299 5020 16300 5060
rect 16340 5020 16341 5060
rect 16299 5011 16341 5020
rect 18315 5060 18357 5069
rect 18315 5020 18316 5060
rect 18356 5020 18357 5060
rect 18315 5011 18357 5020
rect 34635 5060 34677 5069
rect 34635 5020 34636 5060
rect 34676 5020 34677 5060
rect 34635 5011 34677 5020
rect 36939 5060 36981 5069
rect 36939 5020 36940 5060
rect 36980 5020 36981 5060
rect 36939 5011 36981 5020
rect 1315 4976 1373 4977
rect 1315 4936 1324 4976
rect 1364 4936 1373 4976
rect 1315 4935 1373 4936
rect 2563 4976 2621 4977
rect 2563 4936 2572 4976
rect 2612 4936 2621 4976
rect 2563 4935 2621 4936
rect 3051 4976 3093 4985
rect 3051 4936 3052 4976
rect 3092 4936 3093 4976
rect 3051 4927 3093 4936
rect 3243 4976 3285 4985
rect 3243 4936 3244 4976
rect 3284 4936 3285 4976
rect 3243 4927 3285 4936
rect 3331 4976 3389 4977
rect 3331 4936 3340 4976
rect 3380 4936 3389 4976
rect 3331 4935 3389 4936
rect 3915 4976 3957 4985
rect 3915 4936 3916 4976
rect 3956 4936 3957 4976
rect 3915 4927 3957 4936
rect 4195 4976 4253 4977
rect 4195 4936 4204 4976
rect 4244 4936 4253 4976
rect 4195 4935 4253 4936
rect 4587 4976 4629 4985
rect 4587 4936 4588 4976
rect 4628 4936 4629 4976
rect 4587 4927 4629 4936
rect 4683 4976 4725 4985
rect 4683 4936 4684 4976
rect 4724 4936 4725 4976
rect 4683 4927 4725 4936
rect 4779 4976 4821 4985
rect 4779 4936 4780 4976
rect 4820 4936 4821 4976
rect 4779 4927 4821 4936
rect 4875 4976 4917 4985
rect 4875 4936 4876 4976
rect 4916 4936 4917 4976
rect 4875 4927 4917 4936
rect 5059 4976 5117 4977
rect 5059 4936 5068 4976
rect 5108 4936 5117 4976
rect 5059 4935 5117 4936
rect 6307 4976 6365 4977
rect 6307 4936 6316 4976
rect 6356 4936 6365 4976
rect 6307 4935 6365 4936
rect 6795 4976 6837 4985
rect 6795 4936 6796 4976
rect 6836 4936 6837 4976
rect 6795 4927 6837 4936
rect 6891 4976 6933 4985
rect 6891 4936 6892 4976
rect 6932 4936 6933 4976
rect 6891 4927 6933 4936
rect 7275 4976 7317 4985
rect 7275 4936 7276 4976
rect 7316 4936 7317 4976
rect 7275 4927 7317 4936
rect 7371 4976 7413 4985
rect 7371 4936 7372 4976
rect 7412 4936 7413 4976
rect 7371 4927 7413 4936
rect 7843 4976 7901 4977
rect 7843 4936 7852 4976
rect 7892 4936 7901 4976
rect 8899 4976 8957 4977
rect 7843 4935 7901 4936
rect 8331 4962 8373 4971
rect 8331 4922 8332 4962
rect 8372 4922 8373 4962
rect 8899 4936 8908 4976
rect 8948 4936 8957 4976
rect 8899 4935 8957 4936
rect 10147 4976 10205 4977
rect 10147 4936 10156 4976
rect 10196 4936 10205 4976
rect 10147 4935 10205 4936
rect 10435 4976 10493 4977
rect 10435 4936 10444 4976
rect 10484 4936 10493 4976
rect 10435 4935 10493 4936
rect 11683 4976 11741 4977
rect 11683 4936 11692 4976
rect 11732 4936 11741 4976
rect 11683 4935 11741 4936
rect 12075 4976 12117 4985
rect 12075 4936 12076 4976
rect 12116 4936 12117 4976
rect 12075 4927 12117 4936
rect 12171 4976 12213 4985
rect 12171 4936 12172 4976
rect 12212 4936 12213 4976
rect 12171 4927 12213 4936
rect 12267 4976 12309 4985
rect 12267 4936 12268 4976
rect 12308 4936 12309 4976
rect 12267 4927 12309 4936
rect 12363 4976 12405 4985
rect 12363 4936 12364 4976
rect 12404 4936 12405 4976
rect 12363 4927 12405 4936
rect 12547 4976 12605 4977
rect 12547 4936 12556 4976
rect 12596 4936 12605 4976
rect 12547 4935 12605 4936
rect 13795 4976 13853 4977
rect 13795 4936 13804 4976
rect 13844 4936 13853 4976
rect 13795 4935 13853 4936
rect 14851 4976 14909 4977
rect 14851 4936 14860 4976
rect 14900 4936 14909 4976
rect 14851 4935 14909 4936
rect 16099 4976 16157 4977
rect 16099 4936 16108 4976
rect 16148 4936 16157 4976
rect 16099 4935 16157 4936
rect 16587 4976 16629 4985
rect 16587 4936 16588 4976
rect 16628 4936 16629 4976
rect 16587 4927 16629 4936
rect 16683 4976 16725 4985
rect 16683 4936 16684 4976
rect 16724 4936 16725 4976
rect 16683 4927 16725 4936
rect 17067 4976 17109 4985
rect 17067 4936 17068 4976
rect 17108 4936 17109 4976
rect 17067 4927 17109 4936
rect 17163 4976 17205 4985
rect 17163 4936 17164 4976
rect 17204 4936 17205 4976
rect 17163 4927 17205 4936
rect 17635 4976 17693 4977
rect 17635 4936 17644 4976
rect 17684 4936 17693 4976
rect 17635 4935 17693 4936
rect 18123 4971 18165 4980
rect 18123 4931 18124 4971
rect 18164 4931 18165 4971
rect 22051 4976 22109 4977
rect 22051 4936 22060 4976
rect 22100 4936 22109 4976
rect 22051 4935 22109 4936
rect 23299 4976 23357 4977
rect 23299 4936 23308 4976
rect 23348 4936 23357 4976
rect 23299 4935 23357 4936
rect 24547 4976 24605 4977
rect 24547 4936 24556 4976
rect 24596 4936 24605 4976
rect 24547 4935 24605 4936
rect 25795 4976 25853 4977
rect 25795 4936 25804 4976
rect 25844 4936 25853 4976
rect 25795 4935 25853 4936
rect 26947 4976 27005 4977
rect 26947 4936 26956 4976
rect 26996 4936 27005 4976
rect 26947 4935 27005 4936
rect 28195 4976 28253 4977
rect 28195 4936 28204 4976
rect 28244 4936 28253 4976
rect 28195 4935 28253 4936
rect 29635 4976 29693 4977
rect 29635 4936 29644 4976
rect 29684 4936 29693 4976
rect 29635 4935 29693 4936
rect 30883 4976 30941 4977
rect 30883 4936 30892 4976
rect 30932 4936 30941 4976
rect 30883 4935 30941 4936
rect 31267 4976 31325 4977
rect 31267 4936 31276 4976
rect 31316 4936 31325 4976
rect 31267 4935 31325 4936
rect 32515 4976 32573 4977
rect 32515 4936 32524 4976
rect 32564 4936 32573 4976
rect 32515 4935 32573 4936
rect 33187 4976 33245 4977
rect 33187 4936 33196 4976
rect 33236 4936 33245 4976
rect 33187 4935 33245 4936
rect 34435 4976 34493 4977
rect 34435 4936 34444 4976
rect 34484 4936 34493 4976
rect 34435 4935 34493 4936
rect 35779 4976 35837 4977
rect 35779 4936 35788 4976
rect 35828 4936 35837 4976
rect 35779 4935 35837 4936
rect 37123 4976 37181 4977
rect 37123 4936 37132 4976
rect 37172 4936 37181 4976
rect 37123 4935 37181 4936
rect 38371 4976 38429 4977
rect 38371 4936 38380 4976
rect 38420 4936 38429 4976
rect 38371 4935 38429 4936
rect 38755 4976 38813 4977
rect 38755 4936 38764 4976
rect 38804 4936 38813 4976
rect 38755 4935 38813 4936
rect 40003 4976 40061 4977
rect 40003 4936 40012 4976
rect 40052 4936 40061 4976
rect 40003 4935 40061 4936
rect 18123 4922 18165 4931
rect 8331 4913 8373 4922
rect 20227 4892 20285 4893
rect 20227 4852 20236 4892
rect 20276 4852 20285 4892
rect 20227 4851 20285 4852
rect 20995 4892 21053 4893
rect 20995 4852 21004 4892
rect 21044 4852 21053 4892
rect 20995 4851 21053 4852
rect 26563 4892 26621 4893
rect 26563 4852 26572 4892
rect 26612 4852 26621 4892
rect 26563 4851 26621 4852
rect 28771 4892 28829 4893
rect 28771 4852 28780 4892
rect 28820 4852 28829 4892
rect 28771 4851 28829 4852
rect 29443 4892 29501 4893
rect 29443 4852 29452 4892
rect 29492 4852 29501 4892
rect 29443 4851 29501 4852
rect 35011 4892 35069 4893
rect 35011 4852 35020 4892
rect 35060 4852 35069 4892
rect 35011 4851 35069 4852
rect 35395 4892 35453 4893
rect 35395 4852 35404 4892
rect 35444 4852 35453 4892
rect 35395 4851 35453 4852
rect 40483 4892 40541 4893
rect 40483 4852 40492 4892
rect 40532 4852 40541 4892
rect 40483 4851 40541 4852
rect 40867 4892 40925 4893
rect 40867 4852 40876 4892
rect 40916 4852 40925 4892
rect 40867 4851 40925 4852
rect 41251 4892 41309 4893
rect 41251 4852 41260 4892
rect 41300 4852 41309 4892
rect 41251 4851 41309 4852
rect 2763 4808 2805 4817
rect 2763 4768 2764 4808
rect 2804 4768 2805 4808
rect 2763 4759 2805 4768
rect 35211 4808 35253 4817
rect 35211 4768 35212 4808
rect 35252 4768 35253 4808
rect 35211 4759 35253 4768
rect 40683 4808 40725 4817
rect 40683 4768 40684 4808
rect 40724 4768 40725 4808
rect 40683 4759 40725 4768
rect 41067 4808 41109 4817
rect 41067 4768 41068 4808
rect 41108 4768 41109 4808
rect 41067 4759 41109 4768
rect 41451 4808 41493 4817
rect 41451 4768 41452 4808
rect 41492 4768 41493 4808
rect 41451 4759 41493 4768
rect 11883 4724 11925 4733
rect 11883 4684 11884 4724
rect 11924 4684 11925 4724
rect 11883 4675 11925 4684
rect 20427 4724 20469 4733
rect 20427 4684 20428 4724
rect 20468 4684 20469 4724
rect 20427 4675 20469 4684
rect 21195 4724 21237 4733
rect 21195 4684 21196 4724
rect 21236 4684 21237 4724
rect 21195 4675 21237 4684
rect 23499 4724 23541 4733
rect 23499 4684 23500 4724
rect 23540 4684 23541 4724
rect 23499 4675 23541 4684
rect 25995 4724 26037 4733
rect 25995 4684 25996 4724
rect 26036 4684 26037 4724
rect 25995 4675 26037 4684
rect 26763 4724 26805 4733
rect 26763 4684 26764 4724
rect 26804 4684 26805 4724
rect 26763 4675 26805 4684
rect 28395 4724 28437 4733
rect 28395 4684 28396 4724
rect 28436 4684 28437 4724
rect 28395 4675 28437 4684
rect 28587 4724 28629 4733
rect 28587 4684 28588 4724
rect 28628 4684 28629 4724
rect 28587 4675 28629 4684
rect 29259 4724 29301 4733
rect 29259 4684 29260 4724
rect 29300 4684 29301 4724
rect 29259 4675 29301 4684
rect 32715 4724 32757 4733
rect 32715 4684 32716 4724
rect 32756 4684 32757 4724
rect 32715 4675 32757 4684
rect 34827 4724 34869 4733
rect 34827 4684 34828 4724
rect 34868 4684 34869 4724
rect 34827 4675 34869 4684
rect 38571 4724 38613 4733
rect 38571 4684 38572 4724
rect 38612 4684 38613 4724
rect 38571 4675 38613 4684
rect 1152 4556 41856 4580
rect 1152 4516 3688 4556
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 4056 4516 18808 4556
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 19176 4516 33928 4556
rect 33968 4516 34010 4556
rect 34050 4516 34092 4556
rect 34132 4516 34174 4556
rect 34214 4516 34256 4556
rect 34296 4516 41856 4556
rect 1152 4492 41856 4516
rect 8995 4388 9053 4389
rect 8995 4348 9004 4388
rect 9044 4348 9053 4388
rect 8995 4347 9053 4348
rect 37227 4388 37269 4397
rect 37227 4348 37228 4388
rect 37268 4348 37269 4388
rect 37227 4339 37269 4348
rect 39243 4388 39285 4397
rect 39243 4348 39244 4388
rect 39284 4348 39285 4388
rect 39243 4339 39285 4348
rect 41067 4388 41109 4397
rect 41067 4348 41068 4388
rect 41108 4348 41109 4388
rect 41067 4339 41109 4348
rect 40299 4304 40341 4313
rect 40299 4264 40300 4304
rect 40340 4264 40341 4304
rect 40299 4255 40341 4264
rect 4203 4220 4245 4229
rect 4203 4180 4204 4220
rect 4244 4180 4245 4220
rect 4203 4171 4245 4180
rect 4299 4220 4341 4229
rect 4299 4180 4300 4220
rect 4340 4180 4341 4220
rect 4299 4171 4341 4180
rect 6699 4220 6741 4229
rect 6699 4180 6700 4220
rect 6740 4180 6741 4220
rect 18027 4220 18069 4229
rect 6699 4171 6741 4180
rect 15771 4178 15813 4187
rect 3243 4150 3285 4159
rect 1411 4136 1469 4137
rect 1411 4096 1420 4136
rect 1460 4096 1469 4136
rect 1411 4095 1469 4096
rect 2659 4136 2717 4137
rect 2659 4096 2668 4136
rect 2708 4096 2717 4136
rect 3243 4110 3244 4150
rect 3284 4110 3285 4150
rect 7659 4150 7701 4159
rect 3243 4101 3285 4110
rect 3715 4136 3773 4137
rect 2659 4095 2717 4096
rect 3715 4096 3724 4136
rect 3764 4096 3773 4136
rect 3715 4095 3773 4096
rect 4683 4136 4725 4145
rect 4683 4096 4684 4136
rect 4724 4096 4725 4136
rect 4683 4087 4725 4096
rect 4779 4136 4821 4145
rect 4779 4096 4780 4136
rect 4820 4096 4821 4136
rect 4779 4087 4821 4096
rect 5067 4136 5109 4145
rect 5067 4096 5068 4136
rect 5108 4096 5109 4136
rect 5067 4087 5109 4096
rect 5163 4136 5205 4145
rect 5163 4096 5164 4136
rect 5204 4096 5205 4136
rect 5163 4087 5205 4096
rect 5355 4136 5397 4145
rect 5355 4096 5356 4136
rect 5396 4096 5397 4136
rect 5355 4087 5397 4096
rect 5547 4136 5589 4145
rect 5547 4096 5548 4136
rect 5588 4096 5589 4136
rect 5547 4087 5589 4096
rect 5643 4136 5685 4145
rect 5643 4096 5644 4136
rect 5684 4096 5685 4136
rect 5643 4087 5685 4096
rect 5739 4136 5781 4145
rect 5739 4096 5740 4136
rect 5780 4096 5781 4136
rect 5739 4087 5781 4096
rect 5835 4136 5877 4145
rect 5835 4096 5836 4136
rect 5876 4096 5877 4136
rect 5835 4087 5877 4096
rect 6123 4136 6165 4145
rect 6123 4096 6124 4136
rect 6164 4096 6165 4136
rect 6123 4087 6165 4096
rect 6219 4136 6261 4145
rect 6219 4096 6220 4136
rect 6260 4096 6261 4136
rect 6219 4087 6261 4096
rect 6603 4136 6645 4145
rect 6603 4096 6604 4136
rect 6644 4096 6645 4136
rect 6603 4087 6645 4096
rect 7171 4136 7229 4137
rect 7171 4096 7180 4136
rect 7220 4096 7229 4136
rect 7659 4110 7660 4150
rect 7700 4110 7701 4150
rect 7659 4101 7701 4110
rect 8323 4136 8381 4137
rect 7171 4095 7229 4096
rect 8323 4096 8332 4136
rect 8372 4096 8381 4136
rect 8323 4095 8381 4096
rect 8619 4136 8661 4145
rect 8619 4096 8620 4136
rect 8660 4096 8661 4136
rect 8619 4087 8661 4096
rect 8715 4136 8757 4145
rect 8715 4096 8716 4136
rect 8756 4096 8757 4136
rect 8715 4087 8757 4096
rect 9187 4136 9245 4137
rect 9187 4096 9196 4136
rect 9236 4096 9245 4136
rect 9187 4095 9245 4096
rect 10435 4136 10493 4137
rect 10435 4096 10444 4136
rect 10484 4096 10493 4136
rect 10435 4095 10493 4096
rect 10819 4136 10877 4137
rect 10819 4096 10828 4136
rect 10868 4096 10877 4136
rect 10819 4095 10877 4096
rect 12067 4136 12125 4137
rect 12067 4096 12076 4136
rect 12116 4096 12125 4136
rect 12067 4095 12125 4096
rect 12451 4136 12509 4137
rect 12451 4096 12460 4136
rect 12500 4096 12509 4136
rect 12451 4095 12509 4096
rect 13699 4136 13757 4137
rect 13699 4096 13708 4136
rect 13748 4096 13757 4136
rect 13699 4095 13757 4096
rect 14187 4136 14229 4145
rect 14187 4096 14188 4136
rect 14228 4096 14229 4136
rect 14187 4087 14229 4096
rect 14283 4136 14325 4145
rect 14283 4096 14284 4136
rect 14324 4096 14325 4136
rect 14283 4087 14325 4096
rect 14667 4136 14709 4145
rect 14667 4096 14668 4136
rect 14708 4096 14709 4136
rect 14667 4087 14709 4096
rect 14763 4136 14805 4145
rect 15771 4138 15772 4178
rect 15812 4138 15813 4178
rect 18027 4180 18028 4220
rect 18068 4180 18069 4220
rect 18027 4171 18069 4180
rect 18123 4220 18165 4229
rect 18123 4180 18124 4220
rect 18164 4180 18165 4220
rect 24843 4220 24885 4229
rect 18123 4171 18165 4180
rect 22251 4178 22293 4187
rect 14763 4096 14764 4136
rect 14804 4096 14805 4136
rect 14763 4087 14805 4096
rect 15235 4136 15293 4137
rect 15235 4096 15244 4136
rect 15284 4096 15293 4136
rect 15771 4129 15813 4138
rect 17547 4136 17589 4145
rect 15235 4095 15293 4096
rect 17547 4096 17548 4136
rect 17588 4096 17589 4136
rect 17547 4087 17589 4096
rect 17643 4136 17685 4145
rect 19083 4141 19125 4150
rect 17643 4096 17644 4136
rect 17684 4096 17685 4136
rect 17643 4087 17685 4096
rect 18595 4136 18653 4137
rect 18595 4096 18604 4136
rect 18644 4096 18653 4136
rect 18595 4095 18653 4096
rect 19083 4101 19084 4141
rect 19124 4101 19125 4141
rect 19083 4092 19125 4101
rect 20035 4136 20093 4137
rect 20035 4096 20044 4136
rect 20084 4096 20093 4136
rect 20035 4095 20093 4096
rect 21283 4136 21341 4137
rect 21283 4096 21292 4136
rect 21332 4096 21341 4136
rect 21283 4095 21341 4096
rect 21771 4136 21813 4145
rect 21771 4096 21772 4136
rect 21812 4096 21813 4136
rect 21771 4087 21813 4096
rect 21867 4136 21909 4145
rect 21867 4096 21868 4136
rect 21908 4096 21909 4136
rect 22251 4138 22252 4178
rect 22292 4138 22293 4178
rect 22251 4129 22293 4138
rect 22347 4178 22389 4187
rect 22347 4138 22348 4178
rect 22388 4138 22389 4178
rect 22347 4129 22389 4138
rect 23355 4178 23397 4187
rect 23355 4138 23356 4178
rect 23396 4138 23397 4178
rect 24843 4180 24844 4220
rect 24884 4180 24885 4220
rect 24843 4171 24885 4180
rect 28587 4220 28629 4229
rect 28587 4180 28588 4220
rect 28628 4180 28629 4220
rect 28587 4171 28629 4180
rect 32035 4220 32093 4221
rect 32035 4180 32044 4220
rect 32084 4180 32093 4220
rect 32035 4179 32093 4180
rect 32907 4220 32949 4229
rect 32907 4180 32908 4220
rect 32948 4180 32949 4220
rect 32907 4171 32949 4180
rect 34435 4220 34493 4221
rect 34435 4180 34444 4220
rect 34484 4180 34493 4220
rect 34435 4179 34493 4180
rect 35011 4220 35069 4221
rect 35011 4180 35020 4220
rect 35060 4180 35069 4220
rect 35011 4179 35069 4180
rect 35787 4220 35829 4229
rect 35787 4180 35788 4220
rect 35828 4180 35829 4220
rect 35787 4171 35829 4180
rect 35883 4220 35925 4229
rect 35883 4180 35884 4220
rect 35924 4180 35925 4220
rect 35883 4171 35925 4180
rect 37411 4220 37469 4221
rect 37411 4180 37420 4220
rect 37460 4180 37469 4220
rect 37411 4179 37469 4180
rect 39619 4220 39677 4221
rect 39619 4180 39628 4220
rect 39668 4180 39677 4220
rect 39619 4179 39677 4180
rect 39907 4220 39965 4221
rect 39907 4180 39916 4220
rect 39956 4180 39965 4220
rect 39907 4179 39965 4180
rect 40483 4220 40541 4221
rect 40483 4180 40492 4220
rect 40532 4180 40541 4220
rect 40483 4179 40541 4180
rect 40867 4220 40925 4221
rect 40867 4180 40876 4220
rect 40916 4180 40925 4220
rect 40867 4179 40925 4180
rect 41251 4220 41309 4221
rect 41251 4180 41260 4220
rect 41300 4180 41309 4220
rect 41251 4179 41309 4180
rect 25851 4145 25893 4154
rect 29643 4150 29685 4159
rect 22819 4136 22877 4137
rect 21867 4087 21909 4096
rect 22819 4096 22828 4136
rect 22868 4096 22877 4136
rect 23355 4129 23397 4138
rect 24267 4136 24309 4145
rect 22819 4095 22877 4096
rect 24267 4096 24268 4136
rect 24308 4096 24309 4136
rect 24267 4087 24309 4096
rect 24363 4136 24405 4145
rect 24363 4096 24364 4136
rect 24404 4096 24405 4136
rect 24363 4087 24405 4096
rect 24747 4136 24789 4145
rect 24747 4096 24748 4136
rect 24788 4096 24789 4136
rect 24747 4087 24789 4096
rect 25315 4136 25373 4137
rect 25315 4096 25324 4136
rect 25364 4096 25373 4136
rect 25851 4105 25852 4145
rect 25892 4105 25893 4145
rect 25851 4096 25893 4105
rect 26179 4136 26237 4137
rect 26179 4096 26188 4136
rect 26228 4096 26237 4136
rect 25315 4095 25373 4096
rect 26179 4095 26237 4096
rect 27427 4136 27485 4137
rect 27427 4096 27436 4136
rect 27476 4096 27485 4136
rect 27427 4095 27485 4096
rect 28107 4136 28149 4145
rect 28107 4096 28108 4136
rect 28148 4096 28149 4136
rect 28107 4087 28149 4096
rect 28203 4136 28245 4145
rect 28203 4096 28204 4136
rect 28244 4096 28245 4136
rect 28203 4087 28245 4096
rect 28683 4136 28725 4145
rect 28683 4096 28684 4136
rect 28724 4096 28725 4136
rect 28683 4087 28725 4096
rect 29155 4136 29213 4137
rect 29155 4096 29164 4136
rect 29204 4096 29213 4136
rect 29643 4110 29644 4150
rect 29684 4110 29685 4150
rect 32331 4155 32373 4164
rect 29643 4101 29685 4110
rect 30211 4136 30269 4137
rect 29155 4095 29213 4096
rect 30211 4096 30220 4136
rect 30260 4096 30269 4136
rect 30211 4095 30269 4096
rect 31459 4136 31517 4137
rect 31459 4096 31468 4136
rect 31508 4096 31517 4136
rect 32331 4115 32332 4155
rect 32372 4115 32373 4155
rect 32331 4106 32373 4115
rect 32427 4136 32469 4145
rect 31459 4095 31517 4096
rect 32427 4096 32428 4136
rect 32468 4096 32469 4136
rect 32427 4087 32469 4096
rect 32811 4136 32853 4145
rect 33867 4141 33909 4150
rect 32811 4096 32812 4136
rect 32852 4096 32853 4136
rect 32811 4087 32853 4096
rect 33379 4136 33437 4137
rect 33379 4096 33388 4136
rect 33428 4096 33437 4136
rect 33379 4095 33437 4096
rect 33867 4101 33868 4141
rect 33908 4101 33909 4141
rect 33867 4092 33909 4101
rect 35307 4136 35349 4145
rect 35307 4096 35308 4136
rect 35348 4096 35349 4136
rect 35307 4087 35349 4096
rect 35403 4136 35445 4145
rect 36843 4141 36885 4150
rect 35403 4096 35404 4136
rect 35444 4096 35445 4136
rect 35403 4087 35445 4096
rect 36355 4136 36413 4137
rect 36355 4096 36364 4136
rect 36404 4096 36413 4136
rect 36355 4095 36413 4096
rect 36843 4101 36844 4141
rect 36884 4101 36885 4141
rect 36843 4092 36885 4101
rect 37795 4136 37853 4137
rect 37795 4096 37804 4136
rect 37844 4096 37853 4136
rect 37795 4095 37853 4096
rect 39043 4136 39101 4137
rect 39043 4096 39052 4136
rect 39092 4096 39101 4136
rect 39043 4095 39101 4096
rect 21483 4052 21525 4061
rect 21483 4012 21484 4052
rect 21524 4012 21525 4052
rect 21483 4003 21525 4012
rect 25995 4052 26037 4061
rect 25995 4012 25996 4052
rect 26036 4012 26037 4052
rect 25995 4003 26037 4012
rect 34059 4052 34101 4061
rect 34059 4012 34060 4052
rect 34100 4012 34101 4052
rect 34059 4003 34101 4012
rect 37035 4052 37077 4061
rect 37035 4012 37036 4052
rect 37076 4012 37077 4052
rect 37035 4003 37077 4012
rect 2859 3968 2901 3977
rect 2859 3928 2860 3968
rect 2900 3928 2901 3968
rect 2859 3919 2901 3928
rect 3051 3968 3093 3977
rect 3051 3928 3052 3968
rect 3092 3928 3093 3968
rect 3051 3919 3093 3928
rect 7851 3968 7893 3977
rect 7851 3928 7852 3968
rect 7892 3928 7893 3968
rect 7851 3919 7893 3928
rect 10635 3968 10677 3977
rect 10635 3928 10636 3968
rect 10676 3928 10677 3968
rect 10635 3919 10677 3928
rect 12267 3968 12309 3977
rect 12267 3928 12268 3968
rect 12308 3928 12309 3968
rect 12267 3919 12309 3928
rect 13899 3968 13941 3977
rect 13899 3928 13900 3968
rect 13940 3928 13941 3968
rect 13899 3919 13941 3928
rect 15915 3968 15957 3977
rect 15915 3928 15916 3968
rect 15956 3928 15957 3968
rect 15915 3919 15957 3928
rect 19275 3968 19317 3977
rect 19275 3928 19276 3968
rect 19316 3928 19317 3968
rect 19275 3919 19317 3928
rect 23499 3968 23541 3977
rect 23499 3928 23500 3968
rect 23540 3928 23541 3968
rect 23499 3919 23541 3928
rect 27627 3968 27669 3977
rect 27627 3928 27628 3968
rect 27668 3928 27669 3968
rect 27627 3919 27669 3928
rect 29835 3968 29877 3977
rect 29835 3928 29836 3968
rect 29876 3928 29877 3968
rect 29835 3919 29877 3928
rect 30027 3968 30069 3977
rect 30027 3928 30028 3968
rect 30068 3928 30069 3968
rect 30027 3919 30069 3928
rect 31851 3968 31893 3977
rect 31851 3928 31852 3968
rect 31892 3928 31893 3968
rect 31851 3919 31893 3928
rect 34251 3968 34293 3977
rect 34251 3928 34252 3968
rect 34292 3928 34293 3968
rect 34251 3919 34293 3928
rect 34827 3968 34869 3977
rect 34827 3928 34828 3968
rect 34868 3928 34869 3968
rect 34827 3919 34869 3928
rect 39435 3968 39477 3977
rect 39435 3928 39436 3968
rect 39476 3928 39477 3968
rect 39435 3919 39477 3928
rect 40107 3968 40149 3977
rect 40107 3928 40108 3968
rect 40148 3928 40149 3968
rect 40107 3919 40149 3928
rect 41451 3968 41493 3977
rect 41451 3928 41452 3968
rect 41492 3928 41493 3968
rect 41451 3919 41493 3928
rect 1152 3800 41856 3824
rect 1152 3760 4928 3800
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 5296 3760 20048 3800
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20416 3760 35168 3800
rect 35208 3760 35250 3800
rect 35290 3760 35332 3800
rect 35372 3760 35414 3800
rect 35454 3760 35496 3800
rect 35536 3760 41856 3800
rect 1152 3736 41856 3760
rect 3051 3632 3093 3641
rect 3051 3592 3052 3632
rect 3092 3592 3093 3632
rect 3051 3583 3093 3592
rect 3523 3632 3581 3633
rect 3523 3592 3532 3632
rect 3572 3592 3581 3632
rect 3523 3591 3581 3592
rect 4195 3632 4253 3633
rect 4195 3592 4204 3632
rect 4244 3592 4253 3632
rect 4195 3591 4253 3592
rect 5931 3632 5973 3641
rect 5931 3592 5932 3632
rect 5972 3592 5973 3632
rect 5931 3583 5973 3592
rect 17451 3632 17493 3641
rect 17451 3592 17452 3632
rect 17492 3592 17493 3632
rect 17451 3583 17493 3592
rect 19083 3632 19125 3641
rect 19083 3592 19084 3632
rect 19124 3592 19125 3632
rect 19083 3583 19125 3592
rect 24555 3632 24597 3641
rect 24555 3592 24556 3632
rect 24596 3592 24597 3632
rect 24555 3583 24597 3592
rect 29931 3632 29973 3641
rect 29931 3592 29932 3632
rect 29972 3592 29973 3632
rect 29931 3583 29973 3592
rect 32139 3632 32181 3641
rect 32139 3592 32140 3632
rect 32180 3592 32181 3632
rect 32139 3583 32181 3592
rect 32331 3632 32373 3641
rect 32331 3592 32332 3632
rect 32372 3592 32373 3632
rect 32331 3583 32373 3592
rect 34443 3632 34485 3641
rect 34443 3592 34444 3632
rect 34484 3592 34485 3632
rect 34443 3583 34485 3592
rect 34635 3632 34677 3641
rect 34635 3592 34636 3632
rect 34676 3592 34677 3632
rect 34635 3583 34677 3592
rect 41067 3632 41109 3641
rect 41067 3592 41068 3632
rect 41108 3592 41109 3632
rect 41067 3583 41109 3592
rect 8331 3548 8373 3557
rect 8331 3508 8332 3548
rect 8372 3508 8373 3548
rect 8331 3499 8373 3508
rect 10443 3548 10485 3557
rect 10443 3508 10444 3548
rect 10484 3508 10485 3548
rect 10443 3499 10485 3508
rect 12459 3548 12501 3557
rect 12459 3508 12460 3548
rect 12500 3508 12501 3548
rect 12459 3499 12501 3508
rect 14859 3548 14901 3557
rect 14859 3508 14860 3548
rect 14900 3508 14901 3548
rect 14859 3499 14901 3508
rect 27243 3548 27285 3557
rect 27243 3508 27244 3548
rect 27284 3508 27285 3548
rect 27243 3499 27285 3508
rect 39147 3548 39189 3557
rect 39147 3508 39148 3548
rect 39188 3508 39189 3548
rect 39147 3499 39189 3508
rect 1411 3485 1469 3486
rect 1227 3464 1269 3473
rect 1227 3424 1228 3464
rect 1268 3424 1269 3464
rect 1411 3445 1420 3485
rect 1460 3445 1469 3485
rect 1411 3444 1469 3445
rect 1603 3464 1661 3465
rect 1227 3415 1269 3424
rect 1603 3424 1612 3464
rect 1652 3424 1661 3464
rect 1603 3423 1661 3424
rect 2851 3464 2909 3465
rect 2851 3424 2860 3464
rect 2900 3424 2909 3464
rect 2851 3423 2909 3424
rect 3243 3464 3285 3473
rect 3243 3424 3244 3464
rect 3284 3424 3285 3464
rect 3243 3415 3285 3424
rect 3339 3464 3381 3473
rect 3339 3424 3340 3464
rect 3380 3424 3381 3464
rect 3339 3415 3381 3424
rect 3435 3464 3477 3473
rect 3435 3424 3436 3464
rect 3476 3424 3477 3464
rect 3435 3415 3477 3424
rect 3715 3464 3773 3465
rect 3715 3424 3724 3464
rect 3764 3424 3773 3464
rect 3715 3423 3773 3424
rect 3811 3464 3869 3465
rect 3811 3424 3820 3464
rect 3860 3424 3869 3464
rect 3811 3423 3869 3424
rect 4011 3464 4053 3473
rect 4011 3424 4012 3464
rect 4052 3424 4053 3464
rect 4011 3415 4053 3424
rect 4107 3464 4149 3473
rect 4107 3424 4108 3464
rect 4148 3424 4149 3464
rect 4107 3415 4149 3424
rect 4200 3464 4258 3465
rect 4200 3424 4209 3464
rect 4249 3424 4258 3464
rect 4200 3423 4258 3424
rect 4483 3464 4541 3465
rect 4483 3424 4492 3464
rect 4532 3424 4541 3464
rect 4483 3423 4541 3424
rect 5731 3464 5789 3465
rect 5731 3424 5740 3464
rect 5780 3424 5789 3464
rect 5731 3423 5789 3424
rect 6403 3464 6461 3465
rect 6403 3424 6412 3464
rect 6452 3424 6461 3464
rect 6403 3423 6461 3424
rect 7651 3464 7709 3465
rect 7651 3424 7660 3464
rect 7700 3424 7709 3464
rect 7651 3423 7709 3424
rect 7939 3464 7997 3465
rect 7939 3424 7948 3464
rect 7988 3424 7997 3464
rect 7939 3423 7997 3424
rect 8235 3464 8277 3473
rect 8235 3424 8236 3464
rect 8276 3424 8277 3464
rect 8235 3415 8277 3424
rect 8995 3464 9053 3465
rect 8995 3424 9004 3464
rect 9044 3424 9053 3464
rect 8995 3423 9053 3424
rect 10243 3464 10301 3465
rect 10243 3424 10252 3464
rect 10292 3424 10301 3464
rect 10243 3423 10301 3424
rect 10731 3464 10773 3473
rect 10731 3424 10732 3464
rect 10772 3424 10773 3464
rect 10731 3415 10773 3424
rect 10827 3464 10869 3473
rect 10827 3424 10828 3464
rect 10868 3424 10869 3464
rect 10827 3415 10869 3424
rect 11307 3464 11349 3473
rect 11307 3424 11308 3464
rect 11348 3424 11349 3464
rect 11307 3415 11349 3424
rect 11779 3464 11837 3465
rect 11779 3424 11788 3464
rect 11828 3424 11837 3464
rect 11779 3423 11837 3424
rect 12267 3459 12309 3468
rect 12267 3419 12268 3459
rect 12308 3419 12309 3459
rect 12267 3410 12309 3419
rect 13131 3464 13173 3473
rect 13131 3424 13132 3464
rect 13172 3424 13173 3464
rect 13131 3415 13173 3424
rect 13227 3464 13269 3473
rect 13227 3424 13228 3464
rect 13268 3424 13269 3464
rect 13227 3415 13269 3424
rect 13611 3464 13653 3473
rect 13611 3424 13612 3464
rect 13652 3424 13653 3464
rect 13611 3415 13653 3424
rect 14179 3464 14237 3465
rect 14179 3424 14188 3464
rect 14228 3424 14237 3464
rect 14179 3423 14237 3424
rect 14667 3459 14709 3468
rect 14667 3419 14668 3459
rect 14708 3419 14709 3459
rect 16003 3464 16061 3465
rect 16003 3424 16012 3464
rect 16052 3424 16061 3464
rect 16003 3423 16061 3424
rect 17251 3464 17309 3465
rect 17251 3424 17260 3464
rect 17300 3424 17309 3464
rect 17251 3423 17309 3424
rect 17635 3464 17693 3465
rect 17635 3424 17644 3464
rect 17684 3424 17693 3464
rect 17635 3423 17693 3424
rect 18883 3464 18941 3465
rect 18883 3424 18892 3464
rect 18932 3424 18941 3464
rect 18883 3423 18941 3424
rect 20515 3464 20573 3465
rect 20515 3424 20524 3464
rect 20564 3424 20573 3464
rect 20515 3423 20573 3424
rect 21763 3464 21821 3465
rect 21763 3424 21772 3464
rect 21812 3424 21821 3464
rect 21763 3423 21821 3424
rect 23107 3464 23165 3465
rect 23107 3424 23116 3464
rect 23156 3424 23165 3464
rect 23107 3423 23165 3424
rect 24355 3464 24413 3465
rect 24355 3424 24364 3464
rect 24404 3424 24413 3464
rect 24355 3423 24413 3424
rect 25515 3464 25557 3473
rect 25515 3424 25516 3464
rect 25556 3424 25557 3464
rect 14667 3410 14709 3419
rect 25515 3415 25557 3424
rect 25611 3464 25653 3473
rect 25611 3424 25612 3464
rect 25652 3424 25653 3464
rect 25611 3415 25653 3424
rect 26091 3464 26133 3473
rect 26091 3424 26092 3464
rect 26132 3424 26133 3464
rect 26091 3415 26133 3424
rect 26563 3464 26621 3465
rect 26563 3424 26572 3464
rect 26612 3424 26621 3464
rect 28203 3464 28245 3473
rect 26563 3423 26621 3424
rect 27051 3450 27093 3459
rect 27051 3410 27052 3450
rect 27092 3410 27093 3450
rect 28203 3424 28204 3464
rect 28244 3424 28245 3464
rect 28203 3415 28245 3424
rect 28299 3464 28341 3473
rect 28299 3424 28300 3464
rect 28340 3424 28341 3464
rect 28299 3415 28341 3424
rect 28683 3464 28725 3473
rect 28683 3424 28684 3464
rect 28724 3424 28725 3464
rect 28683 3415 28725 3424
rect 29251 3464 29309 3465
rect 29251 3424 29260 3464
rect 29300 3424 29309 3464
rect 30411 3464 30453 3473
rect 29251 3423 29309 3424
rect 29739 3450 29781 3459
rect 27051 3401 27093 3410
rect 29739 3410 29740 3450
rect 29780 3410 29781 3450
rect 30411 3424 30412 3464
rect 30452 3424 30453 3464
rect 30411 3415 30453 3424
rect 30507 3464 30549 3473
rect 30507 3424 30508 3464
rect 30548 3424 30549 3464
rect 30507 3415 30549 3424
rect 30987 3464 31029 3473
rect 30987 3424 30988 3464
rect 31028 3424 31029 3464
rect 30987 3415 31029 3424
rect 31459 3464 31517 3465
rect 31459 3424 31468 3464
rect 31508 3424 31517 3464
rect 32995 3464 33053 3465
rect 31459 3423 31517 3424
rect 31947 3450 31989 3459
rect 29739 3401 29781 3410
rect 31947 3410 31948 3450
rect 31988 3410 31989 3450
rect 32995 3424 33004 3464
rect 33044 3424 33053 3464
rect 32995 3423 33053 3424
rect 34243 3464 34301 3465
rect 34243 3424 34252 3464
rect 34292 3424 34301 3464
rect 34243 3423 34301 3424
rect 34819 3464 34877 3465
rect 34819 3424 34828 3464
rect 34868 3424 34877 3464
rect 34819 3423 34877 3424
rect 36067 3464 36125 3465
rect 36067 3424 36076 3464
rect 36116 3424 36125 3464
rect 36067 3423 36125 3424
rect 37419 3464 37461 3473
rect 37419 3424 37420 3464
rect 37460 3424 37461 3464
rect 37419 3415 37461 3424
rect 37515 3464 37557 3473
rect 37515 3424 37516 3464
rect 37556 3424 37557 3464
rect 37515 3415 37557 3424
rect 37995 3464 38037 3473
rect 37995 3424 37996 3464
rect 38036 3424 38037 3464
rect 37995 3415 38037 3424
rect 38467 3464 38525 3465
rect 38467 3424 38476 3464
rect 38516 3424 38525 3464
rect 38467 3423 38525 3424
rect 38955 3459 38997 3468
rect 38955 3419 38956 3459
rect 38996 3419 38997 3459
rect 38955 3410 38997 3419
rect 31947 3401 31989 3410
rect 11211 3380 11253 3389
rect 11211 3340 11212 3380
rect 11252 3340 11253 3380
rect 11211 3331 11253 3340
rect 12643 3380 12701 3381
rect 12643 3340 12652 3380
rect 12692 3340 12701 3380
rect 12643 3339 12701 3340
rect 13707 3380 13749 3389
rect 13707 3340 13708 3380
rect 13748 3340 13749 3380
rect 13707 3331 13749 3340
rect 19939 3380 19997 3381
rect 19939 3340 19948 3380
rect 19988 3340 19997 3380
rect 19939 3339 19997 3340
rect 22723 3380 22781 3381
rect 22723 3340 22732 3380
rect 22772 3340 22781 3380
rect 22723 3339 22781 3340
rect 25219 3380 25277 3381
rect 25219 3340 25228 3380
rect 25268 3340 25277 3380
rect 25219 3339 25277 3340
rect 25995 3380 26037 3389
rect 25995 3340 25996 3380
rect 26036 3340 26037 3380
rect 25995 3331 26037 3340
rect 27619 3380 27677 3381
rect 27619 3340 27628 3380
rect 27668 3340 27677 3380
rect 27619 3339 27677 3340
rect 28779 3380 28821 3389
rect 28779 3340 28780 3380
rect 28820 3340 28821 3380
rect 28779 3331 28821 3340
rect 30891 3380 30933 3389
rect 30891 3340 30892 3380
rect 30932 3340 30933 3380
rect 30891 3331 30933 3340
rect 32515 3380 32573 3381
rect 32515 3340 32524 3380
rect 32564 3340 32573 3380
rect 32515 3339 32573 3340
rect 36451 3380 36509 3381
rect 36451 3340 36460 3380
rect 36500 3340 36509 3380
rect 36451 3339 36509 3340
rect 37123 3380 37181 3381
rect 37123 3340 37132 3380
rect 37172 3340 37181 3380
rect 37123 3339 37181 3340
rect 37899 3380 37941 3389
rect 37899 3340 37900 3380
rect 37940 3340 37941 3380
rect 37899 3331 37941 3340
rect 39331 3380 39389 3381
rect 39331 3340 39340 3380
rect 39380 3340 39389 3380
rect 39331 3339 39389 3340
rect 39715 3380 39773 3381
rect 39715 3340 39724 3380
rect 39764 3340 39773 3380
rect 39715 3339 39773 3340
rect 40099 3380 40157 3381
rect 40099 3340 40108 3380
rect 40148 3340 40157 3380
rect 40099 3339 40157 3340
rect 40483 3380 40541 3381
rect 40483 3340 40492 3380
rect 40532 3340 40541 3380
rect 40483 3339 40541 3340
rect 40867 3380 40925 3381
rect 40867 3340 40876 3380
rect 40916 3340 40925 3380
rect 40867 3339 40925 3340
rect 41251 3380 41309 3381
rect 41251 3340 41260 3380
rect 41300 3340 41309 3380
rect 41251 3339 41309 3340
rect 8611 3296 8669 3297
rect 8611 3256 8620 3296
rect 8660 3256 8669 3296
rect 8611 3255 8669 3256
rect 40683 3296 40725 3305
rect 40683 3256 40684 3296
rect 40724 3256 40725 3296
rect 40683 3247 40725 3256
rect 1323 3212 1365 3221
rect 1323 3172 1324 3212
rect 1364 3172 1365 3212
rect 1323 3163 1365 3172
rect 5931 3212 5973 3221
rect 5931 3172 5932 3212
rect 5972 3172 5973 3212
rect 5931 3163 5973 3172
rect 6219 3212 6261 3221
rect 6219 3172 6220 3212
rect 6260 3172 6261 3212
rect 6219 3163 6261 3172
rect 12843 3212 12885 3221
rect 12843 3172 12844 3212
rect 12884 3172 12885 3212
rect 12843 3163 12885 3172
rect 20139 3212 20181 3221
rect 20139 3172 20140 3212
rect 20180 3172 20181 3212
rect 20139 3163 20181 3172
rect 21963 3212 22005 3221
rect 21963 3172 21964 3212
rect 22004 3172 22005 3212
rect 21963 3163 22005 3172
rect 22923 3212 22965 3221
rect 22923 3172 22924 3212
rect 22964 3172 22965 3212
rect 22923 3163 22965 3172
rect 25035 3212 25077 3221
rect 25035 3172 25036 3212
rect 25076 3172 25077 3212
rect 25035 3163 25077 3172
rect 27435 3212 27477 3221
rect 27435 3172 27436 3212
rect 27476 3172 27477 3212
rect 27435 3163 27477 3172
rect 36267 3212 36309 3221
rect 36267 3172 36268 3212
rect 36308 3172 36309 3212
rect 36267 3163 36309 3172
rect 36939 3212 36981 3221
rect 36939 3172 36940 3212
rect 36980 3172 36981 3212
rect 36939 3163 36981 3172
rect 39531 3212 39573 3221
rect 39531 3172 39532 3212
rect 39572 3172 39573 3212
rect 39531 3163 39573 3172
rect 39915 3212 39957 3221
rect 39915 3172 39916 3212
rect 39956 3172 39957 3212
rect 39915 3163 39957 3172
rect 40299 3212 40341 3221
rect 40299 3172 40300 3212
rect 40340 3172 40341 3212
rect 40299 3163 40341 3172
rect 41451 3212 41493 3221
rect 41451 3172 41452 3212
rect 41492 3172 41493 3212
rect 41451 3163 41493 3172
rect 1152 3044 41856 3068
rect 1152 3004 3688 3044
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 4056 3004 18808 3044
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 19176 3004 33928 3044
rect 33968 3004 34010 3044
rect 34050 3004 34092 3044
rect 34132 3004 34174 3044
rect 34214 3004 34256 3044
rect 34296 3004 41856 3044
rect 1152 2980 41856 3004
rect 5067 2876 5109 2885
rect 5067 2836 5068 2876
rect 5108 2836 5109 2876
rect 5067 2827 5109 2836
rect 15051 2876 15093 2885
rect 15051 2836 15052 2876
rect 15092 2836 15093 2876
rect 15051 2827 15093 2836
rect 28107 2876 28149 2885
rect 28107 2836 28108 2876
rect 28148 2836 28149 2876
rect 28107 2827 28149 2836
rect 29739 2876 29781 2885
rect 29739 2836 29740 2876
rect 29780 2836 29781 2876
rect 29739 2827 29781 2836
rect 31371 2876 31413 2885
rect 31371 2836 31372 2876
rect 31412 2836 31413 2876
rect 31371 2827 31413 2836
rect 37995 2876 38037 2885
rect 37995 2836 37996 2876
rect 38036 2836 38037 2876
rect 37995 2827 38037 2836
rect 14571 2792 14613 2801
rect 14571 2752 14572 2792
rect 14612 2752 14613 2792
rect 14571 2743 14613 2752
rect 25707 2792 25749 2801
rect 25707 2752 25708 2792
rect 25748 2752 25749 2792
rect 25707 2743 25749 2752
rect 36363 2792 36405 2801
rect 36363 2752 36364 2792
rect 36404 2752 36405 2792
rect 36363 2743 36405 2752
rect 41643 2792 41685 2801
rect 41643 2752 41644 2792
rect 41684 2752 41685 2792
rect 41643 2743 41685 2752
rect 11019 2708 11061 2717
rect 11019 2668 11020 2708
rect 11060 2668 11061 2708
rect 11019 2659 11061 2668
rect 15523 2708 15581 2709
rect 15523 2668 15532 2708
rect 15572 2668 15581 2708
rect 15523 2667 15581 2668
rect 15907 2708 15965 2709
rect 15907 2668 15916 2708
rect 15956 2668 15965 2708
rect 15907 2667 15965 2668
rect 22443 2708 22485 2717
rect 22443 2668 22444 2708
rect 22484 2668 22485 2708
rect 22443 2659 22485 2668
rect 22539 2708 22581 2717
rect 22539 2668 22540 2708
rect 22580 2668 22581 2708
rect 22539 2659 22581 2668
rect 24067 2708 24125 2709
rect 24067 2668 24076 2708
rect 24116 2668 24125 2708
rect 41443 2708 41501 2709
rect 24067 2667 24125 2668
rect 26763 2666 26805 2675
rect 41443 2668 41452 2708
rect 41492 2668 41501 2708
rect 41443 2667 41501 2668
rect 12075 2638 12117 2647
rect 1323 2624 1365 2633
rect 1323 2584 1324 2624
rect 1364 2584 1365 2624
rect 1323 2575 1365 2584
rect 1419 2624 1461 2633
rect 1419 2584 1420 2624
rect 1460 2584 1461 2624
rect 1419 2575 1461 2584
rect 1515 2624 1557 2633
rect 1515 2584 1516 2624
rect 1556 2584 1557 2624
rect 1515 2575 1557 2584
rect 1611 2624 1653 2633
rect 1611 2584 1612 2624
rect 1652 2584 1653 2624
rect 1611 2575 1653 2584
rect 1795 2624 1853 2625
rect 1795 2584 1804 2624
rect 1844 2584 1853 2624
rect 1795 2583 1853 2584
rect 3043 2624 3101 2625
rect 3043 2584 3052 2624
rect 3092 2584 3101 2624
rect 3043 2583 3101 2584
rect 3427 2624 3485 2625
rect 3427 2584 3436 2624
rect 3476 2584 3485 2624
rect 3427 2583 3485 2584
rect 4675 2624 4733 2625
rect 4675 2584 4684 2624
rect 4724 2584 4733 2624
rect 4675 2583 4733 2584
rect 5059 2624 5117 2625
rect 5059 2584 5068 2624
rect 5108 2584 5117 2624
rect 5059 2583 5117 2584
rect 5259 2624 5301 2633
rect 5259 2584 5260 2624
rect 5300 2584 5301 2624
rect 5259 2575 5301 2584
rect 5347 2624 5405 2625
rect 5347 2584 5356 2624
rect 5396 2584 5405 2624
rect 5347 2583 5405 2584
rect 5539 2624 5597 2625
rect 5539 2584 5548 2624
rect 5588 2584 5597 2624
rect 5539 2583 5597 2584
rect 6787 2624 6845 2625
rect 6787 2584 6796 2624
rect 6836 2584 6845 2624
rect 6787 2583 6845 2584
rect 7171 2624 7229 2625
rect 7171 2584 7180 2624
rect 7220 2584 7229 2624
rect 7171 2583 7229 2584
rect 8419 2624 8477 2625
rect 8419 2584 8428 2624
rect 8468 2584 8477 2624
rect 8419 2583 8477 2584
rect 8803 2624 8861 2625
rect 8803 2584 8812 2624
rect 8852 2584 8861 2624
rect 8803 2583 8861 2584
rect 10051 2624 10109 2625
rect 10051 2584 10060 2624
rect 10100 2584 10109 2624
rect 10051 2583 10109 2584
rect 10539 2624 10581 2633
rect 10539 2584 10540 2624
rect 10580 2584 10581 2624
rect 10539 2575 10581 2584
rect 10635 2624 10677 2633
rect 10635 2584 10636 2624
rect 10676 2584 10677 2624
rect 10635 2575 10677 2584
rect 11115 2624 11157 2633
rect 11115 2584 11116 2624
rect 11156 2584 11157 2624
rect 11115 2575 11157 2584
rect 11587 2624 11645 2625
rect 11587 2584 11596 2624
rect 11636 2584 11645 2624
rect 12075 2598 12076 2638
rect 12116 2598 12117 2638
rect 23547 2633 23589 2642
rect 12075 2589 12117 2598
rect 12451 2624 12509 2625
rect 11587 2583 11645 2584
rect 12451 2584 12460 2624
rect 12500 2584 12509 2624
rect 12451 2583 12509 2584
rect 13699 2624 13757 2625
rect 13699 2584 13708 2624
rect 13748 2584 13757 2624
rect 13699 2583 13757 2584
rect 14187 2624 14229 2633
rect 14187 2584 14188 2624
rect 14228 2584 14229 2624
rect 14187 2575 14229 2584
rect 14283 2624 14325 2633
rect 14283 2584 14284 2624
rect 14324 2584 14325 2624
rect 14283 2575 14325 2584
rect 14379 2624 14421 2633
rect 14379 2584 14380 2624
rect 14420 2584 14421 2624
rect 14379 2575 14421 2584
rect 14571 2624 14613 2633
rect 14571 2584 14572 2624
rect 14612 2584 14613 2624
rect 14571 2575 14613 2584
rect 14859 2624 14901 2633
rect 14859 2584 14860 2624
rect 14900 2584 14901 2624
rect 14859 2575 14901 2584
rect 15051 2624 15093 2633
rect 15051 2584 15052 2624
rect 15092 2584 15093 2624
rect 15051 2575 15093 2584
rect 15243 2624 15285 2633
rect 15243 2584 15244 2624
rect 15284 2584 15285 2624
rect 15243 2575 15285 2584
rect 15331 2624 15389 2625
rect 15331 2584 15340 2624
rect 15380 2584 15389 2624
rect 15331 2583 15389 2584
rect 20035 2624 20093 2625
rect 20035 2584 20044 2624
rect 20084 2584 20093 2624
rect 20035 2583 20093 2584
rect 21283 2624 21341 2625
rect 21283 2584 21292 2624
rect 21332 2584 21341 2624
rect 21283 2583 21341 2584
rect 21963 2624 22005 2633
rect 21963 2584 21964 2624
rect 22004 2584 22005 2624
rect 21963 2575 22005 2584
rect 22059 2624 22101 2633
rect 22059 2584 22060 2624
rect 22100 2584 22101 2624
rect 22059 2575 22101 2584
rect 23011 2624 23069 2625
rect 23011 2584 23020 2624
rect 23060 2584 23069 2624
rect 23547 2593 23548 2633
rect 23588 2593 23589 2633
rect 23547 2584 23589 2593
rect 24259 2624 24317 2625
rect 24259 2584 24268 2624
rect 24308 2584 24317 2624
rect 23011 2583 23069 2584
rect 24259 2583 24317 2584
rect 25507 2624 25565 2625
rect 25507 2584 25516 2624
rect 25556 2584 25565 2624
rect 25507 2583 25565 2584
rect 26187 2624 26229 2633
rect 26187 2584 26188 2624
rect 26228 2584 26229 2624
rect 26187 2575 26229 2584
rect 26283 2624 26325 2633
rect 26283 2584 26284 2624
rect 26324 2584 26325 2624
rect 26283 2575 26325 2584
rect 26667 2624 26709 2633
rect 26667 2584 26668 2624
rect 26708 2584 26709 2624
rect 26763 2626 26764 2666
rect 26804 2626 26805 2666
rect 26763 2617 26805 2626
rect 27723 2633 27765 2642
rect 27235 2624 27293 2625
rect 26667 2575 26709 2584
rect 27235 2584 27244 2624
rect 27284 2584 27293 2624
rect 27723 2593 27724 2633
rect 27764 2593 27765 2633
rect 27723 2584 27765 2593
rect 28291 2624 28349 2625
rect 28291 2584 28300 2624
rect 28340 2584 28349 2624
rect 27235 2583 27293 2584
rect 28291 2583 28349 2584
rect 29539 2624 29597 2625
rect 29539 2584 29548 2624
rect 29588 2584 29597 2624
rect 29539 2583 29597 2584
rect 29923 2624 29981 2625
rect 29923 2584 29932 2624
rect 29972 2584 29981 2624
rect 29923 2583 29981 2584
rect 31171 2624 31229 2625
rect 31171 2584 31180 2624
rect 31220 2584 31229 2624
rect 31171 2583 31229 2584
rect 31555 2624 31613 2625
rect 31555 2584 31564 2624
rect 31604 2584 31613 2624
rect 31555 2583 31613 2584
rect 32803 2624 32861 2625
rect 32803 2584 32812 2624
rect 32852 2584 32861 2624
rect 32803 2583 32861 2584
rect 32995 2624 33053 2625
rect 32995 2584 33004 2624
rect 33044 2584 33053 2624
rect 32995 2583 33053 2584
rect 34243 2624 34301 2625
rect 34243 2584 34252 2624
rect 34292 2584 34301 2624
rect 34243 2583 34301 2584
rect 34915 2624 34973 2625
rect 34915 2584 34924 2624
rect 34964 2584 34973 2624
rect 34915 2583 34973 2584
rect 36163 2624 36221 2625
rect 36163 2584 36172 2624
rect 36212 2584 36221 2624
rect 36163 2583 36221 2584
rect 36547 2624 36605 2625
rect 36547 2584 36556 2624
rect 36596 2584 36605 2624
rect 36547 2583 36605 2584
rect 37795 2624 37853 2625
rect 37795 2584 37804 2624
rect 37844 2584 37853 2624
rect 37795 2583 37853 2584
rect 38371 2624 38429 2625
rect 38371 2584 38380 2624
rect 38420 2584 38429 2624
rect 38371 2583 38429 2584
rect 39619 2624 39677 2625
rect 39619 2584 39628 2624
rect 39668 2584 39677 2624
rect 39619 2583 39677 2584
rect 40003 2624 40061 2625
rect 40003 2584 40012 2624
rect 40052 2584 40061 2624
rect 40003 2583 40061 2584
rect 41251 2624 41309 2625
rect 41251 2584 41260 2624
rect 41300 2584 41309 2624
rect 41251 2583 41309 2584
rect 4875 2540 4917 2549
rect 4875 2500 4876 2540
rect 4916 2500 4917 2540
rect 4875 2491 4917 2500
rect 6987 2540 7029 2549
rect 6987 2500 6988 2540
rect 7028 2500 7029 2540
rect 6987 2491 7029 2500
rect 12267 2540 12309 2549
rect 12267 2500 12268 2540
rect 12308 2500 12309 2540
rect 12267 2491 12309 2500
rect 23691 2540 23733 2549
rect 23691 2500 23692 2540
rect 23732 2500 23733 2540
rect 23691 2491 23733 2500
rect 34443 2540 34485 2549
rect 34443 2500 34444 2540
rect 34484 2500 34485 2540
rect 34443 2491 34485 2500
rect 3243 2456 3285 2465
rect 3243 2416 3244 2456
rect 3284 2416 3285 2456
rect 3243 2407 3285 2416
rect 8619 2456 8661 2465
rect 8619 2416 8620 2456
rect 8660 2416 8661 2456
rect 8619 2407 8661 2416
rect 10251 2456 10293 2465
rect 10251 2416 10252 2456
rect 10292 2416 10293 2456
rect 10251 2407 10293 2416
rect 13899 2456 13941 2465
rect 13899 2416 13900 2456
rect 13940 2416 13941 2456
rect 13899 2407 13941 2416
rect 14083 2456 14141 2457
rect 14083 2416 14092 2456
rect 14132 2416 14141 2456
rect 14083 2415 14141 2416
rect 15723 2456 15765 2465
rect 15723 2416 15724 2456
rect 15764 2416 15765 2456
rect 15723 2407 15765 2416
rect 16107 2456 16149 2465
rect 16107 2416 16108 2456
rect 16148 2416 16149 2456
rect 16107 2407 16149 2416
rect 21483 2456 21525 2465
rect 21483 2416 21484 2456
rect 21524 2416 21525 2456
rect 21483 2407 21525 2416
rect 23883 2456 23925 2465
rect 23883 2416 23884 2456
rect 23924 2416 23925 2456
rect 23883 2407 23925 2416
rect 27915 2456 27957 2465
rect 27915 2416 27916 2456
rect 27956 2416 27957 2456
rect 27915 2407 27957 2416
rect 38187 2456 38229 2465
rect 38187 2416 38188 2456
rect 38228 2416 38229 2456
rect 38187 2407 38229 2416
rect 39819 2456 39861 2465
rect 39819 2416 39820 2456
rect 39860 2416 39861 2456
rect 39819 2407 39861 2416
rect 1152 2288 41856 2312
rect 1152 2248 4928 2288
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 5296 2248 20048 2288
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20416 2248 35168 2288
rect 35208 2248 35250 2288
rect 35290 2248 35332 2288
rect 35372 2248 35414 2288
rect 35454 2248 35496 2288
rect 35536 2248 41856 2288
rect 1152 2224 41856 2248
rect 3243 2120 3285 2129
rect 3243 2080 3244 2120
rect 3284 2080 3285 2120
rect 3243 2071 3285 2080
rect 7267 2120 7325 2121
rect 7267 2080 7276 2120
rect 7316 2080 7325 2120
rect 7267 2079 7325 2080
rect 10243 2120 10301 2121
rect 10243 2080 10252 2120
rect 10292 2080 10301 2120
rect 10243 2079 10301 2080
rect 13227 2120 13269 2129
rect 13227 2080 13228 2120
rect 13268 2080 13269 2120
rect 13227 2071 13269 2080
rect 15627 2120 15669 2129
rect 15627 2080 15628 2120
rect 15668 2080 15669 2120
rect 15627 2071 15669 2080
rect 25995 2120 26037 2129
rect 25995 2080 25996 2120
rect 26036 2080 26037 2120
rect 25995 2071 26037 2080
rect 26187 2120 26229 2129
rect 26187 2080 26188 2120
rect 26228 2080 26229 2120
rect 26187 2071 26229 2080
rect 33963 2120 34005 2129
rect 33963 2080 33964 2120
rect 34004 2080 34005 2120
rect 33963 2071 34005 2080
rect 36075 2120 36117 2129
rect 36075 2080 36076 2120
rect 36116 2080 36117 2120
rect 36075 2071 36117 2080
rect 38475 2120 38517 2129
rect 38475 2080 38476 2120
rect 38516 2080 38517 2120
rect 38475 2071 38517 2080
rect 41259 2120 41301 2129
rect 41259 2080 41260 2120
rect 41300 2080 41301 2120
rect 41259 2071 41301 2080
rect 41643 2120 41685 2129
rect 41643 2080 41644 2120
rect 41684 2080 41685 2120
rect 41643 2071 41685 2080
rect 4875 2036 4917 2045
rect 4875 1996 4876 2036
rect 4916 1996 4917 2036
rect 4875 1987 4917 1996
rect 6891 2036 6933 2045
rect 6891 1996 6892 2036
rect 6932 1996 6933 2036
rect 6891 1987 6933 1996
rect 9579 2036 9621 2045
rect 9579 1996 9580 2036
rect 9620 1996 9621 2036
rect 9579 1987 9621 1996
rect 12555 2036 12597 2045
rect 12555 1996 12556 2036
rect 12596 1996 12597 2036
rect 12555 1987 12597 1996
rect 12747 2036 12789 2045
rect 12747 1996 12748 2036
rect 12788 1996 12789 2036
rect 12747 1987 12789 1996
rect 17835 2036 17877 2045
rect 17835 1996 17836 2036
rect 17876 1996 17877 2036
rect 17835 1987 17877 1996
rect 19851 2036 19893 2045
rect 19851 1996 19852 2036
rect 19892 1996 19893 2036
rect 19851 1987 19893 1996
rect 23115 2036 23157 2045
rect 23115 1996 23116 2036
rect 23156 1996 23157 2036
rect 23115 1987 23157 1996
rect 30699 2036 30741 2045
rect 30699 1996 30700 2036
rect 30740 1996 30741 2036
rect 30699 1987 30741 1996
rect 40491 2036 40533 2045
rect 40491 1996 40492 2036
rect 40532 1996 40533 2036
rect 40491 1987 40533 1996
rect 12843 1973 12885 1982
rect 1323 1952 1365 1961
rect 1323 1912 1324 1952
rect 1364 1912 1365 1952
rect 1323 1903 1365 1912
rect 1419 1952 1461 1961
rect 1419 1912 1420 1952
rect 1460 1912 1461 1952
rect 1419 1903 1461 1912
rect 1515 1952 1557 1961
rect 1515 1912 1516 1952
rect 1556 1912 1557 1952
rect 1515 1903 1557 1912
rect 1611 1952 1653 1961
rect 1611 1912 1612 1952
rect 1652 1912 1653 1952
rect 1611 1903 1653 1912
rect 1795 1952 1853 1953
rect 1795 1912 1804 1952
rect 1844 1912 1853 1952
rect 1795 1911 1853 1912
rect 3043 1952 3101 1953
rect 3043 1912 3052 1952
rect 3092 1912 3101 1952
rect 3043 1911 3101 1912
rect 3427 1952 3485 1953
rect 3427 1912 3436 1952
rect 3476 1912 3485 1952
rect 3427 1911 3485 1912
rect 4675 1952 4733 1953
rect 4675 1912 4684 1952
rect 4724 1912 4733 1952
rect 4675 1911 4733 1912
rect 5163 1952 5205 1961
rect 5163 1912 5164 1952
rect 5204 1912 5205 1952
rect 5163 1903 5205 1912
rect 5259 1952 5301 1961
rect 5259 1912 5260 1952
rect 5300 1912 5301 1952
rect 5259 1903 5301 1912
rect 5739 1952 5781 1961
rect 5739 1912 5740 1952
rect 5780 1912 5781 1952
rect 5739 1903 5781 1912
rect 6211 1952 6269 1953
rect 6211 1912 6220 1952
rect 6260 1912 6269 1952
rect 7371 1952 7413 1961
rect 6211 1911 6269 1912
rect 6699 1938 6741 1947
rect 6699 1898 6700 1938
rect 6740 1898 6741 1938
rect 7371 1912 7372 1952
rect 7412 1912 7413 1952
rect 7371 1903 7413 1912
rect 7467 1952 7509 1961
rect 7467 1912 7468 1952
rect 7508 1912 7509 1952
rect 7467 1903 7509 1912
rect 7563 1952 7605 1961
rect 7563 1912 7564 1952
rect 7604 1912 7605 1952
rect 7563 1903 7605 1912
rect 7851 1952 7893 1961
rect 7851 1912 7852 1952
rect 7892 1912 7893 1952
rect 7851 1903 7893 1912
rect 7947 1952 7989 1961
rect 7947 1912 7948 1952
rect 7988 1912 7989 1952
rect 7947 1903 7989 1912
rect 8899 1952 8957 1953
rect 8899 1912 8908 1952
rect 8948 1912 8957 1952
rect 8899 1911 8957 1912
rect 9387 1947 9429 1956
rect 9387 1907 9388 1947
rect 9428 1907 9429 1947
rect 9387 1898 9429 1907
rect 9771 1952 9813 1961
rect 9771 1912 9772 1952
rect 9812 1912 9813 1952
rect 9771 1903 9813 1912
rect 9867 1952 9909 1961
rect 9867 1912 9868 1952
rect 9908 1912 9909 1952
rect 9867 1903 9909 1912
rect 9963 1952 10005 1961
rect 9963 1912 9964 1952
rect 10004 1912 10005 1952
rect 9963 1903 10005 1912
rect 10059 1952 10101 1961
rect 10059 1912 10060 1952
rect 10100 1912 10101 1952
rect 10059 1903 10101 1912
rect 10443 1952 10485 1961
rect 10443 1912 10444 1952
rect 10484 1912 10485 1952
rect 10443 1903 10485 1912
rect 10539 1952 10581 1961
rect 10539 1912 10540 1952
rect 10580 1912 10581 1952
rect 10539 1903 10581 1912
rect 10827 1952 10869 1961
rect 10827 1912 10828 1952
rect 10868 1912 10869 1952
rect 10827 1903 10869 1912
rect 10923 1952 10965 1961
rect 10923 1912 10924 1952
rect 10964 1912 10965 1952
rect 10923 1903 10965 1912
rect 11403 1952 11445 1961
rect 11403 1912 11404 1952
rect 11444 1912 11445 1952
rect 11403 1903 11445 1912
rect 11875 1952 11933 1953
rect 11875 1912 11884 1952
rect 11924 1912 11933 1952
rect 11875 1911 11933 1912
rect 12363 1938 12405 1947
rect 12363 1898 12364 1938
rect 12404 1898 12405 1938
rect 12843 1933 12844 1973
rect 12884 1933 12885 1973
rect 12843 1924 12885 1933
rect 12939 1952 12981 1961
rect 12939 1912 12940 1952
rect 12980 1912 12981 1952
rect 12939 1903 12981 1912
rect 13035 1952 13077 1961
rect 13035 1912 13036 1952
rect 13076 1912 13077 1952
rect 13035 1903 13077 1912
rect 13419 1952 13461 1961
rect 13419 1912 13420 1952
rect 13460 1912 13461 1952
rect 13419 1903 13461 1912
rect 13899 1952 13941 1961
rect 13899 1912 13900 1952
rect 13940 1912 13941 1952
rect 13899 1903 13941 1912
rect 13995 1952 14037 1961
rect 13995 1912 13996 1952
rect 14036 1912 14037 1952
rect 13995 1903 14037 1912
rect 14475 1952 14517 1961
rect 14475 1912 14476 1952
rect 14516 1912 14517 1952
rect 14475 1903 14517 1912
rect 14947 1952 15005 1953
rect 14947 1912 14956 1952
rect 14996 1912 15005 1952
rect 16387 1952 16445 1953
rect 14947 1911 15005 1912
rect 15435 1938 15477 1947
rect 6699 1889 6741 1898
rect 12363 1889 12405 1898
rect 15435 1898 15436 1938
rect 15476 1898 15477 1938
rect 16387 1912 16396 1952
rect 16436 1912 16445 1952
rect 16387 1911 16445 1912
rect 17635 1952 17693 1953
rect 17635 1912 17644 1952
rect 17684 1912 17693 1952
rect 17635 1911 17693 1912
rect 18123 1952 18165 1961
rect 18123 1912 18124 1952
rect 18164 1912 18165 1952
rect 18123 1903 18165 1912
rect 18219 1952 18261 1961
rect 18219 1912 18220 1952
rect 18260 1912 18261 1952
rect 18219 1903 18261 1912
rect 18603 1952 18645 1961
rect 18603 1912 18604 1952
rect 18644 1912 18645 1952
rect 18603 1903 18645 1912
rect 19171 1952 19229 1953
rect 19171 1912 19180 1952
rect 19220 1912 19229 1952
rect 21387 1952 21429 1961
rect 19171 1911 19229 1912
rect 19659 1938 19701 1947
rect 15435 1889 15477 1898
rect 19659 1898 19660 1938
rect 19700 1898 19701 1938
rect 21387 1912 21388 1952
rect 21428 1912 21429 1952
rect 21387 1903 21429 1912
rect 21483 1952 21525 1961
rect 21483 1912 21484 1952
rect 21524 1912 21525 1952
rect 21483 1903 21525 1912
rect 21867 1952 21909 1961
rect 21867 1912 21868 1952
rect 21908 1912 21909 1952
rect 21867 1903 21909 1912
rect 21963 1952 22005 1961
rect 21963 1912 21964 1952
rect 22004 1912 22005 1952
rect 21963 1903 22005 1912
rect 22435 1952 22493 1953
rect 22435 1912 22444 1952
rect 22484 1912 22493 1952
rect 24267 1952 24309 1961
rect 22435 1911 22493 1912
rect 22971 1910 23013 1919
rect 19659 1889 19701 1898
rect 5643 1868 5685 1877
rect 5643 1828 5644 1868
rect 5684 1828 5685 1868
rect 5643 1819 5685 1828
rect 8331 1868 8373 1877
rect 8331 1828 8332 1868
rect 8372 1828 8373 1868
rect 8331 1819 8373 1828
rect 8427 1868 8469 1877
rect 8427 1828 8428 1868
rect 8468 1828 8469 1868
rect 8427 1819 8469 1828
rect 11307 1868 11349 1877
rect 11307 1828 11308 1868
rect 11348 1828 11349 1868
rect 11307 1819 11349 1828
rect 14379 1868 14421 1877
rect 14379 1828 14380 1868
rect 14420 1828 14421 1868
rect 14379 1819 14421 1828
rect 15811 1868 15869 1869
rect 15811 1828 15820 1868
rect 15860 1828 15869 1868
rect 15811 1827 15869 1828
rect 18699 1868 18741 1877
rect 22971 1870 22972 1910
rect 23012 1870 23013 1910
rect 24267 1912 24268 1952
rect 24308 1912 24309 1952
rect 24267 1903 24309 1912
rect 24363 1952 24405 1961
rect 24363 1912 24364 1952
rect 24404 1912 24405 1952
rect 24363 1903 24405 1912
rect 24747 1952 24789 1961
rect 24747 1912 24748 1952
rect 24788 1912 24789 1952
rect 24747 1903 24789 1912
rect 25315 1952 25373 1953
rect 25315 1912 25324 1952
rect 25364 1912 25373 1952
rect 26371 1952 26429 1953
rect 25315 1911 25373 1912
rect 25803 1938 25845 1947
rect 25803 1898 25804 1938
rect 25844 1898 25845 1938
rect 26371 1912 26380 1952
rect 26420 1912 26429 1952
rect 26371 1911 26429 1912
rect 27619 1952 27677 1953
rect 27619 1912 27628 1952
rect 27668 1912 27677 1952
rect 27619 1911 27677 1912
rect 28971 1952 29013 1961
rect 28971 1912 28972 1952
rect 29012 1912 29013 1952
rect 28971 1903 29013 1912
rect 29067 1952 29109 1961
rect 29067 1912 29068 1952
rect 29108 1912 29109 1952
rect 29067 1903 29109 1912
rect 30019 1952 30077 1953
rect 30019 1912 30028 1952
rect 30068 1912 30077 1952
rect 32235 1952 32277 1961
rect 30019 1911 30077 1912
rect 30507 1938 30549 1947
rect 25803 1889 25845 1898
rect 30507 1898 30508 1938
rect 30548 1898 30549 1938
rect 32235 1912 32236 1952
rect 32276 1912 32277 1952
rect 32235 1903 32277 1912
rect 32331 1952 32373 1961
rect 32331 1912 32332 1952
rect 32372 1912 32373 1952
rect 32331 1903 32373 1912
rect 32715 1952 32757 1961
rect 32715 1912 32716 1952
rect 32756 1912 32757 1952
rect 32715 1903 32757 1912
rect 32811 1952 32853 1961
rect 32811 1912 32812 1952
rect 32852 1912 32853 1952
rect 32811 1903 32853 1912
rect 33283 1952 33341 1953
rect 33283 1912 33292 1952
rect 33332 1912 33341 1952
rect 33283 1911 33341 1912
rect 33771 1947 33813 1956
rect 33771 1907 33772 1947
rect 33812 1907 33813 1947
rect 33771 1898 33813 1907
rect 34347 1952 34389 1961
rect 34347 1912 34348 1952
rect 34388 1912 34389 1952
rect 34347 1903 34389 1912
rect 34443 1952 34485 1961
rect 34443 1912 34444 1952
rect 34484 1912 34485 1952
rect 34443 1903 34485 1912
rect 34923 1952 34965 1961
rect 34923 1912 34924 1952
rect 34964 1912 34965 1952
rect 34923 1903 34965 1912
rect 35395 1952 35453 1953
rect 35395 1912 35404 1952
rect 35444 1912 35453 1952
rect 36747 1952 36789 1961
rect 35395 1911 35453 1912
rect 35883 1938 35925 1947
rect 35883 1898 35884 1938
rect 35924 1898 35925 1938
rect 36747 1912 36748 1952
rect 36788 1912 36789 1952
rect 36747 1903 36789 1912
rect 36843 1952 36885 1961
rect 36843 1912 36844 1952
rect 36884 1912 36885 1952
rect 36843 1903 36885 1912
rect 37227 1952 37269 1961
rect 37227 1912 37228 1952
rect 37268 1912 37269 1952
rect 37227 1903 37269 1912
rect 37323 1952 37365 1961
rect 37323 1912 37324 1952
rect 37364 1912 37365 1952
rect 37323 1903 37365 1912
rect 37795 1952 37853 1953
rect 37795 1912 37804 1952
rect 37844 1912 37853 1952
rect 37795 1911 37853 1912
rect 38283 1947 38325 1956
rect 38283 1907 38284 1947
rect 38324 1907 38325 1947
rect 38283 1898 38325 1907
rect 38763 1952 38805 1961
rect 38763 1912 38764 1952
rect 38804 1912 38805 1952
rect 38763 1903 38805 1912
rect 38859 1952 38901 1961
rect 38859 1912 38860 1952
rect 38900 1912 38901 1952
rect 38859 1903 38901 1912
rect 39339 1952 39381 1961
rect 39339 1912 39340 1952
rect 39380 1912 39381 1952
rect 39339 1903 39381 1912
rect 39811 1952 39869 1953
rect 39811 1912 39820 1952
rect 39860 1912 39869 1952
rect 39811 1911 39869 1912
rect 40299 1947 40341 1956
rect 40299 1907 40300 1947
rect 40340 1907 40341 1947
rect 40299 1898 40341 1907
rect 30507 1889 30549 1898
rect 35883 1889 35925 1898
rect 18699 1828 18700 1868
rect 18740 1828 18741 1868
rect 18699 1819 18741 1828
rect 20899 1868 20957 1869
rect 20899 1828 20908 1868
rect 20948 1828 20957 1868
rect 22971 1861 23013 1870
rect 23299 1868 23357 1869
rect 20899 1827 20957 1828
rect 23299 1828 23308 1868
rect 23348 1828 23357 1868
rect 23299 1827 23357 1828
rect 23875 1868 23933 1869
rect 23875 1828 23884 1868
rect 23924 1828 23933 1868
rect 23875 1827 23933 1828
rect 24843 1868 24885 1877
rect 24843 1828 24844 1868
rect 24884 1828 24885 1868
rect 24843 1819 24885 1828
rect 28003 1868 28061 1869
rect 28003 1828 28012 1868
rect 28052 1828 28061 1868
rect 28003 1827 28061 1828
rect 28387 1868 28445 1869
rect 28387 1828 28396 1868
rect 28436 1828 28445 1868
rect 28387 1827 28445 1828
rect 29451 1868 29493 1877
rect 29451 1828 29452 1868
rect 29492 1828 29493 1868
rect 29451 1819 29493 1828
rect 29547 1868 29589 1877
rect 29547 1828 29548 1868
rect 29588 1828 29589 1868
rect 29547 1819 29589 1828
rect 31075 1868 31133 1869
rect 31075 1828 31084 1868
rect 31124 1828 31133 1868
rect 31075 1827 31133 1828
rect 31459 1868 31517 1869
rect 31459 1828 31468 1868
rect 31508 1828 31517 1868
rect 31459 1827 31517 1828
rect 31939 1868 31997 1869
rect 31939 1828 31948 1868
rect 31988 1828 31997 1868
rect 31939 1827 31997 1828
rect 34827 1868 34869 1877
rect 34827 1828 34828 1868
rect 34868 1828 34869 1868
rect 34827 1819 34869 1828
rect 36451 1868 36509 1869
rect 36451 1828 36460 1868
rect 36500 1828 36509 1868
rect 36451 1827 36509 1828
rect 39243 1868 39285 1877
rect 39243 1828 39244 1868
rect 39284 1828 39285 1868
rect 39243 1819 39285 1828
rect 40867 1868 40925 1869
rect 40867 1828 40876 1868
rect 40916 1828 40925 1868
rect 40867 1827 40925 1828
rect 41059 1868 41117 1869
rect 41059 1828 41068 1868
rect 41108 1828 41117 1868
rect 41059 1827 41117 1828
rect 41443 1868 41501 1869
rect 41443 1828 41452 1868
rect 41492 1828 41501 1868
rect 41443 1827 41501 1828
rect 13419 1784 13461 1793
rect 13419 1744 13420 1784
rect 13460 1744 13461 1784
rect 13419 1735 13461 1744
rect 16011 1700 16053 1709
rect 16011 1660 16012 1700
rect 16052 1660 16053 1700
rect 16011 1651 16053 1660
rect 21099 1700 21141 1709
rect 21099 1660 21100 1700
rect 21140 1660 21141 1700
rect 21099 1651 21141 1660
rect 23499 1700 23541 1709
rect 23499 1660 23500 1700
rect 23540 1660 23541 1700
rect 23499 1651 23541 1660
rect 23691 1700 23733 1709
rect 23691 1660 23692 1700
rect 23732 1660 23733 1700
rect 23691 1651 23733 1660
rect 27819 1700 27861 1709
rect 27819 1660 27820 1700
rect 27860 1660 27861 1700
rect 27819 1651 27861 1660
rect 28203 1700 28245 1709
rect 28203 1660 28204 1700
rect 28244 1660 28245 1700
rect 28203 1651 28245 1660
rect 30891 1700 30933 1709
rect 30891 1660 30892 1700
rect 30932 1660 30933 1700
rect 30891 1651 30933 1660
rect 31275 1700 31317 1709
rect 31275 1660 31276 1700
rect 31316 1660 31317 1700
rect 31275 1651 31317 1660
rect 31755 1700 31797 1709
rect 31755 1660 31756 1700
rect 31796 1660 31797 1700
rect 31755 1651 31797 1660
rect 36267 1700 36309 1709
rect 36267 1660 36268 1700
rect 36308 1660 36309 1700
rect 36267 1651 36309 1660
rect 40683 1700 40725 1709
rect 40683 1660 40684 1700
rect 40724 1660 40725 1700
rect 40683 1651 40725 1660
rect 1152 1532 41856 1556
rect 1152 1492 3688 1532
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 4056 1492 18808 1532
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 19176 1492 33928 1532
rect 33968 1492 34010 1532
rect 34050 1492 34092 1532
rect 34132 1492 34174 1532
rect 34214 1492 34256 1532
rect 34296 1492 41856 1532
rect 1152 1468 41856 1492
rect 19563 1364 19605 1373
rect 19563 1324 19564 1364
rect 19604 1324 19605 1364
rect 19563 1315 19605 1324
rect 22155 1364 22197 1373
rect 22155 1324 22156 1364
rect 22196 1324 22197 1364
rect 22155 1315 22197 1324
rect 23979 1364 24021 1373
rect 23979 1324 23980 1364
rect 24020 1324 24021 1364
rect 23979 1315 24021 1324
rect 25611 1364 25653 1373
rect 25611 1324 25612 1364
rect 25652 1324 25653 1364
rect 25611 1315 25653 1324
rect 30507 1364 30549 1373
rect 30507 1324 30508 1364
rect 30548 1324 30549 1364
rect 30507 1315 30549 1324
rect 32139 1364 32181 1373
rect 32139 1324 32140 1364
rect 32180 1324 32181 1364
rect 32139 1315 32181 1324
rect 35403 1364 35445 1373
rect 35403 1324 35404 1364
rect 35444 1324 35445 1364
rect 35403 1315 35445 1324
rect 37035 1364 37077 1373
rect 37035 1324 37036 1364
rect 37076 1324 37077 1364
rect 37035 1315 37077 1324
rect 38667 1364 38709 1373
rect 38667 1324 38668 1364
rect 38708 1324 38709 1364
rect 38667 1315 38709 1324
rect 1611 1280 1653 1289
rect 1611 1240 1612 1280
rect 1652 1240 1653 1280
rect 1611 1231 1653 1240
rect 4003 1280 4061 1281
rect 4003 1240 4012 1280
rect 4052 1240 4061 1280
rect 4003 1239 4061 1240
rect 7747 1280 7805 1281
rect 7747 1240 7756 1280
rect 7796 1240 7805 1280
rect 7747 1239 7805 1240
rect 14859 1280 14901 1289
rect 14859 1240 14860 1280
rect 14900 1240 14901 1280
rect 14859 1231 14901 1240
rect 27243 1280 27285 1289
rect 27243 1240 27244 1280
rect 27284 1240 27285 1280
rect 27243 1231 27285 1240
rect 28875 1280 28917 1289
rect 28875 1240 28876 1280
rect 28916 1240 28917 1280
rect 28875 1231 28917 1240
rect 33771 1280 33813 1289
rect 33771 1240 33772 1280
rect 33812 1240 33813 1280
rect 33771 1231 33813 1240
rect 41067 1280 41109 1289
rect 41067 1240 41068 1280
rect 41108 1240 41109 1280
rect 41067 1231 41109 1240
rect 5547 1196 5589 1205
rect 5547 1156 5548 1196
rect 5588 1156 5589 1196
rect 5547 1147 5589 1156
rect 10251 1196 10293 1205
rect 10251 1156 10252 1196
rect 10292 1156 10293 1196
rect 10251 1147 10293 1156
rect 15523 1196 15581 1197
rect 15523 1156 15532 1196
rect 15572 1156 15581 1196
rect 15523 1155 15581 1156
rect 40483 1196 40541 1197
rect 40483 1156 40492 1196
rect 40532 1156 40541 1196
rect 40483 1155 40541 1156
rect 40867 1196 40925 1197
rect 40867 1156 40876 1196
rect 40916 1156 40925 1196
rect 40867 1155 40925 1156
rect 41251 1196 41309 1197
rect 41251 1156 41260 1196
rect 41300 1156 41309 1196
rect 41251 1155 41309 1156
rect 11211 1126 11253 1135
rect 1315 1112 1373 1113
rect 1315 1072 1324 1112
rect 1364 1072 1373 1112
rect 1315 1071 1373 1072
rect 1419 1112 1461 1121
rect 1419 1072 1420 1112
rect 1460 1072 1461 1112
rect 1419 1063 1461 1072
rect 1611 1112 1653 1121
rect 1611 1072 1612 1112
rect 1652 1072 1653 1112
rect 1611 1063 1653 1072
rect 1795 1112 1853 1113
rect 1795 1072 1804 1112
rect 1844 1072 1853 1112
rect 1795 1071 1853 1072
rect 3043 1112 3101 1113
rect 3043 1072 3052 1112
rect 3092 1072 3101 1112
rect 3043 1071 3101 1072
rect 3523 1112 3581 1113
rect 3523 1072 3532 1112
rect 3572 1072 3581 1112
rect 3523 1071 3581 1072
rect 3723 1112 3765 1121
rect 3723 1072 3724 1112
rect 3764 1072 3765 1112
rect 3723 1063 3765 1072
rect 3811 1112 3869 1113
rect 3811 1072 3820 1112
rect 3860 1072 3869 1112
rect 3811 1071 3869 1072
rect 4299 1112 4341 1121
rect 4299 1072 4300 1112
rect 4340 1072 4341 1112
rect 4299 1063 4341 1072
rect 4395 1112 4437 1121
rect 4395 1072 4396 1112
rect 4436 1072 4437 1112
rect 4395 1063 4437 1072
rect 4675 1112 4733 1113
rect 4675 1072 4684 1112
rect 4724 1072 4733 1112
rect 4675 1071 4733 1072
rect 5067 1112 5109 1121
rect 5067 1072 5068 1112
rect 5108 1072 5109 1112
rect 5067 1063 5109 1072
rect 5163 1112 5205 1121
rect 5163 1072 5164 1112
rect 5204 1072 5205 1112
rect 5163 1063 5205 1072
rect 5643 1112 5685 1121
rect 6603 1117 6645 1126
rect 5643 1072 5644 1112
rect 5684 1072 5685 1112
rect 5643 1063 5685 1072
rect 6115 1112 6173 1113
rect 6115 1072 6124 1112
rect 6164 1072 6173 1112
rect 6115 1071 6173 1072
rect 6603 1077 6604 1117
rect 6644 1077 6645 1117
rect 6603 1068 6645 1077
rect 7075 1112 7133 1113
rect 7075 1072 7084 1112
rect 7124 1072 7133 1112
rect 7075 1071 7133 1072
rect 7371 1112 7413 1121
rect 7371 1072 7372 1112
rect 7412 1072 7413 1112
rect 7371 1063 7413 1072
rect 7939 1112 7997 1113
rect 7939 1072 7948 1112
rect 7988 1072 7997 1112
rect 7939 1071 7997 1072
rect 9187 1112 9245 1113
rect 9187 1072 9196 1112
rect 9236 1072 9245 1112
rect 9187 1071 9245 1072
rect 9675 1112 9717 1121
rect 9675 1072 9676 1112
rect 9716 1072 9717 1112
rect 9675 1063 9717 1072
rect 9771 1112 9813 1121
rect 9771 1072 9772 1112
rect 9812 1072 9813 1112
rect 9771 1063 9813 1072
rect 10155 1112 10197 1121
rect 10155 1072 10156 1112
rect 10196 1072 10197 1112
rect 10155 1063 10197 1072
rect 10723 1112 10781 1113
rect 10723 1072 10732 1112
rect 10772 1072 10781 1112
rect 11211 1086 11212 1126
rect 11252 1086 11253 1126
rect 11211 1077 11253 1086
rect 11587 1112 11645 1113
rect 10723 1071 10781 1072
rect 11587 1072 11596 1112
rect 11636 1072 11645 1112
rect 11587 1071 11645 1072
rect 12835 1112 12893 1113
rect 12835 1072 12844 1112
rect 12884 1072 12893 1112
rect 12835 1071 12893 1072
rect 14659 1112 14717 1113
rect 14659 1072 14668 1112
rect 14708 1072 14717 1112
rect 14659 1071 14717 1072
rect 15051 1112 15093 1121
rect 15051 1072 15052 1112
rect 15092 1072 15093 1112
rect 13411 1070 13469 1071
rect 7467 1028 7509 1037
rect 7467 988 7468 1028
rect 7508 988 7509 1028
rect 7467 979 7509 988
rect 9387 1028 9429 1037
rect 9387 988 9388 1028
rect 9428 988 9429 1028
rect 9387 979 9429 988
rect 11403 1028 11445 1037
rect 11403 988 11404 1028
rect 11444 988 11445 1028
rect 11403 979 11445 988
rect 13035 1028 13077 1037
rect 13411 1030 13420 1070
rect 13460 1030 13469 1070
rect 15051 1063 15093 1072
rect 15147 1112 15189 1121
rect 15147 1072 15148 1112
rect 15188 1072 15189 1112
rect 15147 1063 15189 1072
rect 18115 1112 18173 1113
rect 18115 1072 18124 1112
rect 18164 1072 18173 1112
rect 18115 1071 18173 1072
rect 19363 1112 19421 1113
rect 19363 1072 19372 1112
rect 19412 1072 19421 1112
rect 19363 1071 19421 1072
rect 20707 1112 20765 1113
rect 20707 1072 20716 1112
rect 20756 1072 20765 1112
rect 20707 1071 20765 1072
rect 21955 1112 22013 1113
rect 21955 1072 21964 1112
rect 22004 1072 22013 1112
rect 21955 1071 22013 1072
rect 22339 1112 22397 1113
rect 22339 1072 22348 1112
rect 22388 1072 22397 1112
rect 22339 1071 22397 1072
rect 23587 1112 23645 1113
rect 23587 1072 23596 1112
rect 23636 1072 23645 1112
rect 23587 1071 23645 1072
rect 24163 1112 24221 1113
rect 24163 1072 24172 1112
rect 24212 1072 24221 1112
rect 24163 1071 24221 1072
rect 25795 1112 25853 1113
rect 25795 1072 25804 1112
rect 25844 1072 25853 1112
rect 25795 1071 25853 1072
rect 27043 1112 27101 1113
rect 27043 1072 27052 1112
rect 27092 1072 27101 1112
rect 27043 1071 27101 1072
rect 27427 1112 27485 1113
rect 27427 1072 27436 1112
rect 27476 1072 27485 1112
rect 27427 1071 27485 1072
rect 28675 1112 28733 1113
rect 28675 1072 28684 1112
rect 28724 1072 28733 1112
rect 28675 1071 28733 1072
rect 29059 1112 29117 1113
rect 29059 1072 29068 1112
rect 29108 1072 29117 1112
rect 29059 1071 29117 1072
rect 30307 1112 30365 1113
rect 30307 1072 30316 1112
rect 30356 1072 30365 1112
rect 30307 1071 30365 1072
rect 30691 1112 30749 1113
rect 30691 1072 30700 1112
rect 30740 1072 30749 1112
rect 30691 1071 30749 1072
rect 31939 1112 31997 1113
rect 31939 1072 31948 1112
rect 31988 1072 31997 1112
rect 31939 1071 31997 1072
rect 32323 1112 32381 1113
rect 32323 1072 32332 1112
rect 32372 1072 32381 1112
rect 32323 1071 32381 1072
rect 33571 1112 33629 1113
rect 33571 1072 33580 1112
rect 33620 1072 33629 1112
rect 33571 1071 33629 1072
rect 33955 1112 34013 1113
rect 33955 1072 33964 1112
rect 34004 1072 34013 1112
rect 33955 1071 34013 1072
rect 35203 1112 35261 1113
rect 35203 1072 35212 1112
rect 35252 1072 35261 1112
rect 35203 1071 35261 1072
rect 35587 1112 35645 1113
rect 35587 1072 35596 1112
rect 35636 1072 35645 1112
rect 35587 1071 35645 1072
rect 36835 1112 36893 1113
rect 36835 1072 36844 1112
rect 36884 1072 36893 1112
rect 36835 1071 36893 1072
rect 37219 1112 37277 1113
rect 37219 1072 37228 1112
rect 37268 1072 37277 1112
rect 37219 1071 37277 1072
rect 38467 1112 38525 1113
rect 38467 1072 38476 1112
rect 38516 1072 38525 1112
rect 38467 1071 38525 1072
rect 38851 1112 38909 1113
rect 38851 1072 38860 1112
rect 38900 1072 38909 1112
rect 38851 1071 38909 1072
rect 40099 1112 40157 1113
rect 40099 1072 40108 1112
rect 40148 1072 40157 1112
rect 40099 1071 40157 1072
rect 25411 1070 25469 1071
rect 13411 1029 13469 1030
rect 13035 988 13036 1028
rect 13076 988 13077 1028
rect 13035 979 13077 988
rect 23787 1028 23829 1037
rect 25411 1030 25420 1070
rect 25460 1030 25469 1070
rect 25411 1029 25469 1030
rect 23787 988 23788 1028
rect 23828 988 23829 1028
rect 23787 979 23829 988
rect 3243 944 3285 953
rect 3243 904 3244 944
rect 3284 904 3285 944
rect 3243 895 3285 904
rect 3531 944 3573 953
rect 3531 904 3532 944
rect 3572 904 3573 944
rect 3531 895 3573 904
rect 6795 944 6837 953
rect 6795 904 6796 944
rect 6836 904 6837 944
rect 6795 895 6837 904
rect 15331 944 15389 945
rect 15331 904 15340 944
rect 15380 904 15389 944
rect 15331 903 15389 904
rect 15723 944 15765 953
rect 15723 904 15724 944
rect 15764 904 15765 944
rect 15723 895 15765 904
rect 40299 944 40341 953
rect 40299 904 40300 944
rect 40340 904 40341 944
rect 40299 895 40341 904
rect 41451 944 41493 953
rect 41451 904 41452 944
rect 41492 904 41493 944
rect 41451 895 41493 904
rect 1152 776 41856 800
rect 1152 736 4928 776
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 5296 736 20048 776
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20416 736 35168 776
rect 35208 736 35250 776
rect 35290 736 35332 776
rect 35372 736 35414 776
rect 35454 736 35496 776
rect 35536 736 41856 776
rect 1152 712 41856 736
<< via1 >>
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 35168 9808 35208 9848
rect 35250 9808 35290 9848
rect 35332 9808 35372 9848
rect 35414 9808 35454 9848
rect 35496 9808 35536 9848
rect 1420 9640 1460 9680
rect 2188 9640 2228 9680
rect 7468 9640 7508 9680
rect 9388 9640 9428 9680
rect 32236 9640 32276 9680
rect 34540 9640 34580 9680
rect 36556 9640 36596 9680
rect 36940 9640 36980 9680
rect 37324 9640 37364 9680
rect 39340 9640 39380 9680
rect 39724 9640 39764 9680
rect 40108 9640 40148 9680
rect 40684 9640 40724 9680
rect 41068 9640 41108 9680
rect 3820 9556 3860 9596
rect 1516 9472 1556 9512
rect 1612 9472 1652 9512
rect 1708 9472 1748 9512
rect 1900 9472 1940 9512
rect 1996 9472 2036 9512
rect 2380 9472 2420 9512
rect 3628 9472 3668 9512
rect 4295 9472 4335 9512
rect 4396 9472 4436 9512
rect 4492 9472 4532 9512
rect 4684 9472 4724 9512
rect 4780 9472 4820 9512
rect 4972 9472 5012 9512
rect 5452 9472 5492 9512
rect 6700 9472 6740 9512
rect 6988 9472 7028 9512
rect 7180 9472 7220 9512
rect 7276 9472 7316 9512
rect 7660 9472 7700 9512
rect 7756 9472 7796 9512
rect 7852 9472 7892 9512
rect 7948 9472 7988 9512
rect 8332 9472 8372 9512
rect 8620 9472 8660 9512
rect 8716 9472 8756 9512
rect 8812 9472 8852 9512
rect 8908 9472 8948 9512
rect 9100 9472 9140 9512
rect 9196 9472 9236 9512
rect 9868 9472 9908 9512
rect 11116 9472 11156 9512
rect 11500 9472 11540 9512
rect 12748 9472 12788 9512
rect 13132 9472 13172 9512
rect 14380 9472 14420 9512
rect 14764 9472 14804 9512
rect 16012 9472 16052 9512
rect 16396 9472 16436 9512
rect 17644 9472 17684 9512
rect 18124 9472 18164 9512
rect 19372 9472 19412 9512
rect 19756 9472 19796 9512
rect 21004 9472 21044 9512
rect 21388 9472 21428 9512
rect 22636 9472 22676 9512
rect 23212 9472 23252 9512
rect 24460 9472 24500 9512
rect 25036 9472 25076 9512
rect 26284 9472 26324 9512
rect 26668 9472 26708 9512
rect 27916 9472 27956 9512
rect 28300 9472 28340 9512
rect 29548 9472 29588 9512
rect 30700 9472 30740 9512
rect 31852 9472 31892 9512
rect 32908 9472 32948 9512
rect 34156 9472 34196 9512
rect 34924 9472 34964 9512
rect 36172 9472 36212 9512
rect 37708 9472 37748 9512
rect 38956 9472 38996 9512
rect 31084 9388 31124 9428
rect 32428 9388 32468 9428
rect 34732 9388 34772 9428
rect 36748 9388 36788 9428
rect 37132 9388 37172 9428
rect 37516 9388 37556 9428
rect 39532 9388 39572 9428
rect 39916 9388 39956 9428
rect 40300 9388 40340 9428
rect 40492 9388 40532 9428
rect 40876 9388 40916 9428
rect 41260 9388 41300 9428
rect 5260 9304 5300 9344
rect 8332 9304 8372 9344
rect 41452 9304 41492 9344
rect 4780 9220 4820 9260
rect 5068 9220 5108 9260
rect 6892 9220 6932 9260
rect 8140 9220 8180 9260
rect 11308 9220 11348 9260
rect 12940 9220 12980 9260
rect 14572 9220 14612 9260
rect 16204 9220 16244 9260
rect 17836 9220 17876 9260
rect 19564 9220 19604 9260
rect 21196 9220 21236 9260
rect 22828 9220 22868 9260
rect 24652 9220 24692 9260
rect 24844 9220 24884 9260
rect 26476 9220 26516 9260
rect 28108 9220 28148 9260
rect 30220 9220 30260 9260
rect 34348 9220 34388 9260
rect 36364 9220 36404 9260
rect 39148 9220 39188 9260
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 33928 9052 33968 9092
rect 34010 9052 34050 9092
rect 34092 9052 34132 9092
rect 34174 9052 34214 9092
rect 34256 9052 34296 9092
rect 5644 8884 5684 8924
rect 9196 8884 9236 8924
rect 20236 8800 20276 8840
rect 21100 8800 21140 8840
rect 22732 8800 22772 8840
rect 30892 8800 30932 8840
rect 11116 8716 11156 8756
rect 20044 8716 20084 8756
rect 20524 8716 20564 8756
rect 20908 8716 20948 8756
rect 1324 8632 1364 8672
rect 2572 8632 2612 8672
rect 3148 8637 3188 8677
rect 3628 8632 3668 8672
rect 4108 8632 4148 8672
rect 4204 8632 4244 8672
rect 4588 8632 4628 8672
rect 4684 8632 4724 8672
rect 5260 8632 5300 8672
rect 5356 8632 5396 8672
rect 6124 8632 6164 8672
rect 7372 8632 7412 8672
rect 7756 8632 7796 8672
rect 9004 8632 9044 8672
rect 9484 8632 9524 8672
rect 9580 8632 9620 8672
rect 9676 8632 9716 8672
rect 9964 8632 10004 8672
rect 10060 8632 10100 8672
rect 10540 8632 10580 8672
rect 10636 8632 10676 8672
rect 11020 8632 11060 8672
rect 11596 8632 11636 8672
rect 12076 8646 12116 8686
rect 12460 8632 12500 8672
rect 12556 8632 12596 8672
rect 13132 8632 13172 8672
rect 13228 8632 13268 8672
rect 13516 8632 13556 8672
rect 13612 8632 13652 8672
rect 13996 8632 14036 8672
rect 14092 8632 14132 8672
rect 14572 8632 14612 8672
rect 15052 8637 15092 8677
rect 15436 8632 15476 8672
rect 15532 8632 15572 8672
rect 15628 8632 15668 8672
rect 15724 8632 15764 8672
rect 16204 8632 16244 8672
rect 17452 8632 17492 8672
rect 17932 8632 17972 8672
rect 18028 8632 18068 8672
rect 18412 8632 18452 8672
rect 19516 8674 19556 8714
rect 27244 8716 27284 8756
rect 38764 8716 38804 8756
rect 40876 8716 40916 8756
rect 41260 8716 41300 8756
rect 18508 8632 18548 8672
rect 18988 8632 19028 8672
rect 21292 8632 21332 8672
rect 22540 8632 22580 8672
rect 23020 8632 23060 8672
rect 23116 8632 23156 8672
rect 23500 8632 23540 8672
rect 24604 8674 24644 8714
rect 23596 8632 23636 8672
rect 24076 8632 24116 8672
rect 25132 8632 25172 8672
rect 25228 8632 25268 8672
rect 25612 8632 25652 8672
rect 25708 8632 25748 8672
rect 26188 8632 26228 8672
rect 26668 8646 26708 8686
rect 28780 8632 28820 8672
rect 29644 8632 29684 8672
rect 31084 8632 31124 8672
rect 31948 8632 31988 8672
rect 32812 8632 32852 8672
rect 35500 8632 35540 8672
rect 36364 8632 36404 8672
rect 37132 8632 37172 8672
rect 38380 8632 38420 8672
rect 39148 8632 39188 8672
rect 40396 8632 40436 8672
rect 2956 8548 2996 8588
rect 26860 8548 26900 8588
rect 30028 8548 30068 8588
rect 31564 8548 31604 8588
rect 36748 8548 36788 8588
rect 2764 8464 2804 8504
rect 5164 8460 5204 8500
rect 7564 8464 7604 8504
rect 9772 8464 9812 8504
rect 10252 8464 10292 8504
rect 12268 8464 12308 8504
rect 12748 8464 12788 8504
rect 12940 8464 12980 8504
rect 15244 8464 15284 8504
rect 17644 8464 17684 8504
rect 19660 8464 19700 8504
rect 20716 8464 20756 8504
rect 24748 8464 24788 8504
rect 27052 8464 27092 8504
rect 27628 8464 27668 8504
rect 33964 8464 34004 8504
rect 34348 8464 34388 8504
rect 36940 8464 36980 8504
rect 38572 8464 38612 8504
rect 40588 8464 40628 8504
rect 41068 8464 41108 8504
rect 41452 8464 41492 8504
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 35168 8296 35208 8336
rect 35250 8296 35290 8336
rect 35332 8296 35372 8336
rect 35414 8296 35454 8336
rect 35496 8296 35536 8336
rect 2860 8128 2900 8168
rect 3052 8128 3092 8168
rect 8140 8128 8180 8168
rect 9868 8128 9908 8168
rect 10348 8128 10388 8168
rect 13612 8128 13652 8168
rect 15724 8128 15764 8168
rect 18316 8128 18356 8168
rect 22444 8128 22484 8168
rect 38188 8128 38228 8168
rect 40876 8128 40916 8168
rect 26572 8044 26612 8084
rect 28588 8044 28628 8084
rect 40492 8044 40532 8084
rect 1420 7960 1460 8000
rect 2668 7960 2708 8000
rect 3244 7960 3284 8000
rect 4492 7960 4532 8000
rect 4972 7960 5012 8000
rect 5260 7960 5300 8000
rect 5356 7960 5396 8000
rect 5836 7960 5876 8000
rect 7084 7960 7124 8000
rect 7660 7960 7700 8000
rect 7756 7960 7796 8000
rect 7948 7960 7988 8000
rect 8044 7960 8084 8000
rect 8201 7945 8241 7985
rect 8524 7960 8564 8000
rect 8812 7960 8852 8000
rect 8908 7960 8948 8000
rect 9388 7960 9428 8000
rect 9484 7960 9524 8000
rect 9580 7960 9620 8000
rect 9676 7960 9716 8000
rect 9964 7960 10004 8000
rect 10060 7960 10100 8000
rect 10156 7960 10196 8000
rect 10540 7960 10580 8000
rect 11788 7960 11828 8000
rect 12172 7960 12212 8000
rect 13420 7960 13460 8000
rect 13804 7960 13844 8000
rect 15052 7960 15092 8000
rect 15436 7960 15476 8000
rect 15532 7960 15572 8000
rect 15916 7960 15956 8000
rect 16012 7960 16052 8000
rect 16108 7960 16148 8000
rect 16204 7960 16244 8000
rect 16588 7960 16628 8000
rect 16684 7960 16724 8000
rect 17644 7960 17684 8000
rect 18124 7955 18164 7995
rect 18508 7960 18548 8000
rect 19756 7960 19796 8000
rect 20812 7960 20852 8000
rect 22060 7960 22100 8000
rect 23500 7960 23540 8000
rect 24748 7960 24788 8000
rect 25132 7960 25172 8000
rect 26380 7960 26420 8000
rect 26860 7960 26900 8000
rect 26956 7960 26996 8000
rect 27340 7960 27380 8000
rect 27916 7960 27956 8000
rect 28396 7955 28436 7995
rect 28972 7960 29012 8000
rect 30220 7960 30260 8000
rect 30604 7960 30644 8000
rect 31852 7960 31892 8000
rect 32428 7960 32468 8000
rect 33676 7960 33716 8000
rect 35116 7960 35156 8000
rect 35980 7960 36020 8000
rect 36364 7960 36404 8000
rect 36652 7960 36692 8000
rect 38764 7960 38804 8000
rect 38860 7960 38900 8000
rect 39820 7960 39860 8000
rect 40348 7950 40388 7990
rect 17068 7876 17108 7916
rect 17164 7876 17204 7916
rect 20428 7876 20468 7916
rect 22636 7876 22676 7916
rect 27436 7876 27476 7916
rect 38380 7876 38420 7916
rect 39244 7876 39284 7916
rect 39340 7876 39380 7916
rect 40684 7876 40724 7916
rect 41068 7876 41108 7916
rect 41452 7876 41492 7916
rect 9196 7792 9236 7832
rect 37804 7792 37844 7832
rect 41644 7792 41684 7832
rect 5644 7708 5684 7748
rect 7276 7708 7316 7748
rect 15244 7708 15284 7748
rect 19948 7708 19988 7748
rect 20620 7708 20660 7748
rect 22252 7708 22292 7748
rect 24940 7708 24980 7748
rect 30412 7708 30452 7748
rect 32044 7708 32084 7748
rect 32236 7708 32276 7748
rect 33964 7708 34004 7748
rect 36940 7708 36980 7748
rect 41260 7708 41300 7748
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 33928 7540 33968 7580
rect 34010 7540 34050 7580
rect 34092 7540 34132 7580
rect 34174 7540 34214 7580
rect 34256 7540 34296 7580
rect 3532 7372 3572 7412
rect 9004 7372 9044 7412
rect 9868 7372 9908 7412
rect 32332 7372 32372 7412
rect 37804 7372 37844 7412
rect 2956 7288 2996 7328
rect 29548 7288 29588 7328
rect 3244 7204 3284 7244
rect 5452 7204 5492 7244
rect 25228 7204 25268 7244
rect 25612 7204 25652 7244
rect 29356 7204 29396 7244
rect 1324 7120 1364 7160
rect 1516 7120 1556 7160
rect 2764 7120 2804 7160
rect 3148 7120 3188 7160
rect 3340 7120 3380 7160
rect 3916 7120 3956 7160
rect 4204 7120 4244 7160
rect 4492 7120 4532 7160
rect 4684 7120 4724 7160
rect 4972 7120 5012 7160
rect 5068 7120 5108 7160
rect 5548 7120 5588 7160
rect 6028 7120 6068 7160
rect 6508 7125 6548 7165
rect 7084 7120 7124 7160
rect 7180 7120 7220 7160
rect 7564 7120 7604 7160
rect 7660 7120 7700 7160
rect 8140 7120 8180 7160
rect 8620 7125 8660 7165
rect 9004 7120 9044 7160
rect 9292 7120 9332 7160
rect 9484 7120 9524 7160
rect 9580 7120 9620 7160
rect 9676 7120 9716 7160
rect 10060 7120 10100 7160
rect 11308 7120 11348 7160
rect 11884 7120 11924 7160
rect 13132 7120 13172 7160
rect 13516 7120 13556 7160
rect 13708 7120 13748 7160
rect 13804 7120 13844 7160
rect 13996 7120 14036 7160
rect 14092 7120 14132 7160
rect 14188 7120 14228 7160
rect 14284 7120 14324 7160
rect 14476 7120 14516 7160
rect 15724 7120 15764 7160
rect 16108 7120 16148 7160
rect 17356 7120 17396 7160
rect 17740 7120 17780 7160
rect 18988 7120 19028 7160
rect 19372 7120 19412 7160
rect 20620 7120 20660 7160
rect 21388 7120 21428 7160
rect 22636 7120 22676 7160
rect 23116 7120 23156 7160
rect 23212 7120 23252 7160
rect 23596 7120 23636 7160
rect 24700 7162 24740 7202
rect 32140 7204 32180 7244
rect 32524 7204 32564 7244
rect 36460 7204 36500 7244
rect 23692 7120 23732 7160
rect 24172 7120 24212 7160
rect 25900 7120 25940 7160
rect 27148 7120 27188 7160
rect 27532 7120 27572 7160
rect 28780 7120 28820 7160
rect 30028 7120 30068 7160
rect 30124 7120 30164 7160
rect 30508 7120 30548 7160
rect 31612 7162 31652 7202
rect 37996 7204 38036 7244
rect 39052 7204 39092 7244
rect 40684 7204 40724 7244
rect 40876 7204 40916 7244
rect 41260 7204 41300 7244
rect 30604 7120 30644 7160
rect 31084 7120 31124 7160
rect 32908 7120 32948 7160
rect 34156 7120 34196 7160
rect 34540 7120 34580 7160
rect 35500 7120 35540 7160
rect 35884 7120 35924 7160
rect 35980 7120 36020 7160
rect 36364 7120 36404 7160
rect 36940 7120 36980 7160
rect 37420 7134 37460 7174
rect 38572 7120 38612 7160
rect 38668 7120 38708 7160
rect 39148 7120 39188 7160
rect 39628 7120 39668 7160
rect 40108 7125 40148 7165
rect 3820 7036 3860 7076
rect 4588 7036 4628 7076
rect 6700 7036 6740 7076
rect 8812 7036 8852 7076
rect 13612 7036 13652 7076
rect 22828 7036 22868 7076
rect 24844 7036 24884 7076
rect 31756 7036 31796 7076
rect 1228 6952 1268 6992
rect 13324 6952 13364 6992
rect 15916 6952 15956 6992
rect 17548 6952 17588 6992
rect 19180 6952 19220 6992
rect 20812 6952 20852 6992
rect 25036 6952 25076 6992
rect 25420 6952 25460 6992
rect 27340 6952 27380 6992
rect 28972 6952 29012 6992
rect 29164 6952 29204 6992
rect 31948 6952 31988 6992
rect 34348 6952 34388 6992
rect 35020 6952 35060 6992
rect 37612 6952 37652 6992
rect 40300 6952 40340 6992
rect 40492 6952 40532 6992
rect 41068 6952 41108 6992
rect 41452 6952 41492 6992
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 35168 6784 35208 6824
rect 35250 6784 35290 6824
rect 35332 6784 35372 6824
rect 35414 6784 35454 6824
rect 35496 6784 35536 6824
rect 1228 6616 1268 6656
rect 3148 6616 3188 6656
rect 6700 6616 6740 6656
rect 8812 6616 8852 6656
rect 11692 6616 11732 6656
rect 15916 6616 15956 6656
rect 20044 6616 20084 6656
rect 38764 6616 38804 6656
rect 40588 6616 40628 6656
rect 4972 6532 5012 6572
rect 5740 6532 5780 6572
rect 15340 6532 15380 6572
rect 19852 6532 19892 6572
rect 22924 6532 22964 6572
rect 28780 6532 28820 6572
rect 34156 6532 34196 6572
rect 36172 6532 36212 6572
rect 1420 6448 1460 6488
rect 1516 6448 1556 6488
rect 1708 6448 1748 6488
rect 2956 6448 2996 6488
rect 3820 6448 3860 6488
rect 3916 6448 3956 6488
rect 4204 6448 4244 6488
rect 4588 6448 4628 6488
rect 4876 6448 4916 6488
rect 5836 6448 5876 6488
rect 6124 6448 6164 6488
rect 6508 6448 6548 6488
rect 6604 6448 6644 6488
rect 6796 6448 6836 6488
rect 7084 6448 7124 6488
rect 7180 6448 7220 6488
rect 8140 6448 8180 6488
rect 8620 6434 8660 6474
rect 7564 6364 7604 6404
rect 7660 6364 7700 6404
rect 9004 6403 9044 6443
rect 9100 6448 9140 6488
rect 9196 6448 9236 6488
rect 9292 6448 9332 6488
rect 9580 6448 9620 6488
rect 10828 6448 10868 6488
rect 11404 6448 11444 6488
rect 11500 6448 11540 6488
rect 11596 6448 11636 6488
rect 11884 6448 11924 6488
rect 13132 6448 13172 6488
rect 13612 6448 13652 6488
rect 13708 6448 13748 6488
rect 14668 6448 14708 6488
rect 15196 6438 15236 6478
rect 16108 6448 16148 6488
rect 17356 6448 17396 6488
rect 18124 6448 18164 6488
rect 18220 6448 18260 6488
rect 19180 6448 19220 6488
rect 19708 6438 19748 6478
rect 21196 6448 21236 6488
rect 21292 6448 21332 6488
rect 22252 6448 22292 6488
rect 22732 6443 22772 6483
rect 23116 6448 23156 6488
rect 24364 6448 24404 6488
rect 24940 6448 24980 6488
rect 26188 6448 26228 6488
rect 27052 6448 27092 6488
rect 27148 6448 27188 6488
rect 27532 6448 27572 6488
rect 28108 6448 28148 6488
rect 28636 6438 28676 6478
rect 29164 6448 29204 6488
rect 30412 6448 30452 6488
rect 30700 6448 30740 6488
rect 31948 6448 31988 6488
rect 32428 6448 32468 6488
rect 32524 6448 32564 6488
rect 33484 6448 33524 6488
rect 33964 6443 34004 6483
rect 34444 6448 34484 6488
rect 34540 6448 34580 6488
rect 34924 6448 34964 6488
rect 35500 6448 35540 6488
rect 36028 6438 36068 6478
rect 37324 6448 37364 6488
rect 38572 6448 38612 6488
rect 39148 6448 39188 6488
rect 40396 6448 40436 6488
rect 14092 6364 14132 6404
rect 14188 6364 14228 6404
rect 15724 6364 15764 6404
rect 18604 6364 18644 6404
rect 18700 6364 18740 6404
rect 20236 6364 20276 6404
rect 21676 6364 21716 6404
rect 21772 6364 21812 6404
rect 27628 6364 27668 6404
rect 32908 6364 32948 6404
rect 33004 6364 33044 6404
rect 35020 6364 35060 6404
rect 40876 6364 40916 6404
rect 41260 6364 41300 6404
rect 5260 6280 5300 6320
rect 5452 6280 5492 6320
rect 17548 6280 17588 6320
rect 36364 6280 36404 6320
rect 36748 6280 36788 6320
rect 41068 6280 41108 6320
rect 3532 6196 3572 6236
rect 11020 6196 11060 6236
rect 13324 6196 13364 6236
rect 24556 6196 24596 6236
rect 26380 6196 26420 6236
rect 28972 6196 29012 6236
rect 32140 6196 32180 6236
rect 41452 6196 41492 6236
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 33928 6028 33968 6068
rect 34010 6028 34050 6068
rect 34092 6028 34132 6068
rect 34174 6028 34214 6068
rect 34256 6028 34296 6068
rect 3148 5860 3188 5900
rect 5836 5860 5876 5900
rect 8140 5860 8180 5900
rect 31660 5860 31700 5900
rect 34252 5860 34292 5900
rect 36172 5860 36212 5900
rect 41452 5860 41492 5900
rect 3724 5776 3764 5816
rect 4684 5776 4724 5816
rect 10060 5776 10100 5816
rect 41068 5776 41108 5816
rect 6604 5692 6644 5732
rect 13228 5692 13268 5732
rect 21100 5692 21140 5732
rect 22828 5692 22868 5732
rect 23212 5692 23252 5732
rect 23884 5692 23924 5732
rect 26476 5692 26516 5732
rect 27148 5692 27188 5732
rect 29932 5692 29972 5732
rect 1228 5608 1268 5648
rect 1420 5608 1460 5648
rect 1516 5608 1556 5648
rect 1708 5608 1748 5648
rect 2956 5608 2996 5648
rect 3340 5608 3380 5648
rect 3532 5608 3572 5648
rect 4108 5608 4148 5648
rect 4396 5608 4436 5648
rect 4684 5608 4724 5648
rect 4876 5608 4916 5648
rect 5164 5608 5204 5648
rect 5452 5608 5492 5648
rect 6124 5608 6164 5648
rect 6220 5608 6260 5648
rect 6700 5608 6740 5648
rect 7180 5608 7220 5648
rect 7660 5617 7700 5657
rect 8524 5627 8564 5667
rect 8812 5608 8852 5648
rect 9100 5608 9140 5648
rect 9196 5608 9236 5648
rect 9676 5608 9716 5648
rect 9772 5608 9812 5648
rect 9868 5608 9908 5648
rect 10060 5608 10100 5648
rect 10252 5608 10292 5648
rect 10348 5608 10388 5648
rect 10540 5608 10580 5648
rect 10924 5608 10964 5648
rect 12172 5608 12212 5648
rect 12652 5608 12692 5648
rect 12748 5608 12788 5648
rect 13132 5608 13172 5648
rect 13708 5608 13748 5648
rect 14188 5613 14228 5653
rect 16204 5608 16244 5648
rect 17452 5608 17492 5648
rect 17932 5608 17972 5648
rect 18028 5627 18068 5667
rect 18412 5608 18452 5648
rect 18508 5608 18548 5648
rect 18988 5608 19028 5648
rect 19468 5622 19508 5662
rect 20620 5608 20660 5648
rect 20716 5608 20756 5648
rect 21196 5608 21236 5648
rect 21676 5608 21716 5648
rect 22156 5622 22196 5662
rect 24364 5608 24404 5648
rect 24460 5608 24500 5648
rect 24844 5608 24884 5648
rect 25948 5650 25988 5690
rect 31468 5692 31508 5732
rect 31852 5692 31892 5732
rect 32812 5692 32852 5732
rect 34444 5692 34484 5732
rect 36556 5692 36596 5732
rect 37228 5692 37268 5732
rect 40108 5692 40148 5732
rect 40492 5692 40532 5732
rect 40876 5692 40916 5732
rect 41260 5692 41300 5732
rect 24940 5608 24980 5648
rect 25420 5608 25460 5648
rect 27628 5608 27668 5648
rect 28876 5608 28916 5648
rect 29356 5608 29396 5648
rect 29452 5608 29492 5648
rect 29836 5608 29876 5648
rect 30412 5608 30452 5648
rect 30940 5617 30980 5657
rect 32332 5608 32372 5648
rect 32428 5608 32468 5648
rect 32908 5608 32948 5648
rect 33388 5608 33428 5648
rect 33868 5622 33908 5662
rect 34732 5608 34772 5648
rect 35980 5608 36020 5648
rect 37516 5608 37556 5648
rect 37612 5608 37652 5648
rect 37996 5608 38036 5648
rect 38092 5608 38132 5648
rect 38572 5608 38612 5648
rect 39100 5617 39140 5657
rect 3436 5524 3476 5564
rect 4012 5524 4052 5564
rect 5548 5524 5588 5564
rect 8428 5524 8468 5564
rect 12364 5524 12404 5564
rect 22348 5524 22388 5564
rect 26092 5524 26132 5564
rect 29068 5524 29108 5564
rect 31084 5524 31124 5564
rect 1324 5440 1364 5480
rect 3148 5440 3188 5480
rect 7852 5440 7892 5480
rect 9388 5440 9428 5480
rect 9580 5440 9620 5480
rect 10636 5440 10676 5480
rect 14380 5440 14420 5480
rect 17644 5440 17684 5480
rect 19660 5440 19700 5480
rect 22636 5440 22676 5480
rect 23020 5440 23060 5480
rect 24076 5440 24116 5480
rect 26284 5440 26324 5480
rect 27340 5440 27380 5480
rect 31276 5440 31316 5480
rect 34060 5440 34100 5480
rect 36364 5440 36404 5480
rect 37036 5440 37076 5480
rect 39244 5440 39284 5480
rect 39916 5440 39956 5480
rect 40684 5440 40724 5480
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 35168 5272 35208 5312
rect 35250 5272 35290 5312
rect 35332 5272 35372 5312
rect 35414 5272 35454 5312
rect 35496 5272 35536 5312
rect 3532 5146 3572 5186
rect 6508 5104 6548 5144
rect 8716 5104 8756 5144
rect 13996 5104 14036 5144
rect 31084 5104 31124 5144
rect 36268 5104 36308 5144
rect 3148 5020 3188 5060
rect 3820 5020 3860 5060
rect 8524 5020 8564 5060
rect 16300 5020 16340 5060
rect 18316 5020 18356 5060
rect 34636 5020 34676 5060
rect 36940 5020 36980 5060
rect 1324 4936 1364 4976
rect 2572 4936 2612 4976
rect 3052 4936 3092 4976
rect 3244 4936 3284 4976
rect 3340 4936 3380 4976
rect 3916 4936 3956 4976
rect 4204 4936 4244 4976
rect 4588 4936 4628 4976
rect 4684 4936 4724 4976
rect 4780 4936 4820 4976
rect 4876 4936 4916 4976
rect 5068 4936 5108 4976
rect 6316 4936 6356 4976
rect 6796 4936 6836 4976
rect 6892 4936 6932 4976
rect 7276 4936 7316 4976
rect 7372 4936 7412 4976
rect 7852 4936 7892 4976
rect 8332 4922 8372 4962
rect 8908 4936 8948 4976
rect 10156 4936 10196 4976
rect 10444 4936 10484 4976
rect 11692 4936 11732 4976
rect 12076 4936 12116 4976
rect 12172 4936 12212 4976
rect 12268 4936 12308 4976
rect 12364 4936 12404 4976
rect 12556 4936 12596 4976
rect 13804 4936 13844 4976
rect 14860 4936 14900 4976
rect 16108 4936 16148 4976
rect 16588 4936 16628 4976
rect 16684 4936 16724 4976
rect 17068 4936 17108 4976
rect 17164 4936 17204 4976
rect 17644 4936 17684 4976
rect 18124 4931 18164 4971
rect 22060 4936 22100 4976
rect 23308 4936 23348 4976
rect 24556 4936 24596 4976
rect 25804 4936 25844 4976
rect 26956 4936 26996 4976
rect 28204 4936 28244 4976
rect 29644 4936 29684 4976
rect 30892 4936 30932 4976
rect 31276 4936 31316 4976
rect 32524 4936 32564 4976
rect 33196 4936 33236 4976
rect 34444 4936 34484 4976
rect 35788 4936 35828 4976
rect 37132 4936 37172 4976
rect 38380 4936 38420 4976
rect 38764 4936 38804 4976
rect 40012 4936 40052 4976
rect 20236 4852 20276 4892
rect 21004 4852 21044 4892
rect 26572 4852 26612 4892
rect 28780 4852 28820 4892
rect 29452 4852 29492 4892
rect 35020 4852 35060 4892
rect 35404 4852 35444 4892
rect 40492 4852 40532 4892
rect 40876 4852 40916 4892
rect 41260 4852 41300 4892
rect 2764 4768 2804 4808
rect 35212 4768 35252 4808
rect 40684 4768 40724 4808
rect 41068 4768 41108 4808
rect 41452 4768 41492 4808
rect 11884 4684 11924 4724
rect 20428 4684 20468 4724
rect 21196 4684 21236 4724
rect 23500 4684 23540 4724
rect 25996 4684 26036 4724
rect 26764 4684 26804 4724
rect 28396 4684 28436 4724
rect 28588 4684 28628 4724
rect 29260 4684 29300 4724
rect 32716 4684 32756 4724
rect 34828 4684 34868 4724
rect 38572 4684 38612 4724
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 33928 4516 33968 4556
rect 34010 4516 34050 4556
rect 34092 4516 34132 4556
rect 34174 4516 34214 4556
rect 34256 4516 34296 4556
rect 9004 4348 9044 4388
rect 37228 4348 37268 4388
rect 39244 4348 39284 4388
rect 41068 4348 41108 4388
rect 40300 4264 40340 4304
rect 4204 4180 4244 4220
rect 4300 4180 4340 4220
rect 6700 4180 6740 4220
rect 1420 4096 1460 4136
rect 2668 4096 2708 4136
rect 3244 4110 3284 4150
rect 3724 4096 3764 4136
rect 4684 4096 4724 4136
rect 4780 4096 4820 4136
rect 5068 4096 5108 4136
rect 5164 4096 5204 4136
rect 5356 4096 5396 4136
rect 5548 4096 5588 4136
rect 5644 4096 5684 4136
rect 5740 4096 5780 4136
rect 5836 4096 5876 4136
rect 6124 4096 6164 4136
rect 6220 4096 6260 4136
rect 6604 4096 6644 4136
rect 7180 4096 7220 4136
rect 7660 4110 7700 4150
rect 8332 4096 8372 4136
rect 8620 4096 8660 4136
rect 8716 4096 8756 4136
rect 9196 4096 9236 4136
rect 10444 4096 10484 4136
rect 10828 4096 10868 4136
rect 12076 4096 12116 4136
rect 12460 4096 12500 4136
rect 13708 4096 13748 4136
rect 14188 4096 14228 4136
rect 14284 4096 14324 4136
rect 14668 4096 14708 4136
rect 15772 4138 15812 4178
rect 18028 4180 18068 4220
rect 18124 4180 18164 4220
rect 14764 4096 14804 4136
rect 15244 4096 15284 4136
rect 17548 4096 17588 4136
rect 17644 4096 17684 4136
rect 18604 4096 18644 4136
rect 19084 4101 19124 4141
rect 20044 4096 20084 4136
rect 21292 4096 21332 4136
rect 21772 4096 21812 4136
rect 21868 4096 21908 4136
rect 22252 4138 22292 4178
rect 22348 4138 22388 4178
rect 23356 4138 23396 4178
rect 24844 4180 24884 4220
rect 28588 4180 28628 4220
rect 32044 4180 32084 4220
rect 32908 4180 32948 4220
rect 34444 4180 34484 4220
rect 35020 4180 35060 4220
rect 35788 4180 35828 4220
rect 35884 4180 35924 4220
rect 37420 4180 37460 4220
rect 39628 4180 39668 4220
rect 39916 4180 39956 4220
rect 40492 4180 40532 4220
rect 40876 4180 40916 4220
rect 41260 4180 41300 4220
rect 22828 4096 22868 4136
rect 24268 4096 24308 4136
rect 24364 4096 24404 4136
rect 24748 4096 24788 4136
rect 25324 4096 25364 4136
rect 25852 4105 25892 4145
rect 26188 4096 26228 4136
rect 27436 4096 27476 4136
rect 28108 4096 28148 4136
rect 28204 4096 28244 4136
rect 28684 4096 28724 4136
rect 29164 4096 29204 4136
rect 29644 4110 29684 4150
rect 30220 4096 30260 4136
rect 31468 4096 31508 4136
rect 32332 4115 32372 4155
rect 32428 4096 32468 4136
rect 32812 4096 32852 4136
rect 33388 4096 33428 4136
rect 33868 4101 33908 4141
rect 35308 4096 35348 4136
rect 35404 4096 35444 4136
rect 36364 4096 36404 4136
rect 36844 4101 36884 4141
rect 37804 4096 37844 4136
rect 39052 4096 39092 4136
rect 21484 4012 21524 4052
rect 25996 4012 26036 4052
rect 34060 4012 34100 4052
rect 37036 4012 37076 4052
rect 2860 3928 2900 3968
rect 3052 3928 3092 3968
rect 7852 3928 7892 3968
rect 10636 3928 10676 3968
rect 12268 3928 12308 3968
rect 13900 3928 13940 3968
rect 15916 3928 15956 3968
rect 19276 3928 19316 3968
rect 23500 3928 23540 3968
rect 27628 3928 27668 3968
rect 29836 3928 29876 3968
rect 30028 3928 30068 3968
rect 31852 3928 31892 3968
rect 34252 3928 34292 3968
rect 34828 3928 34868 3968
rect 39436 3928 39476 3968
rect 40108 3928 40148 3968
rect 41452 3928 41492 3968
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 35168 3760 35208 3800
rect 35250 3760 35290 3800
rect 35332 3760 35372 3800
rect 35414 3760 35454 3800
rect 35496 3760 35536 3800
rect 3052 3592 3092 3632
rect 3532 3592 3572 3632
rect 4204 3592 4244 3632
rect 5932 3592 5972 3632
rect 17452 3592 17492 3632
rect 19084 3592 19124 3632
rect 24556 3592 24596 3632
rect 29932 3592 29972 3632
rect 32140 3592 32180 3632
rect 32332 3592 32372 3632
rect 34444 3592 34484 3632
rect 34636 3592 34676 3632
rect 41068 3592 41108 3632
rect 8332 3508 8372 3548
rect 10444 3508 10484 3548
rect 12460 3508 12500 3548
rect 14860 3508 14900 3548
rect 27244 3508 27284 3548
rect 39148 3508 39188 3548
rect 1228 3424 1268 3464
rect 1420 3445 1460 3485
rect 1612 3424 1652 3464
rect 2860 3424 2900 3464
rect 3244 3424 3284 3464
rect 3340 3424 3380 3464
rect 3436 3424 3476 3464
rect 3724 3424 3764 3464
rect 3820 3424 3860 3464
rect 4012 3424 4052 3464
rect 4108 3424 4148 3464
rect 4209 3424 4249 3464
rect 4492 3424 4532 3464
rect 5740 3424 5780 3464
rect 6412 3424 6452 3464
rect 7660 3424 7700 3464
rect 7948 3424 7988 3464
rect 8236 3424 8276 3464
rect 9004 3424 9044 3464
rect 10252 3424 10292 3464
rect 10732 3424 10772 3464
rect 10828 3424 10868 3464
rect 11308 3424 11348 3464
rect 11788 3424 11828 3464
rect 12268 3419 12308 3459
rect 13132 3424 13172 3464
rect 13228 3424 13268 3464
rect 13612 3424 13652 3464
rect 14188 3424 14228 3464
rect 14668 3419 14708 3459
rect 16012 3424 16052 3464
rect 17260 3424 17300 3464
rect 17644 3424 17684 3464
rect 18892 3424 18932 3464
rect 20524 3424 20564 3464
rect 21772 3424 21812 3464
rect 23116 3424 23156 3464
rect 24364 3424 24404 3464
rect 25516 3424 25556 3464
rect 25612 3424 25652 3464
rect 26092 3424 26132 3464
rect 26572 3424 26612 3464
rect 27052 3410 27092 3450
rect 28204 3424 28244 3464
rect 28300 3424 28340 3464
rect 28684 3424 28724 3464
rect 29260 3424 29300 3464
rect 29740 3410 29780 3450
rect 30412 3424 30452 3464
rect 30508 3424 30548 3464
rect 30988 3424 31028 3464
rect 31468 3424 31508 3464
rect 31948 3410 31988 3450
rect 33004 3424 33044 3464
rect 34252 3424 34292 3464
rect 34828 3424 34868 3464
rect 36076 3424 36116 3464
rect 37420 3424 37460 3464
rect 37516 3424 37556 3464
rect 37996 3424 38036 3464
rect 38476 3424 38516 3464
rect 38956 3419 38996 3459
rect 11212 3340 11252 3380
rect 12652 3340 12692 3380
rect 13708 3340 13748 3380
rect 19948 3340 19988 3380
rect 22732 3340 22772 3380
rect 25228 3340 25268 3380
rect 25996 3340 26036 3380
rect 27628 3340 27668 3380
rect 28780 3340 28820 3380
rect 30892 3340 30932 3380
rect 32524 3340 32564 3380
rect 36460 3340 36500 3380
rect 37132 3340 37172 3380
rect 37900 3340 37940 3380
rect 39340 3340 39380 3380
rect 39724 3340 39764 3380
rect 40108 3340 40148 3380
rect 40492 3340 40532 3380
rect 40876 3340 40916 3380
rect 41260 3340 41300 3380
rect 8620 3256 8660 3296
rect 40684 3256 40724 3296
rect 1324 3172 1364 3212
rect 5932 3172 5972 3212
rect 6220 3172 6260 3212
rect 12844 3172 12884 3212
rect 20140 3172 20180 3212
rect 21964 3172 22004 3212
rect 22924 3172 22964 3212
rect 25036 3172 25076 3212
rect 27436 3172 27476 3212
rect 36268 3172 36308 3212
rect 36940 3172 36980 3212
rect 39532 3172 39572 3212
rect 39916 3172 39956 3212
rect 40300 3172 40340 3212
rect 41452 3172 41492 3212
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 33928 3004 33968 3044
rect 34010 3004 34050 3044
rect 34092 3004 34132 3044
rect 34174 3004 34214 3044
rect 34256 3004 34296 3044
rect 5068 2836 5108 2876
rect 15052 2836 15092 2876
rect 28108 2836 28148 2876
rect 29740 2836 29780 2876
rect 31372 2836 31412 2876
rect 37996 2836 38036 2876
rect 14572 2752 14612 2792
rect 25708 2752 25748 2792
rect 36364 2752 36404 2792
rect 41644 2752 41684 2792
rect 11020 2668 11060 2708
rect 15532 2668 15572 2708
rect 15916 2668 15956 2708
rect 22444 2668 22484 2708
rect 22540 2668 22580 2708
rect 24076 2668 24116 2708
rect 41452 2668 41492 2708
rect 1324 2584 1364 2624
rect 1420 2584 1460 2624
rect 1516 2584 1556 2624
rect 1612 2584 1652 2624
rect 1804 2584 1844 2624
rect 3052 2584 3092 2624
rect 3436 2584 3476 2624
rect 4684 2584 4724 2624
rect 5068 2584 5108 2624
rect 5260 2584 5300 2624
rect 5356 2584 5396 2624
rect 5548 2584 5588 2624
rect 6796 2584 6836 2624
rect 7180 2584 7220 2624
rect 8428 2584 8468 2624
rect 8812 2584 8852 2624
rect 10060 2584 10100 2624
rect 10540 2584 10580 2624
rect 10636 2584 10676 2624
rect 11116 2584 11156 2624
rect 11596 2584 11636 2624
rect 12076 2598 12116 2638
rect 12460 2584 12500 2624
rect 13708 2584 13748 2624
rect 14188 2584 14228 2624
rect 14284 2584 14324 2624
rect 14380 2584 14420 2624
rect 14572 2584 14612 2624
rect 14860 2584 14900 2624
rect 15052 2584 15092 2624
rect 15244 2584 15284 2624
rect 15340 2584 15380 2624
rect 20044 2584 20084 2624
rect 21292 2584 21332 2624
rect 21964 2584 22004 2624
rect 22060 2584 22100 2624
rect 23020 2584 23060 2624
rect 23548 2593 23588 2633
rect 24268 2584 24308 2624
rect 25516 2584 25556 2624
rect 26188 2584 26228 2624
rect 26284 2584 26324 2624
rect 26668 2584 26708 2624
rect 26764 2626 26804 2666
rect 27244 2584 27284 2624
rect 27724 2593 27764 2633
rect 28300 2584 28340 2624
rect 29548 2584 29588 2624
rect 29932 2584 29972 2624
rect 31180 2584 31220 2624
rect 31564 2584 31604 2624
rect 32812 2584 32852 2624
rect 33004 2584 33044 2624
rect 34252 2584 34292 2624
rect 34924 2584 34964 2624
rect 36172 2584 36212 2624
rect 36556 2584 36596 2624
rect 37804 2584 37844 2624
rect 38380 2584 38420 2624
rect 39628 2584 39668 2624
rect 40012 2584 40052 2624
rect 41260 2584 41300 2624
rect 4876 2500 4916 2540
rect 6988 2500 7028 2540
rect 12268 2500 12308 2540
rect 23692 2500 23732 2540
rect 34444 2500 34484 2540
rect 3244 2416 3284 2456
rect 8620 2416 8660 2456
rect 10252 2416 10292 2456
rect 13900 2416 13940 2456
rect 14092 2416 14132 2456
rect 15724 2416 15764 2456
rect 16108 2416 16148 2456
rect 21484 2416 21524 2456
rect 23884 2416 23924 2456
rect 27916 2416 27956 2456
rect 38188 2416 38228 2456
rect 39820 2416 39860 2456
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 35168 2248 35208 2288
rect 35250 2248 35290 2288
rect 35332 2248 35372 2288
rect 35414 2248 35454 2288
rect 35496 2248 35536 2288
rect 3244 2080 3284 2120
rect 7276 2080 7316 2120
rect 10252 2080 10292 2120
rect 13228 2080 13268 2120
rect 15628 2080 15668 2120
rect 25996 2080 26036 2120
rect 26188 2080 26228 2120
rect 33964 2080 34004 2120
rect 36076 2080 36116 2120
rect 38476 2080 38516 2120
rect 41260 2080 41300 2120
rect 41644 2080 41684 2120
rect 4876 1996 4916 2036
rect 6892 1996 6932 2036
rect 9580 1996 9620 2036
rect 12556 1996 12596 2036
rect 12748 1996 12788 2036
rect 17836 1996 17876 2036
rect 19852 1996 19892 2036
rect 23116 1996 23156 2036
rect 30700 1996 30740 2036
rect 40492 1996 40532 2036
rect 1324 1912 1364 1952
rect 1420 1912 1460 1952
rect 1516 1912 1556 1952
rect 1612 1912 1652 1952
rect 1804 1912 1844 1952
rect 3052 1912 3092 1952
rect 3436 1912 3476 1952
rect 4684 1912 4724 1952
rect 5164 1912 5204 1952
rect 5260 1912 5300 1952
rect 5740 1912 5780 1952
rect 6220 1912 6260 1952
rect 6700 1898 6740 1938
rect 7372 1912 7412 1952
rect 7468 1912 7508 1952
rect 7564 1912 7604 1952
rect 7852 1912 7892 1952
rect 7948 1912 7988 1952
rect 8908 1912 8948 1952
rect 9388 1907 9428 1947
rect 9772 1912 9812 1952
rect 9868 1912 9908 1952
rect 9964 1912 10004 1952
rect 10060 1912 10100 1952
rect 10444 1912 10484 1952
rect 10540 1912 10580 1952
rect 10828 1912 10868 1952
rect 10924 1912 10964 1952
rect 11404 1912 11444 1952
rect 11884 1912 11924 1952
rect 12364 1898 12404 1938
rect 12844 1933 12884 1973
rect 12940 1912 12980 1952
rect 13036 1912 13076 1952
rect 13420 1912 13460 1952
rect 13900 1912 13940 1952
rect 13996 1912 14036 1952
rect 14476 1912 14516 1952
rect 14956 1912 14996 1952
rect 15436 1898 15476 1938
rect 16396 1912 16436 1952
rect 17644 1912 17684 1952
rect 18124 1912 18164 1952
rect 18220 1912 18260 1952
rect 18604 1912 18644 1952
rect 19180 1912 19220 1952
rect 19660 1898 19700 1938
rect 21388 1912 21428 1952
rect 21484 1912 21524 1952
rect 21868 1912 21908 1952
rect 21964 1912 22004 1952
rect 22444 1912 22484 1952
rect 5644 1828 5684 1868
rect 8332 1828 8372 1868
rect 8428 1828 8468 1868
rect 11308 1828 11348 1868
rect 14380 1828 14420 1868
rect 15820 1828 15860 1868
rect 22972 1870 23012 1910
rect 24268 1912 24308 1952
rect 24364 1912 24404 1952
rect 24748 1912 24788 1952
rect 25324 1912 25364 1952
rect 25804 1898 25844 1938
rect 26380 1912 26420 1952
rect 27628 1912 27668 1952
rect 28972 1912 29012 1952
rect 29068 1912 29108 1952
rect 30028 1912 30068 1952
rect 30508 1898 30548 1938
rect 32236 1912 32276 1952
rect 32332 1912 32372 1952
rect 32716 1912 32756 1952
rect 32812 1912 32852 1952
rect 33292 1912 33332 1952
rect 33772 1907 33812 1947
rect 34348 1912 34388 1952
rect 34444 1912 34484 1952
rect 34924 1912 34964 1952
rect 35404 1912 35444 1952
rect 35884 1898 35924 1938
rect 36748 1912 36788 1952
rect 36844 1912 36884 1952
rect 37228 1912 37268 1952
rect 37324 1912 37364 1952
rect 37804 1912 37844 1952
rect 38284 1907 38324 1947
rect 38764 1912 38804 1952
rect 38860 1912 38900 1952
rect 39340 1912 39380 1952
rect 39820 1912 39860 1952
rect 40300 1907 40340 1947
rect 18700 1828 18740 1868
rect 20908 1828 20948 1868
rect 23308 1828 23348 1868
rect 23884 1828 23924 1868
rect 24844 1828 24884 1868
rect 28012 1828 28052 1868
rect 28396 1828 28436 1868
rect 29452 1828 29492 1868
rect 29548 1828 29588 1868
rect 31084 1828 31124 1868
rect 31468 1828 31508 1868
rect 31948 1828 31988 1868
rect 34828 1828 34868 1868
rect 36460 1828 36500 1868
rect 39244 1828 39284 1868
rect 40876 1828 40916 1868
rect 41068 1828 41108 1868
rect 41452 1828 41492 1868
rect 13420 1744 13460 1784
rect 16012 1660 16052 1700
rect 21100 1660 21140 1700
rect 23500 1660 23540 1700
rect 23692 1660 23732 1700
rect 27820 1660 27860 1700
rect 28204 1660 28244 1700
rect 30892 1660 30932 1700
rect 31276 1660 31316 1700
rect 31756 1660 31796 1700
rect 36268 1660 36308 1700
rect 40684 1660 40724 1700
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 33928 1492 33968 1532
rect 34010 1492 34050 1532
rect 34092 1492 34132 1532
rect 34174 1492 34214 1532
rect 34256 1492 34296 1532
rect 19564 1324 19604 1364
rect 22156 1324 22196 1364
rect 23980 1324 24020 1364
rect 25612 1324 25652 1364
rect 30508 1324 30548 1364
rect 32140 1324 32180 1364
rect 35404 1324 35444 1364
rect 37036 1324 37076 1364
rect 38668 1324 38708 1364
rect 1612 1240 1652 1280
rect 4012 1240 4052 1280
rect 7756 1240 7796 1280
rect 14860 1240 14900 1280
rect 27244 1240 27284 1280
rect 28876 1240 28916 1280
rect 33772 1240 33812 1280
rect 41068 1240 41108 1280
rect 5548 1156 5588 1196
rect 10252 1156 10292 1196
rect 15532 1156 15572 1196
rect 40492 1156 40532 1196
rect 40876 1156 40916 1196
rect 41260 1156 41300 1196
rect 1324 1072 1364 1112
rect 1420 1072 1460 1112
rect 1612 1072 1652 1112
rect 1804 1072 1844 1112
rect 3052 1072 3092 1112
rect 3532 1072 3572 1112
rect 3724 1072 3764 1112
rect 3820 1072 3860 1112
rect 4300 1072 4340 1112
rect 4396 1072 4436 1112
rect 4684 1072 4724 1112
rect 5068 1072 5108 1112
rect 5164 1072 5204 1112
rect 5644 1072 5684 1112
rect 6124 1072 6164 1112
rect 6604 1077 6644 1117
rect 7084 1072 7124 1112
rect 7372 1072 7412 1112
rect 7948 1072 7988 1112
rect 9196 1072 9236 1112
rect 9676 1072 9716 1112
rect 9772 1072 9812 1112
rect 10156 1072 10196 1112
rect 10732 1072 10772 1112
rect 11212 1086 11252 1126
rect 11596 1072 11636 1112
rect 12844 1072 12884 1112
rect 14668 1072 14708 1112
rect 15052 1072 15092 1112
rect 7468 988 7508 1028
rect 9388 988 9428 1028
rect 11404 988 11444 1028
rect 13420 1030 13460 1070
rect 15148 1072 15188 1112
rect 18124 1072 18164 1112
rect 19372 1072 19412 1112
rect 20716 1072 20756 1112
rect 21964 1072 22004 1112
rect 22348 1072 22388 1112
rect 23596 1072 23636 1112
rect 24172 1072 24212 1112
rect 25804 1072 25844 1112
rect 27052 1072 27092 1112
rect 27436 1072 27476 1112
rect 28684 1072 28724 1112
rect 29068 1072 29108 1112
rect 30316 1072 30356 1112
rect 30700 1072 30740 1112
rect 31948 1072 31988 1112
rect 32332 1072 32372 1112
rect 33580 1072 33620 1112
rect 33964 1072 34004 1112
rect 35212 1072 35252 1112
rect 35596 1072 35636 1112
rect 36844 1072 36884 1112
rect 37228 1072 37268 1112
rect 38476 1072 38516 1112
rect 38860 1072 38900 1112
rect 40108 1072 40148 1112
rect 13036 988 13076 1028
rect 25420 1030 25460 1070
rect 23788 988 23828 1028
rect 3244 904 3284 944
rect 3532 904 3572 944
rect 6796 904 6836 944
rect 15340 904 15380 944
rect 15724 904 15764 944
rect 40300 904 40340 944
rect 41452 904 41492 944
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 35168 736 35208 776
rect 35250 736 35290 776
rect 35332 736 35372 776
rect 35414 736 35454 776
rect 35496 736 35536 776
<< metal2 >>
rect 2936 10688 3016 10752
rect 3148 10692 3476 10732
rect 3148 10688 3188 10692
rect 2936 10672 3188 10688
rect 2956 10648 3188 10672
rect 1419 10184 1461 10193
rect 1419 10144 1420 10184
rect 1460 10144 1461 10184
rect 1419 10135 1461 10144
rect 1420 9680 1460 10135
rect 2187 9680 2229 9689
rect 1420 9631 1460 9640
rect 1900 9640 2132 9680
rect 1707 9596 1749 9605
rect 1707 9556 1708 9596
rect 1748 9556 1749 9596
rect 1707 9547 1749 9556
rect 1419 9512 1461 9521
rect 1419 9472 1420 9512
rect 1460 9472 1461 9512
rect 1419 9463 1461 9472
rect 1516 9512 1556 9521
rect 1227 9176 1269 9185
rect 1227 9136 1228 9176
rect 1268 9136 1269 9176
rect 1227 9127 1269 9136
rect 1228 8765 1268 9127
rect 1420 8933 1460 9463
rect 1419 8924 1461 8933
rect 1419 8884 1420 8924
rect 1460 8884 1461 8924
rect 1419 8875 1461 8884
rect 1227 8756 1269 8765
rect 1227 8716 1228 8756
rect 1268 8716 1269 8756
rect 1227 8707 1269 8716
rect 1323 8672 1365 8681
rect 1323 8632 1324 8672
rect 1364 8632 1365 8672
rect 1323 8623 1365 8632
rect 1324 8538 1364 8623
rect 1420 8000 1460 8009
rect 1420 7169 1460 7960
rect 1516 7832 1556 9472
rect 1611 9512 1653 9521
rect 1611 9472 1612 9512
rect 1652 9472 1653 9512
rect 1611 9463 1653 9472
rect 1708 9512 1748 9547
rect 1612 9378 1652 9463
rect 1708 9461 1748 9472
rect 1900 9512 1940 9640
rect 1900 9463 1940 9472
rect 1996 9512 2036 9521
rect 1516 7792 1940 7832
rect 1611 7664 1653 7673
rect 1611 7624 1612 7664
rect 1652 7624 1653 7664
rect 1611 7615 1653 7624
rect 1324 7160 1364 7169
rect 1228 6992 1268 7001
rect 1132 6952 1228 6992
rect 1132 5648 1172 6952
rect 1228 6943 1268 6952
rect 1324 6917 1364 7120
rect 1419 7160 1461 7169
rect 1419 7120 1420 7160
rect 1460 7120 1461 7160
rect 1419 7111 1461 7120
rect 1516 7160 1556 7171
rect 1516 7085 1556 7120
rect 1515 7076 1557 7085
rect 1515 7036 1516 7076
rect 1556 7036 1557 7076
rect 1515 7027 1557 7036
rect 1323 6908 1365 6917
rect 1323 6868 1324 6908
rect 1364 6868 1365 6908
rect 1323 6859 1365 6868
rect 1228 6656 1268 6665
rect 1228 6236 1268 6616
rect 1515 6656 1557 6665
rect 1515 6616 1516 6656
rect 1556 6616 1557 6656
rect 1515 6607 1557 6616
rect 1420 6488 1460 6497
rect 1323 6236 1365 6245
rect 1228 6196 1324 6236
rect 1364 6196 1365 6236
rect 1323 6187 1365 6196
rect 1420 6068 1460 6448
rect 1324 6028 1460 6068
rect 1516 6488 1556 6607
rect 1324 5657 1364 6028
rect 1516 5984 1556 6448
rect 1420 5944 1556 5984
rect 1228 5648 1268 5657
rect 1132 5608 1228 5648
rect 1228 5599 1268 5608
rect 1323 5648 1365 5657
rect 1323 5608 1324 5648
rect 1364 5608 1365 5648
rect 1323 5599 1365 5608
rect 1420 5648 1460 5944
rect 1420 5599 1460 5608
rect 1515 5648 1557 5657
rect 1515 5608 1516 5648
rect 1556 5608 1557 5648
rect 1515 5599 1557 5608
rect 1516 5514 1556 5599
rect 1324 5480 1364 5489
rect 1324 5396 1364 5440
rect 1612 5396 1652 7615
rect 1803 7580 1845 7589
rect 1803 7540 1804 7580
rect 1844 7540 1845 7580
rect 1803 7531 1845 7540
rect 1804 7160 1844 7531
rect 1900 7244 1940 7792
rect 1996 7421 2036 9472
rect 2092 9428 2132 9640
rect 2187 9640 2188 9680
rect 2228 9640 2229 9680
rect 2187 9631 2229 9640
rect 2188 9546 2228 9631
rect 2475 9596 2517 9605
rect 2475 9556 2476 9596
rect 2516 9556 2517 9596
rect 2475 9547 2517 9556
rect 2380 9512 2420 9521
rect 2092 9388 2324 9428
rect 2187 7916 2229 7925
rect 2187 7876 2188 7916
rect 2228 7876 2229 7916
rect 2187 7867 2229 7876
rect 1995 7412 2037 7421
rect 1995 7372 1996 7412
rect 2036 7372 2037 7412
rect 1995 7363 2037 7372
rect 1900 7204 2132 7244
rect 1804 7120 1940 7160
rect 1707 6488 1749 6497
rect 1707 6448 1708 6488
rect 1748 6448 1749 6488
rect 1707 6439 1749 6448
rect 1708 6354 1748 6439
rect 1803 6320 1845 6329
rect 1803 6280 1804 6320
rect 1844 6280 1845 6320
rect 1803 6271 1845 6280
rect 1708 5648 1748 5657
rect 1804 5648 1844 6271
rect 1748 5608 1844 5648
rect 1708 5599 1748 5608
rect 1900 5489 1940 7120
rect 1995 6824 2037 6833
rect 1995 6784 1996 6824
rect 2036 6784 2037 6824
rect 1995 6775 2037 6784
rect 1899 5480 1941 5489
rect 1899 5440 1900 5480
rect 1940 5440 1941 5480
rect 1899 5431 1941 5440
rect 1324 5356 1652 5396
rect 1323 4976 1365 4985
rect 1323 4936 1324 4976
rect 1364 4936 1365 4976
rect 1323 4927 1365 4936
rect 1324 4842 1364 4927
rect 1996 4892 2036 6775
rect 1516 4852 2036 4892
rect 1323 4724 1365 4733
rect 1323 4684 1324 4724
rect 1364 4684 1365 4724
rect 1323 4675 1365 4684
rect 1228 3464 1268 3473
rect 1228 1205 1268 3424
rect 1324 3380 1364 4675
rect 1420 4136 1460 4145
rect 1420 3725 1460 4096
rect 1419 3716 1461 3725
rect 1419 3676 1420 3716
rect 1460 3676 1461 3716
rect 1419 3667 1461 3676
rect 1516 3548 1556 4852
rect 1707 4472 1749 4481
rect 1707 4432 1708 4472
rect 1748 4432 1749 4472
rect 1707 4423 1749 4432
rect 1611 3716 1653 3725
rect 1611 3676 1612 3716
rect 1652 3676 1653 3716
rect 1611 3667 1653 3676
rect 1420 3508 1556 3548
rect 1420 3485 1460 3508
rect 1420 3436 1460 3445
rect 1612 3464 1652 3667
rect 1324 3340 1455 3380
rect 1415 3296 1455 3340
rect 1515 3296 1557 3305
rect 1415 3256 1460 3296
rect 1324 3212 1364 3221
rect 1324 2801 1364 3172
rect 1323 2792 1365 2801
rect 1323 2752 1324 2792
rect 1364 2752 1365 2792
rect 1323 2743 1365 2752
rect 1323 2624 1365 2633
rect 1323 2584 1324 2624
rect 1364 2584 1365 2624
rect 1323 2575 1365 2584
rect 1420 2624 1460 3256
rect 1515 3256 1516 3296
rect 1556 3256 1557 3296
rect 1515 3247 1557 3256
rect 1420 2575 1460 2584
rect 1516 2624 1556 3247
rect 1612 3137 1652 3424
rect 1611 3128 1653 3137
rect 1611 3088 1612 3128
rect 1652 3088 1653 3128
rect 1611 3079 1653 3088
rect 1611 2960 1653 2969
rect 1611 2920 1612 2960
rect 1652 2920 1653 2960
rect 1611 2911 1653 2920
rect 1516 2575 1556 2584
rect 1612 2624 1652 2911
rect 1612 2575 1652 2584
rect 1324 2490 1364 2575
rect 1419 2288 1461 2297
rect 1419 2248 1420 2288
rect 1460 2248 1461 2288
rect 1419 2239 1461 2248
rect 1324 1952 1364 1961
rect 1324 1289 1364 1912
rect 1420 1952 1460 2239
rect 1515 2204 1557 2213
rect 1515 2164 1516 2204
rect 1556 2164 1557 2204
rect 1515 2155 1557 2164
rect 1420 1903 1460 1912
rect 1516 1952 1556 2155
rect 1516 1903 1556 1912
rect 1612 1952 1652 1961
rect 1708 1952 1748 4423
rect 1803 3968 1845 3977
rect 1803 3928 1804 3968
rect 1844 3928 1845 3968
rect 1803 3919 1845 3928
rect 1804 3305 1844 3919
rect 1899 3464 1941 3473
rect 1899 3424 1900 3464
rect 1940 3424 1941 3464
rect 1899 3415 1941 3424
rect 1803 3296 1845 3305
rect 1803 3256 1804 3296
rect 1844 3256 1845 3296
rect 1803 3247 1845 3256
rect 1803 2876 1845 2885
rect 1803 2836 1804 2876
rect 1844 2836 1845 2876
rect 1803 2827 1845 2836
rect 1804 2624 1844 2827
rect 1804 2575 1844 2584
rect 1804 1961 1844 2046
rect 1652 1912 1748 1952
rect 1803 1952 1845 1961
rect 1803 1912 1804 1952
rect 1844 1912 1845 1952
rect 1612 1903 1652 1912
rect 1803 1903 1845 1912
rect 1419 1784 1461 1793
rect 1419 1744 1420 1784
rect 1460 1744 1461 1784
rect 1419 1735 1461 1744
rect 1323 1280 1365 1289
rect 1323 1240 1324 1280
rect 1364 1240 1365 1280
rect 1323 1231 1365 1240
rect 1227 1196 1269 1205
rect 1227 1156 1228 1196
rect 1268 1156 1269 1196
rect 1227 1147 1269 1156
rect 1228 1028 1268 1147
rect 1324 1112 1364 1121
rect 1324 1028 1364 1072
rect 1420 1112 1460 1735
rect 1803 1700 1845 1709
rect 1803 1660 1804 1700
rect 1844 1660 1845 1700
rect 1803 1651 1845 1660
rect 1611 1532 1653 1541
rect 1611 1492 1612 1532
rect 1652 1492 1653 1532
rect 1611 1483 1653 1492
rect 1612 1280 1652 1483
rect 1612 1231 1652 1240
rect 1420 1063 1460 1072
rect 1612 1112 1652 1121
rect 1228 988 1364 1028
rect 1612 869 1652 1072
rect 1804 1112 1844 1651
rect 1900 1541 1940 3415
rect 1899 1532 1941 1541
rect 1899 1492 1900 1532
rect 1940 1492 1941 1532
rect 1899 1483 1941 1492
rect 1611 860 1653 869
rect 1611 820 1612 860
rect 1652 820 1653 860
rect 1611 811 1653 820
rect 1804 617 1844 1072
rect 2092 953 2132 7204
rect 2188 2297 2228 7867
rect 2284 6665 2324 9388
rect 2380 8681 2420 9472
rect 2379 8672 2421 8681
rect 2379 8632 2380 8672
rect 2420 8632 2421 8672
rect 2379 8623 2421 8632
rect 2476 7916 2516 9547
rect 2955 9512 2997 9521
rect 2955 9472 2956 9512
rect 2996 9472 2997 9512
rect 2955 9463 2997 9472
rect 3243 9512 3285 9521
rect 3243 9472 3244 9512
rect 3284 9472 3285 9512
rect 3243 9463 3285 9472
rect 2572 8672 2612 8681
rect 2612 8632 2708 8672
rect 2572 8623 2612 8632
rect 2668 8000 2708 8632
rect 2956 8588 2996 9463
rect 2956 8539 2996 8548
rect 3148 8677 3188 8686
rect 2764 8504 2804 8515
rect 2764 8429 2804 8464
rect 2859 8504 2901 8513
rect 2859 8464 2860 8504
rect 2900 8464 2901 8504
rect 2859 8455 2901 8464
rect 2763 8420 2805 8429
rect 2763 8380 2764 8420
rect 2804 8380 2805 8420
rect 2763 8371 2805 8380
rect 2860 8168 2900 8455
rect 3148 8429 3188 8637
rect 3147 8420 3189 8429
rect 3147 8380 3148 8420
rect 3188 8380 3189 8420
rect 3147 8371 3189 8380
rect 2860 8119 2900 8128
rect 3051 8168 3093 8177
rect 3051 8128 3052 8168
rect 3092 8128 3093 8168
rect 3051 8119 3093 8128
rect 2763 8000 2805 8009
rect 2708 7960 2764 8000
rect 2804 7960 2805 8000
rect 2668 7951 2708 7960
rect 2763 7951 2805 7960
rect 2476 7876 2612 7916
rect 2572 7832 2612 7876
rect 2572 7792 2708 7832
rect 2475 7160 2517 7169
rect 2475 7120 2476 7160
rect 2516 7120 2517 7160
rect 2475 7111 2517 7120
rect 2476 6749 2516 7111
rect 2475 6740 2517 6749
rect 2475 6700 2476 6740
rect 2516 6700 2517 6740
rect 2475 6691 2517 6700
rect 2283 6656 2325 6665
rect 2283 6616 2284 6656
rect 2324 6616 2325 6656
rect 2283 6607 2325 6616
rect 2283 6152 2325 6161
rect 2283 6112 2284 6152
rect 2324 6112 2325 6152
rect 2283 6103 2325 6112
rect 2187 2288 2229 2297
rect 2187 2248 2188 2288
rect 2228 2248 2229 2288
rect 2187 2239 2229 2248
rect 2284 1793 2324 6103
rect 2571 5732 2613 5741
rect 2571 5692 2572 5732
rect 2612 5692 2613 5732
rect 2571 5683 2613 5692
rect 2572 4976 2612 5683
rect 2572 4136 2612 4936
rect 2668 4556 2708 7792
rect 2764 7160 2804 7951
rect 3052 7925 3092 8119
rect 3051 7916 3093 7925
rect 3051 7876 3052 7916
rect 3092 7876 3093 7916
rect 3051 7867 3093 7876
rect 2956 7337 2996 7422
rect 2955 7328 2997 7337
rect 2955 7288 2956 7328
rect 2996 7288 2997 7328
rect 2955 7279 2997 7288
rect 3148 7160 3188 8371
rect 3244 8009 3284 9463
rect 3339 8168 3381 8177
rect 3339 8128 3340 8168
rect 3380 8128 3381 8168
rect 3339 8119 3381 8128
rect 3243 8000 3285 8009
rect 3243 7960 3244 8000
rect 3284 7960 3285 8000
rect 3243 7951 3285 7960
rect 3244 7866 3284 7951
rect 3243 7244 3285 7253
rect 3243 7204 3244 7244
rect 3284 7204 3285 7244
rect 3243 7195 3285 7204
rect 2804 7120 2996 7160
rect 2764 7111 2804 7120
rect 2859 6656 2901 6665
rect 2859 6616 2860 6656
rect 2900 6616 2901 6656
rect 2859 6607 2901 6616
rect 2860 4985 2900 6607
rect 2956 6488 2996 7120
rect 2956 5741 2996 6448
rect 3052 7120 3148 7160
rect 2955 5732 2997 5741
rect 2955 5692 2956 5732
rect 2996 5692 2997 5732
rect 2955 5683 2997 5692
rect 2956 5648 2996 5683
rect 2956 5598 2996 5608
rect 3052 5480 3092 7120
rect 3148 7111 3188 7120
rect 3244 7110 3284 7195
rect 3340 7160 3380 8119
rect 3340 7111 3380 7120
rect 3339 6992 3381 7001
rect 3339 6952 3340 6992
rect 3380 6952 3381 6992
rect 3339 6943 3381 6952
rect 3147 6656 3189 6665
rect 3147 6616 3148 6656
rect 3188 6616 3189 6656
rect 3147 6607 3189 6616
rect 3148 6522 3188 6607
rect 3243 6320 3285 6329
rect 3243 6280 3244 6320
rect 3284 6280 3285 6320
rect 3243 6271 3285 6280
rect 3147 5984 3189 5993
rect 3147 5944 3148 5984
rect 3188 5944 3189 5984
rect 3147 5935 3189 5944
rect 3148 5900 3188 5935
rect 3148 5849 3188 5860
rect 2956 5440 3092 5480
rect 3148 5480 3188 5489
rect 2859 4976 2901 4985
rect 2859 4936 2860 4976
rect 2900 4936 2901 4976
rect 2859 4927 2901 4936
rect 2763 4808 2805 4817
rect 2763 4768 2764 4808
rect 2804 4768 2805 4808
rect 2763 4759 2805 4768
rect 2764 4674 2804 4759
rect 2668 4516 2804 4556
rect 2668 4136 2708 4145
rect 2572 4096 2668 4136
rect 2668 3725 2708 4096
rect 2667 3716 2709 3725
rect 2667 3676 2668 3716
rect 2708 3676 2709 3716
rect 2667 3667 2709 3676
rect 2668 3557 2708 3667
rect 2667 3548 2709 3557
rect 2667 3508 2668 3548
rect 2708 3508 2709 3548
rect 2667 3499 2709 3508
rect 2764 3305 2804 4516
rect 2956 4481 2996 5440
rect 3148 5396 3188 5440
rect 3052 5356 3188 5396
rect 3052 4976 3092 5356
rect 3244 5144 3284 6271
rect 3340 5993 3380 6943
rect 3436 6581 3476 10692
rect 4088 10672 4168 10752
rect 5240 10672 5320 10752
rect 6392 10672 6472 10752
rect 7544 10672 7624 10752
rect 7756 10692 8276 10732
rect 3819 9596 3861 9605
rect 3819 9556 3820 9596
rect 3860 9556 3861 9596
rect 3819 9547 3861 9556
rect 3627 9512 3669 9521
rect 3627 9472 3628 9512
rect 3668 9472 3669 9512
rect 3627 9463 3669 9472
rect 3628 9378 3668 9463
rect 3820 9462 3860 9547
rect 3688 9092 4056 9101
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 3688 9043 4056 9052
rect 4011 8840 4053 8849
rect 4108 8840 4148 10672
rect 5260 10016 5300 10672
rect 5643 10100 5685 10109
rect 5643 10060 5644 10100
rect 5684 10060 5685 10100
rect 5643 10051 5685 10060
rect 5260 9976 5588 10016
rect 4928 9848 5296 9857
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 4928 9799 5296 9808
rect 4491 9680 4533 9689
rect 4491 9640 4492 9680
rect 4532 9640 4533 9680
rect 4491 9631 4533 9640
rect 4295 9512 4335 9521
rect 4396 9512 4436 9521
rect 4335 9472 4340 9512
rect 4295 9463 4340 9472
rect 4203 9176 4245 9185
rect 4203 9136 4204 9176
rect 4244 9136 4245 9176
rect 4203 9127 4245 9136
rect 4204 8849 4244 9127
rect 4011 8800 4012 8840
rect 4052 8800 4148 8840
rect 4203 8840 4245 8849
rect 4203 8800 4204 8840
rect 4244 8800 4245 8840
rect 4011 8791 4053 8800
rect 4203 8791 4245 8800
rect 3628 8672 3668 8681
rect 3628 8429 3668 8632
rect 4108 8672 4148 8681
rect 4204 8672 4244 8681
rect 3627 8420 3669 8429
rect 3627 8380 3628 8420
rect 3668 8380 3669 8420
rect 3627 8371 3669 8380
rect 4108 8345 4148 8632
rect 4196 8632 4204 8672
rect 4196 8623 4244 8632
rect 4196 8504 4236 8623
rect 4196 8464 4244 8504
rect 4107 8336 4149 8345
rect 4107 8296 4108 8336
rect 4148 8296 4149 8336
rect 4107 8287 4149 8296
rect 3688 7580 4056 7589
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 3688 7531 4056 7540
rect 3531 7412 3573 7421
rect 3531 7372 3532 7412
rect 3572 7372 3573 7412
rect 3531 7363 3573 7372
rect 3532 7278 3572 7363
rect 3915 7160 3957 7169
rect 3915 7120 3916 7160
rect 3956 7120 3957 7160
rect 3915 7111 3957 7120
rect 3820 7076 3860 7085
rect 3820 6917 3860 7036
rect 3916 7026 3956 7111
rect 3819 6908 3861 6917
rect 3819 6868 3820 6908
rect 3860 6868 3861 6908
rect 3819 6859 3861 6868
rect 3435 6572 3477 6581
rect 3435 6532 3436 6572
rect 3476 6532 3477 6572
rect 3435 6523 3477 6532
rect 3820 6488 3860 6497
rect 3820 6404 3860 6448
rect 3915 6488 3957 6497
rect 3915 6448 3916 6488
rect 3956 6448 3957 6488
rect 3915 6439 3957 6448
rect 3436 6364 3860 6404
rect 3339 5984 3381 5993
rect 3339 5944 3340 5984
rect 3380 5944 3381 5984
rect 3339 5935 3381 5944
rect 3339 5816 3381 5825
rect 3339 5776 3340 5816
rect 3380 5776 3381 5816
rect 3339 5767 3381 5776
rect 3340 5648 3380 5767
rect 3436 5732 3476 6364
rect 3916 6354 3956 6439
rect 3532 6236 3572 6245
rect 3532 5816 3572 6196
rect 3688 6068 4056 6077
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 3688 6019 4056 6028
rect 4108 5900 4148 8287
rect 4204 7841 4244 8464
rect 4203 7832 4245 7841
rect 4203 7792 4204 7832
rect 4244 7792 4245 7832
rect 4203 7783 4245 7792
rect 4203 7328 4245 7337
rect 4203 7288 4204 7328
rect 4244 7288 4245 7328
rect 4203 7279 4245 7288
rect 4204 7160 4244 7279
rect 4204 6497 4244 7120
rect 4203 6488 4245 6497
rect 4203 6448 4204 6488
rect 4244 6448 4245 6488
rect 4203 6439 4245 6448
rect 3916 5860 4148 5900
rect 3724 5816 3764 5825
rect 3532 5776 3668 5816
rect 3436 5692 3572 5732
rect 3340 5599 3380 5608
rect 3532 5648 3572 5692
rect 3532 5573 3572 5608
rect 3436 5564 3476 5573
rect 3436 5153 3476 5524
rect 3531 5564 3573 5573
rect 3531 5524 3532 5564
rect 3572 5524 3573 5564
rect 3531 5515 3573 5524
rect 3531 5396 3573 5405
rect 3531 5356 3532 5396
rect 3572 5356 3573 5396
rect 3531 5347 3573 5356
rect 3532 5186 3572 5347
rect 3148 5104 3284 5144
rect 3435 5144 3477 5153
rect 3435 5104 3436 5144
rect 3476 5104 3477 5144
rect 3532 5137 3572 5146
rect 3148 5060 3188 5104
rect 3435 5095 3477 5104
rect 3148 5011 3188 5020
rect 3052 4927 3092 4936
rect 3243 4976 3285 4985
rect 3243 4936 3244 4976
rect 3284 4936 3285 4976
rect 3243 4927 3285 4936
rect 3340 4976 3380 4985
rect 3628 4976 3668 5776
rect 3724 5657 3764 5776
rect 3916 5657 3956 5860
rect 3723 5648 3765 5657
rect 3723 5608 3724 5648
rect 3764 5608 3765 5648
rect 3723 5599 3765 5608
rect 3915 5648 3957 5657
rect 3915 5608 3916 5648
rect 3956 5608 3957 5648
rect 3915 5599 3957 5608
rect 4108 5648 4148 5657
rect 3819 5060 3861 5069
rect 3819 5020 3820 5060
rect 3860 5020 3861 5060
rect 3819 5011 3861 5020
rect 3380 4936 3668 4976
rect 3340 4927 3380 4936
rect 3244 4842 3284 4927
rect 3820 4926 3860 5011
rect 3916 4976 3956 5599
rect 4011 5564 4053 5573
rect 4011 5524 4012 5564
rect 4052 5524 4053 5564
rect 4011 5515 4053 5524
rect 4012 5430 4052 5515
rect 4011 5060 4053 5069
rect 4011 5020 4012 5060
rect 4052 5020 4053 5060
rect 4011 5011 4053 5020
rect 3916 4733 3956 4936
rect 4012 4808 4052 5011
rect 4108 4985 4148 5608
rect 4204 5648 4244 6439
rect 4300 6329 4340 9463
rect 4299 6320 4341 6329
rect 4299 6280 4300 6320
rect 4340 6280 4341 6320
rect 4299 6271 4341 6280
rect 4396 6245 4436 9472
rect 4492 9512 4532 9631
rect 4492 9463 4532 9472
rect 4684 9512 4724 9521
rect 4684 8840 4724 9472
rect 4780 9512 4820 9523
rect 4780 9437 4820 9472
rect 4972 9512 5012 9521
rect 4779 9428 4821 9437
rect 4779 9388 4780 9428
rect 4820 9388 4821 9428
rect 4779 9379 4821 9388
rect 4779 9260 4821 9269
rect 4779 9220 4780 9260
rect 4820 9220 4821 9260
rect 4779 9211 4821 9220
rect 4780 9126 4820 9211
rect 4684 8800 4820 8840
rect 4588 8672 4628 8681
rect 4491 8000 4533 8009
rect 4491 7960 4492 8000
rect 4532 7960 4533 8000
rect 4491 7951 4533 7960
rect 4492 7866 4532 7951
rect 4588 7925 4628 8632
rect 4684 8672 4724 8681
rect 4684 8177 4724 8632
rect 4683 8168 4725 8177
rect 4683 8128 4684 8168
rect 4724 8128 4725 8168
rect 4683 8119 4725 8128
rect 4587 7916 4629 7925
rect 4587 7876 4588 7916
rect 4628 7876 4629 7916
rect 4587 7867 4629 7876
rect 4780 7673 4820 8800
rect 4972 8513 5012 9472
rect 5451 9512 5493 9521
rect 5451 9472 5452 9512
rect 5492 9472 5493 9512
rect 5451 9463 5493 9472
rect 5067 9428 5109 9437
rect 5067 9388 5068 9428
rect 5108 9388 5109 9428
rect 5067 9379 5109 9388
rect 5068 9260 5108 9379
rect 5259 9344 5301 9353
rect 5259 9304 5260 9344
rect 5300 9304 5301 9344
rect 5259 9295 5301 9304
rect 5068 9092 5108 9220
rect 5260 9210 5300 9295
rect 5355 9260 5397 9269
rect 5355 9220 5356 9260
rect 5396 9220 5397 9260
rect 5355 9211 5397 9220
rect 5068 9052 5300 9092
rect 5260 8672 5300 9052
rect 5260 8623 5300 8632
rect 5356 8672 5396 9211
rect 5452 9101 5492 9463
rect 5451 9092 5493 9101
rect 5451 9052 5452 9092
rect 5492 9052 5493 9092
rect 5451 9043 5493 9052
rect 5356 8623 5396 8632
rect 5164 8513 5204 8595
rect 4971 8504 5013 8513
rect 4971 8464 4972 8504
rect 5012 8464 5013 8504
rect 4971 8455 5013 8464
rect 5163 8504 5205 8513
rect 5163 8460 5164 8504
rect 5204 8460 5205 8504
rect 5163 8455 5205 8460
rect 5164 8451 5204 8455
rect 4928 8336 5296 8345
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 4928 8287 5296 8296
rect 4972 8000 5012 8009
rect 4779 7664 4821 7673
rect 4779 7624 4780 7664
rect 4820 7624 4821 7664
rect 4779 7615 4821 7624
rect 4972 7337 5012 7960
rect 5260 8000 5300 8011
rect 5260 7925 5300 7960
rect 5356 8000 5396 8009
rect 5259 7916 5301 7925
rect 5259 7876 5260 7916
rect 5300 7876 5301 7916
rect 5259 7867 5301 7876
rect 5356 7841 5396 7960
rect 5355 7832 5397 7841
rect 5355 7792 5356 7832
rect 5396 7792 5397 7832
rect 5355 7783 5397 7792
rect 5548 7496 5588 9976
rect 5644 8924 5684 10051
rect 5835 9008 5877 9017
rect 5835 8968 5836 9008
rect 5876 8968 5877 9008
rect 5835 8959 5877 8968
rect 5644 8875 5684 8884
rect 5836 8000 5876 8959
rect 6123 8672 6165 8681
rect 6123 8632 6124 8672
rect 6164 8632 6165 8672
rect 6123 8623 6165 8632
rect 6124 8538 6164 8623
rect 5836 7951 5876 7960
rect 5644 7748 5684 7757
rect 5684 7708 6068 7748
rect 5644 7699 5684 7708
rect 5548 7456 5972 7496
rect 4971 7328 5013 7337
rect 4971 7288 4972 7328
rect 5012 7288 5013 7328
rect 4971 7279 5013 7288
rect 5452 7288 5684 7328
rect 4491 7244 4533 7253
rect 4491 7204 4492 7244
rect 4532 7204 4533 7244
rect 4491 7195 4533 7204
rect 5452 7244 5492 7288
rect 5452 7195 5492 7204
rect 4492 7160 4532 7195
rect 4492 7109 4532 7120
rect 4684 7160 4724 7169
rect 4587 7076 4629 7085
rect 4587 7036 4588 7076
rect 4628 7036 4629 7076
rect 4587 7027 4629 7036
rect 4588 6942 4628 7027
rect 4684 6917 4724 7120
rect 4972 7160 5012 7169
rect 4779 7076 4821 7085
rect 4779 7036 4780 7076
rect 4820 7036 4821 7076
rect 4779 7027 4821 7036
rect 4683 6908 4725 6917
rect 4683 6868 4684 6908
rect 4724 6868 4725 6908
rect 4683 6859 4725 6868
rect 4780 6656 4820 7027
rect 4972 7001 5012 7120
rect 5068 7160 5108 7169
rect 5548 7160 5588 7169
rect 5108 7120 5396 7160
rect 5068 7111 5108 7120
rect 4971 6992 5013 7001
rect 4971 6952 4972 6992
rect 5012 6952 5013 6992
rect 4971 6943 5013 6952
rect 4928 6824 5296 6833
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 4928 6775 5296 6784
rect 4780 6616 5012 6656
rect 4972 6572 5012 6616
rect 4972 6523 5012 6532
rect 4587 6488 4629 6497
rect 4587 6448 4588 6488
rect 4628 6448 4629 6488
rect 4587 6439 4629 6448
rect 4876 6488 4916 6497
rect 4588 6354 4628 6439
rect 4876 6329 4916 6448
rect 5163 6488 5205 6497
rect 5163 6448 5164 6488
rect 5204 6448 5205 6488
rect 5163 6439 5205 6448
rect 4875 6320 4917 6329
rect 4875 6280 4876 6320
rect 4916 6280 4917 6320
rect 4875 6271 4917 6280
rect 4395 6236 4437 6245
rect 4395 6196 4396 6236
rect 4436 6196 4437 6236
rect 4395 6187 4437 6196
rect 4684 5825 4724 5910
rect 4683 5816 4725 5825
rect 4683 5776 4684 5816
rect 4724 5776 4725 5816
rect 4683 5767 4725 5776
rect 4396 5648 4436 5657
rect 4684 5648 4724 5657
rect 4876 5648 4916 5657
rect 4204 5608 4396 5648
rect 4107 4976 4149 4985
rect 4107 4936 4108 4976
rect 4148 4936 4149 4976
rect 4107 4927 4149 4936
rect 4204 4976 4244 5608
rect 4396 5599 4436 5608
rect 4492 5608 4684 5648
rect 4204 4927 4244 4936
rect 4012 4768 4148 4808
rect 3915 4724 3957 4733
rect 3915 4684 3916 4724
rect 3956 4684 3957 4724
rect 3915 4675 3957 4684
rect 3688 4556 4056 4565
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 3688 4507 4056 4516
rect 2955 4472 2997 4481
rect 2955 4432 2956 4472
rect 2996 4432 2997 4472
rect 2955 4423 2997 4432
rect 4108 4388 4148 4768
rect 4299 4724 4341 4733
rect 4299 4684 4300 4724
rect 4340 4684 4341 4724
rect 4299 4675 4341 4684
rect 4203 4388 4245 4397
rect 4108 4348 4204 4388
rect 4244 4348 4245 4388
rect 4203 4339 4245 4348
rect 3723 4304 3765 4313
rect 3723 4264 3724 4304
rect 3764 4264 3765 4304
rect 3723 4255 3765 4264
rect 2955 4220 2997 4229
rect 2955 4180 2956 4220
rect 2996 4180 2997 4220
rect 2955 4171 2997 4180
rect 3243 4220 3285 4229
rect 3243 4180 3244 4220
rect 3284 4180 3285 4220
rect 3243 4171 3285 4180
rect 2860 3968 2900 3977
rect 2860 3809 2900 3928
rect 2859 3800 2901 3809
rect 2859 3760 2860 3800
rect 2900 3760 2901 3800
rect 2859 3751 2901 3760
rect 2956 3632 2996 4171
rect 3244 4150 3284 4171
rect 3244 4085 3284 4110
rect 3724 4136 3764 4255
rect 4204 4220 4244 4339
rect 4204 4171 4244 4180
rect 4300 4220 4340 4675
rect 4492 4229 4532 5608
rect 4684 5599 4724 5608
rect 4780 5608 4876 5648
rect 4683 5480 4725 5489
rect 4683 5440 4684 5480
rect 4724 5440 4725 5480
rect 4683 5431 4725 5440
rect 4587 4976 4629 4985
rect 4587 4936 4588 4976
rect 4628 4936 4629 4976
rect 4587 4927 4629 4936
rect 4684 4976 4724 5431
rect 4780 5144 4820 5608
rect 4876 5599 4916 5608
rect 5164 5648 5204 6439
rect 5260 6320 5300 6329
rect 5356 6320 5396 7120
rect 5300 6280 5396 6320
rect 5452 6320 5492 6329
rect 5548 6320 5588 7120
rect 5492 6280 5588 6320
rect 5260 6271 5300 6280
rect 5452 6271 5492 6280
rect 5644 5900 5684 7288
rect 5739 6572 5781 6581
rect 5739 6532 5740 6572
rect 5780 6532 5781 6572
rect 5739 6523 5781 6532
rect 5740 6438 5780 6523
rect 5835 6488 5877 6497
rect 5835 6448 5836 6488
rect 5876 6448 5877 6488
rect 5835 6439 5877 6448
rect 5836 6354 5876 6439
rect 5836 5900 5876 5909
rect 5644 5860 5836 5900
rect 5836 5851 5876 5860
rect 5451 5816 5493 5825
rect 5451 5776 5452 5816
rect 5492 5776 5493 5816
rect 5451 5767 5493 5776
rect 5164 5599 5204 5608
rect 5452 5648 5492 5767
rect 5452 5599 5492 5608
rect 5355 5564 5397 5573
rect 5355 5524 5356 5564
rect 5396 5524 5397 5564
rect 5355 5515 5397 5524
rect 5548 5564 5588 5573
rect 4928 5312 5296 5321
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 4928 5263 5296 5272
rect 4780 5104 5012 5144
rect 4684 4927 4724 4936
rect 4780 4976 4820 4985
rect 4588 4842 4628 4927
rect 4780 4733 4820 4936
rect 4875 4976 4917 4985
rect 4875 4936 4876 4976
rect 4916 4936 4917 4976
rect 4875 4927 4917 4936
rect 4876 4842 4916 4927
rect 4972 4817 5012 5104
rect 5067 4976 5109 4985
rect 5067 4936 5068 4976
rect 5108 4936 5109 4976
rect 5067 4927 5109 4936
rect 5068 4842 5108 4927
rect 4971 4808 5013 4817
rect 4971 4768 4972 4808
rect 5012 4768 5013 4808
rect 4971 4759 5013 4768
rect 4779 4724 4821 4733
rect 4779 4684 4780 4724
rect 4820 4684 4821 4724
rect 4779 4675 4821 4684
rect 4300 4171 4340 4180
rect 4491 4220 4533 4229
rect 4491 4180 4492 4220
rect 4532 4180 4533 4220
rect 4491 4171 4533 4180
rect 4683 4220 4725 4229
rect 4683 4180 4684 4220
rect 4724 4180 4725 4220
rect 4683 4171 4725 4180
rect 3724 4087 3764 4096
rect 4684 4136 4724 4171
rect 4684 4061 4724 4096
rect 4780 4136 4820 4145
rect 4972 4136 5012 4759
rect 5356 4649 5396 5515
rect 5451 5144 5493 5153
rect 5451 5104 5452 5144
rect 5492 5104 5493 5144
rect 5451 5095 5493 5104
rect 5067 4640 5109 4649
rect 5067 4600 5068 4640
rect 5108 4600 5109 4640
rect 5067 4591 5109 4600
rect 5355 4640 5397 4649
rect 5355 4600 5356 4640
rect 5396 4600 5397 4640
rect 5355 4591 5397 4600
rect 4820 4096 5012 4136
rect 5068 4136 5108 4591
rect 5355 4220 5397 4229
rect 5355 4180 5356 4220
rect 5396 4180 5397 4220
rect 5355 4171 5397 4180
rect 4780 4087 4820 4096
rect 5068 4087 5108 4096
rect 5164 4136 5204 4145
rect 5259 4136 5301 4145
rect 5204 4096 5260 4136
rect 5300 4096 5301 4136
rect 5164 4087 5204 4096
rect 5259 4087 5301 4096
rect 5356 4136 5396 4171
rect 5356 4085 5396 4096
rect 4683 4052 4725 4061
rect 4683 4012 4684 4052
rect 4724 4012 4725 4052
rect 4683 4003 4725 4012
rect 3052 3968 3092 3977
rect 3531 3968 3573 3977
rect 4684 3972 4724 4003
rect 3092 3928 3380 3968
rect 3052 3919 3092 3928
rect 3243 3800 3285 3809
rect 3243 3760 3244 3800
rect 3284 3760 3285 3800
rect 3243 3751 3285 3760
rect 3052 3632 3092 3641
rect 2956 3592 3052 3632
rect 2859 3548 2901 3557
rect 2859 3508 2860 3548
rect 2900 3508 2901 3548
rect 2859 3499 2901 3508
rect 2860 3464 2900 3499
rect 2763 3296 2805 3305
rect 2763 3256 2764 3296
rect 2804 3256 2805 3296
rect 2763 3247 2805 3256
rect 2860 2624 2900 3424
rect 2956 2969 2996 3592
rect 3052 3583 3092 3592
rect 3244 3464 3284 3751
rect 3147 3212 3189 3221
rect 3147 3172 3148 3212
rect 3188 3172 3189 3212
rect 3147 3163 3189 3172
rect 2955 2960 2997 2969
rect 2955 2920 2956 2960
rect 2996 2920 2997 2960
rect 2955 2911 2997 2920
rect 3148 2801 3188 3163
rect 3147 2792 3189 2801
rect 3147 2752 3148 2792
rect 3188 2752 3189 2792
rect 3147 2743 3189 2752
rect 3052 2624 3092 2633
rect 2860 2584 3052 2624
rect 3052 1952 3092 2584
rect 3148 2120 3188 2743
rect 3244 2717 3284 3424
rect 3340 3464 3380 3928
rect 3531 3928 3532 3968
rect 3572 3928 3573 3968
rect 3531 3919 3573 3928
rect 3532 3632 3572 3919
rect 4491 3884 4533 3893
rect 4491 3844 4492 3884
rect 4532 3844 4533 3884
rect 4491 3835 4533 3844
rect 3532 3583 3572 3592
rect 4204 3632 4244 3641
rect 4244 3592 4340 3632
rect 4204 3583 4244 3592
rect 3340 3415 3380 3424
rect 3436 3464 3476 3475
rect 3436 3389 3476 3424
rect 3724 3464 3764 3473
rect 3435 3380 3477 3389
rect 3435 3340 3436 3380
rect 3476 3340 3477 3380
rect 3435 3331 3477 3340
rect 3531 3296 3573 3305
rect 3531 3256 3532 3296
rect 3572 3256 3573 3296
rect 3531 3247 3573 3256
rect 3243 2708 3285 2717
rect 3243 2668 3244 2708
rect 3284 2668 3285 2708
rect 3243 2659 3285 2668
rect 3436 2624 3476 2633
rect 3339 2540 3381 2549
rect 3436 2540 3476 2584
rect 3339 2500 3340 2540
rect 3380 2500 3476 2540
rect 3339 2491 3381 2500
rect 3244 2456 3284 2465
rect 3244 2297 3284 2416
rect 3243 2288 3285 2297
rect 3243 2248 3244 2288
rect 3284 2248 3285 2288
rect 3243 2239 3285 2248
rect 3244 2120 3284 2129
rect 3148 2080 3244 2120
rect 3244 2071 3284 2080
rect 2283 1784 2325 1793
rect 2283 1744 2284 1784
rect 2324 1744 2325 1784
rect 2283 1735 2325 1744
rect 3052 1112 3092 1912
rect 3340 1457 3380 2491
rect 3436 1952 3476 1961
rect 3339 1448 3381 1457
rect 3339 1408 3340 1448
rect 3380 1408 3381 1448
rect 3339 1399 3381 1408
rect 3436 1121 3476 1912
rect 3052 1063 3092 1072
rect 3435 1112 3477 1121
rect 3435 1072 3436 1112
rect 3476 1072 3477 1112
rect 3435 1063 3477 1072
rect 3532 1112 3572 3247
rect 3724 3221 3764 3424
rect 3819 3464 3861 3473
rect 3819 3424 3820 3464
rect 3860 3424 3861 3464
rect 3819 3415 3861 3424
rect 4011 3464 4053 3473
rect 4011 3424 4012 3464
rect 4052 3424 4053 3464
rect 4011 3415 4053 3424
rect 4108 3464 4148 3473
rect 4209 3464 4249 3473
rect 3820 3330 3860 3415
rect 4012 3330 4052 3415
rect 3723 3212 3765 3221
rect 3723 3172 3724 3212
rect 3764 3172 3765 3212
rect 3723 3163 3765 3172
rect 3688 3044 4056 3053
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 3688 2995 4056 3004
rect 4108 1709 4148 3424
rect 4204 3424 4209 3464
rect 4204 3415 4249 3424
rect 4107 1700 4149 1709
rect 4107 1660 4108 1700
rect 4148 1660 4149 1700
rect 4107 1651 4149 1660
rect 3688 1532 4056 1541
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 3688 1483 4056 1492
rect 3723 1280 3765 1289
rect 3723 1240 3724 1280
rect 3764 1240 3765 1280
rect 3723 1231 3765 1240
rect 4012 1280 4052 1289
rect 4204 1280 4244 3415
rect 4300 2381 4340 3592
rect 4492 3464 4532 3835
rect 4928 3800 5296 3809
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 4928 3751 5296 3760
rect 4683 3716 4725 3725
rect 4683 3676 4684 3716
rect 4724 3676 4725 3716
rect 4683 3667 4725 3676
rect 4492 2969 4532 3424
rect 4491 2960 4533 2969
rect 4491 2920 4492 2960
rect 4532 2920 4533 2960
rect 4491 2911 4533 2920
rect 4684 2624 4724 3667
rect 5067 3380 5109 3389
rect 5067 3340 5068 3380
rect 5108 3340 5109 3380
rect 5067 3331 5109 3340
rect 5068 2876 5108 3331
rect 5068 2827 5108 2836
rect 4971 2708 5013 2717
rect 4971 2668 4972 2708
rect 5012 2668 5108 2708
rect 4971 2659 5013 2668
rect 4299 2372 4341 2381
rect 4299 2332 4300 2372
rect 4340 2332 4341 2372
rect 4299 2323 4341 2332
rect 4684 1952 4724 2584
rect 5068 2624 5108 2668
rect 5260 2633 5300 2718
rect 5068 2575 5108 2584
rect 5259 2624 5301 2633
rect 5259 2584 5260 2624
rect 5300 2584 5301 2624
rect 5259 2575 5301 2584
rect 5356 2624 5396 2633
rect 5452 2624 5492 5095
rect 5548 4985 5588 5524
rect 5547 4976 5589 4985
rect 5547 4936 5548 4976
rect 5588 4936 5589 4976
rect 5547 4927 5589 4936
rect 5547 4136 5589 4145
rect 5547 4096 5548 4136
rect 5588 4096 5589 4136
rect 5547 4087 5589 4096
rect 5644 4136 5684 4145
rect 5548 4002 5588 4087
rect 5547 3800 5589 3809
rect 5547 3760 5548 3800
rect 5588 3760 5589 3800
rect 5547 3751 5589 3760
rect 5548 3128 5588 3751
rect 5644 3305 5684 4096
rect 5740 4136 5780 4145
rect 5740 3884 5780 4096
rect 5835 4136 5877 4145
rect 5835 4096 5836 4136
rect 5876 4096 5877 4136
rect 5835 4087 5877 4096
rect 5836 4002 5876 4087
rect 5932 3977 5972 7456
rect 6028 7160 6068 7708
rect 6412 7673 6452 10672
rect 7564 10604 7604 10672
rect 7756 10604 7796 10692
rect 7564 10564 7796 10604
rect 7468 9680 7508 9689
rect 6700 9512 6740 9521
rect 6700 9437 6740 9472
rect 6988 9512 7028 9521
rect 6699 9428 6741 9437
rect 6699 9388 6700 9428
rect 6740 9388 6741 9428
rect 6699 9379 6741 9388
rect 6700 8681 6740 9379
rect 6892 9260 6932 9269
rect 6699 8672 6741 8681
rect 6699 8632 6700 8672
rect 6740 8632 6741 8672
rect 6699 8623 6741 8632
rect 6699 8504 6741 8513
rect 6699 8464 6700 8504
rect 6740 8464 6741 8504
rect 6699 8455 6741 8464
rect 6411 7664 6453 7673
rect 6411 7624 6412 7664
rect 6452 7624 6453 7664
rect 6411 7615 6453 7624
rect 6028 7111 6068 7120
rect 6508 7165 6548 7174
rect 6027 6992 6069 7001
rect 6027 6952 6028 6992
rect 6068 6952 6069 6992
rect 6027 6943 6069 6952
rect 6028 6329 6068 6943
rect 6508 6665 6548 7125
rect 6700 7076 6740 8455
rect 6795 7580 6837 7589
rect 6795 7540 6796 7580
rect 6836 7540 6837 7580
rect 6795 7531 6837 7540
rect 6700 7027 6740 7036
rect 6507 6656 6549 6665
rect 6507 6616 6508 6656
rect 6548 6616 6549 6656
rect 6507 6607 6549 6616
rect 6700 6656 6740 6665
rect 6796 6656 6836 7531
rect 6740 6616 6836 6656
rect 6700 6607 6740 6616
rect 6124 6488 6164 6499
rect 6124 6413 6164 6448
rect 6508 6488 6548 6497
rect 6123 6404 6165 6413
rect 6123 6364 6124 6404
rect 6164 6364 6165 6404
rect 6123 6355 6165 6364
rect 6411 6404 6453 6413
rect 6411 6364 6412 6404
rect 6452 6364 6453 6404
rect 6411 6355 6453 6364
rect 6027 6320 6069 6329
rect 6027 6280 6028 6320
rect 6068 6280 6069 6320
rect 6027 6271 6069 6280
rect 6028 5816 6068 6271
rect 6315 5816 6357 5825
rect 6028 5776 6260 5816
rect 5931 3968 5973 3977
rect 5931 3928 5932 3968
rect 5972 3928 5973 3968
rect 5931 3919 5973 3928
rect 5740 3844 5876 3884
rect 5739 3716 5781 3725
rect 5739 3676 5740 3716
rect 5780 3676 5781 3716
rect 5739 3667 5781 3676
rect 5740 3464 5780 3667
rect 5740 3415 5780 3424
rect 5643 3296 5685 3305
rect 5643 3256 5644 3296
rect 5684 3256 5685 3296
rect 5643 3247 5685 3256
rect 5836 3137 5876 3844
rect 6028 3809 6068 5776
rect 6124 5648 6164 5657
rect 6124 4229 6164 5608
rect 6220 5648 6260 5776
rect 6315 5776 6316 5816
rect 6356 5776 6357 5816
rect 6315 5767 6357 5776
rect 6220 5599 6260 5608
rect 6316 5144 6356 5767
rect 6220 5104 6356 5144
rect 6123 4220 6165 4229
rect 6123 4180 6124 4220
rect 6164 4180 6165 4220
rect 6123 4171 6165 4180
rect 6124 4136 6164 4171
rect 6027 3800 6069 3809
rect 6027 3760 6028 3800
rect 6068 3760 6069 3800
rect 6027 3751 6069 3760
rect 5932 3632 5972 3641
rect 6124 3632 6164 4096
rect 5972 3592 6164 3632
rect 6220 4136 6260 5104
rect 6316 4976 6356 4985
rect 6316 4556 6356 4936
rect 6412 4733 6452 6355
rect 6508 6329 6548 6448
rect 6604 6488 6644 6497
rect 6507 6320 6549 6329
rect 6507 6280 6508 6320
rect 6548 6280 6549 6320
rect 6507 6271 6549 6280
rect 6508 5489 6548 6271
rect 6604 6161 6644 6448
rect 6699 6488 6741 6497
rect 6699 6448 6700 6488
rect 6740 6448 6741 6488
rect 6699 6439 6741 6448
rect 6796 6488 6836 6499
rect 6603 6152 6645 6161
rect 6603 6112 6604 6152
rect 6644 6112 6645 6152
rect 6603 6103 6645 6112
rect 6603 5900 6645 5909
rect 6603 5860 6604 5900
rect 6644 5860 6645 5900
rect 6603 5851 6645 5860
rect 6604 5732 6644 5851
rect 6507 5480 6549 5489
rect 6507 5440 6508 5480
rect 6548 5440 6549 5480
rect 6507 5431 6549 5440
rect 6507 5312 6549 5321
rect 6507 5272 6508 5312
rect 6548 5272 6549 5312
rect 6507 5263 6549 5272
rect 6508 5144 6548 5263
rect 6508 5095 6548 5104
rect 6604 4892 6644 5692
rect 6508 4852 6644 4892
rect 6700 5648 6740 6439
rect 6796 6413 6836 6448
rect 6795 6404 6837 6413
rect 6795 6364 6796 6404
rect 6836 6364 6837 6404
rect 6795 6355 6837 6364
rect 6892 6161 6932 9220
rect 6988 8513 7028 9472
rect 7180 9512 7220 9521
rect 7180 9353 7220 9472
rect 7276 9512 7316 9521
rect 7179 9344 7221 9353
rect 7179 9304 7180 9344
rect 7220 9304 7221 9344
rect 7179 9295 7221 9304
rect 7083 9092 7125 9101
rect 7083 9052 7084 9092
rect 7124 9052 7125 9092
rect 7083 9043 7125 9052
rect 6987 8504 7029 8513
rect 6987 8464 6988 8504
rect 7028 8464 7029 8504
rect 6987 8455 7029 8464
rect 7084 8000 7124 9043
rect 7084 7951 7124 7960
rect 7180 7832 7220 9295
rect 7276 8429 7316 9472
rect 7371 9092 7413 9101
rect 7371 9052 7372 9092
rect 7412 9052 7413 9092
rect 7371 9043 7413 9052
rect 7372 8672 7412 9043
rect 7468 8933 7508 9640
rect 7564 9640 7892 9680
rect 7467 8924 7509 8933
rect 7467 8884 7468 8924
rect 7508 8884 7509 8924
rect 7467 8875 7509 8884
rect 7564 8672 7604 9640
rect 7659 9512 7701 9521
rect 7659 9472 7660 9512
rect 7700 9472 7701 9512
rect 7659 9463 7701 9472
rect 7756 9512 7796 9521
rect 7660 9378 7700 9463
rect 7756 8840 7796 9472
rect 7852 9512 7892 9640
rect 7852 9463 7892 9472
rect 7948 9512 7988 9521
rect 7948 9344 7988 9472
rect 7372 8623 7412 8632
rect 7468 8632 7604 8672
rect 7660 8800 7796 8840
rect 7852 9304 7988 9344
rect 7371 8504 7413 8513
rect 7371 8464 7372 8504
rect 7412 8464 7413 8504
rect 7371 8455 7413 8464
rect 7275 8420 7317 8429
rect 7275 8380 7276 8420
rect 7316 8380 7317 8420
rect 7275 8371 7317 8380
rect 7084 7792 7220 7832
rect 7084 7160 7124 7792
rect 7276 7748 7316 7757
rect 7276 7337 7316 7708
rect 7275 7328 7317 7337
rect 7275 7288 7276 7328
rect 7316 7288 7317 7328
rect 7275 7279 7317 7288
rect 6987 6572 7029 6581
rect 6987 6532 6988 6572
rect 7028 6532 7029 6572
rect 6987 6523 7029 6532
rect 6891 6152 6933 6161
rect 6891 6112 6892 6152
rect 6932 6112 6933 6152
rect 6891 6103 6933 6112
rect 6411 4724 6453 4733
rect 6411 4684 6412 4724
rect 6452 4684 6453 4724
rect 6411 4675 6453 4684
rect 6316 4516 6452 4556
rect 5932 3583 5972 3592
rect 6220 3380 6260 4096
rect 6315 4052 6357 4061
rect 6315 4012 6316 4052
rect 6356 4012 6357 4052
rect 6315 4003 6357 4012
rect 6028 3340 6260 3380
rect 5931 3212 5973 3221
rect 5931 3172 5932 3212
rect 5972 3172 5973 3212
rect 5931 3163 5973 3172
rect 5835 3128 5877 3137
rect 5548 3088 5684 3128
rect 5396 2584 5492 2624
rect 5548 2624 5588 2633
rect 5356 2575 5396 2584
rect 4876 2540 4916 2549
rect 5548 2540 5588 2584
rect 4684 1903 4724 1912
rect 4780 2500 4876 2540
rect 4491 1700 4533 1709
rect 4491 1660 4492 1700
rect 4532 1660 4533 1700
rect 4491 1651 4533 1660
rect 4299 1532 4341 1541
rect 4299 1492 4300 1532
rect 4340 1492 4341 1532
rect 4299 1483 4341 1492
rect 4052 1240 4244 1280
rect 4012 1231 4052 1240
rect 3532 1063 3572 1072
rect 3724 1112 3764 1231
rect 3724 1063 3764 1072
rect 3819 1112 3861 1121
rect 3819 1072 3820 1112
rect 3860 1072 3861 1112
rect 3819 1063 3861 1072
rect 4300 1112 4340 1483
rect 4300 1063 4340 1072
rect 4395 1112 4437 1121
rect 4395 1072 4396 1112
rect 4436 1072 4437 1112
rect 4395 1063 4437 1072
rect 3820 978 3860 1063
rect 4396 978 4436 1063
rect 2091 944 2133 953
rect 2091 904 2092 944
rect 2132 904 2133 944
rect 2091 895 2133 904
rect 3244 944 3284 955
rect 3244 869 3284 904
rect 3531 944 3573 953
rect 3531 904 3532 944
rect 3572 904 3573 944
rect 3531 895 3573 904
rect 3243 860 3285 869
rect 3243 820 3244 860
rect 3284 820 3285 860
rect 3243 811 3285 820
rect 3532 810 3572 895
rect 4492 869 4532 1651
rect 4683 1280 4725 1289
rect 4780 1280 4820 2500
rect 4876 2491 4916 2500
rect 5452 2500 5588 2540
rect 5644 2540 5684 3088
rect 5835 3088 5836 3128
rect 5876 3088 5877 3128
rect 5835 3079 5877 3088
rect 5932 3078 5972 3163
rect 6028 2540 6068 3340
rect 6220 3212 6260 3223
rect 6220 3137 6260 3172
rect 6219 3128 6261 3137
rect 6219 3088 6220 3128
rect 6260 3088 6261 3128
rect 6219 3079 6261 3088
rect 5644 2500 5876 2540
rect 4928 2288 5296 2297
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 4928 2239 5296 2248
rect 4875 2036 4917 2045
rect 4875 1996 4876 2036
rect 4916 1996 4917 2036
rect 4875 1987 4917 1996
rect 4876 1902 4916 1987
rect 5164 1952 5204 1961
rect 5164 1625 5204 1912
rect 5259 1952 5301 1961
rect 5259 1912 5260 1952
rect 5300 1912 5301 1952
rect 5259 1903 5301 1912
rect 5260 1818 5300 1903
rect 5355 1784 5397 1793
rect 5355 1744 5356 1784
rect 5396 1744 5397 1784
rect 5355 1735 5397 1744
rect 5163 1616 5205 1625
rect 5068 1576 5164 1616
rect 5204 1576 5205 1616
rect 5068 1289 5108 1576
rect 5163 1567 5205 1576
rect 4683 1240 4684 1280
rect 4724 1240 4820 1280
rect 5067 1280 5109 1289
rect 5067 1240 5068 1280
rect 5108 1240 5109 1280
rect 4683 1231 4725 1240
rect 5067 1231 5109 1240
rect 4684 1112 4724 1231
rect 4684 1063 4724 1072
rect 5068 1112 5108 1231
rect 5068 1063 5108 1072
rect 5163 1112 5205 1121
rect 5163 1072 5164 1112
rect 5204 1072 5205 1112
rect 5163 1063 5205 1072
rect 5164 978 5204 1063
rect 4491 860 4533 869
rect 4491 820 4492 860
rect 4532 820 4533 860
rect 4491 811 4533 820
rect 4928 776 5296 785
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 4928 727 5296 736
rect 1803 608 1845 617
rect 1803 568 1804 608
rect 1844 568 1845 608
rect 1803 559 1845 568
rect 5356 113 5396 1735
rect 5452 1205 5492 2500
rect 5739 2288 5781 2297
rect 5739 2248 5740 2288
rect 5780 2248 5781 2288
rect 5739 2239 5781 2248
rect 5740 1952 5780 2239
rect 5836 1961 5876 2500
rect 5932 2500 6068 2540
rect 5740 1903 5780 1912
rect 5835 1952 5877 1961
rect 5835 1912 5836 1952
rect 5876 1912 5877 1952
rect 5835 1903 5877 1912
rect 5644 1868 5684 1877
rect 5644 1709 5684 1828
rect 5643 1700 5685 1709
rect 5643 1660 5644 1700
rect 5684 1660 5685 1700
rect 5643 1651 5685 1660
rect 5547 1532 5589 1541
rect 5547 1492 5548 1532
rect 5588 1492 5589 1532
rect 5547 1483 5589 1492
rect 5451 1196 5493 1205
rect 5451 1156 5452 1196
rect 5492 1156 5493 1196
rect 5451 1147 5493 1156
rect 5548 1196 5588 1483
rect 5836 1457 5876 1903
rect 5835 1448 5877 1457
rect 5835 1408 5836 1448
rect 5876 1408 5877 1448
rect 5835 1399 5877 1408
rect 5548 1147 5588 1156
rect 5452 701 5492 1147
rect 5932 1121 5972 2500
rect 6220 1952 6260 1963
rect 6220 1877 6260 1912
rect 6219 1868 6261 1877
rect 6219 1828 6220 1868
rect 6260 1828 6261 1868
rect 6219 1819 6261 1828
rect 5644 1112 5684 1121
rect 5451 692 5493 701
rect 5451 652 5452 692
rect 5492 652 5493 692
rect 5451 643 5493 652
rect 5644 113 5684 1072
rect 5931 1112 5973 1121
rect 5931 1072 5932 1112
rect 5972 1072 5973 1112
rect 5931 1063 5973 1072
rect 6124 1112 6164 1121
rect 6316 1112 6356 4003
rect 6412 3725 6452 4516
rect 6411 3716 6453 3725
rect 6411 3676 6412 3716
rect 6452 3676 6453 3716
rect 6411 3667 6453 3676
rect 6412 3464 6452 3667
rect 6412 3415 6452 3424
rect 6508 1709 6548 4852
rect 6603 4724 6645 4733
rect 6603 4684 6604 4724
rect 6644 4684 6645 4724
rect 6700 4724 6740 5608
rect 6891 5648 6933 5657
rect 6891 5608 6892 5648
rect 6932 5608 6933 5648
rect 6988 5648 7028 6523
rect 7084 6488 7124 7120
rect 7180 7160 7220 7169
rect 7180 7001 7220 7120
rect 7179 6992 7221 7001
rect 7179 6952 7180 6992
rect 7220 6952 7221 6992
rect 7179 6943 7221 6952
rect 7084 6329 7124 6448
rect 7180 6488 7220 6497
rect 7083 6320 7125 6329
rect 7083 6280 7084 6320
rect 7124 6280 7125 6320
rect 7083 6271 7125 6280
rect 7180 5825 7220 6448
rect 7276 6413 7316 7279
rect 7275 6404 7317 6413
rect 7275 6364 7276 6404
rect 7316 6364 7317 6404
rect 7275 6355 7317 6364
rect 7275 6236 7317 6245
rect 7275 6196 7276 6236
rect 7316 6196 7317 6236
rect 7275 6187 7317 6196
rect 7179 5816 7221 5825
rect 7179 5776 7180 5816
rect 7220 5776 7221 5816
rect 7179 5767 7221 5776
rect 7180 5648 7220 5657
rect 6988 5608 7180 5648
rect 6891 5599 6933 5608
rect 6795 5312 6837 5321
rect 6795 5272 6796 5312
rect 6836 5272 6837 5312
rect 6795 5263 6837 5272
rect 6796 4976 6836 5263
rect 6796 4901 6836 4936
rect 6892 4976 6932 5599
rect 6892 4927 6932 4936
rect 6795 4892 6837 4901
rect 6795 4852 6796 4892
rect 6836 4852 6837 4892
rect 6795 4843 6837 4852
rect 6700 4684 6932 4724
rect 6603 4675 6645 4684
rect 6604 4136 6644 4675
rect 6699 4472 6741 4481
rect 6699 4432 6700 4472
rect 6740 4432 6741 4472
rect 6699 4423 6741 4432
rect 6604 3977 6644 4096
rect 6700 4220 6740 4423
rect 6603 3968 6645 3977
rect 6603 3928 6604 3968
rect 6644 3928 6645 3968
rect 6603 3919 6645 3928
rect 6700 2540 6740 4180
rect 6795 3716 6837 3725
rect 6795 3676 6796 3716
rect 6836 3676 6837 3716
rect 6795 3667 6837 3676
rect 6796 2624 6836 3667
rect 6796 2575 6836 2584
rect 6604 2500 6740 2540
rect 6507 1700 6549 1709
rect 6507 1660 6508 1700
rect 6548 1660 6549 1700
rect 6507 1651 6549 1660
rect 6604 1280 6644 2500
rect 6892 2297 6932 4684
rect 7084 3389 7124 5608
rect 7180 5599 7220 5608
rect 7276 5153 7316 6187
rect 7372 6077 7412 8455
rect 7468 8336 7508 8632
rect 7564 8504 7604 8513
rect 7660 8504 7700 8800
rect 7755 8672 7797 8681
rect 7755 8632 7756 8672
rect 7796 8632 7797 8672
rect 7755 8623 7797 8632
rect 7756 8538 7796 8623
rect 7604 8464 7700 8504
rect 7564 8455 7604 8464
rect 7468 8296 7604 8336
rect 7564 7328 7604 8296
rect 7660 8009 7700 8464
rect 7659 8000 7701 8009
rect 7659 7960 7660 8000
rect 7700 7960 7701 8000
rect 7659 7951 7701 7960
rect 7756 8000 7796 8009
rect 7660 7866 7700 7951
rect 7756 7589 7796 7960
rect 7755 7580 7797 7589
rect 7755 7540 7756 7580
rect 7796 7540 7797 7580
rect 7755 7531 7797 7540
rect 7852 7421 7892 9304
rect 8140 9260 8180 9269
rect 7948 9220 8140 9260
rect 7948 8000 7988 9220
rect 8140 9211 8180 9220
rect 8140 8177 8180 8262
rect 8139 8168 8181 8177
rect 8139 8128 8140 8168
rect 8180 8128 8181 8168
rect 8139 8119 8181 8128
rect 8236 8084 8276 10692
rect 8696 10672 8776 10752
rect 9848 10672 9928 10752
rect 11000 10672 11080 10752
rect 12152 10732 12232 10752
rect 11788 10692 12232 10732
rect 8716 10193 8756 10672
rect 8715 10184 8757 10193
rect 8715 10144 8716 10184
rect 8756 10144 8757 10184
rect 8715 10135 8757 10144
rect 8812 9892 9140 9932
rect 8619 9680 8661 9689
rect 8619 9640 8620 9680
rect 8660 9640 8661 9680
rect 8619 9631 8661 9640
rect 8332 9512 8372 9521
rect 8620 9512 8660 9631
rect 8372 9472 8468 9512
rect 8332 9463 8372 9472
rect 8331 9344 8373 9353
rect 8331 9304 8332 9344
rect 8372 9304 8373 9344
rect 8331 9295 8373 9304
rect 8332 9210 8372 9295
rect 8428 9185 8468 9472
rect 8620 9463 8660 9472
rect 8715 9512 8757 9521
rect 8715 9472 8716 9512
rect 8756 9472 8757 9512
rect 8715 9463 8757 9472
rect 8812 9512 8852 9892
rect 9003 9764 9045 9773
rect 9003 9724 9004 9764
rect 9044 9724 9045 9764
rect 9003 9715 9045 9724
rect 8812 9463 8852 9472
rect 8908 9512 8948 9521
rect 8716 9378 8756 9463
rect 8427 9176 8469 9185
rect 8427 9136 8428 9176
rect 8468 9136 8469 9176
rect 8427 9127 8469 9136
rect 8811 9092 8853 9101
rect 8811 9052 8812 9092
rect 8852 9052 8853 9092
rect 8811 9043 8853 9052
rect 8812 8597 8852 9043
rect 8811 8588 8853 8597
rect 8811 8548 8812 8588
rect 8852 8548 8853 8588
rect 8811 8539 8853 8548
rect 8619 8504 8661 8513
rect 8619 8464 8620 8504
rect 8660 8464 8661 8504
rect 8619 8455 8661 8464
rect 8236 8044 8372 8084
rect 7948 7951 7988 7960
rect 8044 8000 8084 8009
rect 7851 7412 7893 7421
rect 7851 7372 7852 7412
rect 7892 7372 7893 7412
rect 7851 7363 7893 7372
rect 8044 7337 8084 7960
rect 8201 7985 8241 7994
rect 8201 7664 8241 7945
rect 8201 7624 8276 7664
rect 8043 7328 8085 7337
rect 7564 7288 7796 7328
rect 7564 7160 7604 7171
rect 7564 7085 7604 7120
rect 7660 7160 7700 7169
rect 7563 7076 7605 7085
rect 7468 7036 7564 7076
rect 7604 7036 7605 7076
rect 7371 6068 7413 6077
rect 7371 6028 7372 6068
rect 7412 6028 7413 6068
rect 7371 6019 7413 6028
rect 7275 5144 7317 5153
rect 7275 5104 7276 5144
rect 7316 5104 7317 5144
rect 7275 5095 7317 5104
rect 7275 4976 7317 4985
rect 7180 4936 7276 4976
rect 7316 4936 7317 4976
rect 7180 4313 7220 4936
rect 7275 4927 7317 4936
rect 7372 4976 7412 6019
rect 7468 5909 7508 7036
rect 7563 7027 7605 7036
rect 7660 6581 7700 7120
rect 7659 6572 7701 6581
rect 7659 6532 7660 6572
rect 7700 6532 7701 6572
rect 7659 6523 7701 6532
rect 7564 6404 7604 6413
rect 7467 5900 7509 5909
rect 7467 5860 7468 5900
rect 7508 5860 7509 5900
rect 7467 5851 7509 5860
rect 7564 5732 7604 6364
rect 7660 6404 7700 6413
rect 7660 6245 7700 6364
rect 7659 6236 7701 6245
rect 7659 6196 7660 6236
rect 7700 6196 7701 6236
rect 7659 6187 7701 6196
rect 7276 4842 7316 4927
rect 7372 4397 7412 4936
rect 7468 5692 7604 5732
rect 7371 4388 7413 4397
rect 7371 4348 7372 4388
rect 7412 4348 7413 4388
rect 7371 4339 7413 4348
rect 7179 4304 7221 4313
rect 7179 4264 7180 4304
rect 7220 4264 7221 4304
rect 7179 4255 7221 4264
rect 7468 4220 7508 5692
rect 7660 5657 7700 5666
rect 7564 5617 7660 5648
rect 7564 5608 7700 5617
rect 7564 4901 7604 5608
rect 7756 5564 7796 7288
rect 8043 7288 8044 7328
rect 8084 7288 8085 7328
rect 8043 7279 8085 7288
rect 8140 7160 8180 7169
rect 8140 6665 8180 7120
rect 8139 6656 8181 6665
rect 8139 6616 8140 6656
rect 8180 6616 8181 6656
rect 8139 6607 8181 6616
rect 8139 6488 8181 6497
rect 8139 6448 8140 6488
rect 8180 6448 8181 6488
rect 8139 6439 8181 6448
rect 8140 6354 8180 6439
rect 8140 5900 8180 5909
rect 8236 5900 8276 7624
rect 8180 5860 8276 5900
rect 8140 5851 8180 5860
rect 8235 5732 8277 5741
rect 8235 5692 8236 5732
rect 8276 5692 8277 5732
rect 8235 5683 8277 5692
rect 7660 5524 7796 5564
rect 7660 5069 7700 5524
rect 7852 5480 7892 5489
rect 7756 5440 7852 5480
rect 7659 5060 7701 5069
rect 7659 5020 7660 5060
rect 7700 5020 7701 5060
rect 7659 5011 7701 5020
rect 7563 4892 7605 4901
rect 7563 4852 7564 4892
rect 7604 4852 7700 4892
rect 7563 4843 7605 4852
rect 7372 4180 7508 4220
rect 7180 4136 7220 4147
rect 7180 4061 7220 4096
rect 7179 4052 7221 4061
rect 7179 4012 7180 4052
rect 7220 4012 7221 4052
rect 7179 4003 7221 4012
rect 7372 3977 7412 4180
rect 7660 4150 7700 4852
rect 7660 4052 7700 4110
rect 7468 4012 7700 4052
rect 7371 3968 7413 3977
rect 7371 3928 7372 3968
rect 7412 3928 7413 3968
rect 7371 3919 7413 3928
rect 7468 3800 7508 4012
rect 7563 3884 7605 3893
rect 7563 3844 7564 3884
rect 7604 3844 7605 3884
rect 7563 3835 7605 3844
rect 7372 3760 7508 3800
rect 7083 3380 7125 3389
rect 7083 3340 7084 3380
rect 7124 3340 7125 3380
rect 7083 3331 7125 3340
rect 7275 3296 7317 3305
rect 7275 3256 7276 3296
rect 7316 3256 7317 3296
rect 7275 3247 7317 3256
rect 7083 3044 7125 3053
rect 7083 3004 7084 3044
rect 7124 3004 7125 3044
rect 7083 2995 7125 3004
rect 7084 2801 7124 2995
rect 7083 2792 7125 2801
rect 7083 2752 7084 2792
rect 7124 2752 7125 2792
rect 7083 2743 7125 2752
rect 6988 2549 7028 2634
rect 6987 2540 7029 2549
rect 6987 2500 6988 2540
rect 7028 2500 7029 2540
rect 6987 2491 7029 2500
rect 6891 2288 6933 2297
rect 6891 2248 6892 2288
rect 6932 2248 6933 2288
rect 6891 2239 6933 2248
rect 6892 2036 6932 2045
rect 6164 1072 6356 1112
rect 6508 1240 6644 1280
rect 6700 1938 6740 1947
rect 6124 1063 6164 1072
rect 6508 113 6548 1240
rect 6700 1196 6740 1898
rect 6604 1156 6740 1196
rect 6604 1117 6644 1156
rect 6892 1121 6932 1996
rect 6604 785 6644 1077
rect 6891 1112 6933 1121
rect 6891 1072 6892 1112
rect 6932 1072 6933 1112
rect 6891 1063 6933 1072
rect 7084 1112 7124 2743
rect 7180 2624 7220 2633
rect 7180 2549 7220 2584
rect 7179 2540 7221 2549
rect 7179 2500 7180 2540
rect 7220 2500 7221 2540
rect 7179 2491 7221 2500
rect 7180 1793 7220 2491
rect 7276 2120 7316 3247
rect 7276 2071 7316 2080
rect 7372 1952 7412 3760
rect 7467 3212 7509 3221
rect 7467 3172 7468 3212
rect 7508 3172 7509 3212
rect 7467 3163 7509 3172
rect 7372 1903 7412 1912
rect 7468 1952 7508 3163
rect 7564 2129 7604 3835
rect 7659 3800 7701 3809
rect 7659 3760 7660 3800
rect 7700 3760 7701 3800
rect 7756 3800 7796 5440
rect 7852 5431 7892 5440
rect 7851 5228 7893 5237
rect 7851 5188 7852 5228
rect 7892 5188 7893 5228
rect 7851 5179 7893 5188
rect 7852 4976 7892 5179
rect 8236 5060 8276 5683
rect 8332 5489 8372 8044
rect 8523 8000 8565 8009
rect 8523 7960 8524 8000
rect 8564 7960 8565 8000
rect 8523 7951 8565 7960
rect 8524 7866 8564 7951
rect 8620 7925 8660 8455
rect 8908 8177 8948 9472
rect 9004 8840 9044 9715
rect 9100 9512 9140 9892
rect 9388 9680 9428 9689
rect 9868 9680 9908 10672
rect 11020 10109 11060 10672
rect 11019 10100 11061 10109
rect 11019 10060 11020 10100
rect 11060 10060 11061 10100
rect 11019 10051 11061 10060
rect 11499 9764 11541 9773
rect 11499 9724 11500 9764
rect 11540 9724 11541 9764
rect 11499 9715 11541 9724
rect 9100 8924 9140 9472
rect 9196 9512 9236 9521
rect 9236 9472 9332 9512
rect 9196 9463 9236 9472
rect 9196 8924 9236 8933
rect 9100 8884 9196 8924
rect 9196 8875 9236 8884
rect 9004 8800 9140 8840
rect 9004 8672 9044 8683
rect 9004 8597 9044 8632
rect 9003 8588 9045 8597
rect 9003 8548 9004 8588
rect 9044 8548 9045 8588
rect 9003 8539 9045 8548
rect 8907 8168 8949 8177
rect 8907 8128 8908 8168
rect 8948 8128 8949 8168
rect 8907 8119 8949 8128
rect 8812 8000 8852 8009
rect 8619 7916 8661 7925
rect 8619 7876 8620 7916
rect 8660 7876 8661 7916
rect 8619 7867 8661 7876
rect 8620 7496 8660 7867
rect 8524 7456 8660 7496
rect 8427 6908 8469 6917
rect 8427 6868 8428 6908
rect 8468 6868 8469 6908
rect 8427 6859 8469 6868
rect 8428 5741 8468 6859
rect 8524 6245 8564 7456
rect 8619 7328 8661 7337
rect 8619 7288 8620 7328
rect 8660 7288 8661 7328
rect 8619 7279 8661 7288
rect 8620 7165 8660 7279
rect 8620 6474 8660 7125
rect 8812 7076 8852 7960
rect 8812 7027 8852 7036
rect 8908 8000 8948 8009
rect 8715 6656 8757 6665
rect 8715 6616 8716 6656
rect 8756 6616 8757 6656
rect 8715 6607 8757 6616
rect 8812 6656 8852 6665
rect 8908 6656 8948 7960
rect 9003 7412 9045 7421
rect 9003 7372 9004 7412
rect 9044 7372 9045 7412
rect 9003 7363 9045 7372
rect 9004 7278 9044 7363
rect 8852 6616 8948 6656
rect 9004 7160 9044 7169
rect 8812 6607 8852 6616
rect 8620 6413 8660 6434
rect 8619 6404 8661 6413
rect 8619 6364 8620 6404
rect 8660 6364 8661 6404
rect 8619 6355 8661 6364
rect 8523 6236 8565 6245
rect 8523 6196 8524 6236
rect 8564 6196 8565 6236
rect 8523 6187 8565 6196
rect 8716 6161 8756 6607
rect 9004 6572 9044 7120
rect 9100 6833 9140 8800
rect 9196 7832 9236 7841
rect 9292 7832 9332 9472
rect 9388 8504 9428 9640
rect 9772 9640 9908 9680
rect 9483 8756 9525 8765
rect 9483 8716 9484 8756
rect 9524 8716 9525 8756
rect 9483 8707 9525 8716
rect 9484 8672 9524 8707
rect 9580 8681 9620 8766
rect 9772 8681 9812 9640
rect 9868 9512 9908 9521
rect 9868 9353 9908 9472
rect 10731 9512 10773 9521
rect 10731 9472 10732 9512
rect 10772 9472 10773 9512
rect 10731 9463 10773 9472
rect 11115 9512 11157 9521
rect 11115 9472 11116 9512
rect 11156 9472 11157 9512
rect 11115 9463 11157 9472
rect 11500 9512 11540 9715
rect 9867 9344 9909 9353
rect 9867 9304 9868 9344
rect 9908 9304 9909 9344
rect 9867 9295 9909 9304
rect 9484 8621 9524 8632
rect 9579 8672 9621 8681
rect 9579 8632 9580 8672
rect 9620 8632 9621 8672
rect 9579 8623 9621 8632
rect 9676 8672 9716 8681
rect 9676 8504 9716 8632
rect 9771 8672 9813 8681
rect 9771 8632 9772 8672
rect 9812 8632 9813 8672
rect 9771 8623 9813 8632
rect 9388 8464 9620 8504
rect 9483 8168 9525 8177
rect 9483 8128 9484 8168
rect 9524 8128 9525 8168
rect 9483 8119 9525 8128
rect 9387 8084 9429 8093
rect 9387 8044 9388 8084
rect 9428 8044 9429 8084
rect 9387 8035 9429 8044
rect 9388 8000 9428 8035
rect 9388 7949 9428 7960
rect 9484 8000 9524 8119
rect 9484 7951 9524 7960
rect 9580 8000 9620 8464
rect 9675 8464 9716 8504
rect 9772 8504 9812 8515
rect 9675 8336 9715 8464
rect 9772 8429 9812 8464
rect 9771 8420 9813 8429
rect 9771 8380 9772 8420
rect 9812 8380 9813 8420
rect 9771 8371 9813 8380
rect 9868 8345 9908 9295
rect 10732 9101 10772 9463
rect 11116 9378 11156 9463
rect 11308 9260 11348 9269
rect 11115 9176 11157 9185
rect 11115 9136 11116 9176
rect 11156 9136 11157 9176
rect 11115 9127 11157 9136
rect 10731 9092 10773 9101
rect 10731 9052 10732 9092
rect 10772 9052 10773 9092
rect 10731 9043 10773 9052
rect 10347 8840 10389 8849
rect 10347 8800 10348 8840
rect 10388 8800 10389 8840
rect 10347 8791 10389 8800
rect 9964 8672 10004 8681
rect 9867 8336 9909 8345
rect 9675 8296 9716 8336
rect 9676 8177 9716 8296
rect 9867 8296 9868 8336
rect 9908 8296 9909 8336
rect 9867 8287 9909 8296
rect 9675 8168 9717 8177
rect 9675 8128 9676 8168
rect 9716 8128 9717 8168
rect 9675 8119 9717 8128
rect 9868 8168 9908 8177
rect 9964 8168 10004 8632
rect 10060 8672 10100 8681
rect 10060 8429 10100 8632
rect 10155 8588 10197 8597
rect 10155 8548 10156 8588
rect 10196 8548 10197 8588
rect 10155 8539 10197 8548
rect 10059 8420 10101 8429
rect 10059 8380 10060 8420
rect 10100 8380 10101 8420
rect 10059 8371 10101 8380
rect 10059 8252 10101 8261
rect 10059 8212 10060 8252
rect 10100 8212 10101 8252
rect 10059 8203 10101 8212
rect 9908 8128 10004 8168
rect 9868 8119 9908 8128
rect 9580 7951 9620 7960
rect 9676 8000 9716 8009
rect 9676 7841 9716 7960
rect 9963 8000 10005 8009
rect 9963 7960 9964 8000
rect 10004 7960 10005 8000
rect 9963 7951 10005 7960
rect 10060 8000 10100 8203
rect 10156 8177 10196 8539
rect 10252 8504 10292 8513
rect 10155 8168 10197 8177
rect 10155 8128 10156 8168
rect 10196 8128 10197 8168
rect 10155 8119 10197 8128
rect 10060 7951 10100 7960
rect 10156 8000 10196 8119
rect 9964 7866 10004 7951
rect 9236 7792 9332 7832
rect 9675 7832 9717 7841
rect 10156 7832 10196 7960
rect 9675 7792 9676 7832
rect 9716 7792 9717 7832
rect 9196 7783 9236 7792
rect 9675 7783 9717 7792
rect 10060 7792 10196 7832
rect 9675 7664 9717 7673
rect 9675 7624 9676 7664
rect 9716 7624 9717 7664
rect 9675 7615 9717 7624
rect 9292 7160 9332 7169
rect 9484 7160 9524 7169
rect 9332 7120 9484 7160
rect 9099 6824 9141 6833
rect 9099 6784 9100 6824
rect 9140 6784 9141 6824
rect 9099 6775 9141 6784
rect 9292 6665 9332 7120
rect 9484 7111 9524 7120
rect 9579 7160 9621 7169
rect 9579 7120 9580 7160
rect 9620 7120 9621 7160
rect 9579 7111 9621 7120
rect 9676 7160 9716 7615
rect 9868 7412 9908 7421
rect 10060 7412 10100 7792
rect 10252 7589 10292 8464
rect 10348 8345 10388 8791
rect 10443 8672 10485 8681
rect 10443 8632 10444 8672
rect 10484 8632 10485 8672
rect 10443 8623 10485 8632
rect 10540 8672 10580 8683
rect 10347 8336 10389 8345
rect 10347 8296 10348 8336
rect 10388 8296 10389 8336
rect 10347 8287 10389 8296
rect 10348 8168 10388 8177
rect 10444 8168 10484 8623
rect 10540 8597 10580 8632
rect 10636 8672 10676 8681
rect 10539 8588 10581 8597
rect 10539 8548 10540 8588
rect 10580 8548 10581 8588
rect 10539 8539 10581 8548
rect 10636 8513 10676 8632
rect 10635 8504 10677 8513
rect 10635 8464 10636 8504
rect 10676 8464 10677 8504
rect 10635 8455 10677 8464
rect 10732 8252 10772 9043
rect 11020 8765 11060 8796
rect 11019 8756 11061 8765
rect 11019 8716 11020 8756
rect 11060 8716 11061 8756
rect 11019 8707 11061 8716
rect 11116 8756 11156 9127
rect 11308 8840 11348 9220
rect 11308 8800 11444 8840
rect 11116 8707 11156 8716
rect 11020 8672 11060 8707
rect 11020 8597 11060 8632
rect 11019 8588 11061 8597
rect 11019 8548 11020 8588
rect 11060 8548 11061 8588
rect 11019 8539 11061 8548
rect 10388 8128 10484 8168
rect 10540 8212 10772 8252
rect 10348 8119 10388 8128
rect 10540 8000 10580 8212
rect 10635 8084 10677 8093
rect 10635 8044 10636 8084
rect 10676 8044 10677 8084
rect 10635 8035 10677 8044
rect 10444 7960 10540 8000
rect 10444 7832 10484 7960
rect 10540 7951 10580 7960
rect 10347 7792 10484 7832
rect 10347 7664 10387 7792
rect 10636 7664 10676 8035
rect 11404 8009 11444 8800
rect 11403 8000 11445 8009
rect 11403 7960 11404 8000
rect 11444 7960 11445 8000
rect 11403 7951 11445 7960
rect 10347 7624 10388 7664
rect 10251 7580 10293 7589
rect 10251 7540 10252 7580
rect 10292 7540 10293 7580
rect 10251 7531 10293 7540
rect 10348 7412 10388 7624
rect 9908 7372 10100 7412
rect 10156 7372 10388 7412
rect 10444 7624 10676 7664
rect 9868 7363 9908 7372
rect 10156 7328 10196 7372
rect 9580 7026 9620 7111
rect 9676 6917 9716 7120
rect 10060 7288 10196 7328
rect 10060 7160 10100 7288
rect 10060 7111 10100 7120
rect 9675 6908 9717 6917
rect 9675 6868 9676 6908
rect 9716 6868 9717 6908
rect 9675 6859 9717 6868
rect 9579 6824 9621 6833
rect 9579 6784 9580 6824
rect 9620 6784 9621 6824
rect 9579 6775 9621 6784
rect 9291 6656 9333 6665
rect 9291 6616 9292 6656
rect 9332 6616 9333 6656
rect 9291 6607 9333 6616
rect 8908 6532 9044 6572
rect 8811 6320 8853 6329
rect 8811 6280 8812 6320
rect 8852 6280 8853 6320
rect 8811 6271 8853 6280
rect 8715 6152 8757 6161
rect 8715 6112 8716 6152
rect 8756 6112 8757 6152
rect 8715 6103 8757 6112
rect 8427 5732 8469 5741
rect 8427 5692 8428 5732
rect 8468 5692 8469 5732
rect 8427 5683 8469 5692
rect 8524 5667 8564 5676
rect 8715 5648 8757 5657
rect 8564 5627 8660 5648
rect 8524 5608 8660 5627
rect 8428 5564 8468 5573
rect 8331 5480 8373 5489
rect 8331 5440 8332 5480
rect 8372 5440 8373 5480
rect 8331 5431 8373 5440
rect 8428 5237 8468 5524
rect 8427 5228 8469 5237
rect 8427 5188 8428 5228
rect 8468 5188 8469 5228
rect 8427 5179 8469 5188
rect 8523 5060 8565 5069
rect 8236 5020 8468 5060
rect 7852 4927 7892 4936
rect 8332 4962 8372 4971
rect 8332 4136 8372 4922
rect 8428 4304 8468 5020
rect 8523 5020 8524 5060
rect 8564 5020 8565 5060
rect 8523 5011 8565 5020
rect 8524 4926 8564 5011
rect 8620 4985 8660 5608
rect 8715 5608 8716 5648
rect 8756 5608 8757 5648
rect 8715 5599 8757 5608
rect 8812 5648 8852 6271
rect 8812 5599 8852 5608
rect 8716 5144 8756 5599
rect 8908 5153 8948 6532
rect 9100 6488 9140 6497
rect 9004 6443 9044 6452
rect 9004 5993 9044 6403
rect 9003 5984 9045 5993
rect 9003 5944 9004 5984
rect 9044 5944 9045 5984
rect 9003 5935 9045 5944
rect 9100 5816 9140 6448
rect 9196 6488 9236 6497
rect 9196 5825 9236 6448
rect 9292 6488 9332 6497
rect 9580 6488 9620 6775
rect 9332 6448 9524 6488
rect 9292 6439 9332 6448
rect 9484 6068 9524 6448
rect 9580 6439 9620 6448
rect 9484 6028 9812 6068
rect 9291 5984 9333 5993
rect 9291 5944 9292 5984
rect 9332 5944 9333 5984
rect 9291 5935 9333 5944
rect 9004 5776 9140 5816
rect 9195 5816 9237 5825
rect 9195 5776 9196 5816
rect 9236 5776 9237 5816
rect 8716 5095 8756 5104
rect 8907 5144 8949 5153
rect 8907 5104 8908 5144
rect 8948 5104 8949 5144
rect 8907 5095 8949 5104
rect 9004 5069 9044 5776
rect 9195 5767 9237 5776
rect 9099 5648 9141 5657
rect 9099 5608 9100 5648
rect 9140 5608 9141 5648
rect 9099 5599 9141 5608
rect 9196 5648 9236 5657
rect 9100 5514 9140 5599
rect 9003 5060 9045 5069
rect 9003 5020 9004 5060
rect 9044 5020 9045 5060
rect 9003 5011 9045 5020
rect 8619 4976 8661 4985
rect 8619 4936 8620 4976
rect 8660 4936 8661 4976
rect 8619 4927 8661 4936
rect 8908 4976 8948 4985
rect 8620 4481 8660 4927
rect 8619 4472 8661 4481
rect 8619 4432 8620 4472
rect 8660 4432 8661 4472
rect 8619 4423 8661 4432
rect 8428 4264 8756 4304
rect 8620 4136 8660 4147
rect 8372 4096 8468 4136
rect 8332 4087 8372 4096
rect 7852 3968 7892 3977
rect 7892 3928 8372 3968
rect 7852 3919 7892 3928
rect 7756 3760 8276 3800
rect 7659 3751 7701 3760
rect 7660 3464 7700 3751
rect 7947 3548 7989 3557
rect 7947 3508 7948 3548
rect 7988 3508 7989 3548
rect 7947 3499 7989 3508
rect 7660 3415 7700 3424
rect 7948 3464 7988 3499
rect 7948 3137 7988 3424
rect 8236 3464 8276 3760
rect 8332 3548 8372 3928
rect 8332 3499 8372 3508
rect 8236 3415 8276 3424
rect 8428 3221 8468 4096
rect 8620 4061 8660 4096
rect 8716 4136 8756 4264
rect 8716 4087 8756 4096
rect 8619 4052 8661 4061
rect 8619 4012 8620 4052
rect 8660 4012 8661 4052
rect 8619 4003 8661 4012
rect 8523 3968 8565 3977
rect 8523 3928 8524 3968
rect 8564 3928 8565 3968
rect 8523 3919 8565 3928
rect 8427 3212 8469 3221
rect 8427 3172 8428 3212
rect 8468 3172 8469 3212
rect 8427 3163 8469 3172
rect 7947 3128 7989 3137
rect 7947 3088 7948 3128
rect 7988 3088 7989 3128
rect 7947 3079 7989 3088
rect 8427 2708 8469 2717
rect 8427 2668 8428 2708
rect 8468 2668 8469 2708
rect 8427 2659 8469 2668
rect 8428 2624 8468 2659
rect 8428 2573 8468 2584
rect 8524 2372 8564 3919
rect 8908 3725 8948 4936
rect 9196 4472 9236 5608
rect 9100 4432 9236 4472
rect 9003 4388 9045 4397
rect 9003 4348 9004 4388
rect 9044 4348 9045 4388
rect 9003 4339 9045 4348
rect 9004 4254 9044 4339
rect 9003 3800 9045 3809
rect 9003 3760 9004 3800
rect 9044 3760 9045 3800
rect 9003 3751 9045 3760
rect 8907 3716 8949 3725
rect 8907 3676 8908 3716
rect 8948 3676 8949 3716
rect 8907 3667 8949 3676
rect 9004 3464 9044 3751
rect 9004 3415 9044 3424
rect 9100 3305 9140 4432
rect 9195 4304 9237 4313
rect 9195 4264 9196 4304
rect 9236 4264 9237 4304
rect 9195 4255 9237 4264
rect 9196 4136 9236 4255
rect 9196 4087 9236 4096
rect 9292 3557 9332 5935
rect 9676 5648 9716 5657
rect 9388 5608 9676 5648
rect 9388 5480 9428 5608
rect 9676 5599 9716 5608
rect 9772 5648 9812 6028
rect 10060 5816 10100 5825
rect 9772 5599 9812 5608
rect 9868 5776 10060 5816
rect 9868 5648 9908 5776
rect 10060 5767 10100 5776
rect 10156 5776 10388 5816
rect 10060 5648 10100 5657
rect 9868 5599 9908 5608
rect 9964 5608 10060 5648
rect 9388 5431 9428 5440
rect 9579 5480 9621 5489
rect 9579 5440 9580 5480
rect 9620 5440 9621 5480
rect 9579 5431 9621 5440
rect 9580 5346 9620 5431
rect 9483 5228 9525 5237
rect 9483 5188 9484 5228
rect 9524 5188 9525 5228
rect 9483 5179 9525 5188
rect 9387 5060 9429 5069
rect 9387 5020 9388 5060
rect 9428 5020 9429 5060
rect 9387 5011 9429 5020
rect 9388 4649 9428 5011
rect 9387 4640 9429 4649
rect 9387 4600 9388 4640
rect 9428 4600 9429 4640
rect 9387 4591 9429 4600
rect 9291 3548 9333 3557
rect 9291 3508 9292 3548
rect 9332 3508 9333 3548
rect 9291 3499 9333 3508
rect 8619 3296 8661 3305
rect 8619 3256 8620 3296
rect 8660 3256 8661 3296
rect 8619 3247 8661 3256
rect 9099 3296 9141 3305
rect 9099 3256 9100 3296
rect 9140 3256 9141 3296
rect 9099 3247 9141 3256
rect 8620 3162 8660 3247
rect 9484 3128 9524 5179
rect 9579 5060 9621 5069
rect 9579 5020 9580 5060
rect 9620 5020 9621 5060
rect 9579 5011 9621 5020
rect 9580 3893 9620 5011
rect 9771 4724 9813 4733
rect 9771 4684 9772 4724
rect 9812 4684 9813 4724
rect 9771 4675 9813 4684
rect 9579 3884 9621 3893
rect 9579 3844 9580 3884
rect 9620 3844 9621 3884
rect 9579 3835 9621 3844
rect 8908 3088 9524 3128
rect 8812 2633 8852 2718
rect 8811 2624 8853 2633
rect 8811 2584 8812 2624
rect 8852 2584 8853 2624
rect 8811 2575 8853 2584
rect 8332 2332 8564 2372
rect 8620 2456 8660 2465
rect 7563 2120 7605 2129
rect 7563 2080 7564 2120
rect 7604 2080 7605 2120
rect 7563 2071 7605 2080
rect 7468 1903 7508 1912
rect 7564 1952 7604 2071
rect 7851 2036 7893 2045
rect 7851 1996 7852 2036
rect 7892 1996 7893 2036
rect 7851 1987 7893 1996
rect 7564 1903 7604 1912
rect 7852 1952 7892 1987
rect 7852 1901 7892 1912
rect 7948 1952 7988 1961
rect 7179 1784 7221 1793
rect 7179 1744 7180 1784
rect 7220 1744 7221 1784
rect 7179 1735 7221 1744
rect 7948 1709 7988 1912
rect 8332 1868 8372 2332
rect 7947 1700 7989 1709
rect 7947 1660 7948 1700
rect 7988 1660 7989 1700
rect 7947 1651 7989 1660
rect 8332 1541 8372 1828
rect 8427 1868 8469 1877
rect 8427 1828 8428 1868
rect 8468 1828 8469 1868
rect 8427 1819 8469 1828
rect 8428 1734 8468 1819
rect 8331 1532 8373 1541
rect 8331 1492 8332 1532
rect 8372 1492 8373 1532
rect 8331 1483 8373 1492
rect 7755 1280 7797 1289
rect 7755 1240 7756 1280
rect 7796 1240 7797 1280
rect 7755 1231 7797 1240
rect 7372 1121 7412 1206
rect 7756 1146 7796 1231
rect 8620 1121 8660 2416
rect 8908 1952 8948 3088
rect 9675 2708 9717 2717
rect 9675 2668 9676 2708
rect 9716 2668 9717 2708
rect 9675 2659 9717 2668
rect 9195 2624 9237 2633
rect 9195 2584 9196 2624
rect 9236 2584 9237 2624
rect 9195 2575 9237 2584
rect 8908 1205 8948 1912
rect 8907 1196 8949 1205
rect 8907 1156 8908 1196
rect 8948 1156 8949 1196
rect 8907 1147 8949 1156
rect 7084 1063 7124 1072
rect 7371 1112 7413 1121
rect 7371 1072 7372 1112
rect 7412 1072 7413 1112
rect 7371 1063 7413 1072
rect 7947 1112 7989 1121
rect 7947 1072 7948 1112
rect 7988 1072 7989 1112
rect 7947 1063 7989 1072
rect 8619 1112 8661 1121
rect 8619 1072 8620 1112
rect 8660 1072 8661 1112
rect 8619 1063 8661 1072
rect 9196 1112 9236 2575
rect 9387 2456 9429 2465
rect 9387 2416 9388 2456
rect 9428 2416 9429 2456
rect 9387 2407 9429 2416
rect 9388 1947 9428 2407
rect 9579 2036 9621 2045
rect 9579 1996 9580 2036
rect 9620 1996 9621 2036
rect 9579 1987 9621 1996
rect 9388 1898 9428 1907
rect 9580 1902 9620 1987
rect 9676 1616 9716 2659
rect 9772 2540 9812 4675
rect 9964 4145 10004 5608
rect 10060 5599 10100 5608
rect 10156 5480 10196 5776
rect 10252 5648 10292 5657
rect 10252 5489 10292 5608
rect 10348 5648 10388 5776
rect 10348 5599 10388 5608
rect 10060 5440 10196 5480
rect 10251 5480 10293 5489
rect 10251 5440 10252 5480
rect 10292 5440 10293 5480
rect 10060 4397 10100 5440
rect 10251 5431 10293 5440
rect 10156 4976 10196 4985
rect 10156 4817 10196 4936
rect 10347 4976 10389 4985
rect 10347 4936 10348 4976
rect 10388 4936 10389 4976
rect 10347 4927 10389 4936
rect 10444 4976 10484 7624
rect 10923 7496 10965 7505
rect 10923 7456 10924 7496
rect 10964 7456 10965 7496
rect 10923 7447 10965 7456
rect 10924 7001 10964 7447
rect 11308 7160 11348 7169
rect 11308 7001 11348 7120
rect 10923 6992 10965 7001
rect 10923 6952 10924 6992
rect 10964 6952 10965 6992
rect 10923 6943 10965 6952
rect 11307 6992 11349 7001
rect 11307 6952 11308 6992
rect 11348 6952 11349 6992
rect 11307 6943 11349 6952
rect 10828 6488 10868 6499
rect 10828 6413 10868 6448
rect 11404 6488 11444 7951
rect 11500 7505 11540 9472
rect 11595 8672 11637 8681
rect 11595 8632 11596 8672
rect 11636 8632 11637 8672
rect 11595 8623 11637 8632
rect 11596 8538 11636 8623
rect 11788 8420 11828 10692
rect 12124 10672 12232 10692
rect 13304 10672 13384 10752
rect 14456 10672 14536 10752
rect 15608 10672 15688 10752
rect 16760 10688 16840 10752
rect 16760 10672 16780 10688
rect 12124 10648 12212 10672
rect 12843 10520 12885 10529
rect 12843 10480 12844 10520
rect 12884 10480 12885 10520
rect 12843 10471 12885 10480
rect 12747 9512 12789 9521
rect 12747 9472 12748 9512
rect 12788 9472 12789 9512
rect 12747 9463 12789 9472
rect 12748 9378 12788 9463
rect 12844 9428 12884 10471
rect 13132 9512 13172 9521
rect 13132 9428 13172 9472
rect 12844 9388 13172 9428
rect 12747 8840 12789 8849
rect 12747 8800 12748 8840
rect 12788 8800 12789 8840
rect 12747 8791 12789 8800
rect 12075 8756 12117 8765
rect 12075 8716 12076 8756
rect 12116 8716 12117 8756
rect 12075 8707 12117 8716
rect 12459 8756 12501 8765
rect 12459 8716 12460 8756
rect 12500 8716 12501 8756
rect 12459 8707 12501 8716
rect 12651 8756 12693 8765
rect 12651 8716 12652 8756
rect 12692 8716 12693 8756
rect 12651 8707 12693 8716
rect 12076 8686 12116 8707
rect 11883 8672 11925 8681
rect 11883 8632 11884 8672
rect 11924 8632 11925 8672
rect 11883 8623 11925 8632
rect 11692 8380 11828 8420
rect 11595 8336 11637 8345
rect 11595 8296 11596 8336
rect 11636 8296 11637 8336
rect 11595 8287 11637 8296
rect 11596 7757 11636 8287
rect 11595 7748 11637 7757
rect 11595 7708 11596 7748
rect 11636 7708 11637 7748
rect 11595 7699 11637 7708
rect 11595 7580 11637 7589
rect 11595 7540 11596 7580
rect 11636 7540 11637 7580
rect 11595 7531 11637 7540
rect 11499 7496 11541 7505
rect 11499 7456 11500 7496
rect 11540 7456 11541 7496
rect 11499 7447 11541 7456
rect 11499 7244 11541 7253
rect 11499 7204 11500 7244
rect 11540 7204 11541 7244
rect 11499 7195 11541 7204
rect 11500 7085 11540 7195
rect 11499 7076 11541 7085
rect 11499 7036 11500 7076
rect 11540 7036 11541 7076
rect 11499 7027 11541 7036
rect 11404 6439 11444 6448
rect 11499 6488 11541 6497
rect 11499 6448 11500 6488
rect 11540 6448 11541 6488
rect 11499 6439 11541 6448
rect 11596 6488 11636 7531
rect 11692 6656 11732 8380
rect 11788 8000 11828 8009
rect 11788 7757 11828 7960
rect 11787 7748 11829 7757
rect 11787 7708 11788 7748
rect 11828 7708 11829 7748
rect 11787 7699 11829 7708
rect 11884 7421 11924 8623
rect 12076 8621 12116 8646
rect 12460 8672 12500 8707
rect 12460 8621 12500 8632
rect 12556 8672 12596 8681
rect 12268 8504 12308 8513
rect 12075 8000 12117 8009
rect 12172 8000 12212 8009
rect 12075 7960 12076 8000
rect 12116 7960 12172 8000
rect 12075 7951 12117 7960
rect 12172 7951 12212 7960
rect 11883 7412 11925 7421
rect 11883 7372 11884 7412
rect 11924 7372 11925 7412
rect 11883 7363 11925 7372
rect 11884 7160 11924 7171
rect 11884 7085 11924 7120
rect 11883 7076 11925 7085
rect 11883 7036 11884 7076
rect 11924 7036 11925 7076
rect 11883 7027 11925 7036
rect 11883 6908 11925 6917
rect 11883 6868 11884 6908
rect 11924 6868 11925 6908
rect 11883 6859 11925 6868
rect 11787 6824 11829 6833
rect 11787 6784 11788 6824
rect 11828 6784 11829 6824
rect 11787 6775 11829 6784
rect 11692 6607 11732 6616
rect 11596 6439 11636 6448
rect 10827 6404 10869 6413
rect 10827 6364 10828 6404
rect 10868 6364 10869 6404
rect 10827 6355 10869 6364
rect 11307 6404 11349 6413
rect 11307 6364 11308 6404
rect 11348 6364 11349 6404
rect 11307 6355 11349 6364
rect 11020 6236 11060 6245
rect 10444 4927 10484 4936
rect 10540 5648 10580 5657
rect 10155 4808 10197 4817
rect 10155 4768 10156 4808
rect 10196 4768 10197 4808
rect 10155 4759 10197 4768
rect 10059 4388 10101 4397
rect 10059 4348 10060 4388
rect 10100 4348 10101 4388
rect 10059 4339 10101 4348
rect 9963 4136 10005 4145
rect 9963 4096 9964 4136
rect 10004 4096 10005 4136
rect 9963 4087 10005 4096
rect 10348 4136 10388 4927
rect 10540 4901 10580 5608
rect 10924 5648 10964 5657
rect 10635 5480 10677 5489
rect 10635 5440 10636 5480
rect 10676 5440 10677 5480
rect 10635 5431 10677 5440
rect 10636 5346 10676 5431
rect 10539 4892 10581 4901
rect 10539 4852 10540 4892
rect 10580 4852 10581 4892
rect 10539 4843 10581 4852
rect 10924 4817 10964 5608
rect 10923 4808 10965 4817
rect 10923 4768 10924 4808
rect 10964 4768 10965 4808
rect 10923 4759 10965 4768
rect 10924 4565 10964 4759
rect 10923 4556 10965 4565
rect 10923 4516 10924 4556
rect 10964 4516 10965 4556
rect 10923 4507 10965 4516
rect 10444 4136 10484 4145
rect 10348 4096 10444 4136
rect 10252 3464 10292 3473
rect 10348 3464 10388 4096
rect 10444 4087 10484 4096
rect 10827 4136 10869 4145
rect 10827 4096 10828 4136
rect 10868 4096 10869 4136
rect 10827 4087 10869 4096
rect 10828 4002 10868 4087
rect 10636 3968 10676 3977
rect 10636 3725 10676 3928
rect 10635 3716 10677 3725
rect 10635 3676 10636 3716
rect 10676 3676 10677 3716
rect 10635 3667 10677 3676
rect 10444 3548 10484 3557
rect 10484 3508 10772 3548
rect 10444 3499 10484 3508
rect 10292 3424 10388 3464
rect 10732 3464 10772 3508
rect 10252 3415 10292 3424
rect 10732 3415 10772 3424
rect 10828 3464 10868 3473
rect 10059 3044 10101 3053
rect 10059 3004 10060 3044
rect 10100 3004 10101 3044
rect 10059 2995 10101 3004
rect 10060 2633 10100 2995
rect 10828 2960 10868 3424
rect 10156 2920 10868 2960
rect 10059 2624 10101 2633
rect 10059 2584 10060 2624
rect 10100 2584 10101 2624
rect 10059 2575 10101 2584
rect 9772 2500 10004 2540
rect 9771 2372 9813 2381
rect 9771 2332 9772 2372
rect 9812 2332 9813 2372
rect 9771 2323 9813 2332
rect 9772 1952 9812 2323
rect 9964 2288 10004 2500
rect 9964 2248 10100 2288
rect 9963 2120 10005 2129
rect 9963 2080 9964 2120
rect 10004 2080 10005 2120
rect 9963 2071 10005 2080
rect 9772 1903 9812 1912
rect 9867 1952 9909 1961
rect 9867 1912 9868 1952
rect 9908 1912 9909 1952
rect 9867 1903 9909 1912
rect 9964 1952 10004 2071
rect 9964 1903 10004 1912
rect 10060 1952 10100 2248
rect 10060 1903 10100 1912
rect 9868 1818 9908 1903
rect 10059 1784 10101 1793
rect 10059 1744 10060 1784
rect 10100 1744 10101 1784
rect 10059 1735 10101 1744
rect 9676 1576 9908 1616
rect 9483 1448 9525 1457
rect 9483 1408 9484 1448
rect 9524 1408 9525 1448
rect 9483 1399 9525 1408
rect 9771 1448 9813 1457
rect 9771 1408 9772 1448
rect 9812 1408 9813 1448
rect 9771 1399 9813 1408
rect 9196 1063 9236 1072
rect 7468 1028 7508 1037
rect 6796 944 6836 953
rect 7468 944 7508 988
rect 7948 978 7988 1063
rect 9387 1028 9429 1037
rect 9387 988 9388 1028
rect 9428 988 9429 1028
rect 9387 979 9429 988
rect 6836 904 7508 944
rect 6796 895 6836 904
rect 9388 894 9428 979
rect 6603 776 6645 785
rect 6603 736 6604 776
rect 6644 736 6645 776
rect 6603 727 6645 736
rect 5355 104 5397 113
rect 5355 64 5356 104
rect 5396 64 5397 104
rect 5355 55 5397 64
rect 5643 104 5685 113
rect 5643 64 5644 104
rect 5684 64 5685 104
rect 5643 55 5685 64
rect 6507 104 6549 113
rect 6507 64 6508 104
rect 6548 64 6549 104
rect 9484 80 9524 1399
rect 9675 1112 9717 1121
rect 9675 1072 9676 1112
rect 9716 1072 9717 1112
rect 9675 1063 9717 1072
rect 9772 1112 9812 1399
rect 9772 1063 9812 1072
rect 9676 978 9716 1063
rect 9675 860 9717 869
rect 9675 820 9676 860
rect 9716 820 9717 860
rect 9675 811 9717 820
rect 9676 80 9716 811
rect 9868 80 9908 1576
rect 10060 80 10100 1735
rect 10156 1112 10196 2920
rect 11020 2876 11060 6196
rect 11115 6236 11157 6245
rect 11115 6196 11116 6236
rect 11156 6196 11157 6236
rect 11115 6187 11157 6196
rect 10540 2836 11060 2876
rect 10540 2624 10580 2836
rect 11116 2801 11156 6187
rect 11308 4985 11348 6355
rect 11500 6354 11540 6439
rect 11595 5732 11637 5741
rect 11595 5692 11596 5732
rect 11636 5692 11637 5732
rect 11595 5683 11637 5692
rect 11499 5144 11541 5153
rect 11499 5104 11500 5144
rect 11540 5104 11541 5144
rect 11499 5095 11541 5104
rect 11403 5060 11445 5069
rect 11403 5020 11404 5060
rect 11444 5020 11445 5060
rect 11403 5011 11445 5020
rect 11307 4976 11349 4985
rect 11307 4936 11308 4976
rect 11348 4936 11349 4976
rect 11307 4927 11349 4936
rect 11404 4901 11444 5011
rect 11403 4892 11445 4901
rect 11403 4852 11404 4892
rect 11444 4852 11445 4892
rect 11403 4843 11445 4852
rect 11308 3464 11348 3492
rect 11403 3464 11445 3473
rect 11348 3424 11404 3464
rect 11444 3424 11445 3464
rect 11308 3415 11348 3424
rect 11403 3415 11445 3424
rect 11212 3380 11252 3389
rect 11115 2792 11157 2801
rect 11020 2752 11116 2792
rect 11156 2752 11157 2792
rect 10635 2708 10677 2717
rect 10635 2668 10636 2708
rect 10676 2668 10677 2708
rect 10635 2659 10677 2668
rect 11020 2708 11060 2752
rect 11115 2743 11157 2752
rect 11212 2717 11252 3340
rect 11403 3044 11445 3053
rect 11403 3004 11404 3044
rect 11444 3004 11445 3044
rect 11403 2995 11445 3004
rect 11020 2659 11060 2668
rect 11211 2708 11253 2717
rect 11211 2668 11212 2708
rect 11252 2668 11253 2708
rect 11211 2659 11253 2668
rect 10540 2575 10580 2584
rect 10636 2624 10676 2659
rect 11404 2633 11444 2995
rect 10636 2573 10676 2584
rect 11116 2624 11156 2633
rect 11116 2540 11156 2584
rect 11403 2624 11445 2633
rect 11403 2584 11404 2624
rect 11444 2584 11445 2624
rect 11403 2575 11445 2584
rect 11116 2500 11348 2540
rect 10252 2456 10292 2465
rect 10292 2416 11252 2456
rect 10252 2407 10292 2416
rect 10539 2204 10581 2213
rect 10539 2164 10540 2204
rect 10580 2164 10581 2204
rect 10539 2155 10581 2164
rect 10251 2120 10293 2129
rect 10251 2080 10252 2120
rect 10292 2080 10293 2120
rect 10251 2071 10293 2080
rect 10252 1986 10292 2071
rect 10444 1952 10484 1961
rect 10347 1700 10389 1709
rect 10347 1660 10348 1700
rect 10388 1660 10389 1700
rect 10347 1651 10389 1660
rect 10251 1196 10293 1205
rect 10251 1156 10252 1196
rect 10292 1156 10293 1196
rect 10251 1147 10293 1156
rect 10156 869 10196 1072
rect 10252 1062 10292 1147
rect 10348 1112 10388 1651
rect 10444 1289 10484 1912
rect 10540 1952 10580 2155
rect 10540 1903 10580 1912
rect 10828 1952 10868 1961
rect 10635 1868 10677 1877
rect 10635 1828 10636 1868
rect 10676 1828 10677 1868
rect 10635 1819 10677 1828
rect 10539 1700 10581 1709
rect 10539 1660 10540 1700
rect 10580 1660 10581 1700
rect 10539 1651 10581 1660
rect 10443 1280 10485 1289
rect 10443 1240 10444 1280
rect 10484 1240 10485 1280
rect 10443 1231 10485 1240
rect 10348 1072 10484 1112
rect 10155 860 10197 869
rect 10155 820 10156 860
rect 10196 820 10197 860
rect 10155 811 10197 820
rect 10251 608 10293 617
rect 10251 568 10252 608
rect 10292 568 10293 608
rect 10251 559 10293 568
rect 10252 80 10292 559
rect 10444 80 10484 1072
rect 10540 776 10580 1651
rect 10636 860 10676 1819
rect 10731 1112 10773 1121
rect 10731 1072 10732 1112
rect 10772 1072 10773 1112
rect 10731 1063 10773 1072
rect 10732 978 10772 1063
rect 10828 1037 10868 1912
rect 10924 1952 10964 1961
rect 10924 1457 10964 1912
rect 11115 1532 11157 1541
rect 11115 1492 11116 1532
rect 11156 1492 11157 1532
rect 11115 1483 11157 1492
rect 10923 1448 10965 1457
rect 10923 1408 10924 1448
rect 10964 1408 10965 1448
rect 10923 1399 10965 1408
rect 10923 1280 10965 1289
rect 10923 1240 10924 1280
rect 10964 1240 10965 1280
rect 10923 1231 10965 1240
rect 10827 1028 10869 1037
rect 10827 988 10828 1028
rect 10868 988 10869 1028
rect 10827 979 10869 988
rect 10636 820 10868 860
rect 10540 736 10676 776
rect 10636 80 10676 736
rect 10828 80 10868 820
rect 10924 785 10964 1231
rect 11116 1028 11156 1483
rect 11212 1126 11252 2416
rect 11308 1868 11348 2500
rect 11404 1952 11444 1961
rect 11500 1952 11540 5095
rect 11596 4640 11636 5683
rect 11691 4976 11733 4985
rect 11691 4936 11692 4976
rect 11732 4936 11733 4976
rect 11691 4927 11733 4936
rect 11692 4842 11732 4927
rect 11596 4600 11732 4640
rect 11595 3212 11637 3221
rect 11595 3172 11596 3212
rect 11636 3172 11637 3212
rect 11595 3163 11637 3172
rect 11596 2624 11636 3163
rect 11596 2575 11636 2584
rect 11444 1912 11540 1952
rect 11692 1952 11732 4600
rect 11788 3464 11828 6775
rect 11884 6749 11924 6859
rect 11883 6740 11925 6749
rect 11883 6700 11884 6740
rect 11924 6700 11925 6740
rect 11883 6691 11925 6700
rect 11884 6488 11924 6691
rect 11884 6439 11924 6448
rect 12076 6320 12116 7951
rect 12268 6497 12308 8464
rect 12556 8345 12596 8632
rect 12652 8513 12692 8707
rect 12651 8504 12693 8513
rect 12651 8464 12652 8504
rect 12692 8464 12693 8504
rect 12651 8455 12693 8464
rect 12748 8504 12788 8791
rect 12748 8455 12788 8464
rect 12555 8336 12597 8345
rect 12555 8296 12556 8336
rect 12596 8296 12597 8336
rect 12555 8287 12597 8296
rect 12363 7412 12405 7421
rect 12363 7372 12364 7412
rect 12404 7372 12405 7412
rect 12363 7363 12405 7372
rect 12267 6488 12309 6497
rect 12267 6448 12268 6488
rect 12308 6448 12309 6488
rect 12267 6439 12309 6448
rect 11884 6280 12116 6320
rect 12171 6320 12213 6329
rect 12171 6280 12172 6320
rect 12212 6280 12213 6320
rect 11884 5069 11924 6280
rect 12171 6271 12213 6280
rect 12172 5648 12212 6271
rect 12364 5732 12404 7363
rect 12747 6068 12789 6077
rect 12747 6028 12748 6068
rect 12788 6028 12789 6068
rect 12747 6019 12789 6028
rect 11980 5608 12172 5648
rect 11883 5060 11925 5069
rect 11883 5020 11884 5060
rect 11924 5020 11925 5060
rect 11883 5011 11925 5020
rect 11980 4808 12020 5608
rect 12172 5599 12212 5608
rect 12268 5692 12404 5732
rect 12268 5321 12308 5692
rect 12652 5648 12692 5657
rect 12364 5564 12404 5573
rect 12652 5564 12692 5608
rect 12404 5524 12692 5564
rect 12748 5648 12788 6019
rect 12364 5515 12404 5524
rect 12555 5396 12597 5405
rect 12555 5356 12556 5396
rect 12596 5356 12597 5396
rect 12555 5347 12597 5356
rect 12267 5312 12309 5321
rect 12267 5272 12268 5312
rect 12308 5272 12309 5312
rect 12267 5263 12309 5272
rect 12459 5312 12501 5321
rect 12459 5272 12460 5312
rect 12500 5272 12501 5312
rect 12459 5263 12501 5272
rect 12076 4985 12116 5070
rect 12075 4976 12117 4985
rect 12075 4936 12076 4976
rect 12116 4936 12117 4976
rect 12075 4927 12117 4936
rect 12172 4976 12212 4985
rect 11980 4768 12116 4808
rect 11884 4724 11924 4733
rect 11924 4684 12020 4724
rect 11884 4675 11924 4684
rect 11883 4472 11925 4481
rect 11883 4432 11884 4472
rect 11924 4432 11925 4472
rect 11883 4423 11925 4432
rect 11788 3415 11828 3424
rect 11787 3044 11829 3053
rect 11787 3004 11788 3044
rect 11828 3004 11829 3044
rect 11787 2995 11829 3004
rect 11788 2717 11828 2995
rect 11884 2792 11924 4423
rect 11980 3716 12020 4684
rect 12076 4136 12116 4768
rect 12076 4087 12116 4096
rect 11980 3676 12116 3716
rect 11979 2792 12021 2801
rect 11884 2752 11980 2792
rect 12020 2752 12021 2792
rect 11979 2743 12021 2752
rect 11787 2708 11829 2717
rect 11787 2668 11788 2708
rect 11828 2668 11829 2708
rect 11787 2659 11829 2668
rect 11884 1952 11924 1961
rect 11692 1912 11884 1952
rect 11404 1903 11444 1912
rect 11884 1903 11924 1912
rect 11308 1793 11348 1828
rect 11307 1784 11349 1793
rect 11307 1744 11308 1784
rect 11348 1744 11349 1784
rect 11307 1735 11349 1744
rect 11691 1784 11733 1793
rect 11691 1744 11692 1784
rect 11732 1744 11733 1784
rect 11691 1735 11733 1744
rect 11212 1077 11252 1086
rect 11595 1112 11637 1121
rect 11595 1072 11596 1112
rect 11636 1072 11637 1112
rect 11595 1063 11637 1072
rect 11403 1028 11445 1037
rect 11116 988 11252 1028
rect 11019 944 11061 953
rect 11019 904 11020 944
rect 11060 904 11061 944
rect 11019 895 11061 904
rect 10923 776 10965 785
rect 10923 736 10924 776
rect 10964 736 10965 776
rect 10923 727 10965 736
rect 11020 80 11060 895
rect 11212 80 11252 988
rect 11403 988 11404 1028
rect 11444 988 11445 1028
rect 11403 979 11445 988
rect 11404 894 11444 979
rect 11596 978 11636 1063
rect 11692 860 11732 1735
rect 11787 1532 11829 1541
rect 11787 1492 11788 1532
rect 11828 1492 11829 1532
rect 11787 1483 11829 1492
rect 11596 820 11732 860
rect 11403 104 11445 113
rect 11403 80 11404 104
rect 6507 55 6549 64
rect 9464 0 9544 80
rect 9656 0 9736 80
rect 9848 0 9928 80
rect 10040 0 10120 80
rect 10232 0 10312 80
rect 10424 0 10504 80
rect 10616 0 10696 80
rect 10808 0 10888 80
rect 11000 0 11080 80
rect 11192 0 11272 80
rect 11384 64 11404 80
rect 11444 80 11445 104
rect 11596 80 11636 820
rect 11788 80 11828 1483
rect 11980 1289 12020 2743
rect 12076 2638 12116 3676
rect 12076 2589 12116 2598
rect 12075 2120 12117 2129
rect 12075 2080 12076 2120
rect 12116 2080 12117 2120
rect 12075 2071 12117 2080
rect 11979 1280 12021 1289
rect 11979 1240 11980 1280
rect 12020 1240 12021 1280
rect 11979 1231 12021 1240
rect 12076 1126 12116 2071
rect 12172 1625 12212 4936
rect 12268 4976 12308 4985
rect 12268 4481 12308 4936
rect 12364 4976 12404 4985
rect 12267 4472 12309 4481
rect 12267 4432 12268 4472
rect 12308 4432 12309 4472
rect 12267 4423 12309 4432
rect 12267 3968 12309 3977
rect 12267 3928 12268 3968
rect 12308 3928 12309 3968
rect 12267 3919 12309 3928
rect 12268 3834 12308 3919
rect 12364 3809 12404 4936
rect 12460 4724 12500 5263
rect 12556 4985 12596 5347
rect 12555 4976 12597 4985
rect 12555 4936 12556 4976
rect 12596 4936 12597 4976
rect 12555 4927 12597 4936
rect 12556 4842 12596 4927
rect 12460 4684 12596 4724
rect 12460 4136 12500 4145
rect 12363 3800 12405 3809
rect 12363 3760 12364 3800
rect 12404 3760 12405 3800
rect 12363 3751 12405 3760
rect 12460 3725 12500 4096
rect 12267 3716 12309 3725
rect 12267 3676 12268 3716
rect 12308 3676 12309 3716
rect 12267 3667 12309 3676
rect 12459 3716 12501 3725
rect 12459 3676 12460 3716
rect 12500 3676 12501 3716
rect 12459 3667 12501 3676
rect 12268 3459 12308 3667
rect 12268 3410 12308 3419
rect 12460 3548 12500 3557
rect 12460 3389 12500 3508
rect 12459 3380 12501 3389
rect 12459 3340 12460 3380
rect 12500 3340 12501 3380
rect 12459 3331 12501 3340
rect 12267 2708 12309 2717
rect 12267 2668 12268 2708
rect 12308 2668 12309 2708
rect 12267 2659 12309 2668
rect 12268 2540 12308 2659
rect 12460 2633 12500 2718
rect 12459 2624 12501 2633
rect 12459 2584 12460 2624
rect 12500 2584 12501 2624
rect 12459 2575 12501 2584
rect 12268 2491 12308 2500
rect 12556 2204 12596 4684
rect 12651 3380 12693 3389
rect 12651 3340 12652 3380
rect 12692 3340 12693 3380
rect 12651 3331 12693 3340
rect 12652 3246 12692 3331
rect 12748 2381 12788 5608
rect 12844 4313 12884 9388
rect 12940 9260 12980 9269
rect 12980 9220 13076 9260
rect 12940 9211 12980 9220
rect 12939 8840 12981 8849
rect 12939 8800 12940 8840
rect 12980 8800 12981 8840
rect 12939 8791 12981 8800
rect 12940 8504 12980 8791
rect 13036 8681 13076 9220
rect 13035 8672 13077 8681
rect 13035 8632 13036 8672
rect 13076 8632 13077 8672
rect 13035 8623 13077 8632
rect 13132 8672 13172 8681
rect 12940 8455 12980 8464
rect 13132 8345 13172 8632
rect 13228 8672 13268 8683
rect 13228 8597 13268 8632
rect 13227 8588 13269 8597
rect 13227 8548 13228 8588
rect 13268 8548 13269 8588
rect 13227 8539 13269 8548
rect 12939 8336 12981 8345
rect 12939 8296 12940 8336
rect 12980 8296 12981 8336
rect 12939 8287 12981 8296
rect 13131 8336 13173 8345
rect 13131 8296 13132 8336
rect 13172 8296 13173 8336
rect 13131 8287 13173 8296
rect 12940 5825 12980 8287
rect 13132 7160 13172 7169
rect 13324 7160 13364 10672
rect 13419 9680 13461 9689
rect 13419 9640 13420 9680
rect 13460 9640 13461 9680
rect 13419 9631 13461 9640
rect 13420 8336 13460 9631
rect 14283 9512 14325 9521
rect 14380 9512 14420 9521
rect 14283 9472 14284 9512
rect 14324 9472 14380 9512
rect 14283 9463 14325 9472
rect 14380 9463 14420 9472
rect 14091 9176 14133 9185
rect 14091 9136 14092 9176
rect 14132 9136 14133 9176
rect 14091 9127 14133 9136
rect 13707 8924 13749 8933
rect 13707 8884 13708 8924
rect 13748 8884 13749 8924
rect 13707 8875 13749 8884
rect 13611 8756 13653 8765
rect 13611 8716 13612 8756
rect 13652 8716 13653 8756
rect 13611 8707 13653 8716
rect 13515 8672 13557 8681
rect 13515 8632 13516 8672
rect 13556 8632 13557 8672
rect 13515 8623 13557 8632
rect 13612 8672 13652 8707
rect 13516 8538 13556 8623
rect 13612 8621 13652 8632
rect 13611 8504 13653 8513
rect 13611 8464 13612 8504
rect 13652 8464 13653 8504
rect 13611 8455 13653 8464
rect 13420 8296 13556 8336
rect 13419 8168 13461 8177
rect 13419 8128 13420 8168
rect 13460 8128 13461 8168
rect 13419 8119 13461 8128
rect 13420 8000 13460 8119
rect 13516 8000 13556 8296
rect 13612 8168 13652 8455
rect 13612 8119 13652 8128
rect 13516 7960 13652 8000
rect 13420 7951 13460 7960
rect 13515 7328 13557 7337
rect 13515 7288 13516 7328
rect 13556 7288 13557 7328
rect 13515 7279 13557 7288
rect 13132 6749 13172 7120
rect 13228 7120 13364 7160
rect 13516 7160 13556 7279
rect 13228 6824 13268 7120
rect 13516 7111 13556 7120
rect 13612 7076 13652 7960
rect 13708 7832 13748 8875
rect 13899 8672 13941 8681
rect 13899 8632 13900 8672
rect 13940 8632 13941 8672
rect 13899 8623 13941 8632
rect 13996 8672 14036 8681
rect 13804 8009 13844 8094
rect 13803 8000 13845 8009
rect 13803 7960 13804 8000
rect 13844 7960 13845 8000
rect 13803 7951 13845 7960
rect 13900 7925 13940 8623
rect 13996 8429 14036 8632
rect 14092 8672 14132 9127
rect 14187 8840 14229 8849
rect 14187 8800 14188 8840
rect 14228 8800 14229 8840
rect 14187 8791 14229 8800
rect 14092 8513 14132 8632
rect 14091 8504 14133 8513
rect 14091 8464 14092 8504
rect 14132 8464 14133 8504
rect 14091 8455 14133 8464
rect 13995 8420 14037 8429
rect 13995 8380 13996 8420
rect 14036 8380 14037 8420
rect 13995 8371 14037 8380
rect 13899 7916 13941 7925
rect 13899 7876 13900 7916
rect 13940 7876 13941 7916
rect 13899 7867 13941 7876
rect 13708 7792 13844 7832
rect 13707 7160 13749 7169
rect 13707 7120 13708 7160
rect 13748 7120 13749 7160
rect 13707 7111 13749 7120
rect 13804 7160 13844 7792
rect 13900 7160 13940 7867
rect 13996 7421 14036 8371
rect 14188 7832 14228 8791
rect 14284 8177 14324 9463
rect 14476 9344 14516 10672
rect 15628 9596 15668 10672
rect 16779 10648 16780 10672
rect 16820 10672 16840 10688
rect 17912 10672 17992 10752
rect 19064 10732 19144 10752
rect 19064 10692 19988 10732
rect 19064 10672 19172 10692
rect 16820 10648 16821 10672
rect 16779 10639 16821 10648
rect 15628 9556 15764 9596
rect 14763 9512 14805 9521
rect 14763 9472 14764 9512
rect 14804 9472 14805 9512
rect 14763 9463 14805 9472
rect 14764 9378 14804 9463
rect 14380 9304 14516 9344
rect 14283 8168 14325 8177
rect 14283 8128 14284 8168
rect 14324 8128 14325 8168
rect 14283 8119 14325 8128
rect 14283 8000 14325 8009
rect 14283 7960 14284 8000
rect 14324 7960 14325 8000
rect 14283 7951 14325 7960
rect 14092 7792 14228 7832
rect 13995 7412 14037 7421
rect 13995 7372 13996 7412
rect 14036 7372 14037 7412
rect 13995 7363 14037 7372
rect 13996 7160 14036 7169
rect 13900 7120 13996 7160
rect 13804 7111 13844 7120
rect 13996 7111 14036 7120
rect 14092 7160 14132 7792
rect 14187 7580 14229 7589
rect 14187 7540 14188 7580
rect 14228 7540 14229 7580
rect 14187 7531 14229 7540
rect 14092 7111 14132 7120
rect 14188 7160 14228 7531
rect 14188 7111 14228 7120
rect 14284 7160 14324 7951
rect 14380 7841 14420 9304
rect 14572 9260 14612 9269
rect 14476 9220 14572 9260
rect 14476 8681 14516 9220
rect 14572 9211 14612 9220
rect 14475 8672 14517 8681
rect 14475 8632 14476 8672
rect 14516 8632 14517 8672
rect 14475 8623 14517 8632
rect 14572 8672 14612 8681
rect 15052 8677 15092 8686
rect 15436 8681 15476 8766
rect 14612 8632 14708 8672
rect 14572 8623 14612 8632
rect 14379 7832 14421 7841
rect 14379 7792 14380 7832
rect 14420 7792 14421 7832
rect 14379 7783 14421 7792
rect 14476 7589 14516 8623
rect 14571 8504 14613 8513
rect 14571 8464 14572 8504
rect 14612 8464 14613 8504
rect 14571 8455 14613 8464
rect 14475 7580 14517 7589
rect 14475 7540 14476 7580
rect 14516 7540 14517 7580
rect 14475 7531 14517 7540
rect 14379 7412 14421 7421
rect 14379 7372 14380 7412
rect 14420 7372 14421 7412
rect 14379 7363 14421 7372
rect 14284 7111 14324 7120
rect 13612 7027 13652 7036
rect 13708 7026 13748 7111
rect 13324 6992 13364 7001
rect 13364 6952 13556 6992
rect 13324 6943 13364 6952
rect 13228 6784 13460 6824
rect 13131 6740 13173 6749
rect 13036 6700 13132 6740
rect 13172 6700 13173 6740
rect 13036 6329 13076 6700
rect 13131 6691 13173 6700
rect 13132 6581 13172 6612
rect 13131 6572 13173 6581
rect 13131 6532 13132 6572
rect 13172 6532 13173 6572
rect 13131 6523 13173 6532
rect 13132 6488 13172 6523
rect 13035 6320 13077 6329
rect 13035 6280 13036 6320
rect 13076 6280 13077 6320
rect 13035 6271 13077 6280
rect 13132 6152 13172 6448
rect 13323 6236 13365 6245
rect 13323 6196 13324 6236
rect 13364 6196 13365 6236
rect 13323 6187 13365 6196
rect 13036 6112 13172 6152
rect 12939 5816 12981 5825
rect 12939 5776 12940 5816
rect 12980 5776 12981 5816
rect 12939 5767 12981 5776
rect 12843 4304 12885 4313
rect 12843 4264 12844 4304
rect 12884 4264 12885 4304
rect 12843 4255 12885 4264
rect 13036 3725 13076 6112
rect 13324 6102 13364 6187
rect 13227 5816 13269 5825
rect 13227 5776 13228 5816
rect 13268 5776 13269 5816
rect 13227 5767 13269 5776
rect 13228 5732 13268 5767
rect 13132 5648 13172 5657
rect 13132 5405 13172 5608
rect 13131 5396 13173 5405
rect 13131 5356 13132 5396
rect 13172 5356 13173 5396
rect 13131 5347 13173 5356
rect 13228 4976 13268 5692
rect 13420 5237 13460 6784
rect 13516 6488 13556 6952
rect 13803 6740 13845 6749
rect 13803 6700 13804 6740
rect 13844 6700 13845 6740
rect 13803 6691 13845 6700
rect 13612 6488 13652 6497
rect 13516 6448 13612 6488
rect 13612 6439 13652 6448
rect 13708 6488 13748 6497
rect 13708 6161 13748 6448
rect 13707 6152 13749 6161
rect 13707 6112 13708 6152
rect 13748 6112 13749 6152
rect 13707 6103 13749 6112
rect 13708 5900 13748 6103
rect 13612 5860 13748 5900
rect 13419 5228 13461 5237
rect 13419 5188 13420 5228
rect 13460 5188 13461 5228
rect 13419 5179 13461 5188
rect 13228 4936 13364 4976
rect 13227 4808 13269 4817
rect 13227 4768 13228 4808
rect 13268 4768 13269 4808
rect 13227 4759 13269 4768
rect 13131 3968 13173 3977
rect 13131 3928 13132 3968
rect 13172 3928 13173 3968
rect 13131 3919 13173 3928
rect 13035 3716 13077 3725
rect 13035 3676 13036 3716
rect 13076 3676 13077 3716
rect 13035 3667 13077 3676
rect 12939 3296 12981 3305
rect 12939 3256 12940 3296
rect 12980 3256 12981 3296
rect 12939 3247 12981 3256
rect 12844 3212 12884 3221
rect 12844 2465 12884 3172
rect 12940 2885 12980 3247
rect 12939 2876 12981 2885
rect 12939 2836 12940 2876
rect 12980 2836 12981 2876
rect 12939 2827 12981 2836
rect 13036 2633 13076 3667
rect 13132 3464 13172 3919
rect 13132 3415 13172 3424
rect 13228 3464 13268 4759
rect 13268 3424 13273 3464
rect 13228 3415 13273 3424
rect 13233 3296 13273 3415
rect 13132 3256 13273 3296
rect 13035 2624 13077 2633
rect 13035 2584 13036 2624
rect 13076 2584 13077 2624
rect 13035 2575 13077 2584
rect 12843 2456 12885 2465
rect 12843 2416 12844 2456
rect 12884 2416 12885 2456
rect 12843 2407 12885 2416
rect 12747 2372 12789 2381
rect 12747 2332 12748 2372
rect 12788 2332 12789 2372
rect 12747 2323 12789 2332
rect 12843 2288 12885 2297
rect 12843 2248 12844 2288
rect 12884 2248 12885 2288
rect 12843 2239 12885 2248
rect 13035 2288 13077 2297
rect 13035 2248 13036 2288
rect 13076 2248 13077 2288
rect 13035 2239 13077 2248
rect 12460 2164 12596 2204
rect 12364 1938 12404 1947
rect 12171 1616 12213 1625
rect 12171 1576 12172 1616
rect 12212 1576 12213 1616
rect 12171 1567 12213 1576
rect 12364 1289 12404 1898
rect 12171 1280 12213 1289
rect 12171 1240 12172 1280
rect 12212 1240 12213 1280
rect 12171 1231 12213 1240
rect 12363 1280 12405 1289
rect 12363 1240 12364 1280
rect 12404 1240 12405 1280
rect 12363 1231 12405 1240
rect 11980 1086 12116 1126
rect 11980 80 12020 1086
rect 12172 80 12212 1231
rect 12460 1126 12500 2164
rect 12748 2045 12788 2130
rect 12556 2036 12596 2045
rect 12747 2036 12789 2045
rect 12596 1996 12692 2036
rect 12556 1987 12596 1996
rect 12652 1877 12692 1996
rect 12747 1996 12748 2036
rect 12788 1996 12789 2036
rect 12747 1987 12789 1996
rect 12844 1973 12884 2239
rect 12844 1924 12884 1933
rect 12939 1952 12981 1961
rect 12939 1912 12940 1952
rect 12980 1912 12981 1952
rect 12939 1903 12981 1912
rect 13036 1952 13076 2239
rect 13036 1903 13076 1912
rect 12651 1868 12693 1877
rect 12651 1828 12652 1868
rect 12692 1828 12693 1868
rect 12651 1819 12693 1828
rect 12940 1818 12980 1903
rect 12747 1364 12789 1373
rect 12747 1324 12748 1364
rect 12788 1324 12789 1364
rect 12747 1315 12789 1324
rect 12364 1086 12500 1126
rect 12364 80 12404 1086
rect 12555 608 12597 617
rect 12555 568 12556 608
rect 12596 568 12597 608
rect 12555 559 12597 568
rect 12556 80 12596 559
rect 12748 80 12788 1315
rect 13132 1280 13172 3256
rect 13227 2876 13269 2885
rect 13227 2836 13228 2876
rect 13268 2836 13269 2876
rect 13227 2827 13269 2836
rect 13228 2120 13268 2827
rect 13228 2071 13268 2080
rect 13324 1373 13364 4936
rect 13612 4901 13652 5860
rect 13707 5732 13749 5741
rect 13707 5692 13708 5732
rect 13748 5692 13749 5732
rect 13707 5683 13749 5692
rect 13708 5648 13748 5683
rect 13708 5597 13748 5608
rect 13804 4976 13844 6691
rect 14092 6404 14132 6413
rect 13611 4892 13653 4901
rect 13611 4852 13612 4892
rect 13652 4852 13653 4892
rect 13611 4843 13653 4852
rect 13611 4640 13653 4649
rect 13611 4600 13612 4640
rect 13652 4600 13653 4640
rect 13611 4591 13653 4600
rect 13612 3464 13652 4591
rect 13708 4136 13748 4145
rect 13804 4136 13844 4936
rect 13900 6364 14092 6404
rect 13900 4145 13940 6364
rect 14092 6355 14132 6364
rect 14188 6404 14228 6413
rect 14380 6404 14420 7363
rect 14475 7160 14517 7169
rect 14475 7120 14476 7160
rect 14516 7120 14517 7160
rect 14475 7111 14517 7120
rect 14476 7026 14516 7111
rect 14228 6364 14420 6404
rect 14188 6355 14228 6364
rect 14188 5653 14228 5662
rect 14188 5312 14228 5613
rect 14188 5272 14231 5312
rect 14191 5228 14231 5272
rect 14188 5188 14231 5228
rect 13996 5144 14036 5153
rect 14188 5144 14228 5188
rect 14036 5104 14228 5144
rect 13996 5095 14036 5104
rect 14284 4985 14324 6364
rect 14475 6236 14517 6245
rect 14475 6196 14476 6236
rect 14516 6196 14517 6236
rect 14475 6187 14517 6196
rect 14380 5480 14420 5489
rect 13995 4976 14037 4985
rect 13995 4936 13996 4976
rect 14036 4936 14037 4976
rect 13995 4927 14037 4936
rect 14283 4976 14325 4985
rect 14283 4936 14284 4976
rect 14324 4936 14325 4976
rect 14283 4927 14325 4936
rect 13748 4096 13844 4136
rect 13899 4136 13941 4145
rect 13899 4096 13900 4136
rect 13940 4096 13941 4136
rect 13708 4087 13748 4096
rect 13899 4087 13941 4096
rect 13899 3968 13941 3977
rect 13899 3928 13900 3968
rect 13940 3928 13941 3968
rect 13899 3919 13941 3928
rect 13900 3834 13940 3919
rect 13612 2465 13652 3424
rect 13708 3380 13748 3389
rect 13748 3340 13844 3380
rect 13708 3331 13748 3340
rect 13708 2633 13748 2719
rect 13707 2624 13749 2633
rect 13707 2584 13708 2624
rect 13748 2584 13749 2624
rect 13707 2575 13749 2584
rect 13611 2456 13653 2465
rect 13611 2416 13612 2456
rect 13652 2416 13653 2456
rect 13611 2407 13653 2416
rect 13419 2372 13461 2381
rect 13419 2332 13420 2372
rect 13460 2332 13461 2372
rect 13419 2323 13461 2332
rect 13420 1952 13460 2323
rect 13420 1903 13460 1912
rect 13420 1784 13460 1793
rect 13420 1625 13460 1744
rect 13419 1616 13461 1625
rect 13419 1576 13420 1616
rect 13460 1576 13461 1616
rect 13419 1567 13461 1576
rect 13420 1457 13460 1567
rect 13419 1448 13461 1457
rect 13419 1408 13420 1448
rect 13460 1408 13461 1448
rect 13419 1399 13461 1408
rect 13323 1364 13365 1373
rect 13323 1324 13324 1364
rect 13364 1324 13365 1364
rect 13323 1315 13365 1324
rect 12940 1240 13172 1280
rect 13227 1280 13269 1289
rect 13227 1240 13228 1280
rect 13268 1240 13269 1280
rect 12843 1112 12885 1121
rect 12843 1072 12844 1112
rect 12884 1072 12885 1112
rect 12843 1063 12885 1072
rect 12844 978 12884 1063
rect 12940 80 12980 1240
rect 13227 1231 13269 1240
rect 13036 1028 13076 1037
rect 13228 1028 13268 1231
rect 13612 1196 13652 2407
rect 13076 988 13268 1028
rect 13324 1156 13652 1196
rect 13036 979 13076 988
rect 13324 944 13364 1156
rect 13708 1121 13748 2575
rect 13804 2129 13844 3340
rect 13899 2792 13941 2801
rect 13899 2752 13900 2792
rect 13940 2752 13941 2792
rect 13899 2743 13941 2752
rect 13900 2633 13940 2743
rect 13899 2624 13941 2633
rect 13899 2584 13900 2624
rect 13940 2584 13941 2624
rect 13899 2575 13941 2584
rect 13900 2456 13940 2465
rect 13803 2120 13845 2129
rect 13803 2080 13804 2120
rect 13844 2080 13845 2120
rect 13803 2071 13845 2080
rect 13804 1784 13844 2071
rect 13900 1952 13940 2416
rect 13900 1903 13940 1912
rect 13996 1952 14036 4927
rect 14283 4640 14325 4649
rect 14283 4600 14284 4640
rect 14324 4600 14325 4640
rect 14283 4591 14325 4600
rect 14188 4136 14228 4145
rect 14188 3968 14228 4096
rect 14284 4136 14324 4591
rect 14380 4229 14420 5440
rect 14379 4220 14421 4229
rect 14379 4180 14380 4220
rect 14420 4180 14421 4220
rect 14379 4171 14421 4180
rect 14284 4087 14324 4096
rect 14476 3968 14516 6187
rect 14572 4313 14612 8455
rect 14668 7337 14708 8632
rect 15052 8597 15092 8637
rect 15435 8672 15477 8681
rect 15435 8632 15436 8672
rect 15476 8632 15477 8672
rect 15435 8623 15477 8632
rect 15532 8672 15572 8681
rect 15051 8588 15093 8597
rect 15051 8548 15052 8588
rect 15092 8548 15093 8588
rect 15051 8539 15093 8548
rect 15244 8504 15284 8513
rect 15532 8504 15572 8632
rect 15284 8464 15572 8504
rect 15628 8672 15668 8681
rect 15244 8455 15284 8464
rect 15339 8168 15381 8177
rect 15339 8128 15340 8168
rect 15380 8128 15381 8168
rect 15628 8168 15668 8632
rect 15724 8672 15764 9556
rect 16011 9512 16053 9521
rect 16011 9472 16012 9512
rect 16052 9472 16053 9512
rect 16011 9463 16053 9472
rect 16396 9512 16436 9523
rect 16012 9378 16052 9463
rect 16396 9437 16436 9472
rect 17451 9512 17493 9521
rect 17451 9472 17452 9512
rect 17492 9472 17493 9512
rect 17451 9463 17493 9472
rect 17643 9512 17685 9521
rect 17643 9472 17644 9512
rect 17684 9472 17685 9512
rect 17643 9463 17685 9472
rect 16395 9428 16437 9437
rect 16395 9388 16396 9428
rect 16436 9388 16437 9428
rect 16395 9379 16437 9388
rect 16203 9260 16245 9269
rect 16203 9220 16204 9260
rect 16244 9220 16245 9260
rect 16203 9211 16245 9220
rect 16587 9260 16629 9269
rect 16587 9220 16588 9260
rect 16628 9220 16629 9260
rect 16587 9211 16629 9220
rect 16204 9126 16244 9211
rect 16299 8840 16341 8849
rect 16299 8800 16300 8840
rect 16340 8800 16341 8840
rect 16299 8791 16341 8800
rect 15724 8623 15764 8632
rect 16203 8672 16245 8681
rect 16203 8632 16204 8672
rect 16244 8632 16245 8672
rect 16203 8623 16245 8632
rect 16107 8588 16149 8597
rect 16107 8548 16108 8588
rect 16148 8548 16149 8588
rect 16107 8539 16149 8548
rect 15724 8168 15764 8177
rect 15628 8128 15724 8168
rect 15339 8119 15381 8128
rect 15724 8119 15764 8128
rect 15052 8000 15092 8009
rect 14667 7328 14709 7337
rect 14667 7288 14668 7328
rect 14708 7288 14709 7328
rect 14667 7279 14709 7288
rect 14955 7328 14997 7337
rect 14955 7288 14956 7328
rect 14996 7288 14997 7328
rect 14955 7279 14997 7288
rect 14668 6488 14708 6497
rect 14668 5321 14708 6448
rect 14956 6329 14996 7279
rect 15052 6749 15092 7960
rect 15244 7748 15284 7757
rect 15340 7748 15380 8119
rect 15435 8000 15477 8009
rect 15435 7960 15436 8000
rect 15476 7960 15477 8000
rect 15435 7951 15477 7960
rect 15532 8000 15572 8009
rect 15916 8000 15956 8009
rect 15572 7960 15916 8000
rect 15532 7951 15572 7960
rect 15916 7951 15956 7960
rect 16012 8000 16052 8011
rect 15436 7866 15476 7951
rect 16012 7925 16052 7960
rect 16108 8000 16148 8539
rect 16204 8538 16244 8623
rect 16108 7951 16148 7960
rect 16204 8000 16244 8009
rect 16011 7916 16053 7925
rect 16011 7876 16012 7916
rect 16052 7876 16053 7916
rect 16011 7867 16053 7876
rect 15340 7708 15476 7748
rect 15051 6740 15093 6749
rect 15051 6700 15052 6740
rect 15092 6700 15093 6740
rect 15051 6691 15093 6700
rect 15244 6488 15284 7708
rect 15339 6572 15381 6581
rect 15339 6532 15340 6572
rect 15380 6532 15381 6572
rect 15339 6523 15381 6532
rect 15196 6478 15284 6488
rect 15236 6448 15284 6478
rect 15340 6438 15380 6523
rect 15196 6429 15236 6438
rect 14955 6320 14997 6329
rect 14955 6280 14956 6320
rect 14996 6280 14997 6320
rect 14955 6271 14997 6280
rect 15436 6245 15476 7708
rect 16107 7412 16149 7421
rect 16107 7372 16108 7412
rect 16148 7372 16149 7412
rect 16107 7363 16149 7372
rect 15724 7160 15764 7169
rect 15724 7085 15764 7120
rect 16108 7160 16148 7363
rect 15723 7076 15765 7085
rect 15723 7036 15724 7076
rect 15764 7036 15765 7076
rect 15723 7027 15765 7036
rect 15627 6992 15669 7001
rect 15627 6952 15628 6992
rect 15668 6952 15669 6992
rect 15627 6943 15669 6952
rect 15435 6236 15477 6245
rect 15435 6196 15436 6236
rect 15476 6196 15477 6236
rect 15435 6187 15477 6196
rect 14667 5312 14709 5321
rect 14667 5272 14668 5312
rect 14708 5272 14709 5312
rect 14667 5263 14709 5272
rect 14859 4976 14901 4985
rect 14859 4936 14860 4976
rect 14900 4936 14901 4976
rect 14859 4927 14901 4936
rect 14860 4397 14900 4927
rect 15628 4817 15668 6943
rect 15724 6665 15764 7027
rect 15916 6992 15956 7001
rect 15820 6952 15916 6992
rect 15723 6656 15765 6665
rect 15723 6616 15724 6656
rect 15764 6616 15765 6656
rect 15723 6607 15765 6616
rect 15724 6404 15764 6413
rect 15724 6245 15764 6364
rect 15723 6236 15765 6245
rect 15723 6196 15724 6236
rect 15764 6196 15765 6236
rect 15723 6187 15765 6196
rect 15627 4808 15669 4817
rect 15627 4768 15628 4808
rect 15668 4768 15669 4808
rect 15627 4759 15669 4768
rect 14859 4388 14901 4397
rect 14859 4348 14860 4388
rect 14900 4348 14901 4388
rect 14859 4339 14901 4348
rect 14571 4304 14613 4313
rect 14571 4264 14572 4304
rect 14612 4264 14613 4304
rect 14571 4255 14613 4264
rect 15820 4220 15860 6952
rect 15916 6943 15956 6952
rect 16108 6917 16148 7120
rect 16204 7001 16244 7960
rect 16203 6992 16245 7001
rect 16203 6952 16204 6992
rect 16244 6952 16245 6992
rect 16203 6943 16245 6952
rect 16107 6908 16149 6917
rect 16107 6868 16108 6908
rect 16148 6868 16149 6908
rect 16107 6859 16149 6868
rect 16300 6740 16340 8791
rect 16588 8000 16628 9211
rect 17452 8672 17492 9463
rect 17644 9378 17684 9463
rect 17836 9260 17876 9269
rect 17836 8672 17876 9220
rect 17932 8849 17972 10672
rect 19084 10648 19172 10672
rect 18124 9512 18164 9521
rect 18124 9353 18164 9472
rect 19371 9512 19413 9521
rect 19371 9472 19372 9512
rect 19412 9472 19413 9512
rect 19371 9463 19413 9472
rect 19755 9512 19797 9521
rect 19755 9472 19756 9512
rect 19796 9472 19797 9512
rect 19755 9463 19797 9472
rect 19372 9378 19412 9463
rect 19756 9378 19796 9463
rect 18123 9344 18165 9353
rect 18123 9304 18124 9344
rect 18164 9304 18165 9344
rect 18123 9295 18165 9304
rect 18124 8849 18164 9295
rect 19564 9260 19604 9269
rect 19371 9176 19413 9185
rect 19371 9136 19372 9176
rect 19412 9136 19413 9176
rect 19371 9127 19413 9136
rect 18808 9092 19176 9101
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 18808 9043 19176 9052
rect 17931 8840 17973 8849
rect 17931 8800 17932 8840
rect 17972 8800 17973 8840
rect 17931 8791 17973 8800
rect 18123 8840 18165 8849
rect 18123 8800 18124 8840
rect 18164 8800 18165 8840
rect 18123 8791 18165 8800
rect 18028 8681 18068 8766
rect 17932 8672 17972 8681
rect 17836 8632 17932 8672
rect 16588 7951 16628 7960
rect 16684 8000 16724 8009
rect 16684 7253 16724 7960
rect 17355 8000 17397 8009
rect 17355 7960 17356 8000
rect 17396 7960 17397 8000
rect 17355 7951 17397 7960
rect 17068 7916 17108 7925
rect 16780 7876 17068 7916
rect 16683 7244 16725 7253
rect 16683 7204 16684 7244
rect 16724 7204 16725 7244
rect 16683 7195 16725 7204
rect 15916 6700 16340 6740
rect 15916 6656 15956 6700
rect 16395 6656 16437 6665
rect 15916 6607 15956 6616
rect 16300 6616 16396 6656
rect 16436 6616 16437 6656
rect 16107 6488 16149 6497
rect 16107 6448 16108 6488
rect 16148 6448 16149 6488
rect 16107 6439 16149 6448
rect 16108 6354 16148 6439
rect 16203 5648 16245 5657
rect 16203 5608 16204 5648
rect 16244 5608 16245 5648
rect 16203 5599 16245 5608
rect 16204 5514 16244 5599
rect 16300 5228 16340 6616
rect 16395 6607 16437 6616
rect 16204 5188 16340 5228
rect 15772 4180 15860 4220
rect 16108 4976 16148 4985
rect 15772 4178 15812 4180
rect 14668 4136 14708 4145
rect 14188 3928 14516 3968
rect 14572 4096 14668 4136
rect 14283 3800 14325 3809
rect 14283 3760 14284 3800
rect 14324 3760 14325 3800
rect 14283 3751 14325 3760
rect 14187 3632 14229 3641
rect 14187 3592 14188 3632
rect 14228 3592 14229 3632
rect 14187 3583 14229 3592
rect 14188 3473 14228 3583
rect 14187 3464 14229 3473
rect 14187 3424 14188 3464
rect 14228 3424 14229 3464
rect 14187 3415 14229 3424
rect 14188 3330 14228 3415
rect 14187 3128 14229 3137
rect 14187 3088 14188 3128
rect 14228 3088 14229 3128
rect 14187 3079 14229 3088
rect 14188 2624 14228 3079
rect 14188 2575 14228 2584
rect 14284 2624 14324 3751
rect 14572 3137 14612 4096
rect 14668 4087 14708 4096
rect 14764 4136 14804 4145
rect 15244 4136 15284 4145
rect 14667 3968 14709 3977
rect 14667 3928 14668 3968
rect 14708 3928 14709 3968
rect 14667 3919 14709 3928
rect 14668 3459 14708 3919
rect 14668 3410 14708 3419
rect 14667 3296 14709 3305
rect 14764 3296 14804 4096
rect 15148 4096 15244 4136
rect 15772 4129 15812 4138
rect 14859 3548 14901 3557
rect 14859 3508 14860 3548
rect 14900 3508 14901 3548
rect 14859 3499 14901 3508
rect 14860 3414 14900 3499
rect 14667 3256 14668 3296
rect 14708 3256 14804 3296
rect 14667 3247 14709 3256
rect 14571 3128 14613 3137
rect 14571 3088 14572 3128
rect 14612 3088 14613 3128
rect 14571 3079 14613 3088
rect 14572 2792 14612 2801
rect 14284 2575 14324 2584
rect 14380 2752 14572 2792
rect 14380 2624 14420 2752
rect 14572 2743 14612 2752
rect 14380 2575 14420 2584
rect 14572 2624 14612 2633
rect 14475 2540 14517 2549
rect 14475 2500 14476 2540
rect 14516 2500 14517 2540
rect 14475 2491 14517 2500
rect 14092 2456 14132 2465
rect 14092 1961 14132 2416
rect 14283 2204 14325 2213
rect 14283 2164 14284 2204
rect 14324 2164 14325 2204
rect 14283 2155 14325 2164
rect 13996 1793 14036 1912
rect 14091 1952 14133 1961
rect 14091 1912 14092 1952
rect 14132 1912 14133 1952
rect 14091 1903 14133 1912
rect 13995 1784 14037 1793
rect 13804 1744 13940 1784
rect 13803 1616 13845 1625
rect 13803 1576 13804 1616
rect 13844 1576 13845 1616
rect 13803 1567 13845 1576
rect 13707 1112 13749 1121
rect 13132 904 13364 944
rect 13420 1070 13460 1079
rect 13707 1072 13708 1112
rect 13748 1072 13749 1112
rect 13707 1063 13749 1072
rect 13132 80 13172 904
rect 13323 776 13365 785
rect 13323 736 13324 776
rect 13364 736 13365 776
rect 13323 727 13365 736
rect 13324 80 13364 727
rect 13420 281 13460 1030
rect 13515 860 13557 869
rect 13515 820 13516 860
rect 13556 820 13557 860
rect 13515 811 13557 820
rect 13419 272 13461 281
rect 13419 232 13420 272
rect 13460 232 13461 272
rect 13419 223 13461 232
rect 13516 80 13556 811
rect 13804 785 13844 1567
rect 13900 869 13940 1744
rect 13995 1744 13996 1784
rect 14036 1744 14037 1784
rect 13995 1735 14037 1744
rect 13899 860 13941 869
rect 13899 820 13900 860
rect 13940 820 13941 860
rect 13899 811 13941 820
rect 13803 776 13845 785
rect 13803 736 13804 776
rect 13844 736 13845 776
rect 13803 727 13845 736
rect 13899 692 13941 701
rect 13899 652 13900 692
rect 13940 652 13941 692
rect 13899 643 13941 652
rect 13707 104 13749 113
rect 13707 80 13708 104
rect 11444 64 11464 80
rect 11384 0 11464 64
rect 11576 0 11656 80
rect 11768 0 11848 80
rect 11960 0 12040 80
rect 12152 0 12232 80
rect 12344 0 12424 80
rect 12536 0 12616 80
rect 12728 0 12808 80
rect 12920 0 13000 80
rect 13112 0 13192 80
rect 13304 0 13384 80
rect 13496 0 13576 80
rect 13688 64 13708 80
rect 13748 80 13749 104
rect 13900 80 13940 643
rect 14091 440 14133 449
rect 14091 400 14092 440
rect 14132 400 14133 440
rect 14091 391 14133 400
rect 14092 80 14132 391
rect 14284 80 14324 2155
rect 14476 1952 14516 2491
rect 14572 2465 14612 2584
rect 14571 2456 14613 2465
rect 14571 2416 14572 2456
rect 14612 2416 14613 2456
rect 14571 2407 14613 2416
rect 14476 1903 14516 1912
rect 14380 1868 14420 1877
rect 14380 1784 14420 1828
rect 14668 1784 14708 3247
rect 15052 2876 15092 2885
rect 14956 2836 15052 2876
rect 14860 2624 14900 2633
rect 14860 2540 14900 2584
rect 14380 1744 14708 1784
rect 14764 2500 14900 2540
rect 14380 944 14420 1744
rect 14764 1700 14804 2500
rect 14956 2297 14996 2836
rect 15052 2827 15092 2836
rect 15052 2633 15092 2718
rect 15051 2624 15093 2633
rect 15051 2584 15052 2624
rect 15092 2584 15093 2624
rect 15051 2575 15093 2584
rect 14955 2288 14997 2297
rect 14955 2248 14956 2288
rect 14996 2248 14997 2288
rect 14955 2239 14997 2248
rect 14956 1952 14996 1961
rect 14956 1793 14996 1912
rect 15148 1793 15188 4096
rect 15244 4087 15284 4096
rect 15915 3968 15957 3977
rect 15915 3928 15916 3968
rect 15956 3928 15957 3968
rect 15915 3919 15957 3928
rect 15916 3834 15956 3919
rect 16108 3809 16148 4936
rect 16107 3800 16149 3809
rect 16107 3760 16108 3800
rect 16148 3760 16149 3800
rect 16107 3751 16149 3760
rect 16011 3464 16053 3473
rect 16011 3424 16012 3464
rect 16052 3424 16053 3464
rect 16011 3415 16053 3424
rect 15819 3380 15861 3389
rect 15819 3340 15820 3380
rect 15860 3340 15861 3380
rect 15819 3331 15861 3340
rect 15244 2633 15284 2718
rect 15531 2708 15573 2717
rect 15531 2668 15532 2708
rect 15572 2668 15573 2708
rect 15531 2659 15573 2668
rect 15243 2624 15285 2633
rect 15243 2584 15244 2624
rect 15284 2584 15285 2624
rect 15243 2575 15285 2584
rect 15340 2624 15380 2633
rect 15243 2372 15285 2381
rect 15243 2332 15244 2372
rect 15284 2332 15285 2372
rect 15243 2323 15285 2332
rect 14955 1784 14997 1793
rect 14955 1744 14956 1784
rect 14996 1744 14997 1784
rect 14955 1735 14997 1744
rect 15147 1784 15189 1793
rect 15147 1744 15148 1784
rect 15188 1744 15189 1784
rect 15147 1735 15189 1744
rect 14668 1660 14804 1700
rect 14668 1457 14708 1660
rect 14667 1448 14709 1457
rect 14667 1408 14668 1448
rect 14708 1408 14709 1448
rect 14667 1399 14709 1408
rect 15051 1448 15093 1457
rect 15051 1408 15052 1448
rect 15092 1408 15093 1448
rect 15051 1399 15093 1408
rect 14859 1280 14901 1289
rect 14859 1240 14860 1280
rect 14900 1240 14901 1280
rect 14859 1231 14901 1240
rect 14668 1121 14708 1206
rect 14860 1146 14900 1231
rect 14667 1112 14709 1121
rect 14667 1072 14668 1112
rect 14708 1072 14709 1112
rect 14667 1063 14709 1072
rect 15052 1112 15092 1399
rect 15148 1205 15188 1236
rect 15147 1196 15189 1205
rect 15147 1156 15148 1196
rect 15188 1156 15189 1196
rect 15147 1147 15189 1156
rect 15052 1063 15092 1072
rect 15148 1112 15188 1147
rect 14380 904 14708 944
rect 14475 776 14517 785
rect 14475 736 14476 776
rect 14516 736 14517 776
rect 14475 727 14517 736
rect 14476 80 14516 727
rect 14668 80 14708 904
rect 15051 860 15093 869
rect 15051 820 15052 860
rect 15092 820 15093 860
rect 15051 811 15093 820
rect 14859 188 14901 197
rect 14859 148 14860 188
rect 14900 148 14901 188
rect 14859 139 14901 148
rect 14860 80 14900 139
rect 15052 80 15092 811
rect 15148 617 15188 1072
rect 15147 608 15189 617
rect 15147 568 15148 608
rect 15188 568 15189 608
rect 15147 559 15189 568
rect 15244 80 15284 2323
rect 15340 944 15380 2584
rect 15532 2574 15572 2659
rect 15820 2549 15860 3331
rect 16012 3330 16052 3415
rect 15916 2708 15956 2717
rect 15819 2540 15861 2549
rect 15819 2500 15820 2540
rect 15860 2500 15861 2540
rect 15819 2491 15861 2500
rect 15724 2456 15764 2465
rect 15724 2288 15764 2416
rect 15532 2248 15764 2288
rect 15532 1952 15572 2248
rect 15916 2204 15956 2668
rect 15628 2164 15956 2204
rect 16108 2456 16148 2465
rect 15628 2120 15668 2164
rect 15628 2071 15668 2080
rect 15436 1938 15476 1947
rect 15532 1912 15668 1952
rect 15436 1289 15476 1898
rect 15435 1280 15477 1289
rect 15435 1240 15436 1280
rect 15476 1240 15477 1280
rect 15435 1231 15477 1240
rect 15628 1205 15668 1912
rect 15819 1868 15861 1877
rect 15819 1828 15820 1868
rect 15860 1828 15861 1868
rect 15819 1819 15861 1828
rect 15820 1734 15860 1819
rect 16012 1700 16052 1709
rect 15532 1196 15572 1205
rect 15435 1112 15477 1121
rect 15435 1072 15436 1112
rect 15476 1072 15477 1112
rect 15435 1063 15477 1072
rect 15340 895 15380 904
rect 15436 80 15476 1063
rect 15532 1037 15572 1156
rect 15627 1196 15669 1205
rect 15627 1156 15628 1196
rect 15668 1156 15669 1196
rect 15627 1147 15669 1156
rect 15531 1028 15573 1037
rect 15531 988 15532 1028
rect 15572 988 15573 1028
rect 15531 979 15573 988
rect 15724 944 15764 953
rect 15627 776 15669 785
rect 15627 736 15628 776
rect 15668 736 15669 776
rect 15627 727 15669 736
rect 15628 80 15668 727
rect 15724 533 15764 904
rect 16012 617 16052 1660
rect 16108 1457 16148 2416
rect 16107 1448 16149 1457
rect 16107 1408 16108 1448
rect 16148 1408 16149 1448
rect 16107 1399 16149 1408
rect 16204 944 16244 5188
rect 16300 5060 16340 5069
rect 16340 5020 16628 5060
rect 16300 5011 16340 5020
rect 16588 4976 16628 5020
rect 16588 4927 16628 4936
rect 16683 4976 16725 4985
rect 16683 4936 16684 4976
rect 16724 4936 16725 4976
rect 16683 4927 16725 4936
rect 16684 4842 16724 4927
rect 16299 2876 16341 2885
rect 16299 2836 16300 2876
rect 16340 2836 16341 2876
rect 16299 2827 16341 2836
rect 16300 1121 16340 2827
rect 16780 2465 16820 7876
rect 17068 7867 17108 7876
rect 17164 7916 17204 7925
rect 17204 7876 17300 7916
rect 17164 7867 17204 7876
rect 17163 5480 17205 5489
rect 17163 5440 17164 5480
rect 17204 5440 17205 5480
rect 17163 5431 17205 5440
rect 17067 5144 17109 5153
rect 17067 5104 17068 5144
rect 17108 5104 17109 5144
rect 17067 5095 17109 5104
rect 17068 4976 17108 5095
rect 16876 4936 17068 4976
rect 16779 2456 16821 2465
rect 16779 2416 16780 2456
rect 16820 2416 16821 2456
rect 16779 2407 16821 2416
rect 16587 2204 16629 2213
rect 16587 2164 16588 2204
rect 16628 2164 16629 2204
rect 16587 2155 16629 2164
rect 16491 2036 16533 2045
rect 16491 1996 16492 2036
rect 16532 1996 16533 2036
rect 16491 1987 16533 1996
rect 16395 1952 16437 1961
rect 16395 1912 16396 1952
rect 16436 1912 16437 1952
rect 16395 1903 16437 1912
rect 16299 1112 16341 1121
rect 16299 1072 16300 1112
rect 16340 1072 16341 1112
rect 16299 1063 16341 1072
rect 16108 904 16244 944
rect 16011 608 16053 617
rect 16011 568 16012 608
rect 16052 568 16053 608
rect 16011 559 16053 568
rect 15723 524 15765 533
rect 15723 484 15724 524
rect 15764 484 15765 524
rect 15723 475 15765 484
rect 16108 440 16148 904
rect 16203 776 16245 785
rect 16203 736 16204 776
rect 16244 736 16245 776
rect 16203 727 16245 736
rect 15820 400 16148 440
rect 15820 80 15860 400
rect 16011 272 16053 281
rect 16011 232 16012 272
rect 16052 232 16053 272
rect 16011 223 16053 232
rect 16012 80 16052 223
rect 16204 80 16244 727
rect 16396 524 16436 1903
rect 16492 1373 16532 1987
rect 16491 1364 16533 1373
rect 16491 1324 16492 1364
rect 16532 1324 16533 1364
rect 16491 1315 16533 1324
rect 16396 484 16532 524
rect 16395 356 16437 365
rect 16395 316 16396 356
rect 16436 316 16437 356
rect 16395 307 16437 316
rect 16396 80 16436 307
rect 16492 197 16532 484
rect 16491 188 16533 197
rect 16491 148 16492 188
rect 16532 148 16533 188
rect 16491 139 16533 148
rect 16588 80 16628 2155
rect 16780 2129 16820 2407
rect 16779 2120 16821 2129
rect 16779 2080 16780 2120
rect 16820 2080 16821 2120
rect 16779 2071 16821 2080
rect 16779 860 16821 869
rect 16779 820 16780 860
rect 16820 820 16821 860
rect 16779 811 16821 820
rect 16780 80 16820 811
rect 16876 701 16916 4936
rect 17068 4927 17108 4936
rect 17164 4976 17204 5431
rect 17164 4808 17204 4936
rect 16972 4768 17204 4808
rect 16875 692 16917 701
rect 16875 652 16876 692
rect 16916 652 16917 692
rect 16875 643 16917 652
rect 16972 80 17012 4768
rect 17260 4724 17300 7876
rect 17356 7160 17396 7951
rect 17356 7111 17396 7120
rect 17452 7085 17492 8632
rect 17932 8623 17972 8632
rect 18027 8672 18069 8681
rect 18027 8632 18028 8672
rect 18068 8632 18069 8672
rect 18027 8623 18069 8632
rect 18412 8672 18452 8681
rect 18412 8513 18452 8632
rect 18508 8672 18548 8683
rect 18508 8597 18548 8632
rect 18988 8672 19028 8681
rect 18507 8588 18549 8597
rect 18507 8548 18508 8588
rect 18548 8548 18644 8588
rect 18507 8539 18549 8548
rect 17644 8504 17684 8513
rect 18411 8504 18453 8513
rect 17684 8464 18164 8504
rect 17644 8455 17684 8464
rect 17643 8252 17685 8261
rect 17643 8212 17644 8252
rect 17684 8212 17685 8252
rect 17643 8203 17685 8212
rect 17644 8000 17684 8203
rect 17451 7076 17493 7085
rect 17451 7036 17452 7076
rect 17492 7036 17493 7076
rect 17451 7027 17493 7036
rect 17356 6488 17396 6497
rect 17452 6488 17492 7027
rect 17548 6992 17588 7001
rect 17548 6497 17588 6952
rect 17396 6448 17492 6488
rect 17356 6439 17396 6448
rect 17355 5648 17397 5657
rect 17355 5608 17356 5648
rect 17396 5608 17397 5648
rect 17355 5599 17397 5608
rect 17452 5648 17492 6448
rect 17547 6488 17589 6497
rect 17547 6448 17548 6488
rect 17588 6448 17589 6488
rect 17547 6439 17589 6448
rect 17547 6320 17589 6329
rect 17547 6280 17548 6320
rect 17588 6280 17589 6320
rect 17547 6271 17589 6280
rect 17548 6186 17588 6271
rect 17644 6236 17684 7960
rect 18124 7995 18164 8464
rect 18411 8464 18412 8504
rect 18452 8464 18453 8504
rect 18411 8455 18453 8464
rect 18219 8420 18261 8429
rect 18219 8380 18220 8420
rect 18260 8380 18261 8420
rect 18219 8371 18261 8380
rect 18124 7946 18164 7955
rect 17739 7160 17781 7169
rect 17739 7120 17740 7160
rect 17780 7120 17781 7160
rect 17739 7111 17781 7120
rect 17740 7026 17780 7111
rect 18027 6992 18069 7001
rect 18027 6952 18028 6992
rect 18068 6952 18069 6992
rect 18027 6943 18069 6952
rect 17931 6320 17973 6329
rect 17931 6280 17932 6320
rect 17972 6280 17973 6320
rect 17931 6271 17973 6280
rect 17644 6196 17780 6236
rect 17452 5599 17492 5608
rect 17068 4684 17300 4724
rect 17068 2213 17108 4684
rect 17259 3716 17301 3725
rect 17259 3676 17260 3716
rect 17300 3676 17301 3716
rect 17259 3667 17301 3676
rect 17260 3464 17300 3667
rect 17260 3415 17300 3424
rect 17163 2540 17205 2549
rect 17163 2500 17164 2540
rect 17204 2500 17205 2540
rect 17356 2540 17396 5599
rect 17644 5480 17684 5489
rect 17644 5144 17684 5440
rect 17548 5104 17684 5144
rect 17548 4985 17588 5104
rect 17547 4976 17589 4985
rect 17547 4936 17548 4976
rect 17588 4936 17589 4976
rect 17547 4927 17589 4936
rect 17644 4976 17684 4985
rect 17644 4733 17684 4936
rect 17643 4724 17685 4733
rect 17643 4684 17644 4724
rect 17684 4684 17685 4724
rect 17643 4675 17685 4684
rect 17548 4136 17588 4145
rect 17452 3632 17492 3641
rect 17548 3632 17588 4096
rect 17643 4136 17685 4145
rect 17643 4096 17644 4136
rect 17684 4096 17685 4136
rect 17643 4087 17685 4096
rect 17644 4002 17684 4087
rect 17492 3592 17588 3632
rect 17452 3583 17492 3592
rect 17643 3464 17685 3473
rect 17643 3424 17644 3464
rect 17684 3424 17685 3464
rect 17643 3415 17685 3424
rect 17644 3330 17684 3415
rect 17643 2792 17685 2801
rect 17643 2752 17644 2792
rect 17684 2752 17685 2792
rect 17643 2743 17685 2752
rect 17356 2500 17588 2540
rect 17163 2491 17205 2500
rect 17067 2204 17109 2213
rect 17067 2164 17068 2204
rect 17108 2164 17109 2204
rect 17067 2155 17109 2164
rect 17164 80 17204 2491
rect 17355 2288 17397 2297
rect 17355 2248 17356 2288
rect 17396 2248 17397 2288
rect 17355 2239 17397 2248
rect 17356 80 17396 2239
rect 17548 80 17588 2500
rect 17644 2120 17684 2743
rect 17740 2633 17780 6196
rect 17932 5648 17972 6271
rect 18028 5667 18068 6943
rect 18220 6824 18260 8371
rect 18315 8168 18357 8177
rect 18315 8128 18316 8168
rect 18356 8128 18357 8168
rect 18315 8119 18357 8128
rect 18316 8034 18356 8119
rect 18220 6784 18356 6824
rect 18219 6656 18261 6665
rect 18219 6616 18220 6656
rect 18260 6616 18261 6656
rect 18219 6607 18261 6616
rect 18123 6488 18165 6497
rect 18123 6448 18124 6488
rect 18164 6448 18165 6488
rect 18123 6439 18165 6448
rect 18220 6488 18260 6607
rect 18220 6439 18260 6448
rect 18124 6354 18164 6439
rect 18316 6329 18356 6784
rect 18315 6320 18357 6329
rect 18315 6280 18316 6320
rect 18356 6280 18357 6320
rect 18315 6271 18357 6280
rect 18316 6068 18356 6271
rect 18028 5618 18068 5627
rect 18124 6028 18356 6068
rect 17932 5599 17972 5608
rect 18124 5312 18164 6028
rect 18412 5984 18452 8455
rect 18508 8000 18548 8011
rect 18508 7925 18548 7960
rect 18507 7916 18549 7925
rect 18507 7876 18508 7916
rect 18548 7876 18549 7916
rect 18507 7867 18549 7876
rect 18604 6572 18644 8548
rect 18988 7748 19028 8632
rect 17836 5272 18164 5312
rect 18220 5944 18452 5984
rect 18508 6532 18644 6572
rect 18700 7708 19028 7748
rect 17836 3641 17876 5272
rect 18123 4976 18165 4985
rect 18123 4931 18124 4976
rect 18164 4931 18165 4976
rect 18123 4927 18165 4931
rect 18027 4892 18069 4901
rect 18027 4852 18028 4892
rect 18068 4852 18069 4892
rect 18027 4843 18069 4852
rect 18028 4220 18068 4843
rect 18124 4841 18164 4927
rect 17931 4052 17973 4061
rect 17931 4012 17932 4052
rect 17972 4012 17973 4052
rect 17931 4003 17973 4012
rect 17835 3632 17877 3641
rect 17835 3592 17836 3632
rect 17876 3592 17877 3632
rect 17835 3583 17877 3592
rect 17739 2624 17781 2633
rect 17739 2584 17740 2624
rect 17780 2584 17781 2624
rect 17739 2575 17781 2584
rect 17932 2120 17972 4003
rect 18028 2381 18068 4180
rect 18124 4220 18164 4229
rect 18220 4220 18260 5944
rect 18508 5816 18548 6532
rect 18604 6404 18644 6415
rect 18604 6329 18644 6364
rect 18700 6404 18740 7708
rect 18808 7580 19176 7589
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 18808 7531 19176 7540
rect 19372 7505 19412 9127
rect 19564 8756 19604 9220
rect 19516 8716 19604 8756
rect 19755 8756 19797 8765
rect 19755 8716 19756 8756
rect 19796 8716 19797 8756
rect 19516 8714 19556 8716
rect 19755 8707 19797 8716
rect 19516 8665 19556 8674
rect 19660 8504 19700 8513
rect 19660 7925 19700 8464
rect 19756 8009 19796 8707
rect 19948 8168 19988 10692
rect 20216 10672 20296 10752
rect 21368 10672 21448 10752
rect 22520 10672 22600 10752
rect 23672 10672 23752 10752
rect 24824 10672 24904 10752
rect 25976 10672 26056 10752
rect 27128 10672 27208 10752
rect 28280 10672 28360 10752
rect 29432 10672 29512 10752
rect 30584 10672 30664 10752
rect 31736 10672 31816 10752
rect 32235 10688 32277 10697
rect 20236 10016 20276 10672
rect 20236 9976 20564 10016
rect 20048 9848 20416 9857
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20048 9799 20416 9808
rect 20524 8924 20564 9976
rect 21388 9680 21428 10672
rect 21100 9640 21428 9680
rect 21483 9680 21525 9689
rect 21483 9640 21484 9680
rect 21524 9640 21525 9680
rect 21004 9605 21044 9636
rect 21003 9596 21045 9605
rect 21003 9556 21004 9596
rect 21044 9556 21045 9596
rect 21003 9547 21045 9556
rect 20236 8884 20564 8924
rect 21004 9512 21044 9547
rect 20236 8840 20276 8884
rect 20236 8791 20276 8800
rect 20043 8756 20085 8765
rect 20043 8716 20044 8756
rect 20084 8716 20085 8756
rect 20043 8707 20085 8716
rect 20524 8756 20564 8765
rect 20044 8622 20084 8707
rect 20048 8336 20416 8345
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20048 8287 20416 8296
rect 20524 8177 20564 8716
rect 20908 8756 20948 8765
rect 21004 8756 21044 9472
rect 21100 8840 21140 9640
rect 21483 9631 21525 9640
rect 21388 9512 21428 9521
rect 21484 9512 21524 9631
rect 21428 9472 21524 9512
rect 21388 9463 21428 9472
rect 21100 8791 21140 8800
rect 21196 9260 21236 9269
rect 20948 8716 21044 8756
rect 20908 8707 20948 8716
rect 20716 8504 20756 8513
rect 20756 8464 20948 8504
rect 20716 8455 20756 8464
rect 20523 8168 20565 8177
rect 19948 8128 20084 8168
rect 19755 8000 19797 8009
rect 19755 7960 19756 8000
rect 19796 7960 19797 8000
rect 19755 7951 19797 7960
rect 19659 7916 19701 7925
rect 19659 7876 19660 7916
rect 19700 7876 19701 7916
rect 19659 7867 19701 7876
rect 19756 7866 19796 7951
rect 19948 7748 19988 7757
rect 19756 7708 19948 7748
rect 19371 7496 19413 7505
rect 19371 7456 19372 7496
rect 19412 7456 19413 7496
rect 19371 7447 19413 7456
rect 18795 7328 18837 7337
rect 18795 7288 18796 7328
rect 18836 7288 18837 7328
rect 18795 7279 18837 7288
rect 18796 6497 18836 7279
rect 18987 7160 19029 7169
rect 18987 7120 18988 7160
rect 19028 7120 19029 7160
rect 18987 7111 19029 7120
rect 19372 7160 19412 7447
rect 19372 7111 19412 7120
rect 18988 7026 19028 7111
rect 19180 6992 19220 7001
rect 19220 6952 19508 6992
rect 19180 6943 19220 6952
rect 19179 6824 19221 6833
rect 19179 6784 19180 6824
rect 19220 6784 19221 6824
rect 19179 6775 19221 6784
rect 18795 6488 18837 6497
rect 18795 6448 18796 6488
rect 18836 6448 18837 6488
rect 18795 6439 18837 6448
rect 19180 6488 19220 6775
rect 19180 6439 19220 6448
rect 18603 6320 18645 6329
rect 18603 6280 18604 6320
rect 18644 6280 18645 6320
rect 18603 6271 18645 6280
rect 18316 5776 18548 5816
rect 18603 5816 18645 5825
rect 18603 5776 18604 5816
rect 18644 5776 18645 5816
rect 18316 5228 18356 5776
rect 18603 5767 18645 5776
rect 18411 5648 18453 5657
rect 18411 5608 18412 5648
rect 18452 5608 18453 5648
rect 18411 5599 18453 5608
rect 18508 5648 18548 5659
rect 18412 5514 18452 5599
rect 18508 5573 18548 5608
rect 18507 5564 18549 5573
rect 18507 5524 18508 5564
rect 18548 5524 18549 5564
rect 18507 5515 18549 5524
rect 18316 5188 18452 5228
rect 18316 5060 18356 5069
rect 18316 4901 18356 5020
rect 18412 4985 18452 5188
rect 18411 4976 18453 4985
rect 18411 4936 18412 4976
rect 18452 4936 18453 4976
rect 18411 4927 18453 4936
rect 18315 4892 18357 4901
rect 18315 4852 18316 4892
rect 18356 4852 18357 4892
rect 18315 4843 18357 4852
rect 18411 4724 18453 4733
rect 18411 4684 18412 4724
rect 18452 4684 18453 4724
rect 18411 4675 18453 4684
rect 18164 4180 18260 4220
rect 18027 2372 18069 2381
rect 18027 2332 18028 2372
rect 18068 2332 18069 2372
rect 18027 2323 18069 2332
rect 18124 2297 18164 4180
rect 18315 3044 18357 3053
rect 18315 3004 18316 3044
rect 18356 3004 18357 3044
rect 18315 2995 18357 3004
rect 18316 2633 18356 2995
rect 18412 2792 18452 4675
rect 18604 4304 18644 5767
rect 18508 4264 18644 4304
rect 18508 2876 18548 4264
rect 18604 4136 18644 4145
rect 18700 4136 18740 6364
rect 18808 6068 19176 6077
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 18808 6019 19176 6028
rect 19468 5662 19508 6952
rect 19756 6488 19796 7708
rect 19948 7699 19988 7708
rect 20044 6992 20084 8128
rect 20523 8128 20524 8168
rect 20564 8128 20565 8168
rect 20523 8119 20565 8128
rect 20811 8084 20853 8093
rect 20811 8044 20812 8084
rect 20852 8044 20853 8084
rect 20811 8035 20853 8044
rect 20812 8000 20852 8035
rect 20812 7949 20852 7960
rect 20427 7916 20469 7925
rect 20427 7876 20428 7916
rect 20468 7876 20469 7916
rect 20427 7867 20469 7876
rect 20428 7782 20468 7867
rect 20620 7748 20660 7757
rect 19948 6952 20084 6992
rect 20524 7708 20620 7748
rect 19948 6656 19988 6952
rect 20048 6824 20416 6833
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20048 6775 20416 6784
rect 20044 6656 20084 6665
rect 19948 6616 20044 6656
rect 20044 6607 20084 6616
rect 20235 6656 20277 6665
rect 20235 6616 20236 6656
rect 20276 6616 20277 6656
rect 20235 6607 20277 6616
rect 19851 6572 19893 6581
rect 19851 6532 19852 6572
rect 19892 6532 19893 6572
rect 19851 6523 19893 6532
rect 19708 6478 19796 6488
rect 19748 6448 19796 6478
rect 19852 6438 19892 6523
rect 19708 6429 19748 6438
rect 20236 6404 20276 6607
rect 20236 6355 20276 6364
rect 18988 5648 19028 5657
rect 19028 5608 19316 5648
rect 19468 5613 19508 5622
rect 18988 5599 19028 5608
rect 18808 4556 19176 4565
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 18808 4507 19176 4516
rect 19084 4141 19124 4150
rect 18644 4096 19028 4136
rect 18604 4087 18644 4096
rect 18891 3716 18933 3725
rect 18891 3676 18892 3716
rect 18932 3676 18933 3716
rect 18891 3667 18933 3676
rect 18892 3464 18932 3667
rect 18988 3464 19028 4096
rect 19276 4136 19316 5608
rect 19660 5480 19700 5489
rect 19660 4985 19700 5440
rect 20048 5312 20416 5321
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20048 5263 20416 5272
rect 19659 4976 19701 4985
rect 19659 4936 19660 4976
rect 19700 4936 19701 4976
rect 19659 4927 19701 4936
rect 20524 4901 20564 7708
rect 20620 7699 20660 7708
rect 20620 7169 20660 7254
rect 20619 7160 20661 7169
rect 20619 7120 20620 7160
rect 20660 7120 20661 7160
rect 20619 7111 20661 7120
rect 20812 6992 20852 7001
rect 20620 6952 20812 6992
rect 20620 5648 20660 6952
rect 20812 6943 20852 6952
rect 20620 5599 20660 5608
rect 20716 5648 20756 5657
rect 20716 5405 20756 5608
rect 20715 5396 20757 5405
rect 20715 5356 20716 5396
rect 20756 5356 20757 5396
rect 20715 5347 20757 5356
rect 20619 5312 20661 5321
rect 20619 5272 20620 5312
rect 20660 5272 20661 5312
rect 20619 5263 20661 5272
rect 20620 5153 20660 5263
rect 20619 5144 20661 5153
rect 20619 5104 20620 5144
rect 20660 5104 20661 5144
rect 20619 5095 20661 5104
rect 20908 5069 20948 8464
rect 21004 7589 21044 8716
rect 21003 7580 21045 7589
rect 21003 7540 21004 7580
rect 21044 7540 21045 7580
rect 21003 7531 21045 7540
rect 21004 7169 21044 7531
rect 21003 7160 21045 7169
rect 21003 7120 21004 7160
rect 21044 7120 21045 7160
rect 21003 7111 21045 7120
rect 21003 6656 21045 6665
rect 21003 6616 21004 6656
rect 21044 6616 21045 6656
rect 21003 6607 21045 6616
rect 21004 6413 21044 6607
rect 21196 6488 21236 9220
rect 21484 9017 21524 9472
rect 22540 9260 22580 10672
rect 23692 10445 23732 10672
rect 23691 10436 23733 10445
rect 23691 10396 23692 10436
rect 23732 10396 23733 10436
rect 23691 10387 23733 10396
rect 22635 9596 22677 9605
rect 22635 9556 22636 9596
rect 22676 9556 22677 9596
rect 22635 9547 22677 9556
rect 22636 9512 22676 9547
rect 22636 9461 22676 9472
rect 23212 9512 23252 9523
rect 23212 9437 23252 9472
rect 24459 9512 24501 9521
rect 24459 9472 24460 9512
rect 24500 9472 24501 9512
rect 24459 9463 24501 9472
rect 23211 9428 23253 9437
rect 23211 9388 23212 9428
rect 23252 9388 23253 9428
rect 23211 9379 23253 9388
rect 22444 9220 22580 9260
rect 22828 9260 22868 9269
rect 21483 9008 21525 9017
rect 21483 8968 21484 9008
rect 21524 8968 21525 9008
rect 21483 8959 21525 8968
rect 21291 8840 21333 8849
rect 21291 8800 21292 8840
rect 21332 8800 21333 8840
rect 21291 8791 21333 8800
rect 21292 8681 21332 8791
rect 21291 8672 21333 8681
rect 21291 8632 21292 8672
rect 21332 8632 21333 8672
rect 21291 8623 21333 8632
rect 21292 8538 21332 8623
rect 22444 8168 22484 9220
rect 22731 8840 22773 8849
rect 22731 8800 22732 8840
rect 22772 8800 22773 8840
rect 22731 8791 22773 8800
rect 22539 8756 22581 8765
rect 22539 8716 22540 8756
rect 22580 8716 22581 8756
rect 22539 8707 22581 8716
rect 22444 8119 22484 8128
rect 22540 8672 22580 8707
rect 22732 8706 22772 8791
rect 22060 8000 22100 8009
rect 22060 7589 22100 7960
rect 22252 7748 22292 7757
rect 22156 7708 22252 7748
rect 22059 7580 22101 7589
rect 22059 7540 22060 7580
rect 22100 7540 22101 7580
rect 22059 7531 22101 7540
rect 21388 7160 21428 7169
rect 21483 7160 21525 7169
rect 21428 7120 21484 7160
rect 21524 7120 21525 7160
rect 21388 7111 21428 7120
rect 21483 7111 21525 7120
rect 21387 6908 21429 6917
rect 21387 6868 21388 6908
rect 21428 6868 21429 6908
rect 21387 6859 21429 6868
rect 21196 6439 21236 6448
rect 21292 6488 21332 6499
rect 21292 6413 21332 6448
rect 21003 6404 21045 6413
rect 21003 6364 21004 6404
rect 21044 6364 21045 6404
rect 21003 6355 21045 6364
rect 21291 6404 21333 6413
rect 21291 6364 21292 6404
rect 21332 6364 21333 6404
rect 21291 6355 21333 6364
rect 21099 6320 21141 6329
rect 21099 6280 21100 6320
rect 21140 6280 21141 6320
rect 21099 6271 21141 6280
rect 21100 5732 21140 6271
rect 21100 5489 21140 5692
rect 21196 5648 21236 5657
rect 21388 5648 21428 6859
rect 21676 6404 21716 6413
rect 21676 5816 21716 6364
rect 21772 6404 21812 6413
rect 21772 5993 21812 6364
rect 21771 5984 21813 5993
rect 21771 5944 21772 5984
rect 21812 5944 21813 5984
rect 21771 5935 21813 5944
rect 21676 5776 21812 5816
rect 21236 5608 21428 5648
rect 21676 5648 21716 5657
rect 21099 5480 21141 5489
rect 21099 5440 21100 5480
rect 21140 5440 21141 5480
rect 21099 5431 21141 5440
rect 21196 5321 21236 5608
rect 21195 5312 21237 5321
rect 21195 5272 21196 5312
rect 21236 5272 21237 5312
rect 21195 5263 21237 5272
rect 21676 5069 21716 5608
rect 21772 5321 21812 5776
rect 22156 5662 22196 7708
rect 22252 7699 22292 7708
rect 22540 7589 22580 8632
rect 22636 7916 22676 7925
rect 22539 7580 22581 7589
rect 22539 7540 22540 7580
rect 22580 7540 22581 7580
rect 22539 7531 22581 7540
rect 22443 7496 22485 7505
rect 22443 7456 22444 7496
rect 22484 7456 22485 7496
rect 22443 7447 22485 7456
rect 22444 6665 22484 7447
rect 22540 7160 22580 7531
rect 22636 7505 22676 7876
rect 22828 7832 22868 9220
rect 23019 8840 23061 8849
rect 23019 8800 23020 8840
rect 23060 8800 23061 8840
rect 23019 8791 23061 8800
rect 23020 8672 23060 8791
rect 23020 8623 23060 8632
rect 23116 8672 23156 8681
rect 23500 8672 23540 8681
rect 23156 8632 23348 8672
rect 23116 8623 23156 8632
rect 22732 7792 22868 7832
rect 22635 7496 22677 7505
rect 22635 7456 22636 7496
rect 22676 7456 22677 7496
rect 22635 7447 22677 7456
rect 22636 7160 22676 7169
rect 22540 7120 22636 7160
rect 22636 7111 22676 7120
rect 22443 6656 22485 6665
rect 22443 6616 22444 6656
rect 22484 6616 22485 6656
rect 22443 6607 22485 6616
rect 22252 6488 22292 6497
rect 22252 5909 22292 6448
rect 22251 5900 22293 5909
rect 22251 5860 22252 5900
rect 22292 5860 22293 5900
rect 22251 5851 22293 5860
rect 22156 5613 22196 5622
rect 22252 5489 22292 5851
rect 22347 5732 22389 5741
rect 22347 5692 22348 5732
rect 22388 5692 22389 5732
rect 22347 5683 22389 5692
rect 22348 5564 22388 5683
rect 22348 5515 22388 5524
rect 22251 5480 22293 5489
rect 22251 5440 22252 5480
rect 22292 5440 22293 5480
rect 22251 5431 22293 5440
rect 21771 5312 21813 5321
rect 21771 5272 21772 5312
rect 21812 5272 21813 5312
rect 21771 5263 21813 5272
rect 20907 5060 20949 5069
rect 20907 5020 20908 5060
rect 20948 5020 20949 5060
rect 20907 5011 20949 5020
rect 21387 5060 21429 5069
rect 21387 5020 21388 5060
rect 21428 5020 21429 5060
rect 21387 5011 21429 5020
rect 21675 5060 21717 5069
rect 21675 5020 21676 5060
rect 21716 5020 21717 5060
rect 21675 5011 21717 5020
rect 20235 4892 20277 4901
rect 20235 4852 20236 4892
rect 20276 4852 20277 4892
rect 20235 4843 20277 4852
rect 20523 4892 20565 4901
rect 20523 4852 20524 4892
rect 20564 4852 20565 4892
rect 20523 4843 20565 4852
rect 21003 4892 21045 4901
rect 21003 4852 21004 4892
rect 21044 4852 21045 4892
rect 21003 4843 21045 4852
rect 21291 4892 21333 4901
rect 21291 4852 21292 4892
rect 21332 4852 21333 4892
rect 21291 4843 21333 4852
rect 20236 4758 20276 4843
rect 21004 4758 21044 4843
rect 21099 4808 21141 4817
rect 21099 4768 21100 4808
rect 21140 4768 21141 4808
rect 21099 4759 21141 4768
rect 20428 4724 20468 4733
rect 20468 4684 20948 4724
rect 20428 4675 20468 4684
rect 20619 4304 20661 4313
rect 20619 4264 20620 4304
rect 20660 4264 20661 4304
rect 20619 4255 20661 4264
rect 19084 3632 19124 4101
rect 19180 4096 19316 4136
rect 20043 4136 20085 4145
rect 20043 4096 20044 4136
rect 20084 4096 20085 4136
rect 19180 3800 19220 4096
rect 20043 4087 20085 4096
rect 20044 4002 20084 4087
rect 20620 4061 20660 4255
rect 20619 4052 20661 4061
rect 20619 4012 20620 4052
rect 20660 4012 20661 4052
rect 20619 4003 20661 4012
rect 19276 3968 19316 3977
rect 20811 3968 20853 3977
rect 19316 3928 19988 3968
rect 19276 3919 19316 3928
rect 19180 3760 19604 3800
rect 19084 3583 19124 3592
rect 18988 3424 19316 3464
rect 18892 3415 18932 3424
rect 18808 3044 19176 3053
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 18808 2995 19176 3004
rect 18508 2836 18836 2876
rect 18412 2752 18548 2792
rect 18315 2624 18357 2633
rect 18315 2584 18316 2624
rect 18356 2584 18357 2624
rect 18315 2575 18357 2584
rect 18411 2540 18453 2549
rect 18411 2500 18412 2540
rect 18452 2500 18453 2540
rect 18411 2491 18453 2500
rect 18123 2288 18165 2297
rect 18123 2248 18124 2288
rect 18164 2248 18165 2288
rect 18123 2239 18165 2248
rect 17644 2080 17780 2120
rect 17932 2080 18356 2120
rect 17643 1952 17685 1961
rect 17643 1912 17644 1952
rect 17684 1912 17685 1952
rect 17643 1903 17685 1912
rect 17644 1818 17684 1903
rect 17740 80 17780 2080
rect 17836 2036 17876 2045
rect 17876 1996 18164 2036
rect 17836 1987 17876 1996
rect 18124 1952 18164 1996
rect 18124 1903 18164 1912
rect 18220 1952 18260 1961
rect 18027 1532 18069 1541
rect 18027 1492 18028 1532
rect 18068 1492 18069 1532
rect 18027 1483 18069 1492
rect 18028 944 18068 1483
rect 18124 1121 18164 1206
rect 18123 1112 18165 1121
rect 18123 1072 18124 1112
rect 18164 1072 18165 1112
rect 18123 1063 18165 1072
rect 18028 904 18164 944
rect 17931 692 17973 701
rect 17931 652 17932 692
rect 17972 652 17973 692
rect 17931 643 17973 652
rect 17932 80 17972 643
rect 18124 80 18164 904
rect 18220 785 18260 1912
rect 18219 776 18261 785
rect 18219 736 18220 776
rect 18260 736 18261 776
rect 18219 727 18261 736
rect 18316 80 18356 2080
rect 18412 2045 18452 2491
rect 18411 2036 18453 2045
rect 18411 1996 18412 2036
rect 18452 1996 18453 2036
rect 18411 1987 18453 1996
rect 18412 1541 18452 1987
rect 18411 1532 18453 1541
rect 18411 1492 18412 1532
rect 18452 1492 18453 1532
rect 18411 1483 18453 1492
rect 18508 80 18548 2752
rect 18603 2624 18645 2633
rect 18603 2584 18604 2624
rect 18644 2584 18645 2624
rect 18603 2575 18645 2584
rect 18604 1952 18644 2575
rect 18604 1903 18644 1912
rect 18700 1868 18740 1877
rect 18603 1784 18645 1793
rect 18700 1784 18740 1828
rect 18603 1744 18604 1784
rect 18644 1744 18740 1784
rect 18603 1735 18645 1744
rect 18604 953 18644 1735
rect 18796 1700 18836 2836
rect 19179 2624 19221 2633
rect 19179 2584 19180 2624
rect 19220 2584 19221 2624
rect 19179 2575 19221 2584
rect 19180 1952 19220 2575
rect 19180 1903 19220 1912
rect 18700 1660 18836 1700
rect 18603 944 18645 953
rect 18603 904 18604 944
rect 18644 904 18645 944
rect 18603 895 18645 904
rect 18700 80 18740 1660
rect 18808 1532 19176 1541
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 18808 1483 19176 1492
rect 19276 1364 19316 3424
rect 19371 3212 19413 3221
rect 19371 3172 19372 3212
rect 19412 3172 19413 3212
rect 19371 3163 19413 3172
rect 19372 2549 19412 3163
rect 19467 3044 19509 3053
rect 19467 3004 19468 3044
rect 19508 3004 19509 3044
rect 19467 2995 19509 3004
rect 19371 2540 19413 2549
rect 19371 2500 19372 2540
rect 19412 2500 19413 2540
rect 19371 2491 19413 2500
rect 19468 1961 19508 2995
rect 19564 2129 19604 3760
rect 19948 3380 19988 3928
rect 20811 3928 20812 3968
rect 20852 3928 20853 3968
rect 20811 3919 20853 3928
rect 20048 3800 20416 3809
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20048 3751 20416 3760
rect 20523 3716 20565 3725
rect 20523 3676 20524 3716
rect 20564 3676 20565 3716
rect 20523 3667 20565 3676
rect 20524 3464 20564 3667
rect 20812 3548 20852 3919
rect 20908 3632 20948 4684
rect 21100 3977 21140 4759
rect 21196 4724 21236 4733
rect 21099 3968 21141 3977
rect 21099 3928 21100 3968
rect 21140 3928 21141 3968
rect 21099 3919 21141 3928
rect 21196 3809 21236 4684
rect 21292 4136 21332 4843
rect 21195 3800 21237 3809
rect 21195 3760 21196 3800
rect 21236 3760 21237 3800
rect 21195 3751 21237 3760
rect 21292 3641 21332 4096
rect 21388 3884 21428 5011
rect 21676 4733 21716 5011
rect 22059 4976 22101 4985
rect 22059 4936 22060 4976
rect 22100 4936 22101 4976
rect 22059 4927 22101 4936
rect 22060 4842 22100 4927
rect 22444 4733 22484 6607
rect 22732 6483 22772 7792
rect 23116 7160 23156 7169
rect 22828 7076 22868 7085
rect 23116 7076 23156 7120
rect 22868 7036 23156 7076
rect 23212 7160 23252 7169
rect 22828 7027 22868 7036
rect 23212 6917 23252 7120
rect 23211 6908 23253 6917
rect 23211 6868 23212 6908
rect 23252 6868 23253 6908
rect 23211 6859 23253 6868
rect 22924 6572 22964 6581
rect 22732 6434 22772 6443
rect 22828 6532 22924 6572
rect 22828 5732 22868 6532
rect 22924 6523 22964 6532
rect 23115 6488 23157 6497
rect 23115 6448 23116 6488
rect 23156 6448 23157 6488
rect 23115 6439 23157 6448
rect 23116 6354 23156 6439
rect 22828 5683 22868 5692
rect 23211 5732 23253 5741
rect 23211 5692 23212 5732
rect 23252 5692 23253 5732
rect 23211 5683 23253 5692
rect 23212 5598 23252 5683
rect 22636 5480 22676 5489
rect 23020 5480 23060 5489
rect 22539 5060 22581 5069
rect 22539 5020 22540 5060
rect 22580 5020 22581 5060
rect 22539 5011 22581 5020
rect 21675 4724 21717 4733
rect 21675 4684 21676 4724
rect 21716 4684 21717 4724
rect 21675 4675 21717 4684
rect 22443 4724 22485 4733
rect 22443 4684 22444 4724
rect 22484 4684 22485 4724
rect 22443 4675 22485 4684
rect 22155 4472 22197 4481
rect 22155 4432 22156 4472
rect 22196 4432 22197 4472
rect 22155 4423 22197 4432
rect 22156 4178 22196 4423
rect 22252 4178 22292 4187
rect 21772 4136 21812 4145
rect 21484 4052 21524 4061
rect 21772 4052 21812 4096
rect 21867 4136 21909 4145
rect 22156 4138 22252 4178
rect 21867 4096 21868 4136
rect 21908 4096 21909 4136
rect 22252 4129 22292 4138
rect 22348 4178 22388 4187
rect 21867 4087 21909 4096
rect 21524 4012 21812 4052
rect 21484 4003 21524 4012
rect 21868 3893 21908 4087
rect 22348 4061 22388 4138
rect 22347 4052 22389 4061
rect 22252 4012 22348 4052
rect 22388 4012 22389 4052
rect 22252 3968 22292 4012
rect 22347 4003 22389 4012
rect 22156 3928 22292 3968
rect 21867 3884 21909 3893
rect 21388 3844 21620 3884
rect 21291 3632 21333 3641
rect 20908 3592 21044 3632
rect 20812 3508 20948 3548
rect 20524 3415 20564 3424
rect 19948 3331 19988 3340
rect 20140 3212 20180 3221
rect 20180 3172 20852 3212
rect 20140 3163 20180 3172
rect 19659 3044 19701 3053
rect 19659 3004 19660 3044
rect 19700 3004 19701 3044
rect 19659 2995 19701 3004
rect 20235 3044 20277 3053
rect 20235 3004 20236 3044
rect 20276 3004 20277 3044
rect 20235 2995 20277 3004
rect 19660 2801 19700 2995
rect 19659 2792 19701 2801
rect 19659 2752 19660 2792
rect 19700 2752 19701 2792
rect 19659 2743 19701 2752
rect 20044 2624 20084 2633
rect 19947 2540 19989 2549
rect 20044 2540 20084 2584
rect 19947 2500 19948 2540
rect 19988 2500 20084 2540
rect 20139 2540 20181 2549
rect 20236 2540 20276 2995
rect 20139 2500 20140 2540
rect 20180 2500 20276 2540
rect 19947 2491 19989 2500
rect 20139 2491 20181 2500
rect 20048 2288 20416 2297
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20048 2239 20416 2248
rect 19563 2120 19605 2129
rect 19563 2080 19564 2120
rect 19604 2080 19605 2120
rect 19563 2071 19605 2080
rect 19467 1952 19509 1961
rect 19467 1912 19468 1952
rect 19508 1912 19509 1952
rect 19467 1903 19509 1912
rect 19371 1532 19413 1541
rect 19371 1492 19372 1532
rect 19412 1492 19413 1532
rect 19371 1483 19413 1492
rect 18892 1324 19316 1364
rect 18892 80 18932 1324
rect 19372 1280 19412 1483
rect 19276 1240 19412 1280
rect 19276 1196 19316 1240
rect 19084 1156 19316 1196
rect 19084 80 19124 1156
rect 19372 1112 19412 1121
rect 19468 1112 19508 1903
rect 19564 1541 19604 2071
rect 19851 2036 19893 2045
rect 19851 1996 19852 2036
rect 19892 1996 19893 2036
rect 19851 1987 19893 1996
rect 19660 1938 19700 1947
rect 19852 1902 19892 1987
rect 19563 1532 19605 1541
rect 19563 1492 19564 1532
rect 19604 1492 19605 1532
rect 19563 1483 19605 1492
rect 19564 1364 19604 1373
rect 19660 1364 19700 1898
rect 19604 1324 19700 1364
rect 19564 1315 19604 1324
rect 20523 1280 20565 1289
rect 20523 1240 20524 1280
rect 20564 1240 20565 1280
rect 20523 1231 20565 1240
rect 19659 1196 19701 1205
rect 19659 1156 19660 1196
rect 19700 1156 19701 1196
rect 19659 1147 19701 1156
rect 19412 1072 19508 1112
rect 19372 1063 19412 1072
rect 19275 944 19317 953
rect 19275 904 19276 944
rect 19316 904 19317 944
rect 19275 895 19317 904
rect 19276 80 19316 895
rect 19660 80 19700 1147
rect 20048 776 20416 785
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20048 727 20416 736
rect 20235 608 20277 617
rect 20524 608 20564 1231
rect 20619 1196 20661 1205
rect 20619 1156 20620 1196
rect 20660 1156 20661 1196
rect 20619 1147 20661 1156
rect 20235 568 20236 608
rect 20276 568 20277 608
rect 20235 559 20277 568
rect 20428 568 20564 608
rect 20043 524 20085 533
rect 20043 484 20044 524
rect 20084 484 20085 524
rect 20043 475 20085 484
rect 19851 272 19893 281
rect 19851 232 19852 272
rect 19892 232 19893 272
rect 19851 223 19893 232
rect 19852 80 19892 223
rect 20044 80 20084 475
rect 20236 80 20276 559
rect 20428 80 20468 568
rect 20620 80 20660 1147
rect 20715 1112 20757 1121
rect 20715 1072 20716 1112
rect 20756 1072 20757 1112
rect 20715 1063 20757 1072
rect 20716 978 20756 1063
rect 20812 80 20852 3172
rect 20908 1868 20948 3508
rect 20908 1819 20948 1828
rect 20907 1028 20949 1037
rect 20907 988 20908 1028
rect 20948 988 20949 1028
rect 20907 979 20949 988
rect 20908 524 20948 979
rect 21004 776 21044 3592
rect 21291 3592 21292 3632
rect 21332 3592 21333 3632
rect 21291 3583 21333 3592
rect 21291 2792 21333 2801
rect 21291 2752 21292 2792
rect 21332 2752 21333 2792
rect 21291 2743 21333 2752
rect 21292 2624 21332 2743
rect 21292 2575 21332 2584
rect 21484 2456 21524 2465
rect 21388 2416 21484 2456
rect 21388 1952 21428 2416
rect 21484 2407 21524 2416
rect 21388 1903 21428 1912
rect 21484 1952 21524 1961
rect 21099 1700 21141 1709
rect 21099 1660 21100 1700
rect 21140 1660 21141 1700
rect 21099 1651 21141 1660
rect 21100 1566 21140 1651
rect 21484 1373 21524 1912
rect 21483 1364 21525 1373
rect 21483 1324 21484 1364
rect 21524 1324 21525 1364
rect 21483 1315 21525 1324
rect 21004 736 21236 776
rect 20908 484 21044 524
rect 21004 80 21044 484
rect 21196 80 21236 736
rect 21387 608 21429 617
rect 21387 568 21388 608
rect 21428 568 21429 608
rect 21387 559 21429 568
rect 21388 80 21428 559
rect 21580 80 21620 3844
rect 21867 3844 21868 3884
rect 21908 3844 21909 3884
rect 21867 3835 21909 3844
rect 21772 3464 21812 3473
rect 21772 2801 21812 3424
rect 21964 3212 22004 3221
rect 21771 2792 21813 2801
rect 21771 2752 21772 2792
rect 21812 2752 21813 2792
rect 21771 2743 21813 2752
rect 21772 1121 21812 2743
rect 21964 2624 22004 3172
rect 22059 2876 22101 2885
rect 22059 2836 22060 2876
rect 22100 2836 22101 2876
rect 22059 2827 22101 2836
rect 21964 2575 22004 2584
rect 22060 2624 22100 2827
rect 22060 2575 22100 2584
rect 22156 2456 22196 3928
rect 22347 3884 22389 3893
rect 22347 3844 22348 3884
rect 22388 3844 22389 3884
rect 22347 3835 22389 3844
rect 22251 3800 22293 3809
rect 22251 3760 22252 3800
rect 22292 3760 22293 3800
rect 22251 3751 22293 3760
rect 22060 2416 22196 2456
rect 21867 2372 21909 2381
rect 21867 2332 21868 2372
rect 21908 2332 21909 2372
rect 21867 2323 21909 2332
rect 21868 2213 21908 2323
rect 21963 2288 22005 2297
rect 21963 2248 21964 2288
rect 22004 2248 22005 2288
rect 21963 2239 22005 2248
rect 21867 2204 21909 2213
rect 21867 2164 21868 2204
rect 21908 2164 21909 2204
rect 21867 2155 21909 2164
rect 21868 1952 21908 2155
rect 21868 1903 21908 1912
rect 21964 1952 22004 2239
rect 21964 1793 22004 1912
rect 21963 1784 22005 1793
rect 21963 1744 21964 1784
rect 22004 1744 22005 1784
rect 21963 1735 22005 1744
rect 21867 1700 21909 1709
rect 21867 1660 21868 1700
rect 21908 1660 21909 1700
rect 21867 1651 21909 1660
rect 21771 1112 21813 1121
rect 21771 1072 21772 1112
rect 21812 1072 21813 1112
rect 21771 1063 21813 1072
rect 21771 944 21813 953
rect 21771 904 21772 944
rect 21812 904 21813 944
rect 21771 895 21813 904
rect 21772 80 21812 895
rect 21868 860 21908 1651
rect 21963 1112 22005 1121
rect 21963 1072 21964 1112
rect 22004 1072 22005 1112
rect 21963 1063 22005 1072
rect 21964 978 22004 1063
rect 22060 869 22100 2416
rect 22155 1364 22197 1373
rect 22155 1324 22156 1364
rect 22196 1324 22197 1364
rect 22155 1315 22197 1324
rect 22156 1230 22196 1315
rect 22252 1112 22292 3751
rect 22348 1280 22388 3835
rect 22443 3632 22485 3641
rect 22443 3592 22444 3632
rect 22484 3592 22485 3632
rect 22443 3583 22485 3592
rect 22444 2717 22484 3583
rect 22443 2708 22485 2717
rect 22443 2668 22444 2708
rect 22484 2668 22485 2708
rect 22443 2659 22485 2668
rect 22540 2708 22580 5011
rect 22540 2659 22580 2668
rect 22444 2574 22484 2659
rect 22636 2456 22676 5440
rect 22924 5440 23020 5480
rect 22827 4304 22869 4313
rect 22827 4264 22828 4304
rect 22868 4264 22869 4304
rect 22827 4255 22869 4264
rect 22828 4136 22868 4255
rect 22828 4087 22868 4096
rect 22731 3800 22773 3809
rect 22731 3760 22732 3800
rect 22772 3760 22773 3800
rect 22731 3751 22773 3760
rect 22732 3380 22772 3751
rect 22924 3380 22964 5440
rect 23020 5431 23060 5440
rect 23308 5144 23348 8632
rect 23500 8261 23540 8632
rect 23596 8672 23636 8681
rect 23596 8429 23636 8632
rect 24076 8672 24116 8681
rect 23595 8420 23637 8429
rect 23595 8380 23596 8420
rect 23636 8380 23637 8420
rect 23595 8371 23637 8380
rect 24076 8345 24116 8632
rect 24075 8336 24117 8345
rect 24075 8296 24076 8336
rect 24116 8296 24117 8336
rect 24075 8287 24117 8296
rect 23499 8252 23541 8261
rect 23499 8212 23500 8252
rect 23540 8212 23541 8252
rect 23499 8203 23541 8212
rect 23500 8000 23540 8009
rect 24460 8000 24500 9463
rect 24844 9428 24884 10672
rect 25996 10613 26036 10672
rect 25995 10604 26037 10613
rect 25995 10564 25996 10604
rect 26036 10564 26037 10604
rect 25995 10555 26037 10564
rect 27148 10529 27188 10672
rect 27147 10520 27189 10529
rect 27147 10480 27148 10520
rect 27188 10480 27189 10520
rect 27147 10471 27189 10480
rect 28300 9857 28340 10672
rect 28299 9848 28341 9857
rect 28299 9808 28300 9848
rect 28340 9808 28341 9848
rect 28299 9799 28341 9808
rect 27915 9764 27957 9773
rect 27915 9724 27916 9764
rect 27956 9724 27957 9764
rect 27915 9715 27957 9724
rect 26283 9596 26325 9605
rect 26283 9556 26284 9596
rect 26324 9556 26325 9596
rect 26283 9547 26325 9556
rect 25035 9512 25077 9521
rect 25035 9472 25036 9512
rect 25076 9472 25077 9512
rect 25035 9463 25077 9472
rect 26284 9512 26324 9547
rect 24748 9388 24884 9428
rect 24652 9260 24692 9269
rect 24652 8756 24692 9220
rect 24748 9092 24788 9388
rect 25036 9378 25076 9463
rect 24844 9260 24884 9269
rect 24884 9220 25172 9260
rect 24844 9211 24884 9220
rect 25035 9092 25077 9101
rect 24748 9052 24884 9092
rect 24604 8716 24692 8756
rect 24604 8714 24644 8716
rect 24604 8665 24644 8674
rect 24747 8504 24789 8513
rect 24747 8464 24748 8504
rect 24788 8464 24789 8504
rect 24747 8455 24789 8464
rect 24748 8370 24788 8455
rect 24844 8009 24884 9052
rect 25035 9052 25036 9092
rect 25076 9052 25077 9092
rect 25035 9043 25077 9052
rect 24748 8000 24788 8009
rect 24460 7960 24748 8000
rect 23500 7841 23540 7960
rect 23499 7832 23541 7841
rect 23499 7792 23500 7832
rect 23540 7792 23541 7832
rect 23499 7783 23541 7792
rect 24652 7589 24692 7960
rect 24748 7951 24788 7960
rect 24843 8000 24885 8009
rect 24843 7960 24844 8000
rect 24884 7960 24885 8000
rect 25036 8000 25076 9043
rect 25132 8672 25172 9220
rect 25899 9008 25941 9017
rect 25899 8968 25900 9008
rect 25940 8968 25941 9008
rect 25899 8959 25941 8968
rect 25612 8681 25652 8766
rect 25132 8623 25172 8632
rect 25227 8672 25269 8681
rect 25227 8632 25228 8672
rect 25268 8632 25269 8672
rect 25227 8623 25269 8632
rect 25611 8672 25653 8681
rect 25611 8632 25612 8672
rect 25652 8632 25653 8672
rect 25611 8623 25653 8632
rect 25708 8672 25748 8681
rect 25228 8538 25268 8623
rect 25611 8504 25653 8513
rect 25611 8464 25612 8504
rect 25652 8464 25653 8504
rect 25611 8455 25653 8464
rect 25515 8336 25557 8345
rect 25515 8296 25516 8336
rect 25556 8296 25557 8336
rect 25515 8287 25557 8296
rect 25132 8000 25172 8009
rect 25036 7960 25132 8000
rect 24843 7951 24885 7960
rect 25132 7951 25172 7960
rect 24940 7748 24980 7757
rect 24748 7708 24940 7748
rect 24363 7580 24405 7589
rect 24363 7540 24364 7580
rect 24404 7540 24405 7580
rect 24363 7531 24405 7540
rect 24651 7580 24693 7589
rect 24651 7540 24652 7580
rect 24692 7540 24693 7580
rect 24651 7531 24693 7540
rect 23596 7160 23636 7169
rect 23596 6329 23636 7120
rect 23692 7160 23732 7169
rect 24172 7160 24212 7169
rect 23692 6749 23732 7120
rect 23980 7120 24172 7160
rect 23691 6740 23733 6749
rect 23691 6700 23692 6740
rect 23732 6700 23733 6740
rect 23691 6691 23733 6700
rect 23883 6572 23925 6581
rect 23883 6532 23884 6572
rect 23924 6532 23925 6572
rect 23883 6523 23925 6532
rect 23595 6320 23637 6329
rect 23595 6280 23596 6320
rect 23636 6280 23637 6320
rect 23595 6271 23637 6280
rect 23884 5732 23924 6523
rect 23884 5683 23924 5692
rect 23212 5104 23348 5144
rect 23212 4565 23252 5104
rect 23308 4976 23348 4985
rect 23308 4817 23348 4936
rect 23307 4808 23349 4817
rect 23307 4768 23308 4808
rect 23348 4768 23349 4808
rect 23307 4759 23349 4768
rect 23500 4724 23540 4733
rect 23404 4684 23500 4724
rect 23211 4556 23253 4565
rect 23211 4516 23212 4556
rect 23252 4516 23253 4556
rect 23211 4507 23253 4516
rect 23115 4388 23157 4397
rect 23115 4348 23116 4388
rect 23156 4348 23157 4388
rect 23115 4339 23157 4348
rect 23019 3464 23061 3473
rect 23019 3424 23020 3464
rect 23060 3424 23061 3464
rect 23019 3415 23061 3424
rect 23116 3464 23156 4339
rect 22732 3331 22772 3340
rect 22828 3340 22964 3380
rect 22828 3212 22868 3340
rect 22540 2416 22676 2456
rect 22732 3172 22868 3212
rect 22924 3212 22964 3221
rect 22443 2120 22485 2129
rect 22443 2080 22444 2120
rect 22484 2080 22485 2120
rect 22443 2071 22485 2080
rect 22444 1952 22484 2071
rect 22444 1903 22484 1912
rect 22348 1240 22484 1280
rect 22156 1072 22292 1112
rect 22348 1112 22388 1121
rect 22059 860 22101 869
rect 21868 820 22004 860
rect 21964 80 22004 820
rect 22059 820 22060 860
rect 22100 820 22101 860
rect 22059 811 22101 820
rect 22156 80 22196 1072
rect 22348 1028 22388 1072
rect 22252 988 22388 1028
rect 22252 869 22292 988
rect 22444 944 22484 1240
rect 22348 904 22484 944
rect 22251 860 22293 869
rect 22251 820 22252 860
rect 22292 820 22293 860
rect 22251 811 22293 820
rect 22348 80 22388 904
rect 22540 80 22580 2416
rect 22635 1364 22677 1373
rect 22635 1324 22636 1364
rect 22676 1324 22677 1364
rect 22635 1315 22677 1324
rect 22636 533 22676 1315
rect 22635 524 22677 533
rect 22635 484 22636 524
rect 22676 484 22677 524
rect 22635 475 22677 484
rect 22732 80 22772 3172
rect 22924 2540 22964 3172
rect 23020 3053 23060 3415
rect 23019 3044 23061 3053
rect 23019 3004 23020 3044
rect 23060 3004 23061 3044
rect 23019 2995 23061 3004
rect 23020 2624 23060 2995
rect 23116 2801 23156 3424
rect 23115 2792 23157 2801
rect 23115 2752 23116 2792
rect 23156 2752 23157 2792
rect 23115 2743 23157 2752
rect 23020 2575 23060 2584
rect 22828 2500 22964 2540
rect 22828 1616 22868 2500
rect 23116 2036 23156 2045
rect 22972 1910 23012 1919
rect 23116 1877 23156 1996
rect 22972 1868 23012 1870
rect 23115 1868 23157 1877
rect 22972 1828 23060 1868
rect 22828 1576 22964 1616
rect 22924 80 22964 1576
rect 23020 1289 23060 1828
rect 23115 1828 23116 1868
rect 23156 1828 23157 1868
rect 23115 1819 23157 1828
rect 23115 1700 23157 1709
rect 23115 1660 23116 1700
rect 23156 1660 23157 1700
rect 23115 1651 23157 1660
rect 23019 1280 23061 1289
rect 23019 1240 23020 1280
rect 23060 1240 23061 1280
rect 23019 1231 23061 1240
rect 23116 80 23156 1651
rect 23212 1205 23252 4507
rect 23404 4220 23444 4684
rect 23500 4675 23540 4684
rect 23356 4180 23444 4220
rect 23356 4178 23396 4180
rect 23356 4129 23396 4138
rect 23500 3968 23540 3977
rect 23500 3809 23540 3928
rect 23499 3800 23541 3809
rect 23499 3760 23500 3800
rect 23540 3760 23541 3800
rect 23499 3751 23541 3760
rect 23980 3473 24020 7120
rect 24172 7111 24212 7120
rect 24364 6581 24404 7531
rect 24748 7244 24788 7708
rect 24940 7699 24980 7708
rect 24700 7204 24788 7244
rect 24843 7244 24885 7253
rect 24843 7204 24844 7244
rect 24884 7204 24885 7244
rect 24700 7202 24740 7204
rect 24843 7195 24885 7204
rect 25227 7244 25269 7253
rect 25227 7204 25228 7244
rect 25268 7204 25269 7244
rect 25227 7195 25269 7204
rect 24700 7153 24740 7162
rect 24844 7076 24884 7195
rect 25228 7110 25268 7195
rect 24844 7027 24884 7036
rect 24939 7076 24981 7085
rect 24939 7036 24940 7076
rect 24980 7036 24981 7076
rect 24939 7027 24981 7036
rect 24940 6665 24980 7027
rect 25516 7001 25556 8287
rect 25612 7244 25652 8455
rect 25708 8429 25748 8632
rect 25707 8420 25749 8429
rect 25707 8380 25708 8420
rect 25748 8380 25749 8420
rect 25707 8371 25749 8380
rect 25612 7195 25652 7204
rect 25803 7244 25845 7253
rect 25803 7204 25804 7244
rect 25844 7204 25845 7244
rect 25803 7195 25845 7204
rect 25036 6992 25076 7001
rect 25420 6992 25460 7001
rect 24939 6656 24981 6665
rect 24939 6616 24940 6656
rect 24980 6616 24981 6656
rect 24939 6607 24981 6616
rect 24363 6572 24405 6581
rect 24363 6532 24364 6572
rect 24404 6532 24405 6572
rect 24363 6523 24405 6532
rect 24364 6488 24404 6523
rect 24364 6438 24404 6448
rect 24940 6488 24980 6607
rect 24940 6439 24980 6448
rect 24556 6236 24596 6245
rect 24364 6196 24556 6236
rect 24364 5648 24404 6196
rect 24556 6187 24596 6196
rect 24364 5599 24404 5608
rect 24459 5648 24501 5657
rect 24459 5608 24460 5648
rect 24500 5608 24501 5648
rect 24459 5599 24501 5608
rect 24844 5648 24884 5657
rect 24460 5514 24500 5599
rect 24076 5480 24116 5489
rect 23979 3464 24021 3473
rect 23979 3424 23980 3464
rect 24020 3424 24021 3464
rect 23979 3415 24021 3424
rect 24076 3053 24116 5440
rect 24844 5153 24884 5608
rect 24940 5648 24980 5657
rect 24940 5489 24980 5608
rect 24939 5480 24981 5489
rect 24939 5440 24940 5480
rect 24980 5440 24981 5480
rect 24939 5431 24981 5440
rect 24843 5144 24885 5153
rect 24843 5104 24844 5144
rect 24884 5104 24885 5144
rect 24843 5095 24885 5104
rect 24555 4976 24597 4985
rect 24555 4936 24556 4976
rect 24596 4936 24597 4976
rect 24555 4927 24597 4936
rect 24556 4842 24596 4927
rect 25036 4808 25076 6952
rect 25324 6952 25420 6992
rect 25131 6404 25173 6413
rect 25131 6364 25132 6404
rect 25172 6364 25173 6404
rect 25131 6355 25173 6364
rect 24652 4768 25076 4808
rect 24459 4472 24501 4481
rect 24459 4432 24460 4472
rect 24500 4432 24501 4472
rect 24459 4423 24501 4432
rect 24172 4264 24404 4304
rect 24075 3044 24117 3053
rect 24075 3004 24076 3044
rect 24116 3004 24117 3044
rect 24075 2995 24117 3004
rect 23691 2708 23733 2717
rect 23691 2668 23692 2708
rect 23732 2668 23733 2708
rect 23691 2659 23733 2668
rect 24075 2708 24117 2717
rect 24075 2668 24076 2708
rect 24116 2668 24117 2708
rect 24075 2659 24117 2668
rect 23548 2633 23588 2642
rect 23588 2593 23636 2624
rect 23548 2584 23636 2593
rect 23307 2036 23349 2045
rect 23307 1996 23308 2036
rect 23348 1996 23349 2036
rect 23307 1987 23349 1996
rect 23308 1868 23348 1987
rect 23308 1819 23348 1828
rect 23500 1700 23540 1709
rect 23307 1364 23349 1373
rect 23307 1324 23308 1364
rect 23348 1324 23349 1364
rect 23307 1315 23349 1324
rect 23211 1196 23253 1205
rect 23211 1156 23212 1196
rect 23252 1156 23253 1196
rect 23211 1147 23253 1156
rect 23308 80 23348 1315
rect 23500 80 23540 1660
rect 23596 1280 23636 2584
rect 23692 2540 23732 2659
rect 24076 2574 24116 2659
rect 23692 2491 23732 2500
rect 23884 2456 23924 2465
rect 23788 2416 23884 2456
rect 24172 2456 24212 4264
rect 24268 4136 24308 4145
rect 24268 3809 24308 4096
rect 24364 4136 24404 4264
rect 24364 4087 24404 4096
rect 24267 3800 24309 3809
rect 24267 3760 24268 3800
rect 24308 3760 24309 3800
rect 24267 3751 24309 3760
rect 24364 3464 24404 3473
rect 24460 3464 24500 4423
rect 24555 3800 24597 3809
rect 24555 3760 24556 3800
rect 24596 3760 24597 3800
rect 24555 3751 24597 3760
rect 24556 3632 24596 3751
rect 24556 3583 24596 3592
rect 24404 3424 24500 3464
rect 24364 3415 24404 3424
rect 24460 3137 24500 3424
rect 24459 3128 24501 3137
rect 24459 3088 24460 3128
rect 24500 3088 24501 3128
rect 24459 3079 24501 3088
rect 24267 2708 24309 2717
rect 24267 2668 24268 2708
rect 24308 2668 24309 2708
rect 24267 2659 24309 2668
rect 24268 2624 24308 2659
rect 24268 2573 24308 2584
rect 24172 2416 24404 2456
rect 23691 1700 23733 1709
rect 23691 1660 23692 1700
rect 23732 1660 23733 1700
rect 23691 1651 23733 1660
rect 23692 1566 23732 1651
rect 23788 1280 23828 2416
rect 23884 2407 23924 2416
rect 24268 1952 24308 1961
rect 23980 1912 24268 1952
rect 23883 1868 23925 1877
rect 23883 1828 23884 1868
rect 23924 1828 23925 1868
rect 23883 1819 23925 1828
rect 23884 1734 23924 1819
rect 23980 1364 24020 1912
rect 24268 1903 24308 1912
rect 24364 1952 24404 2416
rect 24364 1625 24404 1912
rect 24363 1616 24405 1625
rect 24363 1576 24364 1616
rect 24404 1576 24405 1616
rect 24363 1567 24405 1576
rect 23980 1315 24020 1324
rect 23596 1240 23732 1280
rect 23788 1240 23924 1280
rect 23595 1112 23637 1121
rect 23595 1072 23596 1112
rect 23636 1072 23637 1112
rect 23595 1063 23637 1072
rect 23596 978 23636 1063
rect 23692 1028 23732 1240
rect 23788 1028 23828 1037
rect 23692 988 23788 1028
rect 23788 979 23828 988
rect 23691 524 23733 533
rect 23691 484 23692 524
rect 23732 484 23733 524
rect 23691 475 23733 484
rect 23692 80 23732 475
rect 23884 80 23924 1240
rect 24171 1112 24213 1121
rect 24171 1072 24172 1112
rect 24212 1072 24213 1112
rect 24171 1063 24213 1072
rect 24172 978 24212 1063
rect 24267 944 24309 953
rect 24267 904 24268 944
rect 24308 904 24309 944
rect 24267 895 24309 904
rect 24075 860 24117 869
rect 24075 820 24076 860
rect 24116 820 24117 860
rect 24075 811 24117 820
rect 24076 80 24116 811
rect 24268 80 24308 895
rect 24459 104 24501 113
rect 24459 80 24460 104
rect 13748 64 13768 80
rect 13688 0 13768 64
rect 13880 0 13960 80
rect 14072 0 14152 80
rect 14264 0 14344 80
rect 14456 0 14536 80
rect 14648 0 14728 80
rect 14840 0 14920 80
rect 15032 0 15112 80
rect 15224 0 15304 80
rect 15416 0 15496 80
rect 15608 0 15688 80
rect 15800 0 15880 80
rect 15992 0 16072 80
rect 16184 0 16264 80
rect 16376 0 16456 80
rect 16568 0 16648 80
rect 16760 0 16840 80
rect 16952 0 17032 80
rect 17144 0 17224 80
rect 17336 0 17416 80
rect 17528 0 17608 80
rect 17720 0 17800 80
rect 17912 0 17992 80
rect 18104 0 18184 80
rect 18296 0 18376 80
rect 18488 0 18568 80
rect 18680 0 18760 80
rect 18872 0 18952 80
rect 19064 0 19144 80
rect 19256 0 19336 80
rect 19448 0 19528 80
rect 19640 0 19720 80
rect 19832 0 19912 80
rect 20024 0 20104 80
rect 20216 0 20296 80
rect 20408 0 20488 80
rect 20600 0 20680 80
rect 20792 0 20872 80
rect 20984 0 21064 80
rect 21176 0 21256 80
rect 21368 0 21448 80
rect 21560 0 21640 80
rect 21752 0 21832 80
rect 21944 0 22024 80
rect 22136 0 22216 80
rect 22328 0 22408 80
rect 22520 0 22600 80
rect 22712 0 22792 80
rect 22904 0 22984 80
rect 23096 0 23176 80
rect 23288 0 23368 80
rect 23480 0 23560 80
rect 23672 0 23752 80
rect 23864 0 23944 80
rect 24056 0 24136 80
rect 24248 0 24328 80
rect 24440 64 24460 80
rect 24500 80 24501 104
rect 24652 80 24692 4768
rect 24844 4220 24884 4229
rect 25132 4220 25172 6355
rect 25227 6320 25269 6329
rect 25227 6280 25228 6320
rect 25268 6280 25269 6320
rect 25227 6271 25269 6280
rect 24884 4180 25172 4220
rect 24844 4171 24884 4180
rect 24747 4136 24789 4145
rect 24747 4096 24748 4136
rect 24788 4096 24789 4136
rect 24747 4087 24789 4096
rect 24748 4002 24788 4087
rect 25228 3548 25268 6271
rect 25324 4388 25364 6952
rect 25420 6943 25460 6952
rect 25515 6992 25557 7001
rect 25515 6952 25516 6992
rect 25556 6952 25557 6992
rect 25515 6943 25557 6952
rect 25419 5816 25461 5825
rect 25419 5776 25420 5816
rect 25460 5776 25461 5816
rect 25419 5767 25461 5776
rect 25420 5648 25460 5767
rect 25420 5599 25460 5608
rect 25324 4348 25460 4388
rect 25324 4136 25364 4145
rect 25324 3809 25364 4096
rect 25323 3800 25365 3809
rect 25323 3760 25324 3800
rect 25364 3760 25365 3800
rect 25323 3751 25365 3760
rect 25132 3508 25268 3548
rect 25036 3212 25076 3221
rect 24940 3172 25036 3212
rect 24747 1952 24789 1961
rect 24747 1912 24748 1952
rect 24788 1912 24789 1952
rect 24747 1903 24789 1912
rect 24748 1818 24788 1903
rect 24844 1868 24884 1877
rect 24844 1625 24884 1828
rect 24843 1616 24885 1625
rect 24843 1576 24844 1616
rect 24884 1576 24885 1616
rect 24843 1567 24885 1576
rect 24844 365 24884 1567
rect 24940 1373 24980 3172
rect 25036 3163 25076 3172
rect 25035 3044 25077 3053
rect 25035 3004 25036 3044
rect 25076 3004 25077 3044
rect 25035 2995 25077 3004
rect 24939 1364 24981 1373
rect 24939 1324 24940 1364
rect 24980 1324 24981 1364
rect 24939 1315 24981 1324
rect 24939 776 24981 785
rect 24939 736 24940 776
rect 24980 736 24981 776
rect 24939 727 24981 736
rect 24843 356 24885 365
rect 24843 316 24844 356
rect 24884 316 24885 356
rect 24843 307 24885 316
rect 24940 188 24980 727
rect 24844 148 24980 188
rect 24844 80 24884 148
rect 25036 80 25076 2995
rect 25132 2213 25172 3508
rect 25228 3380 25268 3389
rect 25131 2204 25173 2213
rect 25131 2164 25132 2204
rect 25172 2164 25173 2204
rect 25131 2155 25173 2164
rect 25228 2129 25268 3340
rect 25324 3221 25364 3751
rect 25323 3212 25365 3221
rect 25323 3172 25324 3212
rect 25364 3172 25365 3212
rect 25323 3163 25365 3172
rect 25227 2120 25269 2129
rect 25227 2080 25228 2120
rect 25268 2080 25269 2120
rect 25227 2071 25269 2080
rect 25227 1952 25269 1961
rect 25227 1912 25228 1952
rect 25268 1912 25269 1952
rect 25227 1903 25269 1912
rect 25324 1952 25364 1963
rect 25228 80 25268 1903
rect 25324 1877 25364 1912
rect 25323 1868 25365 1877
rect 25323 1828 25324 1868
rect 25364 1828 25365 1868
rect 25323 1819 25365 1828
rect 25420 1448 25460 4348
rect 25516 3809 25556 6943
rect 25804 6833 25844 7195
rect 25900 7160 25940 8959
rect 26188 8672 26228 8681
rect 26188 8597 26228 8632
rect 26187 8588 26229 8597
rect 26187 8548 26188 8588
rect 26228 8548 26229 8588
rect 26187 8539 26229 8548
rect 26188 8345 26228 8539
rect 26187 8336 26229 8345
rect 26187 8296 26188 8336
rect 26228 8296 26229 8336
rect 26187 8287 26229 8296
rect 26284 8093 26324 9472
rect 26667 9512 26709 9521
rect 26667 9472 26668 9512
rect 26708 9472 26709 9512
rect 26667 9463 26709 9472
rect 27916 9512 27956 9715
rect 29452 9689 29492 10672
rect 29259 9680 29301 9689
rect 29259 9640 29260 9680
rect 29300 9640 29301 9680
rect 29259 9631 29301 9640
rect 29451 9680 29493 9689
rect 29451 9640 29452 9680
rect 29492 9640 29493 9680
rect 29451 9631 29493 9640
rect 26668 9378 26708 9463
rect 26476 9260 26516 9269
rect 26516 9220 26708 9260
rect 26476 9211 26516 9220
rect 26668 8686 26708 9220
rect 27916 9101 27956 9472
rect 28300 9512 28340 9521
rect 28340 9472 28532 9512
rect 28300 9463 28340 9472
rect 28108 9260 28148 9269
rect 28148 9220 28436 9260
rect 28108 9211 28148 9220
rect 27915 9092 27957 9101
rect 27915 9052 27916 9092
rect 27956 9052 27957 9092
rect 27915 9043 27957 9052
rect 27244 8756 27284 8765
rect 27244 8672 27284 8716
rect 27339 8756 27381 8765
rect 27339 8716 27340 8756
rect 27380 8716 27381 8756
rect 27339 8707 27381 8716
rect 26668 8637 26708 8646
rect 26956 8632 27284 8672
rect 26860 8588 26900 8597
rect 26956 8588 26996 8632
rect 26900 8548 26996 8588
rect 26860 8539 26900 8548
rect 27052 8504 27092 8513
rect 26475 8420 26517 8429
rect 26475 8380 26476 8420
rect 26516 8380 26517 8420
rect 26475 8371 26517 8380
rect 26283 8084 26325 8093
rect 26283 8044 26284 8084
rect 26324 8044 26325 8084
rect 26283 8035 26325 8044
rect 26380 8000 26420 8009
rect 26380 7253 26420 7960
rect 26379 7244 26421 7253
rect 26379 7204 26380 7244
rect 26420 7204 26421 7244
rect 26379 7195 26421 7204
rect 25803 6824 25845 6833
rect 25803 6784 25804 6824
rect 25844 6784 25845 6824
rect 25803 6775 25845 6784
rect 25611 6740 25653 6749
rect 25611 6700 25612 6740
rect 25652 6700 25653 6740
rect 25611 6691 25653 6700
rect 25515 3800 25557 3809
rect 25515 3760 25516 3800
rect 25556 3760 25557 3800
rect 25515 3751 25557 3760
rect 25612 3641 25652 6691
rect 25804 4976 25844 6775
rect 25900 6665 25940 7120
rect 25899 6656 25941 6665
rect 25899 6616 25900 6656
rect 25940 6616 25941 6656
rect 25899 6607 25941 6616
rect 26187 6572 26229 6581
rect 26187 6532 26188 6572
rect 26228 6532 26229 6572
rect 26187 6523 26229 6532
rect 26188 6488 26228 6523
rect 26188 6437 26228 6448
rect 26380 6236 26420 6245
rect 25996 6196 26380 6236
rect 25996 5732 26036 6196
rect 26380 6187 26420 6196
rect 26476 5900 26516 8371
rect 26572 8084 26612 8093
rect 26612 8044 26900 8084
rect 26572 8035 26612 8044
rect 26860 8000 26900 8044
rect 26860 7951 26900 7960
rect 26956 8000 26996 8009
rect 26859 7076 26901 7085
rect 26859 7036 26860 7076
rect 26900 7036 26901 7076
rect 26859 7027 26901 7036
rect 26860 6497 26900 7027
rect 26859 6488 26901 6497
rect 26859 6448 26860 6488
rect 26900 6448 26901 6488
rect 26859 6439 26901 6448
rect 26956 6329 26996 7960
rect 27052 7589 27092 8464
rect 27340 8084 27380 8707
rect 27628 8504 27668 8515
rect 27628 8429 27668 8464
rect 27627 8420 27669 8429
rect 27627 8380 27628 8420
rect 27668 8380 27669 8420
rect 27627 8371 27669 8380
rect 27915 8420 27957 8429
rect 27915 8380 27916 8420
rect 27956 8380 27957 8420
rect 27915 8371 27957 8380
rect 27340 8044 27668 8084
rect 27340 8000 27380 8044
rect 27340 7951 27380 7960
rect 27436 7916 27476 7925
rect 27051 7580 27093 7589
rect 27051 7540 27052 7580
rect 27092 7540 27093 7580
rect 27051 7531 27093 7540
rect 27147 7244 27189 7253
rect 27147 7204 27148 7244
rect 27188 7204 27189 7244
rect 27147 7195 27189 7204
rect 27148 7160 27188 7195
rect 27148 7109 27188 7120
rect 27340 6992 27380 7001
rect 27052 6952 27340 6992
rect 27052 6488 27092 6952
rect 27340 6943 27380 6952
rect 27436 6917 27476 7876
rect 27532 7160 27572 7171
rect 27532 7085 27572 7120
rect 27531 7076 27573 7085
rect 27531 7036 27532 7076
rect 27572 7036 27573 7076
rect 27531 7027 27573 7036
rect 27435 6908 27477 6917
rect 27628 6908 27668 8044
rect 27916 8000 27956 8371
rect 27916 7951 27956 7960
rect 28396 7995 28436 9220
rect 28396 7946 28436 7955
rect 28492 7925 28532 9472
rect 29260 9353 29300 9631
rect 29547 9596 29589 9605
rect 29547 9556 29548 9596
rect 29588 9556 29589 9596
rect 29547 9547 29589 9556
rect 29548 9512 29588 9547
rect 29548 9461 29588 9472
rect 29259 9344 29301 9353
rect 29259 9304 29260 9344
rect 29300 9304 29301 9344
rect 29259 9295 29301 9304
rect 30220 9260 30260 9269
rect 29739 8756 29781 8765
rect 29739 8716 29740 8756
rect 29780 8716 29781 8756
rect 29739 8707 29781 8716
rect 28779 8672 28821 8681
rect 28779 8632 28780 8672
rect 28820 8632 28821 8672
rect 28779 8623 28821 8632
rect 29644 8672 29684 8681
rect 28780 8538 28820 8623
rect 28587 8084 28629 8093
rect 28587 8044 28588 8084
rect 28628 8044 28629 8084
rect 28587 8035 28629 8044
rect 29355 8084 29397 8093
rect 29355 8044 29356 8084
rect 29396 8044 29397 8084
rect 29355 8035 29397 8044
rect 28588 7950 28628 8035
rect 28972 8000 29012 8009
rect 28491 7916 28533 7925
rect 28491 7876 28492 7916
rect 28532 7876 28533 7916
rect 28491 7867 28533 7876
rect 28779 7916 28821 7925
rect 28779 7876 28780 7916
rect 28820 7876 28821 7916
rect 28779 7867 28821 7876
rect 28780 7253 28820 7867
rect 28972 7841 29012 7960
rect 28971 7832 29013 7841
rect 28971 7792 28972 7832
rect 29012 7792 29013 7832
rect 28971 7783 29013 7792
rect 28203 7244 28245 7253
rect 28203 7204 28204 7244
rect 28244 7204 28245 7244
rect 28203 7195 28245 7204
rect 28779 7244 28821 7253
rect 28779 7204 28780 7244
rect 28820 7204 28821 7244
rect 28779 7195 28821 7204
rect 29356 7244 29396 8035
rect 29548 7328 29588 7337
rect 29644 7328 29684 8632
rect 29588 7288 29684 7328
rect 29548 7279 29588 7288
rect 29356 7195 29396 7204
rect 27819 6992 27861 7001
rect 27819 6952 27820 6992
rect 27860 6952 27861 6992
rect 27819 6943 27861 6952
rect 27435 6868 27436 6908
rect 27476 6868 27477 6908
rect 27435 6859 27477 6868
rect 27532 6868 27668 6908
rect 27147 6824 27189 6833
rect 27147 6784 27148 6824
rect 27188 6784 27189 6824
rect 27147 6775 27189 6784
rect 27052 6439 27092 6448
rect 27148 6488 27188 6775
rect 27435 6656 27477 6665
rect 27435 6616 27436 6656
rect 27476 6616 27477 6656
rect 27435 6607 27477 6616
rect 27148 6439 27188 6448
rect 26955 6320 26997 6329
rect 26955 6280 26956 6320
rect 26996 6280 26997 6320
rect 26955 6271 26997 6280
rect 27147 6236 27189 6245
rect 27147 6196 27148 6236
rect 27188 6196 27189 6236
rect 27147 6187 27189 6196
rect 26476 5860 26708 5900
rect 25948 5692 26036 5732
rect 26091 5732 26133 5741
rect 26091 5692 26092 5732
rect 26132 5692 26133 5732
rect 25948 5690 25988 5692
rect 26091 5683 26133 5692
rect 26475 5732 26517 5741
rect 26475 5692 26476 5732
rect 26516 5692 26517 5732
rect 26475 5683 26517 5692
rect 25948 5641 25988 5650
rect 26092 5564 26132 5683
rect 26476 5598 26516 5683
rect 26092 5515 26132 5524
rect 26284 5480 26324 5489
rect 25804 4481 25844 4936
rect 26187 4976 26229 4985
rect 26187 4936 26188 4976
rect 26228 4936 26229 4976
rect 26187 4927 26229 4936
rect 25996 4724 26036 4733
rect 25803 4472 25845 4481
rect 25803 4432 25804 4472
rect 25844 4432 25845 4472
rect 25803 4423 25845 4432
rect 25707 4388 25749 4397
rect 25707 4348 25708 4388
rect 25748 4348 25749 4388
rect 25707 4339 25749 4348
rect 25708 4061 25748 4339
rect 25996 4304 26036 4684
rect 26188 4481 26228 4927
rect 26187 4472 26229 4481
rect 26187 4432 26188 4472
rect 26228 4432 26229 4472
rect 26187 4423 26229 4432
rect 25852 4264 26036 4304
rect 25852 4145 25892 4264
rect 25852 4096 25892 4105
rect 26188 4136 26228 4423
rect 26188 4087 26228 4096
rect 25707 4052 25749 4061
rect 25707 4012 25708 4052
rect 25748 4012 25749 4052
rect 25707 4003 25749 4012
rect 25996 4052 26036 4061
rect 26091 4052 26133 4061
rect 26036 4012 26092 4052
rect 26132 4012 26133 4052
rect 25996 4003 26036 4012
rect 26091 4003 26133 4012
rect 25707 3800 25749 3809
rect 25707 3760 25708 3800
rect 25748 3760 25749 3800
rect 25707 3751 25749 3760
rect 25611 3632 25653 3641
rect 25611 3592 25612 3632
rect 25652 3592 25653 3632
rect 25611 3583 25653 3592
rect 25516 3464 25556 3473
rect 25516 2801 25556 3424
rect 25612 3464 25652 3473
rect 25612 3305 25652 3424
rect 25611 3296 25653 3305
rect 25611 3256 25612 3296
rect 25652 3256 25653 3296
rect 25611 3247 25653 3256
rect 25708 3044 25748 3751
rect 26091 3632 26133 3641
rect 26091 3592 26092 3632
rect 26132 3592 26133 3632
rect 26091 3583 26133 3592
rect 26092 3464 26132 3583
rect 26092 3415 26132 3424
rect 25612 3004 25748 3044
rect 25996 3380 26036 3389
rect 25515 2792 25557 2801
rect 25515 2752 25516 2792
rect 25556 2752 25557 2792
rect 25515 2743 25557 2752
rect 25516 2624 25556 2633
rect 25612 2624 25652 3004
rect 25707 2792 25749 2801
rect 25707 2752 25708 2792
rect 25748 2752 25749 2792
rect 25707 2743 25749 2752
rect 25708 2658 25748 2743
rect 25996 2633 26036 3340
rect 26284 3296 26324 5440
rect 26572 4892 26612 4901
rect 26572 4229 26612 4852
rect 26668 4556 26708 5860
rect 27148 5732 27188 6187
rect 27148 5683 27188 5692
rect 27340 5480 27380 5489
rect 26956 4976 26996 4987
rect 26956 4901 26996 4936
rect 26955 4892 26997 4901
rect 26955 4852 26956 4892
rect 26996 4852 26997 4892
rect 26955 4843 26997 4852
rect 26764 4724 26804 4733
rect 27051 4724 27093 4733
rect 26804 4684 26996 4724
rect 26764 4675 26804 4684
rect 26668 4516 26804 4556
rect 26571 4220 26613 4229
rect 26571 4180 26572 4220
rect 26612 4180 26613 4220
rect 26571 4171 26613 4180
rect 26379 4052 26421 4061
rect 26379 4012 26380 4052
rect 26420 4012 26421 4052
rect 26379 4003 26421 4012
rect 26667 4052 26709 4061
rect 26667 4012 26668 4052
rect 26708 4012 26709 4052
rect 26667 4003 26709 4012
rect 26092 3256 26324 3296
rect 25556 2584 25652 2624
rect 25995 2624 26037 2633
rect 25995 2584 25996 2624
rect 26036 2584 26037 2624
rect 25516 2575 25556 2584
rect 25995 2575 26037 2584
rect 25995 2120 26037 2129
rect 25995 2080 25996 2120
rect 26036 2080 26037 2120
rect 25995 2071 26037 2080
rect 25996 1986 26036 2071
rect 26092 1961 26132 3256
rect 26188 2624 26228 2633
rect 26188 2120 26228 2584
rect 26284 2624 26324 2633
rect 26284 2213 26324 2584
rect 26380 2381 26420 4003
rect 26572 3473 26612 3558
rect 26571 3464 26613 3473
rect 26571 3424 26572 3464
rect 26612 3424 26613 3464
rect 26571 3415 26613 3424
rect 26668 3296 26708 4003
rect 26572 3256 26708 3296
rect 26475 2792 26517 2801
rect 26475 2752 26476 2792
rect 26516 2752 26517 2792
rect 26475 2743 26517 2752
rect 26379 2372 26421 2381
rect 26379 2332 26380 2372
rect 26420 2332 26421 2372
rect 26379 2323 26421 2332
rect 26283 2204 26325 2213
rect 26283 2164 26284 2204
rect 26324 2164 26325 2204
rect 26283 2155 26325 2164
rect 26188 2071 26228 2080
rect 26380 1961 26420 2046
rect 26091 1952 26133 1961
rect 25324 1408 25460 1448
rect 25804 1938 25844 1947
rect 26091 1912 26092 1952
rect 26132 1912 26133 1952
rect 26091 1903 26133 1912
rect 26379 1952 26421 1961
rect 26379 1912 26380 1952
rect 26420 1912 26421 1952
rect 26379 1903 26421 1912
rect 25324 944 25364 1408
rect 25612 1364 25652 1373
rect 25804 1364 25844 1898
rect 26476 1784 26516 2743
rect 26380 1744 26516 1784
rect 26187 1448 26229 1457
rect 26187 1408 26188 1448
rect 26228 1408 26229 1448
rect 26187 1399 26229 1408
rect 25652 1324 25844 1364
rect 25612 1315 25652 1324
rect 25995 1196 26037 1205
rect 25995 1156 25996 1196
rect 26036 1156 26037 1196
rect 25995 1147 26037 1156
rect 25611 1112 25653 1121
rect 25420 1070 25460 1079
rect 25611 1072 25612 1112
rect 25652 1072 25653 1112
rect 25611 1063 25653 1072
rect 25804 1112 25844 1121
rect 25420 1028 25460 1030
rect 25420 988 25556 1028
rect 25324 904 25460 944
rect 25420 80 25460 904
rect 25516 701 25556 988
rect 25515 692 25557 701
rect 25515 652 25516 692
rect 25556 652 25557 692
rect 25515 643 25557 652
rect 25612 80 25652 1063
rect 25707 1028 25749 1037
rect 25804 1028 25844 1072
rect 25707 988 25708 1028
rect 25748 988 25844 1028
rect 25707 979 25749 988
rect 25803 692 25845 701
rect 25803 652 25804 692
rect 25844 652 25845 692
rect 25803 643 25845 652
rect 25804 80 25844 643
rect 25996 80 26036 1147
rect 26188 80 26228 1399
rect 26380 80 26420 1744
rect 26572 701 26612 3256
rect 26764 2666 26804 4516
rect 26859 4136 26901 4145
rect 26859 4096 26860 4136
rect 26900 4096 26901 4136
rect 26859 4087 26901 4096
rect 26668 2624 26708 2633
rect 26764 2617 26804 2626
rect 26668 1793 26708 2584
rect 26667 1784 26709 1793
rect 26667 1744 26668 1784
rect 26708 1744 26709 1784
rect 26667 1735 26709 1744
rect 26860 1205 26900 4087
rect 26956 2540 26996 4684
rect 27051 4684 27052 4724
rect 27092 4684 27093 4724
rect 27051 4675 27093 4684
rect 27052 4397 27092 4675
rect 27051 4388 27093 4397
rect 27051 4348 27052 4388
rect 27092 4348 27093 4388
rect 27051 4339 27093 4348
rect 27340 4145 27380 5440
rect 27339 4136 27381 4145
rect 27339 4096 27340 4136
rect 27380 4096 27381 4136
rect 27339 4087 27381 4096
rect 27436 4136 27476 6607
rect 27532 6488 27572 6868
rect 27532 6439 27572 6448
rect 27628 6404 27668 6413
rect 27628 6068 27668 6364
rect 27532 6028 27668 6068
rect 27532 4556 27572 6028
rect 27627 5900 27669 5909
rect 27627 5860 27628 5900
rect 27668 5860 27669 5900
rect 27627 5851 27669 5860
rect 27628 5657 27668 5851
rect 27627 5648 27669 5657
rect 27627 5608 27628 5648
rect 27668 5608 27669 5648
rect 27627 5599 27669 5608
rect 27628 5514 27668 5599
rect 27532 4516 27764 4556
rect 27147 3884 27189 3893
rect 27147 3844 27148 3884
rect 27188 3844 27189 3884
rect 27147 3835 27189 3844
rect 27148 3716 27188 3835
rect 27436 3809 27476 4096
rect 27628 3968 27668 3977
rect 27628 3809 27668 3928
rect 27435 3800 27477 3809
rect 27435 3760 27436 3800
rect 27476 3760 27477 3800
rect 27435 3751 27477 3760
rect 27627 3800 27669 3809
rect 27627 3760 27628 3800
rect 27668 3760 27669 3800
rect 27627 3751 27669 3760
rect 27130 3676 27188 3716
rect 27130 3548 27170 3676
rect 27052 3508 27170 3548
rect 27244 3548 27284 3557
rect 27627 3548 27669 3557
rect 27284 3508 27380 3548
rect 27052 3450 27092 3508
rect 27244 3499 27284 3508
rect 27052 3401 27092 3410
rect 27243 3212 27285 3221
rect 27243 3172 27244 3212
rect 27284 3172 27285 3212
rect 27243 3163 27285 3172
rect 27244 2624 27284 3163
rect 27244 2575 27284 2584
rect 26956 2500 27188 2540
rect 26955 1952 26997 1961
rect 26955 1912 26956 1952
rect 26996 1912 26997 1952
rect 26955 1903 26997 1912
rect 26859 1196 26901 1205
rect 26859 1156 26860 1196
rect 26900 1156 26901 1196
rect 26859 1147 26901 1156
rect 26571 692 26613 701
rect 26571 652 26572 692
rect 26612 652 26613 692
rect 26571 643 26613 652
rect 26571 440 26613 449
rect 26571 400 26572 440
rect 26612 400 26613 440
rect 26571 391 26613 400
rect 26572 80 26612 391
rect 26763 104 26805 113
rect 26763 80 26764 104
rect 24500 64 24520 80
rect 24440 0 24520 64
rect 24632 0 24712 80
rect 24824 0 24904 80
rect 25016 0 25096 80
rect 25208 0 25288 80
rect 25400 0 25480 80
rect 25592 0 25672 80
rect 25784 0 25864 80
rect 25976 0 26056 80
rect 26168 0 26248 80
rect 26360 0 26440 80
rect 26552 0 26632 80
rect 26744 64 26764 80
rect 26804 80 26805 104
rect 26956 80 26996 1903
rect 27052 1112 27092 1121
rect 27052 869 27092 1072
rect 27051 860 27093 869
rect 27051 820 27052 860
rect 27092 820 27093 860
rect 27051 811 27093 820
rect 27051 692 27093 701
rect 27051 652 27052 692
rect 27092 652 27093 692
rect 27051 643 27093 652
rect 27052 188 27092 643
rect 27148 365 27188 2500
rect 27340 1877 27380 3508
rect 27627 3508 27628 3548
rect 27668 3508 27669 3548
rect 27627 3499 27669 3508
rect 27628 3380 27668 3499
rect 27628 3331 27668 3340
rect 27724 3305 27764 4516
rect 27723 3296 27765 3305
rect 27723 3256 27724 3296
rect 27764 3256 27765 3296
rect 27723 3247 27765 3256
rect 27436 3212 27476 3221
rect 27436 1961 27476 3172
rect 27724 2633 27764 2642
rect 27532 2593 27724 2624
rect 27532 2584 27764 2593
rect 27435 1952 27477 1961
rect 27435 1912 27436 1952
rect 27476 1912 27477 1952
rect 27435 1903 27477 1912
rect 27339 1868 27381 1877
rect 27339 1828 27340 1868
rect 27380 1828 27381 1868
rect 27339 1819 27381 1828
rect 27339 1700 27381 1709
rect 27339 1660 27340 1700
rect 27380 1660 27381 1700
rect 27339 1651 27381 1660
rect 27243 1280 27285 1289
rect 27243 1240 27244 1280
rect 27284 1240 27285 1280
rect 27243 1231 27285 1240
rect 27244 1146 27284 1231
rect 27147 356 27189 365
rect 27147 316 27148 356
rect 27188 316 27189 356
rect 27147 307 27189 316
rect 27052 148 27188 188
rect 27148 80 27188 148
rect 27340 80 27380 1651
rect 27532 1289 27572 2584
rect 27820 2540 27860 6943
rect 28108 6488 28148 6497
rect 28011 6068 28053 6077
rect 28011 6028 28012 6068
rect 28052 6028 28053 6068
rect 28011 6019 28053 6028
rect 28012 2549 28052 6019
rect 28108 5825 28148 6448
rect 28107 5816 28149 5825
rect 28107 5776 28108 5816
rect 28148 5776 28149 5816
rect 28107 5767 28149 5776
rect 28204 5405 28244 7195
rect 28780 7160 28820 7195
rect 28780 7109 28820 7120
rect 28972 6992 29012 7001
rect 28684 6952 28972 6992
rect 28684 6488 28724 6952
rect 28972 6943 29012 6952
rect 29164 6992 29204 7001
rect 29164 6656 29204 6952
rect 28876 6616 29204 6656
rect 28636 6478 28724 6488
rect 28676 6448 28724 6478
rect 28780 6572 28820 6581
rect 28636 6429 28676 6438
rect 28780 5816 28820 6532
rect 28684 5776 28820 5816
rect 28876 5816 28916 6616
rect 29164 6488 29204 6499
rect 29164 6413 29204 6448
rect 29163 6404 29205 6413
rect 29163 6364 29164 6404
rect 29204 6364 29205 6404
rect 29163 6355 29205 6364
rect 28972 6236 29012 6245
rect 29451 6236 29493 6245
rect 29012 6196 29396 6236
rect 28972 6187 29012 6196
rect 28876 5776 29012 5816
rect 28203 5396 28245 5405
rect 28203 5356 28204 5396
rect 28244 5356 28245 5396
rect 28203 5347 28245 5356
rect 28204 4976 28244 5347
rect 28204 4927 28244 4936
rect 28684 4892 28724 5776
rect 28876 5648 28916 5657
rect 28876 5564 28916 5608
rect 28780 5524 28916 5564
rect 28780 5405 28820 5524
rect 28972 5480 29012 5776
rect 29356 5648 29396 6196
rect 29451 6196 29452 6236
rect 29492 6196 29493 6236
rect 29451 6187 29493 6196
rect 29452 5909 29492 6187
rect 29451 5900 29493 5909
rect 29451 5860 29452 5900
rect 29492 5860 29493 5900
rect 29451 5851 29493 5860
rect 29356 5599 29396 5608
rect 29452 5648 29492 5851
rect 29643 5816 29685 5825
rect 29643 5776 29644 5816
rect 29684 5776 29685 5816
rect 29643 5767 29685 5776
rect 29452 5599 29492 5608
rect 29068 5564 29108 5573
rect 29108 5524 29300 5564
rect 29068 5515 29108 5524
rect 28876 5440 29012 5480
rect 28779 5396 28821 5405
rect 28779 5356 28780 5396
rect 28820 5356 28821 5396
rect 28779 5347 28821 5356
rect 28780 4892 28820 4901
rect 28684 4852 28780 4892
rect 28780 4843 28820 4852
rect 28396 4724 28436 4733
rect 28588 4724 28628 4733
rect 28108 4684 28396 4724
rect 28108 4136 28148 4684
rect 28396 4675 28436 4684
rect 28492 4684 28588 4724
rect 28108 4087 28148 4096
rect 28204 4136 28244 4145
rect 28244 4096 28340 4136
rect 28204 4087 28244 4096
rect 28204 3464 28244 3473
rect 28108 2876 28148 2885
rect 28204 2876 28244 3424
rect 28300 3464 28340 4096
rect 28300 3305 28340 3424
rect 28299 3296 28341 3305
rect 28299 3256 28300 3296
rect 28340 3256 28341 3296
rect 28299 3247 28341 3256
rect 28299 3128 28341 3137
rect 28299 3088 28300 3128
rect 28340 3088 28341 3128
rect 28299 3079 28341 3088
rect 28148 2836 28244 2876
rect 28108 2827 28148 2836
rect 28300 2633 28340 3079
rect 28299 2624 28341 2633
rect 28299 2584 28300 2624
rect 28340 2584 28341 2624
rect 28299 2575 28341 2584
rect 27724 2500 27860 2540
rect 28011 2540 28053 2549
rect 28011 2500 28012 2540
rect 28052 2500 28053 2540
rect 27627 2288 27669 2297
rect 27627 2248 27628 2288
rect 27668 2248 27669 2288
rect 27627 2239 27669 2248
rect 27628 1952 27668 2239
rect 27628 1903 27668 1912
rect 27531 1280 27573 1289
rect 27531 1240 27532 1280
rect 27572 1240 27573 1280
rect 27531 1231 27573 1240
rect 27435 1112 27477 1121
rect 27435 1072 27436 1112
rect 27476 1072 27477 1112
rect 27435 1063 27477 1072
rect 27436 978 27476 1063
rect 27531 356 27573 365
rect 27531 316 27532 356
rect 27572 316 27573 356
rect 27531 307 27573 316
rect 27532 80 27572 307
rect 27724 80 27764 2500
rect 28011 2491 28053 2500
rect 27915 2456 27957 2465
rect 27915 2416 27916 2456
rect 27956 2416 27957 2456
rect 27915 2407 27957 2416
rect 27916 2322 27956 2407
rect 28011 2372 28053 2381
rect 28492 2372 28532 4684
rect 28588 4675 28628 4684
rect 28587 4556 28629 4565
rect 28587 4516 28588 4556
rect 28628 4516 28629 4556
rect 28587 4507 28629 4516
rect 28588 4220 28628 4507
rect 28588 3464 28628 4180
rect 28684 4136 28724 4145
rect 28724 4096 28820 4136
rect 28684 4087 28724 4096
rect 28684 3464 28724 3473
rect 28588 3424 28684 3464
rect 28684 3415 28724 3424
rect 28780 3380 28820 4096
rect 28780 2885 28820 3340
rect 28779 2876 28821 2885
rect 28779 2836 28780 2876
rect 28820 2836 28821 2876
rect 28779 2827 28821 2836
rect 28011 2332 28012 2372
rect 28052 2332 28053 2372
rect 28011 2323 28053 2332
rect 28300 2332 28532 2372
rect 28012 1868 28052 2323
rect 28012 1819 28052 1828
rect 27819 1700 27861 1709
rect 27819 1660 27820 1700
rect 27860 1660 27861 1700
rect 27819 1651 27861 1660
rect 28204 1700 28244 1709
rect 27820 1566 27860 1651
rect 27915 1196 27957 1205
rect 27915 1156 27916 1196
rect 27956 1156 27957 1196
rect 27915 1147 27957 1156
rect 27916 80 27956 1147
rect 28204 953 28244 1660
rect 28203 944 28245 953
rect 28203 904 28204 944
rect 28244 904 28245 944
rect 28203 895 28245 904
rect 28107 272 28149 281
rect 28107 232 28108 272
rect 28148 232 28149 272
rect 28107 223 28149 232
rect 28108 80 28148 223
rect 28300 80 28340 2332
rect 28395 1868 28437 1877
rect 28395 1828 28396 1868
rect 28436 1828 28437 1868
rect 28395 1819 28437 1828
rect 28396 1734 28436 1819
rect 28876 1448 28916 5440
rect 29260 5228 29300 5524
rect 29260 5188 29588 5228
rect 29163 5060 29205 5069
rect 29163 5020 29164 5060
rect 29204 5020 29205 5060
rect 29163 5011 29205 5020
rect 29355 5060 29397 5069
rect 29355 5020 29356 5060
rect 29396 5020 29397 5060
rect 29355 5011 29397 5020
rect 29164 4136 29204 5011
rect 29164 4087 29204 4096
rect 29260 4724 29300 4733
rect 29260 4061 29300 4684
rect 29259 4052 29301 4061
rect 29259 4012 29260 4052
rect 29300 4012 29301 4052
rect 29259 4003 29301 4012
rect 29067 3800 29109 3809
rect 29067 3760 29068 3800
rect 29108 3760 29109 3800
rect 29067 3751 29109 3760
rect 28780 1408 28916 1448
rect 28972 1952 29012 1961
rect 28683 1112 28725 1121
rect 28683 1072 28684 1112
rect 28724 1072 28725 1112
rect 28780 1112 28820 1408
rect 28876 1280 28916 1289
rect 28972 1280 29012 1912
rect 29068 1952 29108 3751
rect 29260 3464 29300 3473
rect 29356 3464 29396 5011
rect 29452 4892 29492 4901
rect 29452 3641 29492 4852
rect 29548 4150 29588 5188
rect 29644 4976 29684 5767
rect 29644 4927 29684 4936
rect 29644 4150 29684 4159
rect 29548 4110 29644 4150
rect 29644 4101 29684 4110
rect 29740 4052 29780 8707
rect 30220 8681 30260 9220
rect 30507 8924 30549 8933
rect 30507 8884 30508 8924
rect 30548 8884 30549 8924
rect 30507 8875 30549 8884
rect 30219 8672 30261 8681
rect 30219 8632 30220 8672
rect 30260 8632 30261 8672
rect 30219 8623 30261 8632
rect 30028 8588 30068 8597
rect 29836 8548 30028 8588
rect 29836 6833 29876 8548
rect 30028 8539 30068 8548
rect 30219 8084 30261 8093
rect 30219 8044 30220 8084
rect 30260 8044 30261 8084
rect 30219 8035 30261 8044
rect 30220 8000 30260 8035
rect 30220 7925 30260 7960
rect 30219 7916 30261 7925
rect 30219 7876 30220 7916
rect 30260 7876 30261 7916
rect 30219 7867 30261 7876
rect 29931 7832 29973 7841
rect 30220 7836 30260 7867
rect 29931 7792 29932 7832
rect 29972 7792 29973 7832
rect 29931 7783 29973 7792
rect 29932 6917 29972 7783
rect 30027 7748 30069 7757
rect 30027 7708 30028 7748
rect 30068 7708 30069 7748
rect 30027 7699 30069 7708
rect 30411 7748 30453 7757
rect 30411 7708 30412 7748
rect 30452 7708 30453 7748
rect 30411 7699 30453 7708
rect 30028 7160 30068 7699
rect 30412 7614 30452 7699
rect 30411 7496 30453 7505
rect 30411 7456 30412 7496
rect 30452 7456 30453 7496
rect 30411 7447 30453 7456
rect 30412 7253 30452 7447
rect 30411 7244 30453 7253
rect 30411 7204 30412 7244
rect 30452 7204 30453 7244
rect 30411 7195 30453 7204
rect 30028 7111 30068 7120
rect 30124 7160 30164 7169
rect 29931 6908 29973 6917
rect 29931 6868 29932 6908
rect 29972 6868 29973 6908
rect 29931 6859 29973 6868
rect 29835 6824 29877 6833
rect 29835 6784 29836 6824
rect 29876 6784 29877 6824
rect 29835 6775 29877 6784
rect 29931 6740 29973 6749
rect 29931 6700 29932 6740
rect 29972 6700 29973 6740
rect 29931 6691 29973 6700
rect 29932 5732 29972 6691
rect 30027 6656 30069 6665
rect 30027 6616 30028 6656
rect 30068 6616 30069 6656
rect 30027 6607 30069 6616
rect 29836 5648 29876 5657
rect 29836 5321 29876 5608
rect 29835 5312 29877 5321
rect 29835 5272 29836 5312
rect 29876 5272 29877 5312
rect 29835 5263 29877 5272
rect 29932 5069 29972 5692
rect 29931 5060 29973 5069
rect 29931 5020 29932 5060
rect 29972 5020 29973 5060
rect 29931 5011 29973 5020
rect 30028 4136 30068 6607
rect 29644 4012 29780 4052
rect 29932 4096 30068 4136
rect 29547 3884 29589 3893
rect 29547 3844 29548 3884
rect 29588 3844 29589 3884
rect 29547 3835 29589 3844
rect 29451 3632 29493 3641
rect 29451 3592 29452 3632
rect 29492 3592 29493 3632
rect 29451 3583 29493 3592
rect 29548 3464 29588 3835
rect 29300 3424 29396 3464
rect 29452 3424 29588 3464
rect 29260 3415 29300 3424
rect 29163 2540 29205 2549
rect 29163 2500 29164 2540
rect 29204 2500 29205 2540
rect 29163 2491 29205 2500
rect 29068 1709 29108 1912
rect 29067 1700 29109 1709
rect 29067 1660 29068 1700
rect 29108 1660 29109 1700
rect 29067 1651 29109 1660
rect 28916 1240 29012 1280
rect 28876 1231 28916 1240
rect 29164 1121 29204 2491
rect 29452 1877 29492 3424
rect 29547 3044 29589 3053
rect 29547 3004 29548 3044
rect 29588 3004 29589 3044
rect 29547 2995 29589 3004
rect 29548 2624 29588 2995
rect 29548 2575 29588 2584
rect 29547 2120 29589 2129
rect 29547 2080 29548 2120
rect 29588 2080 29589 2120
rect 29547 2071 29589 2080
rect 29451 1868 29493 1877
rect 29451 1828 29452 1868
rect 29492 1828 29493 1868
rect 29451 1819 29493 1828
rect 29548 1868 29588 2071
rect 29452 1734 29492 1819
rect 29259 1700 29301 1709
rect 29259 1660 29260 1700
rect 29300 1660 29301 1700
rect 29259 1651 29301 1660
rect 29068 1112 29108 1121
rect 29163 1112 29205 1121
rect 28780 1072 28916 1112
rect 28683 1063 28725 1072
rect 28684 978 28724 1063
rect 28491 692 28533 701
rect 28491 652 28492 692
rect 28532 652 28533 692
rect 28491 643 28533 652
rect 28492 80 28532 643
rect 28683 188 28725 197
rect 28683 148 28684 188
rect 28724 148 28725 188
rect 28683 139 28725 148
rect 28684 80 28724 139
rect 28876 80 28916 1072
rect 29108 1072 29164 1112
rect 29204 1072 29205 1112
rect 29068 1063 29108 1072
rect 29163 1063 29205 1072
rect 29164 978 29204 1063
rect 29067 944 29109 953
rect 29067 904 29068 944
rect 29108 904 29109 944
rect 29067 895 29109 904
rect 29068 80 29108 895
rect 29260 80 29300 1651
rect 29548 1541 29588 1828
rect 29547 1532 29589 1541
rect 29547 1492 29548 1532
rect 29588 1492 29589 1532
rect 29547 1483 29589 1492
rect 29451 1364 29493 1373
rect 29451 1324 29452 1364
rect 29492 1324 29493 1364
rect 29451 1315 29493 1324
rect 29452 80 29492 1315
rect 29644 80 29684 4012
rect 29836 3968 29876 3977
rect 29740 3450 29780 3459
rect 29740 2876 29780 3410
rect 29740 2827 29780 2836
rect 29836 1961 29876 3928
rect 29932 3809 29972 4096
rect 30028 3968 30068 3977
rect 29931 3800 29973 3809
rect 29931 3760 29932 3800
rect 29972 3760 29973 3800
rect 29931 3751 29973 3760
rect 29931 3632 29973 3641
rect 29931 3592 29932 3632
rect 29972 3592 29973 3632
rect 29931 3583 29973 3592
rect 29932 3498 29972 3583
rect 30028 3473 30068 3928
rect 30124 3893 30164 7120
rect 30508 7160 30548 8875
rect 30604 8168 30644 10672
rect 30700 9512 30740 9521
rect 30700 8933 30740 9472
rect 31084 9428 31124 9437
rect 30699 8924 30741 8933
rect 30699 8884 30700 8924
rect 30740 8884 30741 8924
rect 30699 8875 30741 8884
rect 30891 8840 30933 8849
rect 30891 8800 30892 8840
rect 30932 8800 30933 8840
rect 30891 8791 30933 8800
rect 30892 8706 30932 8791
rect 31084 8672 31124 9388
rect 31084 8623 31124 8632
rect 31564 8588 31604 8597
rect 31564 8177 31604 8548
rect 31083 8168 31125 8177
rect 30604 8128 30740 8168
rect 30604 8000 30644 8009
rect 30604 7505 30644 7960
rect 30700 7589 30740 8128
rect 31083 8128 31084 8168
rect 31124 8128 31125 8168
rect 31083 8119 31125 8128
rect 31563 8168 31605 8177
rect 31563 8128 31564 8168
rect 31604 8128 31605 8168
rect 31563 8119 31605 8128
rect 30699 7580 30741 7589
rect 30699 7540 30700 7580
rect 30740 7540 30741 7580
rect 30699 7531 30741 7540
rect 30603 7496 30645 7505
rect 30603 7456 30604 7496
rect 30644 7456 30645 7496
rect 30603 7447 30645 7456
rect 31084 7169 31124 8119
rect 31563 8000 31605 8009
rect 31563 7960 31564 8000
rect 31604 7960 31605 8000
rect 31563 7951 31605 7960
rect 31564 7328 31604 7951
rect 31756 7925 31796 10672
rect 32235 10648 32236 10688
rect 32276 10648 32277 10688
rect 32888 10672 32968 10752
rect 33196 10692 33428 10732
rect 32235 10639 32277 10648
rect 32236 9680 32276 10639
rect 32908 10604 32948 10672
rect 33196 10604 33236 10692
rect 32908 10564 33236 10604
rect 32331 10436 32373 10445
rect 32331 10396 32332 10436
rect 32372 10396 32373 10436
rect 32331 10387 32373 10396
rect 32236 9631 32276 9640
rect 31852 9512 31892 9521
rect 31852 8765 31892 9472
rect 31851 8756 31893 8765
rect 31851 8716 31852 8756
rect 31892 8716 31893 8756
rect 31851 8707 31893 8716
rect 31948 8672 31988 8681
rect 31988 8632 32180 8672
rect 31948 8623 31988 8632
rect 31851 8084 31893 8093
rect 31851 8044 31852 8084
rect 31892 8044 31893 8084
rect 31851 8035 31893 8044
rect 31852 8000 31892 8035
rect 31852 7949 31892 7960
rect 31755 7916 31797 7925
rect 31755 7876 31756 7916
rect 31796 7876 31797 7916
rect 31755 7867 31797 7876
rect 32140 7757 32180 8632
rect 32044 7748 32084 7757
rect 31468 7288 31604 7328
rect 31660 7708 32044 7748
rect 30315 7076 30357 7085
rect 30315 7036 30316 7076
rect 30356 7036 30357 7076
rect 30315 7027 30357 7036
rect 30316 5900 30356 7027
rect 30411 6488 30453 6497
rect 30411 6448 30412 6488
rect 30452 6448 30453 6488
rect 30411 6439 30453 6448
rect 30412 6354 30452 6439
rect 30316 5860 30452 5900
rect 30412 5741 30452 5860
rect 30411 5732 30453 5741
rect 30411 5692 30412 5732
rect 30452 5692 30453 5732
rect 30411 5683 30453 5692
rect 30412 5648 30452 5683
rect 30412 5598 30452 5608
rect 30508 5405 30548 7120
rect 30604 7160 30644 7169
rect 30507 5396 30549 5405
rect 30507 5356 30508 5396
rect 30548 5356 30549 5396
rect 30507 5347 30549 5356
rect 30219 4808 30261 4817
rect 30219 4768 30220 4808
rect 30260 4768 30261 4808
rect 30219 4759 30261 4768
rect 30220 4136 30260 4759
rect 30220 4087 30260 4096
rect 30123 3884 30165 3893
rect 30123 3844 30124 3884
rect 30164 3844 30165 3884
rect 30123 3835 30165 3844
rect 30027 3464 30069 3473
rect 30027 3424 30028 3464
rect 30068 3424 30069 3464
rect 30027 3415 30069 3424
rect 30411 3464 30453 3473
rect 30411 3424 30412 3464
rect 30452 3424 30453 3464
rect 30411 3415 30453 3424
rect 30508 3464 30548 3473
rect 30604 3464 30644 7120
rect 31083 7160 31125 7169
rect 31083 7120 31084 7160
rect 31124 7120 31125 7160
rect 31083 7111 31125 7120
rect 31084 7026 31124 7111
rect 31468 7076 31508 7288
rect 31660 7244 31700 7708
rect 32044 7699 32084 7708
rect 32139 7748 32181 7757
rect 32139 7708 32140 7748
rect 32180 7708 32181 7748
rect 32139 7699 32181 7708
rect 32236 7748 32276 7757
rect 32043 7580 32085 7589
rect 32043 7540 32044 7580
rect 32084 7540 32085 7580
rect 32043 7531 32085 7540
rect 31612 7204 31700 7244
rect 31755 7244 31797 7253
rect 31755 7204 31756 7244
rect 31796 7204 31797 7244
rect 31612 7202 31652 7204
rect 31755 7195 31797 7204
rect 31612 7153 31652 7162
rect 31756 7076 31796 7195
rect 31468 7036 31700 7076
rect 30699 6488 30741 6497
rect 30699 6448 30700 6488
rect 30740 6448 30741 6488
rect 30699 6439 30741 6448
rect 30700 6354 30740 6439
rect 30795 6404 30837 6413
rect 30795 6364 30796 6404
rect 30836 6364 30837 6404
rect 30795 6355 30837 6364
rect 30796 6236 30836 6355
rect 30700 6196 30836 6236
rect 30700 4724 30740 6196
rect 31563 6152 31605 6161
rect 31563 6112 31564 6152
rect 31604 6112 31605 6152
rect 31563 6103 31605 6112
rect 31468 5732 31508 5741
rect 31180 5692 31468 5732
rect 30940 5657 30980 5666
rect 30980 5617 31028 5648
rect 30940 5608 31028 5617
rect 30988 5144 31028 5608
rect 31084 5564 31124 5573
rect 31180 5564 31220 5692
rect 31468 5683 31508 5692
rect 31124 5524 31220 5564
rect 31084 5515 31124 5524
rect 31276 5480 31316 5489
rect 31179 5312 31221 5321
rect 31179 5272 31180 5312
rect 31220 5272 31221 5312
rect 31179 5263 31221 5272
rect 31084 5144 31124 5153
rect 30988 5104 31084 5144
rect 31084 5095 31124 5104
rect 30892 4976 30932 4985
rect 31180 4976 31220 5263
rect 31276 5153 31316 5440
rect 31371 5480 31413 5489
rect 31371 5440 31372 5480
rect 31412 5440 31413 5480
rect 31371 5431 31413 5440
rect 31275 5144 31317 5153
rect 31275 5104 31276 5144
rect 31316 5104 31317 5144
rect 31275 5095 31317 5104
rect 30892 4724 30932 4936
rect 30700 4684 30932 4724
rect 30988 4936 31220 4976
rect 31276 4976 31316 4985
rect 30699 4388 30741 4397
rect 30699 4348 30700 4388
rect 30740 4348 30741 4388
rect 30699 4339 30741 4348
rect 30548 3424 30644 3464
rect 30412 3330 30452 3415
rect 30219 2876 30261 2885
rect 30219 2836 30220 2876
rect 30260 2836 30261 2876
rect 30219 2827 30261 2836
rect 29932 2633 29972 2719
rect 29931 2624 29973 2633
rect 29931 2584 29932 2624
rect 29972 2584 29973 2624
rect 29931 2575 29973 2584
rect 29835 1952 29877 1961
rect 29835 1912 29836 1952
rect 29876 1912 29877 1952
rect 29835 1903 29877 1912
rect 29932 1205 29972 2575
rect 30027 2204 30069 2213
rect 30027 2164 30028 2204
rect 30068 2164 30069 2204
rect 30027 2155 30069 2164
rect 30028 1952 30068 2155
rect 30028 1903 30068 1912
rect 30220 1289 30260 2827
rect 30411 2540 30453 2549
rect 30411 2500 30412 2540
rect 30452 2500 30453 2540
rect 30411 2491 30453 2500
rect 30315 2288 30357 2297
rect 30315 2248 30316 2288
rect 30356 2248 30357 2288
rect 30315 2239 30357 2248
rect 30219 1280 30261 1289
rect 30219 1240 30220 1280
rect 30260 1240 30261 1280
rect 30219 1231 30261 1240
rect 29931 1196 29973 1205
rect 29931 1156 29932 1196
rect 29972 1156 29973 1196
rect 29931 1147 29973 1156
rect 29835 1112 29877 1121
rect 29835 1072 29836 1112
rect 29876 1072 29877 1112
rect 29835 1063 29877 1072
rect 29836 80 29876 1063
rect 29932 449 29972 1147
rect 29931 440 29973 449
rect 29931 400 29932 440
rect 29972 400 30068 440
rect 29931 391 29973 400
rect 30028 80 30068 400
rect 30220 80 30260 1231
rect 30316 1112 30356 2239
rect 30316 617 30356 1072
rect 30315 608 30357 617
rect 30315 568 30316 608
rect 30356 568 30357 608
rect 30315 559 30357 568
rect 30412 80 30452 2491
rect 30508 2129 30548 3424
rect 30700 2540 30740 4339
rect 30796 2885 30836 4684
rect 30988 3464 31028 4936
rect 31276 4817 31316 4936
rect 31275 4808 31317 4817
rect 31275 4768 31276 4808
rect 31316 4768 31317 4808
rect 31275 4759 31317 4768
rect 31275 4388 31317 4397
rect 31275 4348 31276 4388
rect 31316 4348 31317 4388
rect 31275 4339 31317 4348
rect 31083 4220 31125 4229
rect 31083 4180 31084 4220
rect 31124 4180 31125 4220
rect 31083 4171 31125 4180
rect 30988 3415 31028 3424
rect 30892 3380 30932 3389
rect 30892 3221 30932 3340
rect 30891 3212 30933 3221
rect 31084 3212 31124 4171
rect 30891 3172 30892 3212
rect 30932 3172 30933 3212
rect 30891 3163 30933 3172
rect 30988 3172 31124 3212
rect 30795 2876 30837 2885
rect 30795 2836 30796 2876
rect 30836 2836 30837 2876
rect 30795 2827 30837 2836
rect 30604 2500 30740 2540
rect 30507 2120 30549 2129
rect 30507 2080 30508 2120
rect 30548 2080 30549 2120
rect 30507 2071 30549 2080
rect 30508 1938 30548 1947
rect 30508 1364 30548 1898
rect 30508 1315 30548 1324
rect 30604 80 30644 2500
rect 30700 2036 30740 2045
rect 30700 1877 30740 1996
rect 30699 1868 30741 1877
rect 30699 1828 30700 1868
rect 30740 1828 30741 1868
rect 30699 1819 30741 1828
rect 30892 1700 30932 1709
rect 30892 1457 30932 1660
rect 30891 1448 30933 1457
rect 30891 1408 30892 1448
rect 30932 1408 30933 1448
rect 30891 1399 30933 1408
rect 30795 1196 30837 1205
rect 30795 1156 30796 1196
rect 30836 1156 30837 1196
rect 30795 1147 30837 1156
rect 30699 1112 30741 1121
rect 30699 1072 30700 1112
rect 30740 1072 30741 1112
rect 30699 1063 30741 1072
rect 30700 978 30740 1063
rect 30796 80 30836 1147
rect 30988 80 31028 3172
rect 31276 3053 31316 4339
rect 31372 3464 31412 5431
rect 31467 4388 31509 4397
rect 31467 4348 31468 4388
rect 31508 4348 31509 4388
rect 31467 4339 31509 4348
rect 31468 4136 31508 4339
rect 31468 4087 31508 4096
rect 31564 3641 31604 6103
rect 31660 5900 31700 7036
rect 31756 7027 31796 7036
rect 31947 6992 31989 7001
rect 31947 6952 31948 6992
rect 31988 6952 31989 6992
rect 31947 6943 31989 6952
rect 31851 6908 31893 6917
rect 31851 6868 31852 6908
rect 31892 6868 31893 6908
rect 31851 6859 31893 6868
rect 31755 6488 31797 6497
rect 31755 6448 31756 6488
rect 31796 6448 31797 6488
rect 31755 6439 31797 6448
rect 31660 5851 31700 5860
rect 31756 5732 31796 6439
rect 31852 6077 31892 6859
rect 31948 6858 31988 6943
rect 31948 6581 31988 6612
rect 31947 6572 31989 6581
rect 31947 6532 31948 6572
rect 31988 6532 31989 6572
rect 31947 6523 31989 6532
rect 31948 6488 31988 6523
rect 31948 6413 31988 6448
rect 31947 6404 31989 6413
rect 31947 6364 31948 6404
rect 31988 6364 31989 6404
rect 31947 6355 31989 6364
rect 31851 6068 31893 6077
rect 31851 6028 31852 6068
rect 31892 6028 31893 6068
rect 31851 6019 31893 6028
rect 31947 5984 31989 5993
rect 31947 5944 31948 5984
rect 31988 5944 31989 5984
rect 31947 5935 31989 5944
rect 31660 5692 31796 5732
rect 31852 5732 31892 5741
rect 31563 3632 31605 3641
rect 31563 3592 31564 3632
rect 31604 3592 31605 3632
rect 31563 3583 31605 3592
rect 31468 3464 31508 3473
rect 31372 3424 31468 3464
rect 31468 3415 31508 3424
rect 31275 3044 31317 3053
rect 31275 3004 31276 3044
rect 31316 3004 31317 3044
rect 31275 2995 31317 3004
rect 31179 2960 31221 2969
rect 31179 2920 31180 2960
rect 31220 2920 31221 2960
rect 31179 2911 31221 2920
rect 31563 2960 31605 2969
rect 31563 2920 31564 2960
rect 31604 2920 31605 2960
rect 31563 2911 31605 2920
rect 31180 2717 31220 2911
rect 31371 2876 31413 2885
rect 31371 2836 31372 2876
rect 31412 2836 31413 2876
rect 31371 2827 31413 2836
rect 31372 2742 31412 2827
rect 31179 2708 31221 2717
rect 31179 2668 31180 2708
rect 31220 2668 31221 2708
rect 31179 2659 31221 2668
rect 31180 2624 31220 2659
rect 31180 2573 31220 2584
rect 31275 2624 31317 2633
rect 31275 2584 31276 2624
rect 31316 2584 31317 2624
rect 31275 2575 31317 2584
rect 31564 2624 31604 2911
rect 31083 2456 31125 2465
rect 31083 2416 31084 2456
rect 31124 2416 31125 2456
rect 31083 2407 31125 2416
rect 31084 1868 31124 2407
rect 31276 1868 31316 2575
rect 31564 2549 31604 2584
rect 31563 2540 31605 2549
rect 31563 2500 31564 2540
rect 31604 2500 31605 2540
rect 31563 2491 31605 2500
rect 31564 2460 31604 2491
rect 31660 2129 31700 5692
rect 31755 5564 31797 5573
rect 31755 5524 31756 5564
rect 31796 5524 31797 5564
rect 31755 5515 31797 5524
rect 31659 2120 31701 2129
rect 31659 2080 31660 2120
rect 31700 2080 31701 2120
rect 31659 2071 31701 2080
rect 31467 2036 31509 2045
rect 31467 1996 31468 2036
rect 31508 1996 31509 2036
rect 31467 1987 31509 1996
rect 31084 1819 31124 1828
rect 31180 1828 31316 1868
rect 31468 1868 31508 1987
rect 31756 1868 31796 5515
rect 31852 4229 31892 5692
rect 31851 4220 31893 4229
rect 31851 4180 31852 4220
rect 31892 4180 31893 4220
rect 31851 4171 31893 4180
rect 31948 4052 31988 5935
rect 32044 4388 32084 7531
rect 32139 7244 32181 7253
rect 32139 7204 32140 7244
rect 32180 7204 32181 7244
rect 32139 7195 32181 7204
rect 32140 7110 32180 7195
rect 32236 6488 32276 7708
rect 32332 7412 32372 10387
rect 32907 9512 32949 9521
rect 32907 9472 32908 9512
rect 32948 9472 32949 9512
rect 32907 9463 32949 9472
rect 32428 9428 32468 9437
rect 32428 8849 32468 9388
rect 32908 9378 32948 9463
rect 32427 8840 32469 8849
rect 32427 8800 32428 8840
rect 32468 8800 32469 8840
rect 32427 8791 32469 8800
rect 32811 8672 32853 8681
rect 32811 8632 32812 8672
rect 32852 8632 32853 8672
rect 32811 8623 32853 8632
rect 32812 8538 32852 8623
rect 32427 8084 32469 8093
rect 32427 8044 32428 8084
rect 32468 8044 32469 8084
rect 32427 8035 32469 8044
rect 32428 8000 32468 8035
rect 32428 7949 32468 7960
rect 32811 7916 32853 7925
rect 32811 7876 32812 7916
rect 32852 7876 32853 7916
rect 32811 7867 32853 7876
rect 32715 7748 32757 7757
rect 32715 7708 32716 7748
rect 32756 7708 32757 7748
rect 32715 7699 32757 7708
rect 32332 7363 32372 7372
rect 32524 7244 32564 7253
rect 32564 7204 32660 7244
rect 32524 7195 32564 7204
rect 32428 6488 32468 6497
rect 32236 6448 32428 6488
rect 32428 6439 32468 6448
rect 32523 6488 32565 6497
rect 32523 6448 32524 6488
rect 32564 6448 32565 6488
rect 32523 6439 32565 6448
rect 32524 6354 32564 6439
rect 32140 6236 32180 6245
rect 32180 6196 32372 6236
rect 32140 6187 32180 6196
rect 32139 6068 32181 6077
rect 32139 6028 32140 6068
rect 32180 6028 32181 6068
rect 32139 6019 32181 6028
rect 32140 5153 32180 6019
rect 32332 5648 32372 6196
rect 32332 5599 32372 5608
rect 32428 5648 32468 5657
rect 32139 5144 32181 5153
rect 32139 5104 32140 5144
rect 32180 5104 32181 5144
rect 32139 5095 32181 5104
rect 32428 5069 32468 5608
rect 32427 5060 32469 5069
rect 32427 5020 32428 5060
rect 32468 5020 32469 5060
rect 32427 5011 32469 5020
rect 32524 4976 32564 4987
rect 32524 4901 32564 4936
rect 32523 4892 32565 4901
rect 32523 4852 32524 4892
rect 32564 4852 32565 4892
rect 32523 4843 32565 4852
rect 32331 4724 32373 4733
rect 32331 4684 32332 4724
rect 32372 4684 32373 4724
rect 32331 4675 32373 4684
rect 32044 4348 32276 4388
rect 32044 4220 32084 4229
rect 32084 4180 32180 4220
rect 32044 4171 32084 4180
rect 31948 4012 32084 4052
rect 31851 3968 31893 3977
rect 31851 3928 31852 3968
rect 31892 3928 31893 3968
rect 31851 3919 31893 3928
rect 31852 3834 31892 3919
rect 31851 3632 31893 3641
rect 31851 3592 31852 3632
rect 31892 3592 31893 3632
rect 31851 3583 31893 3592
rect 31180 80 31220 1828
rect 31468 1819 31508 1828
rect 31564 1828 31796 1868
rect 31276 1700 31316 1709
rect 31276 1373 31316 1660
rect 31275 1364 31317 1373
rect 31275 1324 31276 1364
rect 31316 1324 31317 1364
rect 31275 1315 31317 1324
rect 31371 1280 31413 1289
rect 31371 1240 31372 1280
rect 31412 1240 31413 1280
rect 31371 1231 31413 1240
rect 31372 80 31412 1231
rect 31564 80 31604 1828
rect 31755 1700 31797 1709
rect 31755 1660 31756 1700
rect 31796 1660 31797 1700
rect 31755 1651 31797 1660
rect 31756 1566 31796 1651
rect 31659 1532 31701 1541
rect 31659 1492 31660 1532
rect 31700 1492 31701 1532
rect 31659 1483 31701 1492
rect 31660 785 31700 1483
rect 31659 776 31701 785
rect 31659 736 31660 776
rect 31700 736 31701 776
rect 31659 727 31701 736
rect 31755 692 31797 701
rect 31755 652 31756 692
rect 31796 652 31797 692
rect 31755 643 31797 652
rect 31756 80 31796 643
rect 31852 197 31892 3583
rect 31948 3450 31988 3459
rect 31948 2885 31988 3410
rect 31947 2876 31989 2885
rect 31947 2836 31948 2876
rect 31988 2836 31989 2876
rect 31947 2827 31989 2836
rect 31947 1868 31989 1877
rect 31947 1828 31948 1868
rect 31988 1828 31989 1868
rect 31947 1819 31989 1828
rect 31948 1734 31988 1819
rect 31947 1112 31989 1121
rect 31947 1072 31948 1112
rect 31988 1072 31989 1112
rect 31947 1063 31989 1072
rect 31948 978 31988 1063
rect 32044 1037 32084 4012
rect 32140 3632 32180 4180
rect 32236 3632 32276 4348
rect 32332 4155 32372 4675
rect 32332 4106 32372 4115
rect 32428 4136 32468 4145
rect 32428 4052 32468 4096
rect 32332 4012 32468 4052
rect 32332 3893 32372 4012
rect 32620 3968 32660 7204
rect 32716 5573 32756 7699
rect 32812 7589 32852 7867
rect 32811 7580 32853 7589
rect 32811 7540 32812 7580
rect 32852 7540 32853 7580
rect 32811 7531 32853 7540
rect 32812 5732 32852 7531
rect 33195 7496 33237 7505
rect 33195 7456 33196 7496
rect 33236 7456 33237 7496
rect 33195 7447 33237 7456
rect 32907 7160 32949 7169
rect 32907 7120 32908 7160
rect 32948 7120 32949 7160
rect 32907 7111 32949 7120
rect 32908 7026 32948 7111
rect 32908 6404 32948 6413
rect 32908 5816 32948 6364
rect 33004 6404 33044 6413
rect 33004 6245 33044 6364
rect 33099 6320 33141 6329
rect 33099 6280 33100 6320
rect 33140 6280 33141 6320
rect 33099 6271 33141 6280
rect 33003 6236 33045 6245
rect 33003 6196 33004 6236
rect 33044 6196 33045 6236
rect 33003 6187 33045 6196
rect 32908 5776 33044 5816
rect 32812 5683 32852 5692
rect 32908 5648 32948 5657
rect 32715 5564 32757 5573
rect 32715 5524 32716 5564
rect 32756 5524 32757 5564
rect 32715 5515 32757 5524
rect 32811 5060 32853 5069
rect 32811 5020 32812 5060
rect 32852 5020 32853 5060
rect 32811 5011 32853 5020
rect 32715 4724 32757 4733
rect 32715 4684 32716 4724
rect 32756 4684 32757 4724
rect 32715 4675 32757 4684
rect 32716 4590 32756 4675
rect 32812 4136 32852 5011
rect 32908 4313 32948 5608
rect 33004 5069 33044 5776
rect 33003 5060 33045 5069
rect 33003 5020 33004 5060
rect 33044 5020 33045 5060
rect 33003 5011 33045 5020
rect 32907 4304 32949 4313
rect 32907 4264 32908 4304
rect 32948 4264 32949 4304
rect 32907 4255 32949 4264
rect 32908 4220 32948 4255
rect 32908 4169 32948 4180
rect 32812 4061 32852 4096
rect 32811 4052 32853 4061
rect 32428 3928 32660 3968
rect 32716 4012 32812 4052
rect 32852 4012 32853 4052
rect 32331 3884 32373 3893
rect 32331 3844 32332 3884
rect 32372 3844 32373 3884
rect 32331 3835 32373 3844
rect 32332 3632 32372 3641
rect 32236 3592 32332 3632
rect 32140 3583 32180 3592
rect 32332 3583 32372 3592
rect 32331 2120 32373 2129
rect 32331 2080 32332 2120
rect 32372 2080 32373 2120
rect 32331 2071 32373 2080
rect 32236 1952 32276 1961
rect 32139 1868 32181 1877
rect 32139 1828 32140 1868
rect 32180 1828 32181 1868
rect 32139 1819 32181 1828
rect 32140 1541 32180 1819
rect 32139 1532 32181 1541
rect 32139 1492 32140 1532
rect 32180 1492 32181 1532
rect 32139 1483 32181 1492
rect 32140 1364 32180 1373
rect 32236 1364 32276 1912
rect 32332 1952 32372 2071
rect 32332 1903 32372 1912
rect 32428 1457 32468 3928
rect 32619 3800 32661 3809
rect 32619 3760 32620 3800
rect 32660 3760 32661 3800
rect 32619 3751 32661 3760
rect 32524 3380 32564 3389
rect 32427 1448 32469 1457
rect 32427 1408 32428 1448
rect 32468 1408 32469 1448
rect 32427 1399 32469 1408
rect 32180 1324 32276 1364
rect 32140 1315 32180 1324
rect 32524 1280 32564 3340
rect 32236 1240 32564 1280
rect 32043 1028 32085 1037
rect 32043 988 32044 1028
rect 32084 988 32085 1028
rect 32043 979 32085 988
rect 32236 440 32276 1240
rect 32332 1112 32372 1121
rect 32372 1072 32468 1112
rect 32332 1063 32372 1072
rect 32331 776 32373 785
rect 32331 736 32332 776
rect 32372 736 32373 776
rect 32331 727 32373 736
rect 32044 400 32276 440
rect 31851 188 31893 197
rect 32044 188 32084 400
rect 31851 148 31852 188
rect 31892 148 31893 188
rect 31851 139 31893 148
rect 31948 148 32084 188
rect 32139 188 32181 197
rect 32139 148 32140 188
rect 32180 148 32181 188
rect 31948 80 31988 148
rect 32139 139 32181 148
rect 32140 80 32180 139
rect 32332 80 32372 727
rect 32428 449 32468 1072
rect 32523 1028 32565 1037
rect 32523 988 32524 1028
rect 32564 988 32565 1028
rect 32523 979 32565 988
rect 32427 440 32469 449
rect 32427 400 32428 440
rect 32468 400 32469 440
rect 32427 391 32469 400
rect 32524 80 32564 979
rect 32620 944 32660 3751
rect 32716 2876 32756 4012
rect 32811 4003 32853 4012
rect 33003 3464 33045 3473
rect 33003 3424 33004 3464
rect 33044 3424 33045 3464
rect 33003 3415 33045 3424
rect 33004 3330 33044 3415
rect 32716 2836 32948 2876
rect 32811 2708 32853 2717
rect 32811 2668 32812 2708
rect 32852 2668 32853 2708
rect 32811 2659 32853 2668
rect 32812 2624 32852 2659
rect 32812 2573 32852 2584
rect 32908 2372 32948 2836
rect 32716 2332 32948 2372
rect 33004 2624 33044 2633
rect 32716 1952 32756 2332
rect 32716 1903 32756 1912
rect 32811 1952 32853 1961
rect 32811 1912 32812 1952
rect 32852 1912 32853 1952
rect 32811 1903 32853 1912
rect 32812 1818 32852 1903
rect 33004 1709 33044 2584
rect 33003 1700 33045 1709
rect 33003 1660 33004 1700
rect 33044 1660 33045 1700
rect 33003 1651 33045 1660
rect 32907 1364 32949 1373
rect 32907 1324 32908 1364
rect 32948 1324 32949 1364
rect 32907 1315 32949 1324
rect 32620 904 32756 944
rect 32716 80 32756 904
rect 32908 80 32948 1315
rect 33004 1037 33044 1651
rect 33003 1028 33045 1037
rect 33003 988 33004 1028
rect 33044 988 33045 1028
rect 33003 979 33045 988
rect 33100 80 33140 6271
rect 33196 5237 33236 7447
rect 33291 7160 33333 7169
rect 33291 7120 33292 7160
rect 33332 7120 33333 7160
rect 33291 7111 33333 7120
rect 33292 6413 33332 7111
rect 33291 6404 33333 6413
rect 33291 6364 33292 6404
rect 33332 6364 33333 6404
rect 33291 6355 33333 6364
rect 33195 5228 33237 5237
rect 33195 5188 33196 5228
rect 33236 5188 33237 5228
rect 33195 5179 33237 5188
rect 33196 4976 33236 4985
rect 33292 4976 33332 6355
rect 33388 5909 33428 10692
rect 34040 10672 34120 10752
rect 35192 10732 35272 10752
rect 34828 10692 35272 10732
rect 34060 9941 34100 10672
rect 34059 9932 34101 9941
rect 34059 9892 34060 9932
rect 34100 9892 34101 9932
rect 34059 9883 34101 9892
rect 34539 9848 34581 9857
rect 34539 9808 34540 9848
rect 34580 9808 34581 9848
rect 34539 9799 34581 9808
rect 34540 9680 34580 9799
rect 34540 9631 34580 9640
rect 34156 9512 34196 9521
rect 34156 9428 34196 9472
rect 34732 9428 34772 9437
rect 34156 9388 34484 9428
rect 33771 9260 33813 9269
rect 33771 9220 33772 9260
rect 33812 9220 33813 9260
rect 33771 9211 33813 9220
rect 34347 9260 34389 9269
rect 34347 9220 34348 9260
rect 34388 9220 34389 9260
rect 34347 9211 34389 9220
rect 33675 8000 33717 8009
rect 33675 7960 33676 8000
rect 33716 7960 33717 8000
rect 33675 7951 33717 7960
rect 33676 7866 33716 7951
rect 33772 7412 33812 9211
rect 34348 9126 34388 9211
rect 33928 9092 34296 9101
rect 33968 9052 34010 9092
rect 34050 9052 34092 9092
rect 34132 9052 34174 9092
rect 34214 9052 34256 9092
rect 33928 9043 34296 9052
rect 34444 8597 34484 9388
rect 34539 8924 34581 8933
rect 34539 8884 34540 8924
rect 34580 8884 34581 8924
rect 34539 8875 34581 8884
rect 33963 8588 34005 8597
rect 33963 8548 33964 8588
rect 34004 8548 34005 8588
rect 33963 8539 34005 8548
rect 34443 8588 34485 8597
rect 34443 8548 34444 8588
rect 34484 8548 34485 8588
rect 34443 8539 34485 8548
rect 33964 8504 34004 8539
rect 33964 8453 34004 8464
rect 34348 8504 34388 8513
rect 34348 7832 34388 8464
rect 34444 8093 34484 8539
rect 34443 8084 34485 8093
rect 34443 8044 34444 8084
rect 34484 8044 34485 8084
rect 34443 8035 34485 8044
rect 34348 7792 34484 7832
rect 33964 7748 34004 7757
rect 34004 7708 34388 7748
rect 33964 7699 34004 7708
rect 33928 7580 34296 7589
rect 33968 7540 34010 7580
rect 34050 7540 34092 7580
rect 34132 7540 34174 7580
rect 34214 7540 34256 7580
rect 33928 7531 34296 7540
rect 33772 7372 34004 7412
rect 33771 6992 33813 7001
rect 33771 6952 33772 6992
rect 33812 6952 33813 6992
rect 33771 6943 33813 6952
rect 33483 6824 33525 6833
rect 33483 6784 33484 6824
rect 33524 6784 33525 6824
rect 33483 6775 33525 6784
rect 33484 6488 33524 6775
rect 33524 6448 33716 6488
rect 33484 6439 33524 6448
rect 33579 6236 33621 6245
rect 33579 6196 33580 6236
rect 33620 6196 33621 6236
rect 33579 6187 33621 6196
rect 33387 5900 33429 5909
rect 33387 5860 33388 5900
rect 33428 5860 33429 5900
rect 33387 5851 33429 5860
rect 33388 5741 33428 5772
rect 33387 5732 33429 5741
rect 33387 5692 33388 5732
rect 33428 5692 33429 5732
rect 33387 5683 33429 5692
rect 33388 5648 33428 5683
rect 33388 5321 33428 5608
rect 33483 5396 33525 5405
rect 33483 5356 33484 5396
rect 33524 5356 33525 5396
rect 33483 5347 33525 5356
rect 33387 5312 33429 5321
rect 33387 5272 33388 5312
rect 33428 5272 33429 5312
rect 33387 5263 33429 5272
rect 33484 5069 33524 5347
rect 33483 5060 33525 5069
rect 33483 5020 33484 5060
rect 33524 5020 33525 5060
rect 33483 5011 33525 5020
rect 33236 4936 33332 4976
rect 33196 4927 33236 4936
rect 33291 4724 33333 4733
rect 33291 4684 33292 4724
rect 33332 4684 33333 4724
rect 33291 4675 33333 4684
rect 33292 1952 33332 4675
rect 33483 4220 33525 4229
rect 33483 4180 33484 4220
rect 33524 4180 33525 4220
rect 33483 4171 33525 4180
rect 33387 4136 33429 4145
rect 33387 4096 33388 4136
rect 33428 4096 33429 4136
rect 33387 4087 33429 4096
rect 33388 4002 33428 4087
rect 33292 1903 33332 1912
rect 33291 1448 33333 1457
rect 33291 1408 33292 1448
rect 33332 1408 33333 1448
rect 33291 1399 33333 1408
rect 33292 80 33332 1399
rect 33484 80 33524 4171
rect 33580 3221 33620 6187
rect 33676 4733 33716 6448
rect 33772 5900 33812 6943
rect 33964 6483 34004 7372
rect 34348 7253 34388 7708
rect 34347 7244 34389 7253
rect 34252 7204 34348 7244
rect 34388 7204 34389 7244
rect 34156 7160 34196 7169
rect 34060 7120 34156 7160
rect 34060 6581 34100 7120
rect 34156 7111 34196 7120
rect 34252 6749 34292 7204
rect 34347 7195 34389 7204
rect 34444 7085 34484 7792
rect 34540 7160 34580 8875
rect 34732 7757 34772 9388
rect 34731 7748 34773 7757
rect 34731 7708 34732 7748
rect 34772 7708 34773 7748
rect 34731 7699 34773 7708
rect 34540 7111 34580 7120
rect 34443 7076 34485 7085
rect 34443 7036 34444 7076
rect 34484 7036 34485 7076
rect 34443 7027 34485 7036
rect 34347 6992 34389 7001
rect 34347 6952 34348 6992
rect 34388 6952 34389 6992
rect 34347 6943 34389 6952
rect 34348 6858 34388 6943
rect 34444 6917 34484 7027
rect 34443 6908 34485 6917
rect 34443 6868 34444 6908
rect 34484 6868 34485 6908
rect 34443 6859 34485 6868
rect 34251 6740 34293 6749
rect 34251 6700 34252 6740
rect 34292 6700 34293 6740
rect 34251 6691 34293 6700
rect 34539 6656 34581 6665
rect 34539 6616 34540 6656
rect 34580 6616 34581 6656
rect 34539 6607 34581 6616
rect 34059 6572 34101 6581
rect 34059 6532 34060 6572
rect 34100 6532 34101 6572
rect 34059 6523 34101 6532
rect 34156 6572 34196 6581
rect 34196 6532 34388 6572
rect 34156 6523 34196 6532
rect 33964 6434 34004 6443
rect 33928 6068 34296 6077
rect 33968 6028 34010 6068
rect 34050 6028 34092 6068
rect 34132 6028 34174 6068
rect 34214 6028 34256 6068
rect 33928 6019 34296 6028
rect 34251 5900 34293 5909
rect 33772 5860 33908 5900
rect 33868 5662 33908 5860
rect 34251 5860 34252 5900
rect 34292 5860 34293 5900
rect 34251 5851 34293 5860
rect 34252 5766 34292 5851
rect 33868 5613 33908 5622
rect 34251 5564 34293 5573
rect 34251 5524 34252 5564
rect 34292 5524 34293 5564
rect 34251 5515 34293 5524
rect 34060 5480 34100 5489
rect 34060 4733 34100 5440
rect 33675 4724 33717 4733
rect 33675 4684 33676 4724
rect 33716 4684 33717 4724
rect 33675 4675 33717 4684
rect 34059 4724 34101 4733
rect 34059 4684 34060 4724
rect 34100 4684 34101 4724
rect 34252 4724 34292 5515
rect 34348 5405 34388 6532
rect 34444 6488 34484 6497
rect 34444 5900 34484 6448
rect 34540 6488 34580 6607
rect 34540 6439 34580 6448
rect 34444 5860 34676 5900
rect 34444 5732 34484 5741
rect 34347 5396 34389 5405
rect 34347 5356 34348 5396
rect 34388 5356 34389 5396
rect 34347 5347 34389 5356
rect 34444 5321 34484 5692
rect 34443 5312 34485 5321
rect 34443 5272 34444 5312
rect 34484 5272 34485 5312
rect 34443 5263 34485 5272
rect 34636 5060 34676 5860
rect 34731 5648 34773 5657
rect 34731 5608 34732 5648
rect 34772 5608 34773 5648
rect 34731 5599 34773 5608
rect 34732 5514 34772 5599
rect 34731 5396 34773 5405
rect 34731 5356 34732 5396
rect 34772 5356 34773 5396
rect 34731 5347 34773 5356
rect 34732 5060 34772 5347
rect 34828 5144 34868 10692
rect 35164 10672 35272 10692
rect 36344 10672 36424 10752
rect 37496 10672 37576 10752
rect 38648 10672 38728 10752
rect 39800 10672 39880 10752
rect 35164 10648 35252 10672
rect 35168 9848 35536 9857
rect 35208 9808 35250 9848
rect 35290 9808 35332 9848
rect 35372 9808 35414 9848
rect 35454 9808 35496 9848
rect 35168 9799 35536 9808
rect 34924 9512 34964 9521
rect 34924 9353 34964 9472
rect 36172 9512 36212 9521
rect 34923 9344 34965 9353
rect 34923 9304 34924 9344
rect 34964 9304 34965 9344
rect 34923 9295 34965 9304
rect 35883 9260 35925 9269
rect 35883 9220 35884 9260
rect 35924 9220 35925 9260
rect 35883 9211 35925 9220
rect 35500 8672 35540 8681
rect 35540 8632 35636 8672
rect 35500 8623 35540 8632
rect 35168 8336 35536 8345
rect 35208 8296 35250 8336
rect 35290 8296 35332 8336
rect 35372 8296 35414 8336
rect 35454 8296 35496 8336
rect 35168 8287 35536 8296
rect 35596 8009 35636 8632
rect 35115 8000 35157 8009
rect 35115 7960 35116 8000
rect 35156 7960 35157 8000
rect 35115 7951 35157 7960
rect 35595 8000 35637 8009
rect 35595 7960 35596 8000
rect 35636 7960 35637 8000
rect 35595 7951 35637 7960
rect 35116 7866 35156 7951
rect 35499 7748 35541 7757
rect 35499 7708 35500 7748
rect 35540 7708 35541 7748
rect 35499 7699 35541 7708
rect 35500 7160 35540 7699
rect 35691 7244 35733 7253
rect 35691 7204 35692 7244
rect 35732 7204 35733 7244
rect 35691 7195 35733 7204
rect 35500 7111 35540 7120
rect 35595 7076 35637 7085
rect 35595 7036 35596 7076
rect 35636 7036 35637 7076
rect 35595 7027 35637 7036
rect 35019 6992 35061 7001
rect 35019 6952 35020 6992
rect 35060 6952 35061 6992
rect 35019 6943 35061 6952
rect 35020 6858 35060 6943
rect 35168 6824 35536 6833
rect 35208 6784 35250 6824
rect 35290 6784 35332 6824
rect 35372 6784 35414 6824
rect 35454 6784 35496 6824
rect 35168 6775 35536 6784
rect 34923 6488 34965 6497
rect 34923 6448 34924 6488
rect 34964 6448 34965 6488
rect 34923 6439 34965 6448
rect 35499 6488 35541 6497
rect 35596 6488 35636 7027
rect 35499 6448 35500 6488
rect 35540 6448 35636 6488
rect 35499 6439 35541 6448
rect 34924 6354 34964 6439
rect 35020 6404 35060 6413
rect 35020 5573 35060 6364
rect 35500 6354 35540 6439
rect 35692 6404 35732 7195
rect 35884 7160 35924 9211
rect 35980 8000 36020 8009
rect 36020 7960 36116 8000
rect 35980 7951 36020 7960
rect 35884 7111 35924 7120
rect 35979 7160 36021 7169
rect 35979 7120 35980 7160
rect 36020 7120 36021 7160
rect 35979 7111 36021 7120
rect 35980 7026 36020 7111
rect 35787 6992 35829 7001
rect 35787 6952 35788 6992
rect 35828 6952 35829 6992
rect 35787 6943 35829 6952
rect 35596 6364 35732 6404
rect 35019 5564 35061 5573
rect 35019 5524 35020 5564
rect 35060 5524 35061 5564
rect 35019 5515 35061 5524
rect 35168 5312 35536 5321
rect 35208 5272 35250 5312
rect 35290 5272 35332 5312
rect 35372 5272 35414 5312
rect 35454 5272 35496 5312
rect 35168 5263 35536 5272
rect 34828 5104 35252 5144
rect 34732 5020 35060 5060
rect 34636 5011 34676 5020
rect 34444 4976 34484 4987
rect 34444 4901 34484 4936
rect 34443 4892 34485 4901
rect 34443 4852 34444 4892
rect 34484 4852 34485 4892
rect 34443 4843 34485 4852
rect 35020 4892 35060 5020
rect 35020 4843 35060 4852
rect 35212 4808 35252 5104
rect 35307 5060 35349 5069
rect 35307 5020 35308 5060
rect 35348 5020 35349 5060
rect 35307 5011 35349 5020
rect 35212 4759 35252 4768
rect 34828 4724 34868 4733
rect 34252 4684 34388 4724
rect 34059 4675 34101 4684
rect 33928 4556 34296 4565
rect 33968 4516 34010 4556
rect 34050 4516 34092 4556
rect 34132 4516 34174 4556
rect 34214 4516 34256 4556
rect 33928 4507 34296 4516
rect 33868 4141 33908 4150
rect 33868 3641 33908 4101
rect 34059 4052 34101 4061
rect 34059 4012 34060 4052
rect 34100 4012 34101 4052
rect 34059 4003 34101 4012
rect 34060 3918 34100 4003
rect 34251 3968 34293 3977
rect 34251 3928 34252 3968
rect 34292 3928 34293 3968
rect 34251 3919 34293 3928
rect 34252 3834 34292 3919
rect 33867 3632 33909 3641
rect 33867 3592 33868 3632
rect 33908 3592 33909 3632
rect 33867 3583 33909 3592
rect 34251 3548 34293 3557
rect 34251 3508 34252 3548
rect 34292 3508 34293 3548
rect 34251 3499 34293 3508
rect 34252 3464 34292 3499
rect 34252 3413 34292 3424
rect 33675 3296 33717 3305
rect 33675 3256 33676 3296
rect 33716 3256 33717 3296
rect 33675 3247 33717 3256
rect 33579 3212 33621 3221
rect 33579 3172 33580 3212
rect 33620 3172 33621 3212
rect 33579 3163 33621 3172
rect 33580 1961 33620 3163
rect 33579 1952 33621 1961
rect 33579 1912 33580 1952
rect 33620 1912 33621 1952
rect 33579 1903 33621 1912
rect 33676 1373 33716 3247
rect 33928 3044 34296 3053
rect 33968 3004 34010 3044
rect 34050 3004 34092 3044
rect 34132 3004 34174 3044
rect 34214 3004 34256 3044
rect 33928 2995 34296 3004
rect 34252 2624 34292 2633
rect 33771 2456 33813 2465
rect 33771 2416 33772 2456
rect 33812 2416 33813 2456
rect 33771 2407 33813 2416
rect 33772 1947 33812 2407
rect 34252 2297 34292 2584
rect 34251 2288 34293 2297
rect 34251 2248 34252 2288
rect 34292 2248 34293 2288
rect 34251 2239 34293 2248
rect 33963 2204 34005 2213
rect 33963 2164 33964 2204
rect 34004 2164 34005 2204
rect 33963 2155 34005 2164
rect 33964 2120 34004 2155
rect 34348 2120 34388 4684
rect 34540 4684 34828 4724
rect 34444 4220 34484 4229
rect 34444 4061 34484 4180
rect 34443 4052 34485 4061
rect 34443 4012 34444 4052
rect 34484 4012 34485 4052
rect 34443 4003 34485 4012
rect 34443 3632 34485 3641
rect 34443 3592 34444 3632
rect 34484 3592 34485 3632
rect 34443 3583 34485 3592
rect 34444 3498 34484 3583
rect 34444 2549 34484 2634
rect 34443 2540 34485 2549
rect 34443 2500 34444 2540
rect 34484 2500 34485 2540
rect 34443 2491 34485 2500
rect 33964 2069 34004 2080
rect 34252 2080 34388 2120
rect 34443 2120 34485 2129
rect 34443 2080 34444 2120
rect 34484 2080 34485 2120
rect 33772 1898 33812 1907
rect 34252 1709 34292 2080
rect 34443 2071 34485 2080
rect 34348 1952 34388 1961
rect 34251 1700 34293 1709
rect 34251 1660 34252 1700
rect 34292 1660 34293 1700
rect 34251 1651 34293 1660
rect 33928 1532 34296 1541
rect 33968 1492 34010 1532
rect 34050 1492 34092 1532
rect 34132 1492 34174 1532
rect 34214 1492 34256 1532
rect 33928 1483 34296 1492
rect 33675 1364 33717 1373
rect 33675 1324 33676 1364
rect 33716 1324 33717 1364
rect 33675 1315 33717 1324
rect 34348 1289 34388 1912
rect 34444 1952 34484 2071
rect 34444 1903 34484 1912
rect 33771 1280 33813 1289
rect 33771 1240 33772 1280
rect 33812 1240 33813 1280
rect 33771 1231 33813 1240
rect 34347 1280 34389 1289
rect 34347 1240 34348 1280
rect 34388 1240 34389 1280
rect 34347 1231 34389 1240
rect 33772 1146 33812 1231
rect 33579 1112 33621 1121
rect 33579 1072 33580 1112
rect 33620 1072 33621 1112
rect 33579 1063 33621 1072
rect 33963 1112 34005 1121
rect 33963 1072 33964 1112
rect 34004 1072 34005 1112
rect 33963 1063 34005 1072
rect 33580 978 33620 1063
rect 33964 449 34004 1063
rect 34540 533 34580 4684
rect 34828 4675 34868 4684
rect 35019 4724 35061 4733
rect 35019 4684 35020 4724
rect 35060 4684 35061 4724
rect 35308 4724 35348 5011
rect 35404 4892 35444 4901
rect 35444 4852 35540 4892
rect 35404 4843 35444 4852
rect 35308 4684 35444 4724
rect 35019 4675 35061 4684
rect 35020 4220 35060 4675
rect 35020 4171 35060 4180
rect 35308 4136 35348 4145
rect 34828 3968 34868 3977
rect 35308 3968 35348 4096
rect 35404 4136 35444 4684
rect 35404 4087 35444 4096
rect 35500 3977 35540 4852
rect 34732 3928 34828 3968
rect 34635 3632 34677 3641
rect 34635 3592 34636 3632
rect 34676 3592 34677 3632
rect 34635 3583 34677 3592
rect 34636 3498 34676 3583
rect 34635 2288 34677 2297
rect 34635 2248 34636 2288
rect 34676 2248 34677 2288
rect 34635 2239 34677 2248
rect 34636 1289 34676 2239
rect 34732 1877 34772 3928
rect 34828 3919 34868 3928
rect 35020 3928 35348 3968
rect 35499 3968 35541 3977
rect 35499 3928 35500 3968
rect 35540 3928 35541 3968
rect 35020 3641 35060 3928
rect 35499 3919 35541 3928
rect 35168 3800 35536 3809
rect 35208 3760 35250 3800
rect 35290 3760 35332 3800
rect 35372 3760 35414 3800
rect 35454 3760 35496 3800
rect 35168 3751 35536 3760
rect 35019 3632 35061 3641
rect 35596 3632 35636 6364
rect 35691 5480 35733 5489
rect 35691 5440 35692 5480
rect 35732 5440 35733 5480
rect 35691 5431 35733 5440
rect 35692 4808 35732 5431
rect 35788 4976 35828 6943
rect 35883 6908 35925 6917
rect 35883 6868 35884 6908
rect 35924 6868 35925 6908
rect 35883 6859 35925 6868
rect 35884 6320 35924 6859
rect 36076 6665 36116 7960
rect 36172 6833 36212 9472
rect 36364 9437 36404 10672
rect 36555 10604 36597 10613
rect 36555 10564 36556 10604
rect 36596 10564 36597 10604
rect 36555 10555 36597 10564
rect 36556 9680 36596 10555
rect 36939 10520 36981 10529
rect 36939 10480 36940 10520
rect 36980 10480 36981 10520
rect 36939 10471 36981 10480
rect 36556 9631 36596 9640
rect 36940 9680 36980 10471
rect 36940 9631 36980 9640
rect 37323 9680 37365 9689
rect 37323 9640 37324 9680
rect 37364 9640 37365 9680
rect 37323 9631 37365 9640
rect 37324 9546 37364 9631
rect 37516 9596 37556 10672
rect 38668 9689 38708 10672
rect 39820 10016 39860 10672
rect 40971 10520 41013 10529
rect 40971 10480 40972 10520
rect 41012 10480 41013 10520
rect 40971 10471 41013 10480
rect 40683 10184 40725 10193
rect 40683 10144 40684 10184
rect 40724 10144 40725 10184
rect 40683 10135 40725 10144
rect 39820 9976 40148 10016
rect 39339 9932 39381 9941
rect 39339 9892 39340 9932
rect 39380 9892 39381 9932
rect 39339 9883 39381 9892
rect 38667 9680 38709 9689
rect 38667 9640 38668 9680
rect 38708 9640 38709 9680
rect 38667 9631 38709 9640
rect 39340 9680 39380 9883
rect 39340 9631 39380 9640
rect 39723 9680 39765 9689
rect 39723 9640 39724 9680
rect 39764 9640 39765 9680
rect 39723 9631 39765 9640
rect 40108 9680 40148 9976
rect 40108 9631 40148 9640
rect 40684 9680 40724 10135
rect 40875 9764 40917 9773
rect 40875 9724 40876 9764
rect 40916 9724 40917 9764
rect 40875 9715 40917 9724
rect 40684 9631 40724 9640
rect 37516 9556 37652 9596
rect 36363 9428 36405 9437
rect 36363 9388 36364 9428
rect 36404 9388 36405 9428
rect 36363 9379 36405 9388
rect 36748 9428 36788 9437
rect 36363 9260 36405 9269
rect 36363 9220 36364 9260
rect 36404 9220 36405 9260
rect 36363 9211 36405 9220
rect 36364 9126 36404 9211
rect 36748 8924 36788 9388
rect 37132 9428 37172 9437
rect 37132 9101 37172 9388
rect 37516 9428 37556 9437
rect 37131 9092 37173 9101
rect 37131 9052 37132 9092
rect 37172 9052 37173 9092
rect 37131 9043 37173 9052
rect 36748 8884 37076 8924
rect 36651 8756 36693 8765
rect 36651 8716 36652 8756
rect 36692 8716 36693 8756
rect 36651 8707 36693 8716
rect 36364 8672 36404 8681
rect 36364 8177 36404 8632
rect 36555 8420 36597 8429
rect 36555 8380 36556 8420
rect 36596 8380 36597 8420
rect 36555 8371 36597 8380
rect 36363 8168 36405 8177
rect 36363 8128 36364 8168
rect 36404 8128 36405 8168
rect 36363 8119 36405 8128
rect 36267 8000 36309 8009
rect 36267 7960 36268 8000
rect 36308 7960 36309 8000
rect 36267 7951 36309 7960
rect 36364 8000 36404 8011
rect 36171 6824 36213 6833
rect 36171 6784 36172 6824
rect 36212 6784 36213 6824
rect 36171 6775 36213 6784
rect 36075 6656 36117 6665
rect 36075 6616 36076 6656
rect 36116 6616 36117 6656
rect 36075 6607 36117 6616
rect 36172 6581 36212 6666
rect 36171 6572 36213 6581
rect 36171 6532 36172 6572
rect 36212 6532 36213 6572
rect 36171 6523 36213 6532
rect 36028 6478 36068 6487
rect 36068 6438 36212 6478
rect 36028 6429 36068 6438
rect 35884 6280 36116 6320
rect 35883 5648 35925 5657
rect 35883 5608 35884 5648
rect 35924 5608 35925 5648
rect 35883 5599 35925 5608
rect 35980 5648 36020 5657
rect 35788 4927 35828 4936
rect 35692 4768 35828 4808
rect 35691 4220 35733 4229
rect 35691 4180 35692 4220
rect 35732 4180 35733 4220
rect 35691 4171 35733 4180
rect 35788 4220 35828 4768
rect 35788 4171 35828 4180
rect 35884 4220 35924 5599
rect 35884 4171 35924 4180
rect 35692 3977 35732 4171
rect 35691 3968 35733 3977
rect 35691 3928 35692 3968
rect 35732 3928 35733 3968
rect 35691 3919 35733 3928
rect 35691 3800 35733 3809
rect 35691 3760 35692 3800
rect 35732 3760 35733 3800
rect 35691 3751 35733 3760
rect 35019 3592 35020 3632
rect 35060 3592 35061 3632
rect 35019 3583 35061 3592
rect 35212 3592 35636 3632
rect 34827 3548 34869 3557
rect 34827 3508 34828 3548
rect 34868 3508 34869 3548
rect 34827 3499 34869 3508
rect 34828 3464 34868 3499
rect 34828 3413 34868 3424
rect 34924 2624 34964 2633
rect 34924 2381 34964 2584
rect 35212 2540 35252 3592
rect 35020 2500 35252 2540
rect 34923 2372 34965 2381
rect 34923 2332 34924 2372
rect 34964 2332 34965 2372
rect 34923 2323 34965 2332
rect 34924 1952 34964 1961
rect 35020 1952 35060 2500
rect 35168 2288 35536 2297
rect 35208 2248 35250 2288
rect 35290 2248 35332 2288
rect 35372 2248 35414 2288
rect 35454 2248 35496 2288
rect 35168 2239 35536 2248
rect 34964 1912 35060 1952
rect 35404 1952 35444 1961
rect 35692 1952 35732 3751
rect 35883 3464 35925 3473
rect 35980 3464 36020 5608
rect 36076 3809 36116 6280
rect 36172 5900 36212 6438
rect 36172 5851 36212 5860
rect 36268 5144 36308 7951
rect 36364 7925 36404 7960
rect 36363 7916 36405 7925
rect 36363 7876 36364 7916
rect 36404 7876 36405 7916
rect 36363 7867 36405 7876
rect 36459 7244 36501 7253
rect 36459 7204 36460 7244
rect 36500 7204 36501 7244
rect 36459 7195 36501 7204
rect 36364 7160 36404 7171
rect 36364 7085 36404 7120
rect 36460 7110 36500 7195
rect 36363 7076 36405 7085
rect 36363 7036 36364 7076
rect 36404 7036 36405 7076
rect 36363 7027 36405 7036
rect 36363 6656 36405 6665
rect 36363 6616 36364 6656
rect 36404 6616 36405 6656
rect 36363 6607 36405 6616
rect 36364 6320 36404 6607
rect 36459 6572 36501 6581
rect 36459 6532 36460 6572
rect 36500 6532 36501 6572
rect 36459 6523 36501 6532
rect 36364 6271 36404 6280
rect 36460 5732 36500 6523
rect 36556 5900 36596 8371
rect 36652 8000 36692 8707
rect 36748 8588 36788 8597
rect 36748 8429 36788 8548
rect 36940 8504 36980 8513
rect 36747 8420 36789 8429
rect 36747 8380 36748 8420
rect 36788 8380 36789 8420
rect 36747 8371 36789 8380
rect 36747 8168 36789 8177
rect 36747 8128 36748 8168
rect 36788 8128 36789 8168
rect 36747 8119 36789 8128
rect 36652 7951 36692 7960
rect 36651 6740 36693 6749
rect 36651 6700 36652 6740
rect 36692 6700 36693 6740
rect 36651 6691 36693 6700
rect 36652 6068 36692 6691
rect 36748 6320 36788 8119
rect 36940 8093 36980 8464
rect 36939 8084 36981 8093
rect 36939 8044 36940 8084
rect 36980 8044 36981 8084
rect 36939 8035 36981 8044
rect 36939 7748 36981 7757
rect 36939 7708 36940 7748
rect 36980 7708 36981 7748
rect 36939 7699 36981 7708
rect 36940 7614 36980 7699
rect 36843 7244 36885 7253
rect 36843 7204 36844 7244
rect 36884 7204 36885 7244
rect 36843 7195 36885 7204
rect 36748 6271 36788 6280
rect 36652 6028 36788 6068
rect 36651 5900 36693 5909
rect 36556 5860 36652 5900
rect 36692 5860 36693 5900
rect 36651 5851 36693 5860
rect 36652 5741 36692 5851
rect 36556 5732 36596 5741
rect 36460 5692 36556 5732
rect 36556 5683 36596 5692
rect 36651 5732 36693 5741
rect 36651 5692 36652 5732
rect 36692 5692 36693 5732
rect 36651 5683 36693 5692
rect 36363 5480 36405 5489
rect 36363 5440 36364 5480
rect 36404 5440 36405 5480
rect 36363 5431 36405 5440
rect 36364 5346 36404 5431
rect 36268 5095 36308 5104
rect 36748 4901 36788 6028
rect 36747 4892 36789 4901
rect 36747 4852 36748 4892
rect 36788 4852 36789 4892
rect 36747 4843 36789 4852
rect 36844 4304 36884 7195
rect 36940 7160 36980 7169
rect 36940 6917 36980 7120
rect 36939 6908 36981 6917
rect 36939 6868 36940 6908
rect 36980 6868 36981 6908
rect 36939 6859 36981 6868
rect 37036 5648 37076 8884
rect 37132 8672 37172 8681
rect 37132 8504 37172 8632
rect 37132 8464 37182 8504
rect 37142 8420 37182 8464
rect 37132 8380 37182 8420
rect 37132 6749 37172 8380
rect 37419 8084 37461 8093
rect 37419 8044 37420 8084
rect 37460 8044 37461 8084
rect 37419 8035 37461 8044
rect 37420 7174 37460 8035
rect 37516 7253 37556 9388
rect 37612 7916 37652 9556
rect 39724 9546 39764 9631
rect 37708 9512 37748 9521
rect 37708 9353 37748 9472
rect 38956 9512 38996 9521
rect 38187 9428 38229 9437
rect 38187 9388 38188 9428
rect 38228 9388 38229 9428
rect 38187 9379 38229 9388
rect 37707 9344 37749 9353
rect 37707 9304 37708 9344
rect 37748 9304 37749 9344
rect 37707 9295 37749 9304
rect 37708 8000 37748 9295
rect 38188 8168 38228 9379
rect 38764 8756 38804 8765
rect 38476 8716 38764 8756
rect 38379 8672 38421 8681
rect 38379 8632 38380 8672
rect 38420 8632 38421 8672
rect 38379 8623 38421 8632
rect 38380 8538 38420 8623
rect 38188 8119 38228 8128
rect 38091 8000 38133 8009
rect 37708 7960 37940 8000
rect 37612 7876 37748 7916
rect 37708 7496 37748 7876
rect 37804 7832 37844 7841
rect 37804 7673 37844 7792
rect 37803 7664 37845 7673
rect 37803 7624 37804 7664
rect 37844 7624 37845 7664
rect 37803 7615 37845 7624
rect 37708 7456 37844 7496
rect 37804 7412 37844 7456
rect 37804 7363 37844 7372
rect 37707 7328 37749 7337
rect 37707 7288 37708 7328
rect 37748 7288 37749 7328
rect 37707 7279 37749 7288
rect 37515 7244 37557 7253
rect 37515 7204 37516 7244
rect 37556 7204 37557 7244
rect 37515 7195 37557 7204
rect 37420 7125 37460 7134
rect 37612 6992 37652 7001
rect 37228 6952 37612 6992
rect 37131 6740 37173 6749
rect 37131 6700 37132 6740
rect 37172 6700 37173 6740
rect 37131 6691 37173 6700
rect 37228 5732 37268 6952
rect 37612 6943 37652 6952
rect 37708 6917 37748 7279
rect 37707 6908 37749 6917
rect 37707 6868 37708 6908
rect 37748 6868 37749 6908
rect 37707 6859 37749 6868
rect 37323 6824 37365 6833
rect 37323 6784 37324 6824
rect 37364 6784 37365 6824
rect 37323 6775 37365 6784
rect 37324 6488 37364 6775
rect 37324 6439 37364 6448
rect 37900 6320 37940 7960
rect 38091 7960 38092 8000
rect 38132 7960 38133 8000
rect 38091 7951 38133 7960
rect 37996 7244 38036 7253
rect 37996 6413 38036 7204
rect 37995 6404 38037 6413
rect 37995 6364 37996 6404
rect 38036 6364 38037 6404
rect 37995 6355 38037 6364
rect 37804 6280 37940 6320
rect 37611 6068 37653 6077
rect 37611 6028 37612 6068
rect 37652 6028 37653 6068
rect 37611 6019 37653 6028
rect 37228 5683 37268 5692
rect 37516 5648 37556 5657
rect 37036 5608 37172 5648
rect 37035 5480 37077 5489
rect 37035 5440 37036 5480
rect 37076 5440 37077 5480
rect 37035 5431 37077 5440
rect 37036 5346 37076 5431
rect 37132 5228 37172 5608
rect 37036 5188 37172 5228
rect 36939 5060 36981 5069
rect 36939 5020 36940 5060
rect 36980 5020 36981 5060
rect 36939 5011 36981 5020
rect 36940 4926 36980 5011
rect 37036 4388 37076 5188
rect 37516 5069 37556 5608
rect 37612 5648 37652 6019
rect 37804 5741 37844 6280
rect 37803 5732 37845 5741
rect 37803 5692 37804 5732
rect 37844 5692 37845 5732
rect 37803 5683 37845 5692
rect 37612 5573 37652 5608
rect 37995 5648 38037 5657
rect 37995 5608 37996 5648
rect 38036 5608 38037 5648
rect 37995 5599 38037 5608
rect 38092 5648 38132 7951
rect 38380 7916 38420 7925
rect 37611 5564 37653 5573
rect 37611 5524 37612 5564
rect 37652 5524 37653 5564
rect 37611 5515 37653 5524
rect 37612 5153 37652 5515
rect 37996 5514 38036 5599
rect 37611 5144 37653 5153
rect 37611 5104 37612 5144
rect 37652 5104 37653 5144
rect 37611 5095 37653 5104
rect 37515 5060 37557 5069
rect 37515 5020 37516 5060
rect 37556 5020 37557 5060
rect 37515 5011 37557 5020
rect 37132 4976 37172 4987
rect 37132 4901 37172 4936
rect 37227 4976 37269 4985
rect 37227 4936 37228 4976
rect 37268 4936 37269 4976
rect 37227 4927 37269 4936
rect 37131 4892 37173 4901
rect 37131 4852 37132 4892
rect 37172 4852 37173 4892
rect 37131 4843 37173 4852
rect 37228 4388 37268 4927
rect 37611 4892 37653 4901
rect 37611 4852 37612 4892
rect 37652 4852 37653 4892
rect 37611 4843 37653 4852
rect 37803 4892 37845 4901
rect 37803 4852 37804 4892
rect 37844 4852 37845 4892
rect 37803 4843 37845 4852
rect 37036 4348 37172 4388
rect 36844 4264 36980 4304
rect 36364 4136 36404 4145
rect 36172 4096 36364 4136
rect 36075 3800 36117 3809
rect 36075 3760 36076 3800
rect 36116 3760 36117 3800
rect 36075 3751 36117 3760
rect 36076 3473 36116 3558
rect 35883 3424 35884 3464
rect 35924 3424 36020 3464
rect 35883 3415 35925 3424
rect 35980 2708 36020 3424
rect 36075 3464 36117 3473
rect 36075 3424 36076 3464
rect 36116 3424 36117 3464
rect 36075 3415 36117 3424
rect 36172 3296 36212 4096
rect 36364 4087 36404 4096
rect 36844 4141 36884 4150
rect 36844 3884 36884 4101
rect 36556 3844 36884 3884
rect 36460 3380 36500 3389
rect 36076 3256 36212 3296
rect 36364 3340 36460 3380
rect 36076 2885 36116 3256
rect 36268 3212 36308 3221
rect 36172 3172 36268 3212
rect 36075 2876 36117 2885
rect 36075 2836 36076 2876
rect 36116 2836 36117 2876
rect 36075 2827 36117 2836
rect 36172 2801 36212 3172
rect 36268 3163 36308 3172
rect 36364 2960 36404 3340
rect 36460 3331 36500 3340
rect 36556 3212 36596 3844
rect 36940 3800 36980 4264
rect 37035 4220 37077 4229
rect 37035 4180 37036 4220
rect 37076 4180 37077 4220
rect 37035 4171 37077 4180
rect 37036 4052 37076 4171
rect 37036 4003 37076 4012
rect 36268 2920 36404 2960
rect 36460 3172 36596 3212
rect 36652 3760 36980 3800
rect 36171 2792 36213 2801
rect 36171 2752 36172 2792
rect 36212 2752 36213 2792
rect 36171 2743 36213 2752
rect 35980 2668 36116 2708
rect 36076 2624 36116 2668
rect 36172 2624 36212 2633
rect 36076 2584 36172 2624
rect 36172 2575 36212 2584
rect 36268 2288 36308 2920
rect 36364 2792 36404 2801
rect 36460 2792 36500 3172
rect 36404 2752 36500 2792
rect 36364 2743 36404 2752
rect 36555 2708 36597 2717
rect 36555 2668 36556 2708
rect 36596 2668 36597 2708
rect 36555 2659 36597 2668
rect 36556 2624 36596 2659
rect 36556 2573 36596 2584
rect 36076 2248 36308 2288
rect 36076 2120 36116 2248
rect 36076 2071 36116 2080
rect 36459 2036 36501 2045
rect 36459 1996 36460 2036
rect 36500 1996 36501 2036
rect 36459 1987 36501 1996
rect 35444 1912 35732 1952
rect 35884 1938 35924 1947
rect 34924 1903 34964 1912
rect 35404 1903 35444 1912
rect 34731 1868 34773 1877
rect 34731 1828 34732 1868
rect 34772 1828 34773 1868
rect 34731 1819 34773 1828
rect 34828 1868 34868 1877
rect 34828 1709 34868 1828
rect 34827 1700 34869 1709
rect 34827 1660 34828 1700
rect 34868 1660 34869 1700
rect 34827 1651 34869 1660
rect 35884 1532 35924 1898
rect 36460 1868 36500 1987
rect 36460 1819 36500 1828
rect 36555 1868 36597 1877
rect 36555 1828 36556 1868
rect 36596 1828 36597 1868
rect 36555 1819 36597 1828
rect 35404 1492 35924 1532
rect 36268 1700 36308 1709
rect 35211 1364 35253 1373
rect 35211 1324 35212 1364
rect 35252 1324 35253 1364
rect 35211 1315 35253 1324
rect 35404 1364 35444 1492
rect 35404 1315 35444 1324
rect 34635 1280 34677 1289
rect 34635 1240 34636 1280
rect 34676 1240 34677 1280
rect 34635 1231 34677 1240
rect 34636 1121 34676 1231
rect 35212 1121 35252 1315
rect 35595 1280 35637 1289
rect 35595 1240 35596 1280
rect 35636 1240 35637 1280
rect 35595 1231 35637 1240
rect 35596 1121 35636 1231
rect 34635 1112 34677 1121
rect 34635 1072 34636 1112
rect 34676 1072 34677 1112
rect 34635 1063 34677 1072
rect 35211 1112 35253 1121
rect 35211 1072 35212 1112
rect 35252 1072 35253 1112
rect 35211 1063 35253 1072
rect 35595 1112 35637 1121
rect 35595 1072 35596 1112
rect 35636 1072 35637 1112
rect 35595 1063 35637 1072
rect 35212 978 35252 1063
rect 35596 978 35636 1063
rect 36268 953 36308 1660
rect 36556 1205 36596 1819
rect 36555 1196 36597 1205
rect 36555 1156 36556 1196
rect 36596 1156 36597 1196
rect 36555 1147 36597 1156
rect 36267 944 36309 953
rect 36267 904 36268 944
rect 36308 904 36309 944
rect 36267 895 36309 904
rect 35168 776 35536 785
rect 35208 736 35250 776
rect 35290 736 35332 776
rect 35372 736 35414 776
rect 35454 736 35496 776
rect 35168 727 35536 736
rect 36652 701 36692 3760
rect 37132 3548 37172 4348
rect 37228 4339 37268 4348
rect 37420 4220 37460 4229
rect 37036 3508 37172 3548
rect 37324 4180 37420 4220
rect 36939 3212 36981 3221
rect 36939 3172 36940 3212
rect 36980 3172 36981 3212
rect 36939 3163 36981 3172
rect 36940 3078 36980 3163
rect 37036 2633 37076 3508
rect 37132 3380 37172 3389
rect 37035 2624 37077 2633
rect 37035 2584 37036 2624
rect 37076 2584 37077 2624
rect 37035 2575 37077 2584
rect 37132 2129 37172 3340
rect 37324 2213 37364 4180
rect 37420 4171 37460 4180
rect 37420 3464 37460 3473
rect 37420 2885 37460 3424
rect 37516 3464 37556 3475
rect 37516 3389 37556 3424
rect 37515 3380 37557 3389
rect 37515 3340 37516 3380
rect 37556 3340 37557 3380
rect 37515 3331 37557 3340
rect 37419 2876 37461 2885
rect 37419 2836 37420 2876
rect 37460 2836 37461 2876
rect 37419 2827 37461 2836
rect 37516 2801 37556 3331
rect 37515 2792 37557 2801
rect 37515 2752 37516 2792
rect 37556 2752 37557 2792
rect 37515 2743 37557 2752
rect 37612 2540 37652 4843
rect 37804 4136 37844 4843
rect 38092 4472 38132 5608
rect 37804 4061 37844 4096
rect 37900 4432 38132 4472
rect 38284 7876 38380 7916
rect 37803 4052 37845 4061
rect 37803 4012 37804 4052
rect 37844 4012 37845 4052
rect 37803 4003 37845 4012
rect 37804 3972 37844 4003
rect 37707 3380 37749 3389
rect 37707 3340 37708 3380
rect 37748 3340 37749 3380
rect 37707 3331 37749 3340
rect 37900 3380 37940 4432
rect 37995 4136 38037 4145
rect 37995 4096 37996 4136
rect 38036 4096 38037 4136
rect 37995 4087 38037 4096
rect 37996 3464 38036 4087
rect 37996 3415 38036 3424
rect 37708 2717 37748 3331
rect 37707 2708 37749 2717
rect 37707 2668 37708 2708
rect 37748 2668 37749 2708
rect 37707 2659 37749 2668
rect 37803 2624 37845 2633
rect 37780 2584 37804 2624
rect 37844 2584 37845 2624
rect 37780 2575 37845 2584
rect 37780 2540 37844 2575
rect 37420 2500 37844 2540
rect 37323 2204 37365 2213
rect 37323 2164 37324 2204
rect 37364 2164 37365 2204
rect 37323 2155 37365 2164
rect 37131 2120 37173 2129
rect 37131 2080 37132 2120
rect 37172 2080 37173 2120
rect 37131 2071 37173 2080
rect 37323 2036 37365 2045
rect 37323 1996 37324 2036
rect 37364 1996 37365 2036
rect 37323 1987 37365 1996
rect 36748 1952 36788 1961
rect 36748 1364 36788 1912
rect 36843 1952 36885 1961
rect 36843 1912 36844 1952
rect 36884 1912 36885 1952
rect 36843 1903 36885 1912
rect 37227 1952 37269 1961
rect 37227 1912 37228 1952
rect 37268 1912 37269 1952
rect 37227 1903 37269 1912
rect 37324 1952 37364 1987
rect 36844 1818 36884 1903
rect 37228 1818 37268 1903
rect 37324 1901 37364 1912
rect 37036 1364 37076 1373
rect 36748 1324 37036 1364
rect 37036 1315 37076 1324
rect 36747 1196 36789 1205
rect 36747 1156 36748 1196
rect 36788 1156 36789 1196
rect 36747 1147 36789 1156
rect 36748 1037 36788 1147
rect 36844 1112 36884 1121
rect 36747 1028 36789 1037
rect 36747 988 36748 1028
rect 36788 988 36789 1028
rect 36747 979 36789 988
rect 36844 869 36884 1072
rect 37228 1112 37268 1121
rect 37420 1112 37460 2500
rect 37804 2490 37844 2500
rect 37803 2288 37845 2297
rect 37803 2248 37804 2288
rect 37844 2248 37845 2288
rect 37803 2239 37845 2248
rect 37804 1952 37844 2239
rect 37900 1961 37940 3340
rect 38284 3305 38324 7876
rect 38380 7867 38420 7876
rect 38379 7160 38421 7169
rect 38379 7120 38380 7160
rect 38420 7120 38421 7160
rect 38379 7111 38421 7120
rect 38380 6077 38420 7111
rect 38476 6161 38516 8716
rect 38764 8707 38804 8716
rect 38956 8597 38996 9472
rect 39532 9428 39572 9437
rect 39148 9260 39188 9269
rect 39052 9220 39148 9260
rect 38955 8588 38997 8597
rect 38955 8548 38956 8588
rect 38996 8548 38997 8588
rect 38955 8539 38997 8548
rect 38572 8504 38612 8513
rect 38572 7841 38612 8464
rect 38763 8420 38805 8429
rect 38763 8380 38764 8420
rect 38804 8380 38805 8420
rect 38763 8371 38805 8380
rect 38764 8000 38804 8371
rect 38764 7951 38804 7960
rect 38860 8000 38900 8009
rect 38571 7832 38613 7841
rect 38571 7792 38572 7832
rect 38612 7792 38613 7832
rect 38571 7783 38613 7792
rect 38572 7160 38612 7169
rect 38572 6656 38612 7120
rect 38667 7160 38709 7169
rect 38860 7160 38900 7960
rect 38956 7589 38996 8539
rect 39052 8429 39092 9220
rect 39148 9211 39188 9220
rect 39147 8672 39189 8681
rect 39147 8632 39148 8672
rect 39188 8632 39189 8672
rect 39147 8623 39189 8632
rect 39051 8420 39093 8429
rect 39051 8380 39052 8420
rect 39092 8380 39093 8420
rect 39051 8371 39093 8380
rect 39148 7757 39188 8623
rect 39244 7916 39284 7925
rect 39147 7748 39189 7757
rect 39147 7708 39148 7748
rect 39188 7708 39189 7748
rect 39147 7699 39189 7708
rect 38955 7580 38997 7589
rect 38955 7540 38956 7580
rect 38996 7540 38997 7580
rect 38955 7531 38997 7540
rect 38667 7120 38668 7160
rect 38708 7120 38900 7160
rect 38667 7111 38709 7120
rect 38668 7026 38708 7111
rect 38764 6656 38804 6665
rect 38572 6616 38764 6656
rect 38764 6607 38804 6616
rect 38956 6572 38996 7531
rect 39244 7253 39284 7876
rect 39340 7916 39380 7925
rect 39051 7244 39093 7253
rect 39051 7204 39052 7244
rect 39092 7204 39093 7244
rect 39051 7195 39093 7204
rect 39243 7244 39285 7253
rect 39243 7204 39244 7244
rect 39284 7204 39285 7244
rect 39243 7195 39285 7204
rect 39052 7110 39092 7195
rect 39147 7160 39189 7169
rect 39147 7120 39148 7160
rect 39188 7120 39189 7160
rect 39147 7111 39189 7120
rect 39148 7026 39188 7111
rect 39147 6908 39189 6917
rect 39147 6868 39148 6908
rect 39188 6868 39189 6908
rect 39147 6859 39189 6868
rect 38860 6532 38996 6572
rect 38572 6488 38612 6497
rect 38860 6488 38900 6532
rect 38612 6448 38900 6488
rect 39148 6488 39188 6859
rect 38572 6439 38612 6448
rect 39148 6439 39188 6448
rect 39244 6320 39284 7195
rect 39340 7169 39380 7876
rect 39339 7160 39381 7169
rect 39339 7120 39340 7160
rect 39380 7120 39381 7160
rect 39339 7111 39381 7120
rect 39244 6280 39380 6320
rect 38475 6152 38517 6161
rect 38475 6112 38476 6152
rect 38516 6112 38517 6152
rect 38475 6103 38517 6112
rect 38379 6068 38421 6077
rect 38379 6028 38380 6068
rect 38420 6028 38421 6068
rect 38379 6019 38421 6028
rect 38571 5900 38613 5909
rect 38571 5860 38572 5900
rect 38612 5860 38613 5900
rect 38571 5851 38613 5860
rect 38572 5648 38612 5851
rect 38476 5608 38572 5648
rect 39100 5657 39140 5666
rect 39140 5617 39188 5648
rect 39100 5608 39188 5617
rect 38380 4976 38420 4985
rect 38380 4817 38420 4936
rect 38379 4808 38421 4817
rect 38379 4768 38380 4808
rect 38420 4768 38421 4808
rect 38379 4759 38421 4768
rect 38476 3464 38516 5608
rect 38572 5599 38612 5608
rect 38859 5144 38901 5153
rect 38859 5104 38860 5144
rect 38900 5104 38901 5144
rect 38859 5095 38901 5104
rect 38763 5060 38805 5069
rect 38763 5020 38764 5060
rect 38804 5020 38805 5060
rect 38763 5011 38805 5020
rect 38764 4976 38804 5011
rect 38764 4925 38804 4936
rect 38571 4724 38613 4733
rect 38571 4684 38572 4724
rect 38612 4684 38613 4724
rect 38571 4675 38613 4684
rect 38572 4590 38612 4675
rect 38283 3296 38325 3305
rect 38283 3256 38284 3296
rect 38324 3256 38325 3296
rect 38283 3247 38325 3256
rect 37995 2876 38037 2885
rect 37995 2836 37996 2876
rect 38036 2836 38037 2876
rect 37995 2827 38037 2836
rect 37996 2742 38036 2827
rect 38380 2633 38420 2718
rect 38379 2624 38421 2633
rect 38379 2584 38380 2624
rect 38420 2584 38421 2624
rect 38379 2575 38421 2584
rect 38188 2456 38228 2465
rect 38379 2456 38421 2465
rect 38228 2416 38324 2456
rect 38188 2407 38228 2416
rect 37804 1903 37844 1912
rect 37899 1952 37941 1961
rect 37899 1912 37900 1952
rect 37940 1912 37941 1952
rect 37899 1903 37941 1912
rect 38284 1947 38324 2416
rect 38379 2416 38380 2456
rect 38420 2416 38421 2456
rect 38379 2407 38421 2416
rect 38284 1898 38324 1907
rect 38380 1289 38420 2407
rect 38476 2297 38516 3424
rect 38571 2708 38613 2717
rect 38571 2668 38572 2708
rect 38612 2668 38613 2708
rect 38571 2659 38613 2668
rect 38475 2288 38517 2297
rect 38475 2248 38476 2288
rect 38516 2248 38517 2288
rect 38475 2239 38517 2248
rect 38475 2120 38517 2129
rect 38475 2080 38476 2120
rect 38516 2080 38517 2120
rect 38475 2071 38517 2080
rect 38476 1986 38516 2071
rect 38572 1373 38612 2659
rect 38764 1952 38804 1961
rect 38571 1364 38613 1373
rect 38571 1324 38572 1364
rect 38612 1324 38613 1364
rect 38571 1315 38613 1324
rect 38668 1364 38708 1373
rect 38764 1364 38804 1912
rect 38860 1952 38900 5095
rect 39051 5060 39093 5069
rect 39051 5020 39052 5060
rect 39092 5020 39093 5060
rect 39051 5011 39093 5020
rect 38955 4724 38997 4733
rect 38955 4684 38956 4724
rect 38996 4684 38997 4724
rect 38955 4675 38997 4684
rect 38956 3459 38996 4675
rect 39052 4136 39092 5011
rect 39148 4388 39188 5608
rect 39244 5480 39284 5489
rect 39244 4565 39284 5440
rect 39243 4556 39285 4565
rect 39243 4516 39244 4556
rect 39284 4516 39285 4556
rect 39243 4507 39285 4516
rect 39244 4388 39284 4397
rect 39148 4348 39244 4388
rect 39244 4339 39284 4348
rect 39340 4220 39380 6280
rect 39532 5993 39572 9388
rect 39916 9428 39956 9437
rect 40300 9428 40340 9437
rect 39627 8504 39669 8513
rect 39627 8464 39628 8504
rect 39668 8464 39669 8504
rect 39627 8455 39669 8464
rect 39628 7160 39668 8455
rect 39819 8000 39861 8009
rect 39819 7960 39820 8000
rect 39860 7960 39861 8000
rect 39819 7951 39861 7960
rect 39820 7866 39860 7951
rect 39628 7111 39668 7120
rect 39819 7160 39861 7169
rect 39819 7120 39820 7160
rect 39860 7120 39861 7160
rect 39819 7111 39861 7120
rect 39531 5984 39573 5993
rect 39531 5944 39532 5984
rect 39572 5944 39573 5984
rect 39531 5935 39573 5944
rect 39820 5825 39860 7111
rect 39819 5816 39861 5825
rect 39819 5776 39820 5816
rect 39860 5776 39861 5816
rect 39819 5767 39861 5776
rect 39916 5648 39956 9388
rect 39724 5608 39956 5648
rect 40012 9388 40300 9428
rect 39627 4556 39669 4565
rect 39627 4516 39628 4556
rect 39668 4516 39669 4556
rect 39627 4507 39669 4516
rect 39052 4087 39092 4096
rect 39148 4180 39380 4220
rect 39628 4220 39668 4507
rect 39148 3968 39188 4180
rect 39628 4171 39668 4180
rect 39436 3968 39476 3977
rect 38956 3410 38996 3419
rect 39052 3928 39188 3968
rect 39244 3928 39436 3968
rect 38860 1903 38900 1912
rect 39052 1793 39092 3928
rect 39148 3548 39188 3557
rect 39148 2549 39188 3508
rect 39147 2540 39189 2549
rect 39147 2500 39148 2540
rect 39188 2500 39189 2540
rect 39147 2491 39189 2500
rect 39244 2045 39284 3928
rect 39436 3919 39476 3928
rect 39627 3548 39669 3557
rect 39627 3508 39628 3548
rect 39668 3508 39669 3548
rect 39724 3548 39764 5608
rect 39915 5480 39957 5489
rect 39915 5440 39916 5480
rect 39956 5440 39957 5480
rect 39915 5431 39957 5440
rect 39916 5346 39956 5431
rect 40012 5144 40052 9388
rect 40300 9379 40340 9388
rect 40491 9428 40533 9437
rect 40491 9388 40492 9428
rect 40532 9388 40533 9428
rect 40491 9379 40533 9388
rect 40876 9428 40916 9715
rect 40876 9379 40916 9388
rect 40492 9294 40532 9379
rect 40779 8924 40821 8933
rect 40779 8884 40780 8924
rect 40820 8884 40821 8924
rect 40779 8875 40821 8884
rect 40396 8681 40436 8766
rect 40395 8672 40437 8681
rect 40395 8632 40396 8672
rect 40436 8632 40437 8672
rect 40395 8623 40437 8632
rect 40588 8504 40628 8513
rect 40396 8464 40588 8504
rect 40396 8000 40436 8464
rect 40588 8455 40628 8464
rect 40492 8084 40532 8093
rect 40532 8044 40628 8084
rect 40492 8035 40532 8044
rect 40348 7990 40436 8000
rect 40388 7960 40436 7990
rect 40348 7941 40388 7950
rect 40395 7580 40437 7589
rect 40395 7540 40396 7580
rect 40436 7540 40437 7580
rect 40395 7531 40437 7540
rect 40108 7165 40148 7174
rect 40108 6665 40148 7125
rect 40300 6992 40340 7001
rect 40107 6656 40149 6665
rect 40107 6616 40108 6656
rect 40148 6616 40149 6656
rect 40107 6607 40149 6616
rect 40300 6320 40340 6952
rect 40396 6488 40436 7531
rect 40588 7244 40628 8044
rect 40684 7916 40724 7925
rect 40684 7421 40724 7876
rect 40683 7412 40725 7421
rect 40683 7372 40684 7412
rect 40724 7372 40725 7412
rect 40683 7363 40725 7372
rect 40684 7244 40724 7253
rect 40588 7204 40684 7244
rect 40684 7195 40724 7204
rect 40491 6992 40533 7001
rect 40491 6952 40492 6992
rect 40532 6952 40533 6992
rect 40491 6943 40533 6952
rect 40492 6858 40532 6943
rect 40587 6656 40629 6665
rect 40587 6616 40588 6656
rect 40628 6616 40629 6656
rect 40587 6607 40629 6616
rect 40588 6522 40628 6607
rect 40396 6439 40436 6448
rect 40108 6280 40340 6320
rect 40108 5732 40148 6280
rect 40780 5909 40820 8875
rect 40875 8756 40917 8765
rect 40875 8716 40876 8756
rect 40916 8716 40917 8756
rect 40875 8707 40917 8716
rect 40876 8622 40916 8707
rect 40876 8168 40916 8177
rect 40972 8168 41012 10471
rect 41067 9848 41109 9857
rect 41067 9808 41068 9848
rect 41108 9808 41109 9848
rect 41067 9799 41109 9808
rect 41068 9680 41108 9799
rect 41068 9631 41108 9640
rect 41259 9596 41301 9605
rect 41259 9556 41260 9596
rect 41300 9556 41301 9596
rect 41259 9547 41301 9556
rect 41260 9428 41300 9547
rect 41451 9512 41493 9521
rect 41451 9472 41452 9512
rect 41492 9472 41493 9512
rect 41451 9463 41493 9472
rect 41260 9379 41300 9388
rect 41452 9344 41492 9463
rect 41452 9295 41492 9304
rect 41355 9176 41397 9185
rect 41355 9136 41356 9176
rect 41396 9136 41397 9176
rect 41355 9127 41397 9136
rect 41163 9008 41205 9017
rect 41163 8968 41164 9008
rect 41204 8968 41205 9008
rect 41163 8959 41205 8968
rect 41068 8504 41108 8513
rect 41068 8177 41108 8464
rect 40916 8128 41012 8168
rect 41067 8168 41109 8177
rect 41067 8128 41068 8168
rect 41108 8128 41109 8168
rect 40876 8119 40916 8128
rect 41067 8119 41109 8128
rect 41068 7916 41108 7925
rect 41164 7916 41204 8959
rect 41259 8756 41301 8765
rect 41259 8716 41260 8756
rect 41300 8716 41301 8756
rect 41259 8707 41301 8716
rect 41260 8622 41300 8707
rect 41108 7876 41204 7916
rect 41068 7867 41108 7876
rect 41163 7748 41205 7757
rect 41163 7708 41164 7748
rect 41204 7708 41205 7748
rect 41163 7699 41205 7708
rect 41260 7748 41300 7757
rect 40971 7412 41013 7421
rect 40971 7372 40972 7412
rect 41012 7372 41013 7412
rect 40971 7363 41013 7372
rect 40876 7244 40916 7253
rect 40876 7085 40916 7204
rect 40875 7076 40917 7085
rect 40875 7036 40876 7076
rect 40916 7036 40917 7076
rect 40875 7027 40917 7036
rect 40875 6572 40917 6581
rect 40875 6532 40876 6572
rect 40916 6532 40917 6572
rect 40875 6523 40917 6532
rect 40876 6404 40916 6523
rect 40876 6355 40916 6364
rect 40972 5993 41012 7363
rect 41068 6992 41108 7001
rect 41068 6833 41108 6952
rect 41067 6824 41109 6833
rect 41067 6784 41068 6824
rect 41108 6784 41109 6824
rect 41067 6775 41109 6784
rect 41067 6488 41109 6497
rect 41067 6448 41068 6488
rect 41108 6448 41109 6488
rect 41067 6439 41109 6448
rect 41068 6320 41108 6439
rect 41068 6271 41108 6280
rect 40971 5984 41013 5993
rect 40971 5944 40972 5984
rect 41012 5944 41013 5984
rect 40971 5935 41013 5944
rect 40779 5900 40821 5909
rect 40779 5860 40780 5900
rect 40820 5860 40821 5900
rect 40779 5851 40821 5860
rect 40203 5816 40245 5825
rect 40203 5776 40204 5816
rect 40244 5776 40245 5816
rect 40203 5767 40245 5776
rect 41067 5816 41109 5825
rect 41067 5776 41068 5816
rect 41108 5776 41109 5816
rect 41067 5767 41109 5776
rect 40108 5683 40148 5692
rect 39820 5104 40052 5144
rect 39820 3977 39860 5104
rect 40012 4976 40052 4985
rect 40012 4397 40052 4936
rect 40011 4388 40053 4397
rect 40011 4348 40012 4388
rect 40052 4348 40053 4388
rect 40011 4339 40053 4348
rect 39916 4220 39956 4229
rect 39819 3968 39861 3977
rect 39819 3928 39820 3968
rect 39860 3928 39861 3968
rect 39819 3919 39861 3928
rect 39916 3893 39956 4180
rect 40108 3968 40148 3977
rect 39915 3884 39957 3893
rect 39915 3844 39916 3884
rect 39956 3844 39957 3884
rect 39915 3835 39957 3844
rect 40108 3557 40148 3928
rect 40107 3548 40149 3557
rect 39724 3508 39860 3548
rect 39627 3499 39669 3508
rect 39340 3380 39380 3389
rect 39380 3340 39476 3380
rect 39340 3331 39380 3340
rect 39339 2792 39381 2801
rect 39339 2752 39340 2792
rect 39380 2752 39381 2792
rect 39339 2743 39381 2752
rect 39243 2036 39285 2045
rect 39243 1996 39244 2036
rect 39284 1996 39285 2036
rect 39243 1987 39285 1996
rect 39340 1952 39380 2743
rect 39340 1903 39380 1912
rect 39244 1868 39284 1879
rect 39244 1793 39284 1828
rect 39051 1784 39093 1793
rect 39051 1744 39052 1784
rect 39092 1744 39093 1784
rect 39051 1735 39093 1744
rect 39243 1784 39285 1793
rect 39243 1744 39244 1784
rect 39284 1744 39285 1784
rect 39243 1735 39285 1744
rect 38708 1324 38804 1364
rect 38668 1315 38708 1324
rect 38379 1280 38421 1289
rect 38379 1240 38380 1280
rect 38420 1240 38421 1280
rect 38379 1231 38421 1240
rect 37268 1072 37460 1112
rect 38380 1112 38420 1231
rect 38476 1112 38516 1121
rect 38380 1072 38476 1112
rect 37228 1063 37268 1072
rect 38476 1063 38516 1072
rect 38859 1112 38901 1121
rect 38859 1072 38860 1112
rect 38900 1072 38901 1112
rect 38859 1063 38901 1072
rect 38860 978 38900 1063
rect 39436 953 39476 3340
rect 39532 3212 39572 3221
rect 39532 2633 39572 3172
rect 39531 2624 39573 2633
rect 39531 2584 39532 2624
rect 39572 2584 39573 2624
rect 39531 2575 39573 2584
rect 39628 2624 39668 3499
rect 39724 3380 39764 3389
rect 39724 2717 39764 3340
rect 39723 2708 39765 2717
rect 39723 2668 39724 2708
rect 39764 2668 39765 2708
rect 39723 2659 39765 2668
rect 39820 2624 39860 3508
rect 40107 3508 40108 3548
rect 40148 3508 40149 3548
rect 40107 3499 40149 3508
rect 40108 3380 40148 3389
rect 39915 3212 39957 3221
rect 39915 3172 39916 3212
rect 39956 3172 39957 3212
rect 39915 3163 39957 3172
rect 39916 3078 39956 3163
rect 40012 2624 40052 2633
rect 39820 2584 39956 2624
rect 39628 1373 39668 2584
rect 39819 2456 39861 2465
rect 39819 2416 39820 2456
rect 39860 2416 39861 2456
rect 39819 2407 39861 2416
rect 39820 2322 39860 2407
rect 39819 1952 39861 1961
rect 39819 1912 39820 1952
rect 39860 1912 39861 1952
rect 39819 1903 39861 1912
rect 39820 1818 39860 1903
rect 39916 1457 39956 2584
rect 39915 1448 39957 1457
rect 39915 1408 39916 1448
rect 39956 1408 39957 1448
rect 39915 1399 39957 1408
rect 39627 1364 39669 1373
rect 39627 1324 39628 1364
rect 39668 1324 39669 1364
rect 39627 1315 39669 1324
rect 40012 1121 40052 2584
rect 40108 1877 40148 3340
rect 40204 2801 40244 5767
rect 40492 5732 40532 5741
rect 40492 5573 40532 5692
rect 40876 5732 40916 5741
rect 40491 5564 40533 5573
rect 40491 5524 40492 5564
rect 40532 5524 40533 5564
rect 40491 5515 40533 5524
rect 40683 5480 40725 5489
rect 40683 5440 40684 5480
rect 40724 5440 40725 5480
rect 40683 5431 40725 5440
rect 40684 5346 40724 5431
rect 40876 5405 40916 5692
rect 41068 5682 41108 5767
rect 40875 5396 40917 5405
rect 40875 5356 40876 5396
rect 40916 5356 40917 5396
rect 40875 5347 40917 5356
rect 41067 5144 41109 5153
rect 41067 5104 41068 5144
rect 41108 5104 41109 5144
rect 41067 5095 41109 5104
rect 40492 4892 40532 4903
rect 40492 4817 40532 4852
rect 40875 4892 40917 4901
rect 40875 4852 40876 4892
rect 40916 4852 40917 4892
rect 40875 4843 40917 4852
rect 40491 4808 40533 4817
rect 40491 4768 40492 4808
rect 40532 4768 40533 4808
rect 40491 4759 40533 4768
rect 40683 4808 40725 4817
rect 40683 4768 40684 4808
rect 40724 4768 40725 4808
rect 40683 4759 40725 4768
rect 40684 4674 40724 4759
rect 40876 4758 40916 4843
rect 41068 4808 41108 5095
rect 41164 4892 41204 7699
rect 41260 7505 41300 7708
rect 41259 7496 41301 7505
rect 41259 7456 41260 7496
rect 41300 7456 41301 7496
rect 41259 7447 41301 7456
rect 41260 7244 41300 7253
rect 41260 6917 41300 7204
rect 41259 6908 41301 6917
rect 41259 6868 41260 6908
rect 41300 6868 41301 6908
rect 41259 6859 41301 6868
rect 41260 6413 41300 6498
rect 41259 6404 41301 6413
rect 41259 6364 41260 6404
rect 41300 6364 41301 6404
rect 41259 6355 41301 6364
rect 41259 5732 41301 5741
rect 41259 5692 41260 5732
rect 41300 5692 41301 5732
rect 41259 5683 41301 5692
rect 41260 5598 41300 5683
rect 41260 4892 41300 4901
rect 41164 4852 41260 4892
rect 41260 4843 41300 4852
rect 41356 4808 41396 9127
rect 41451 8504 41493 8513
rect 41451 8464 41452 8504
rect 41492 8464 41493 8504
rect 41451 8455 41493 8464
rect 41452 8370 41492 8455
rect 41451 7916 41493 7925
rect 41451 7876 41452 7916
rect 41492 7876 41493 7916
rect 41451 7867 41493 7876
rect 41452 7782 41492 7867
rect 41643 7832 41685 7841
rect 41643 7792 41644 7832
rect 41684 7792 41685 7832
rect 41643 7783 41685 7792
rect 41644 7698 41684 7783
rect 41451 7160 41493 7169
rect 41451 7120 41452 7160
rect 41492 7120 41493 7160
rect 41451 7111 41493 7120
rect 41452 6992 41492 7111
rect 41452 6943 41492 6952
rect 41451 6236 41493 6245
rect 41451 6196 41452 6236
rect 41492 6196 41493 6236
rect 41451 6187 41493 6196
rect 41452 6102 41492 6187
rect 41451 5900 41493 5909
rect 41451 5860 41452 5900
rect 41492 5860 41493 5900
rect 41451 5851 41493 5860
rect 41452 5766 41492 5851
rect 41452 4808 41492 4817
rect 41356 4768 41452 4808
rect 41068 4759 41108 4768
rect 41452 4759 41492 4768
rect 41259 4640 41301 4649
rect 41259 4600 41260 4640
rect 41300 4600 41301 4640
rect 41259 4591 41301 4600
rect 40875 4472 40917 4481
rect 40875 4432 40876 4472
rect 40916 4432 40917 4472
rect 40875 4423 40917 4432
rect 41067 4472 41109 4481
rect 41067 4432 41068 4472
rect 41108 4432 41109 4472
rect 41067 4423 41109 4432
rect 40395 4388 40437 4397
rect 40395 4348 40396 4388
rect 40436 4348 40437 4388
rect 40395 4339 40437 4348
rect 40299 4304 40341 4313
rect 40299 4264 40300 4304
rect 40340 4264 40341 4304
rect 40299 4255 40341 4264
rect 40300 4170 40340 4255
rect 40396 3380 40436 4339
rect 40491 4220 40533 4229
rect 40491 4180 40492 4220
rect 40532 4180 40533 4220
rect 40491 4171 40533 4180
rect 40876 4220 40916 4423
rect 41068 4388 41108 4423
rect 41068 4337 41108 4348
rect 40876 4171 40916 4180
rect 41260 4220 41300 4591
rect 41260 4171 41300 4180
rect 40492 4086 40532 4171
rect 41451 4136 41493 4145
rect 41451 4096 41452 4136
rect 41492 4096 41493 4136
rect 41451 4087 41493 4096
rect 41452 3968 41492 4087
rect 41452 3919 41492 3928
rect 41067 3800 41109 3809
rect 41067 3760 41068 3800
rect 41108 3760 41109 3800
rect 41067 3751 41109 3760
rect 41068 3632 41108 3751
rect 41259 3716 41301 3725
rect 41259 3676 41260 3716
rect 41300 3676 41301 3716
rect 41259 3667 41301 3676
rect 41068 3583 41108 3592
rect 40683 3464 40725 3473
rect 40683 3424 40684 3464
rect 40724 3424 40725 3464
rect 40683 3415 40725 3424
rect 40492 3380 40532 3389
rect 40396 3340 40492 3380
rect 40492 3331 40532 3340
rect 40684 3296 40724 3415
rect 40875 3380 40917 3389
rect 40875 3340 40876 3380
rect 40916 3340 40917 3380
rect 40875 3331 40917 3340
rect 41260 3380 41300 3667
rect 41260 3331 41300 3340
rect 40684 3247 40724 3256
rect 40876 3246 40916 3331
rect 40300 3212 40340 3221
rect 40779 3212 40821 3221
rect 40340 3172 40436 3212
rect 40300 3163 40340 3172
rect 40203 2792 40245 2801
rect 40203 2752 40204 2792
rect 40244 2752 40245 2792
rect 40203 2743 40245 2752
rect 40299 2456 40341 2465
rect 40299 2416 40300 2456
rect 40340 2416 40341 2456
rect 40299 2407 40341 2416
rect 40300 1947 40340 2407
rect 40300 1898 40340 1907
rect 40107 1868 40149 1877
rect 40107 1828 40108 1868
rect 40148 1828 40149 1868
rect 40107 1819 40149 1828
rect 40107 1364 40149 1373
rect 40107 1324 40108 1364
rect 40148 1324 40149 1364
rect 40107 1315 40149 1324
rect 40011 1112 40053 1121
rect 40011 1072 40012 1112
rect 40052 1072 40053 1112
rect 40011 1063 40053 1072
rect 40108 1112 40148 1315
rect 40108 1063 40148 1072
rect 39435 944 39477 953
rect 39435 904 39436 944
rect 39476 904 39477 944
rect 39435 895 39477 904
rect 40300 944 40340 953
rect 36843 860 36885 869
rect 36843 820 36844 860
rect 36884 820 36885 860
rect 36843 811 36885 820
rect 36651 692 36693 701
rect 36651 652 36652 692
rect 36692 652 36693 692
rect 36651 643 36693 652
rect 34539 524 34581 533
rect 34539 484 34540 524
rect 34580 484 34581 524
rect 34539 475 34581 484
rect 33963 440 34005 449
rect 33963 400 33964 440
rect 34004 400 34005 440
rect 33963 391 34005 400
rect 40300 113 40340 904
rect 40396 449 40436 3172
rect 40779 3172 40780 3212
rect 40820 3172 40821 3212
rect 40779 3163 40821 3172
rect 41451 3212 41493 3221
rect 41451 3172 41452 3212
rect 41492 3172 41493 3212
rect 41451 3163 41493 3172
rect 40587 2624 40629 2633
rect 40587 2584 40588 2624
rect 40628 2584 40629 2624
rect 40587 2575 40629 2584
rect 40492 2036 40532 2045
rect 40492 1196 40532 1996
rect 40492 1147 40532 1156
rect 40588 1121 40628 2575
rect 40683 1700 40725 1709
rect 40683 1660 40684 1700
rect 40724 1660 40725 1700
rect 40683 1651 40725 1660
rect 40684 1566 40724 1651
rect 40587 1112 40629 1121
rect 40587 1072 40588 1112
rect 40628 1072 40629 1112
rect 40587 1063 40629 1072
rect 40780 785 40820 3163
rect 41452 3078 41492 3163
rect 41643 2792 41685 2801
rect 41643 2752 41644 2792
rect 41684 2752 41685 2792
rect 41643 2743 41685 2752
rect 41451 2708 41493 2717
rect 41451 2668 41452 2708
rect 41492 2668 41493 2708
rect 41451 2659 41493 2668
rect 41260 2624 41300 2633
rect 41164 2584 41260 2624
rect 40875 2540 40917 2549
rect 40875 2500 40876 2540
rect 40916 2500 40917 2540
rect 40875 2491 40917 2500
rect 40876 1868 40916 2491
rect 41068 1868 41108 1877
rect 41164 1868 41204 2584
rect 41260 2575 41300 2584
rect 41452 2574 41492 2659
rect 41644 2658 41684 2743
rect 41259 2456 41301 2465
rect 41259 2416 41260 2456
rect 41300 2416 41301 2456
rect 41259 2407 41301 2416
rect 41260 2120 41300 2407
rect 41260 2071 41300 2080
rect 41643 2120 41685 2129
rect 41643 2080 41644 2120
rect 41684 2080 41685 2120
rect 41643 2071 41685 2080
rect 41644 1986 41684 2071
rect 40876 1819 40916 1828
rect 40972 1828 41068 1868
rect 41108 1828 41204 1868
rect 41452 1868 41492 1877
rect 40972 1289 41012 1828
rect 41068 1819 41108 1828
rect 41067 1700 41109 1709
rect 41067 1660 41068 1700
rect 41108 1660 41109 1700
rect 41067 1651 41109 1660
rect 40971 1280 41013 1289
rect 40971 1240 40972 1280
rect 41012 1240 41013 1280
rect 40971 1231 41013 1240
rect 41068 1280 41108 1651
rect 41452 1373 41492 1828
rect 41451 1364 41493 1373
rect 41451 1324 41452 1364
rect 41492 1324 41493 1364
rect 41451 1315 41493 1324
rect 41068 1231 41108 1240
rect 40875 1196 40917 1205
rect 40875 1156 40876 1196
rect 40916 1156 40917 1196
rect 40875 1147 40917 1156
rect 41260 1196 41300 1205
rect 40876 1062 40916 1147
rect 41260 869 41300 1156
rect 41452 944 41492 953
rect 41259 860 41301 869
rect 41259 820 41260 860
rect 41300 820 41301 860
rect 41259 811 41301 820
rect 40779 776 40821 785
rect 40779 736 40780 776
rect 40820 736 40821 776
rect 40779 727 40821 736
rect 40395 440 40437 449
rect 40395 400 40396 440
rect 40436 400 40437 440
rect 40395 391 40437 400
rect 41452 113 41492 904
rect 40299 104 40341 113
rect 26804 64 26824 80
rect 26744 0 26824 64
rect 26936 0 27016 80
rect 27128 0 27208 80
rect 27320 0 27400 80
rect 27512 0 27592 80
rect 27704 0 27784 80
rect 27896 0 27976 80
rect 28088 0 28168 80
rect 28280 0 28360 80
rect 28472 0 28552 80
rect 28664 0 28744 80
rect 28856 0 28936 80
rect 29048 0 29128 80
rect 29240 0 29320 80
rect 29432 0 29512 80
rect 29624 0 29704 80
rect 29816 0 29896 80
rect 30008 0 30088 80
rect 30200 0 30280 80
rect 30392 0 30472 80
rect 30584 0 30664 80
rect 30776 0 30856 80
rect 30968 0 31048 80
rect 31160 0 31240 80
rect 31352 0 31432 80
rect 31544 0 31624 80
rect 31736 0 31816 80
rect 31928 0 32008 80
rect 32120 0 32200 80
rect 32312 0 32392 80
rect 32504 0 32584 80
rect 32696 0 32776 80
rect 32888 0 32968 80
rect 33080 0 33160 80
rect 33272 0 33352 80
rect 33464 0 33544 80
rect 40299 64 40300 104
rect 40340 64 40341 104
rect 40299 55 40341 64
rect 41451 104 41493 113
rect 41451 64 41452 104
rect 41492 64 41493 104
rect 41451 55 41493 64
<< via2 >>
rect 1420 10144 1460 10184
rect 1708 9556 1748 9596
rect 1420 9472 1460 9512
rect 1228 9136 1268 9176
rect 1420 8884 1460 8924
rect 1228 8716 1268 8756
rect 1324 8632 1364 8672
rect 1612 9472 1652 9512
rect 1612 7624 1652 7664
rect 1420 7120 1460 7160
rect 1516 7036 1556 7076
rect 1324 6868 1364 6908
rect 1516 6616 1556 6656
rect 1324 6196 1364 6236
rect 1324 5608 1364 5648
rect 1516 5608 1556 5648
rect 1804 7540 1844 7580
rect 2188 9640 2228 9680
rect 2476 9556 2516 9596
rect 2188 7876 2228 7916
rect 1996 7372 2036 7412
rect 1708 6448 1748 6488
rect 1804 6280 1844 6320
rect 1996 6784 2036 6824
rect 1900 5440 1940 5480
rect 1324 4936 1364 4976
rect 1324 4684 1364 4724
rect 1420 3676 1460 3716
rect 1708 4432 1748 4472
rect 1612 3676 1652 3716
rect 1324 2752 1364 2792
rect 1324 2584 1364 2624
rect 1516 3256 1556 3296
rect 1612 3088 1652 3128
rect 1612 2920 1652 2960
rect 1420 2248 1460 2288
rect 1516 2164 1556 2204
rect 1804 3928 1844 3968
rect 1900 3424 1940 3464
rect 1804 3256 1844 3296
rect 1804 2836 1844 2876
rect 1804 1912 1844 1952
rect 1420 1744 1460 1784
rect 1324 1240 1364 1280
rect 1228 1156 1268 1196
rect 1804 1660 1844 1700
rect 1612 1492 1652 1532
rect 1900 1492 1940 1532
rect 1612 820 1652 860
rect 2380 8632 2420 8672
rect 2956 9472 2996 9512
rect 3244 9472 3284 9512
rect 2860 8464 2900 8504
rect 2764 8380 2804 8420
rect 3148 8380 3188 8420
rect 3052 8128 3092 8168
rect 2764 7960 2804 8000
rect 2476 7120 2516 7160
rect 2476 6700 2516 6740
rect 2284 6616 2324 6656
rect 2284 6112 2324 6152
rect 2188 2248 2228 2288
rect 2572 5692 2612 5732
rect 3052 7876 3092 7916
rect 2956 7288 2996 7328
rect 3340 8128 3380 8168
rect 3244 7960 3284 8000
rect 3244 7204 3284 7244
rect 2860 6616 2900 6656
rect 2956 5692 2996 5732
rect 3340 6952 3380 6992
rect 3148 6616 3188 6656
rect 3244 6280 3284 6320
rect 3148 5944 3188 5984
rect 2860 4936 2900 4976
rect 2764 4768 2804 4808
rect 2668 3676 2708 3716
rect 2668 3508 2708 3548
rect 3820 9556 3860 9596
rect 3628 9472 3668 9512
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 5644 10060 5684 10100
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 4492 9640 4532 9680
rect 4204 9136 4244 9176
rect 4012 8800 4052 8840
rect 4204 8800 4244 8840
rect 3628 8380 3668 8420
rect 4108 8296 4148 8336
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 3532 7372 3572 7412
rect 3916 7120 3956 7160
rect 3820 6868 3860 6908
rect 3436 6532 3476 6572
rect 3916 6448 3956 6488
rect 3340 5944 3380 5984
rect 3340 5776 3380 5816
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 4204 7792 4244 7832
rect 4204 7288 4244 7328
rect 4204 6448 4244 6488
rect 3532 5524 3572 5564
rect 3532 5356 3572 5396
rect 3436 5104 3476 5144
rect 3244 4936 3284 4976
rect 3724 5608 3764 5648
rect 3916 5608 3956 5648
rect 3820 5020 3860 5060
rect 4012 5524 4052 5564
rect 4012 5020 4052 5060
rect 4300 6280 4340 6320
rect 4780 9388 4820 9428
rect 4780 9220 4820 9260
rect 4492 7960 4532 8000
rect 4684 8128 4724 8168
rect 4588 7876 4628 7916
rect 5452 9472 5492 9512
rect 5068 9388 5108 9428
rect 5260 9304 5300 9344
rect 5356 9220 5396 9260
rect 5452 9052 5492 9092
rect 4972 8464 5012 8504
rect 5164 8500 5204 8504
rect 5164 8464 5204 8500
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 4780 7624 4820 7664
rect 5260 7876 5300 7916
rect 5356 7792 5396 7832
rect 5836 8968 5876 9008
rect 6124 8632 6164 8672
rect 4972 7288 5012 7328
rect 4492 7204 4532 7244
rect 4588 7036 4628 7076
rect 4780 7036 4820 7076
rect 4684 6868 4724 6908
rect 4972 6952 5012 6992
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 4588 6448 4628 6488
rect 5164 6448 5204 6488
rect 4876 6280 4916 6320
rect 4396 6196 4436 6236
rect 4684 5776 4724 5816
rect 4108 4936 4148 4976
rect 3916 4684 3956 4724
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 2956 4432 2996 4472
rect 4300 4684 4340 4724
rect 4204 4348 4244 4388
rect 3724 4264 3764 4304
rect 2956 4180 2996 4220
rect 3244 4180 3284 4220
rect 2860 3760 2900 3800
rect 4684 5440 4724 5480
rect 4588 4936 4628 4976
rect 5740 6532 5780 6572
rect 5836 6448 5876 6488
rect 5452 5776 5492 5816
rect 5356 5524 5396 5564
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 4876 4936 4916 4976
rect 5068 4936 5108 4976
rect 4972 4768 5012 4808
rect 4780 4684 4820 4724
rect 4492 4180 4532 4220
rect 4684 4180 4724 4220
rect 5452 5104 5492 5144
rect 5068 4600 5108 4640
rect 5356 4600 5396 4640
rect 5356 4180 5396 4220
rect 5260 4096 5300 4136
rect 4684 4012 4724 4052
rect 3244 3760 3284 3800
rect 2860 3508 2900 3548
rect 2764 3256 2804 3296
rect 3148 3172 3188 3212
rect 2956 2920 2996 2960
rect 3148 2752 3188 2792
rect 3532 3928 3572 3968
rect 4492 3844 4532 3884
rect 3436 3340 3476 3380
rect 3532 3256 3572 3296
rect 3244 2668 3284 2708
rect 3340 2500 3380 2540
rect 3244 2248 3284 2288
rect 2284 1744 2324 1784
rect 3340 1408 3380 1448
rect 3436 1072 3476 1112
rect 3820 3424 3860 3464
rect 4012 3424 4052 3464
rect 3724 3172 3764 3212
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 4108 1660 4148 1700
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 3724 1240 3764 1280
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 4684 3676 4724 3716
rect 4492 2920 4532 2960
rect 5068 3340 5108 3380
rect 4972 2668 5012 2708
rect 4300 2332 4340 2372
rect 5260 2584 5300 2624
rect 5548 4936 5588 4976
rect 5548 4096 5588 4136
rect 5548 3760 5588 3800
rect 5836 4096 5876 4136
rect 6700 9388 6740 9428
rect 6700 8632 6740 8672
rect 6700 8464 6740 8504
rect 6412 7624 6452 7664
rect 6028 6952 6068 6992
rect 6796 7540 6836 7580
rect 6508 6616 6548 6656
rect 6124 6364 6164 6404
rect 6412 6364 6452 6404
rect 6028 6280 6068 6320
rect 5932 3928 5972 3968
rect 5740 3676 5780 3716
rect 5644 3256 5684 3296
rect 6316 5776 6356 5816
rect 6124 4180 6164 4220
rect 6028 3760 6068 3800
rect 6508 6280 6548 6320
rect 6700 6448 6740 6488
rect 6604 6112 6644 6152
rect 6604 5860 6644 5900
rect 6508 5440 6548 5480
rect 6508 5272 6548 5312
rect 6796 6364 6836 6404
rect 7180 9304 7220 9344
rect 7084 9052 7124 9092
rect 6988 8464 7028 8504
rect 7372 9052 7412 9092
rect 7468 8884 7508 8924
rect 7660 9472 7700 9512
rect 7372 8464 7412 8504
rect 7276 8380 7316 8420
rect 7276 7288 7316 7328
rect 6988 6532 7028 6572
rect 6892 6112 6932 6152
rect 6412 4684 6452 4724
rect 6316 4012 6356 4052
rect 5932 3172 5972 3212
rect 4492 1660 4532 1700
rect 4300 1492 4340 1532
rect 3820 1072 3860 1112
rect 4396 1072 4436 1112
rect 2092 904 2132 944
rect 3532 904 3572 944
rect 3244 820 3284 860
rect 5836 3088 5876 3128
rect 6220 3088 6260 3128
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 4876 1996 4916 2036
rect 5260 1912 5300 1952
rect 5356 1744 5396 1784
rect 5164 1576 5204 1616
rect 4684 1240 4724 1280
rect 5068 1240 5108 1280
rect 5164 1072 5204 1112
rect 4492 820 4532 860
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 1804 568 1844 608
rect 5740 2248 5780 2288
rect 5836 1912 5876 1952
rect 5644 1660 5684 1700
rect 5548 1492 5588 1532
rect 5452 1156 5492 1196
rect 5836 1408 5876 1448
rect 6220 1828 6260 1868
rect 5452 652 5492 692
rect 5932 1072 5972 1112
rect 6412 3676 6452 3716
rect 6604 4684 6644 4724
rect 6892 5608 6932 5648
rect 7180 6952 7220 6992
rect 7084 6280 7124 6320
rect 7276 6364 7316 6404
rect 7276 6196 7316 6236
rect 7180 5776 7220 5816
rect 6796 5272 6836 5312
rect 6796 4852 6836 4892
rect 6700 4432 6740 4472
rect 6604 3928 6644 3968
rect 6796 3676 6836 3716
rect 6508 1660 6548 1700
rect 7756 8632 7796 8672
rect 7660 7960 7700 8000
rect 7756 7540 7796 7580
rect 8140 8128 8180 8168
rect 8716 10144 8756 10184
rect 8620 9640 8660 9680
rect 8332 9304 8372 9344
rect 8716 9472 8756 9512
rect 9004 9724 9044 9764
rect 8428 9136 8468 9176
rect 8812 9052 8852 9092
rect 8812 8548 8852 8588
rect 8620 8464 8660 8504
rect 7852 7372 7892 7412
rect 7564 7036 7604 7076
rect 7372 6028 7412 6068
rect 7276 5104 7316 5144
rect 7276 4936 7316 4976
rect 7660 6532 7700 6572
rect 7468 5860 7508 5900
rect 7660 6196 7700 6236
rect 7372 4348 7412 4388
rect 7180 4264 7220 4304
rect 8044 7288 8084 7328
rect 8140 6616 8180 6656
rect 8140 6448 8180 6488
rect 8236 5692 8276 5732
rect 7660 5020 7700 5060
rect 7564 4852 7604 4892
rect 7180 4012 7220 4052
rect 7372 3928 7412 3968
rect 7564 3844 7604 3884
rect 7084 3340 7124 3380
rect 7276 3256 7316 3296
rect 7084 3004 7124 3044
rect 7084 2752 7124 2792
rect 6988 2500 7028 2540
rect 6892 2248 6932 2288
rect 6892 1072 6932 1112
rect 7180 2500 7220 2540
rect 7468 3172 7508 3212
rect 7660 3760 7700 3800
rect 7852 5188 7892 5228
rect 8524 7960 8564 8000
rect 11020 10060 11060 10100
rect 11500 9724 11540 9764
rect 9004 8548 9044 8588
rect 8908 8128 8948 8168
rect 8620 7876 8660 7916
rect 8428 6868 8468 6908
rect 8620 7288 8660 7328
rect 8716 6616 8756 6656
rect 9004 7372 9044 7412
rect 8620 6364 8660 6404
rect 8524 6196 8564 6236
rect 9484 8716 9524 8756
rect 10732 9472 10772 9512
rect 11116 9472 11156 9512
rect 9868 9304 9908 9344
rect 9580 8632 9620 8672
rect 9772 8632 9812 8672
rect 9484 8128 9524 8168
rect 9388 8044 9428 8084
rect 9772 8380 9812 8420
rect 11116 9136 11156 9176
rect 10732 9052 10772 9092
rect 10348 8800 10388 8840
rect 9868 8296 9908 8336
rect 9676 8128 9716 8168
rect 10156 8548 10196 8588
rect 10060 8380 10100 8420
rect 10060 8212 10100 8252
rect 9964 7960 10004 8000
rect 10156 8128 10196 8168
rect 9676 7792 9716 7832
rect 9676 7624 9716 7664
rect 9100 6784 9140 6824
rect 9580 7120 9620 7160
rect 10444 8632 10484 8672
rect 10348 8296 10388 8336
rect 10540 8548 10580 8588
rect 10636 8464 10676 8504
rect 11020 8716 11060 8756
rect 11020 8548 11060 8588
rect 10636 8044 10676 8084
rect 11404 7960 11444 8000
rect 10252 7540 10292 7580
rect 9676 6868 9716 6908
rect 9580 6784 9620 6824
rect 9292 6616 9332 6656
rect 8812 6280 8852 6320
rect 8716 6112 8756 6152
rect 8428 5692 8468 5732
rect 8332 5440 8372 5480
rect 8428 5188 8468 5228
rect 8524 5020 8564 5060
rect 8716 5608 8756 5648
rect 9004 5944 9044 5984
rect 9292 5944 9332 5984
rect 9196 5776 9236 5816
rect 8908 5104 8948 5144
rect 9100 5608 9140 5648
rect 9004 5020 9044 5060
rect 8620 4936 8660 4976
rect 8620 4432 8660 4472
rect 7948 3508 7988 3548
rect 8620 4012 8660 4052
rect 8524 3928 8564 3968
rect 8428 3172 8468 3212
rect 7948 3088 7988 3128
rect 8428 2668 8468 2708
rect 9004 4348 9044 4388
rect 9004 3760 9044 3800
rect 8908 3676 8948 3716
rect 9196 4264 9236 4304
rect 9580 5440 9620 5480
rect 9484 5188 9524 5228
rect 9388 5020 9428 5060
rect 9388 4600 9428 4640
rect 9292 3508 9332 3548
rect 8620 3256 8660 3296
rect 9100 3256 9140 3296
rect 9580 5020 9620 5060
rect 9772 4684 9812 4724
rect 9580 3844 9620 3884
rect 8812 2584 8852 2624
rect 7564 2080 7604 2120
rect 7852 1996 7892 2036
rect 7180 1744 7220 1784
rect 7948 1660 7988 1700
rect 8428 1828 8468 1868
rect 8332 1492 8372 1532
rect 7756 1240 7796 1280
rect 9676 2668 9716 2708
rect 9196 2584 9236 2624
rect 8908 1156 8948 1196
rect 7372 1072 7412 1112
rect 7948 1072 7988 1112
rect 8620 1072 8660 1112
rect 9388 2416 9428 2456
rect 9580 1996 9620 2036
rect 10252 5440 10292 5480
rect 10348 4936 10388 4976
rect 10924 7456 10964 7496
rect 10924 6952 10964 6992
rect 11308 6952 11348 6992
rect 11596 8632 11636 8672
rect 12844 10480 12884 10520
rect 12748 9472 12788 9512
rect 12748 8800 12788 8840
rect 12076 8716 12116 8756
rect 12460 8716 12500 8756
rect 12652 8716 12692 8756
rect 11884 8632 11924 8672
rect 11596 8296 11636 8336
rect 11596 7708 11636 7748
rect 11596 7540 11636 7580
rect 11500 7456 11540 7496
rect 11500 7204 11540 7244
rect 11500 7036 11540 7076
rect 11500 6448 11540 6488
rect 11788 7708 11828 7748
rect 12076 7960 12116 8000
rect 11884 7372 11924 7412
rect 11884 7036 11924 7076
rect 11884 6868 11924 6908
rect 11788 6784 11828 6824
rect 10828 6364 10868 6404
rect 11308 6364 11348 6404
rect 10156 4768 10196 4808
rect 10060 4348 10100 4388
rect 9964 4096 10004 4136
rect 10636 5440 10676 5480
rect 10540 4852 10580 4892
rect 10924 4768 10964 4808
rect 10924 4516 10964 4556
rect 10828 4096 10868 4136
rect 10636 3676 10676 3716
rect 10060 3004 10100 3044
rect 10060 2584 10100 2624
rect 9772 2332 9812 2372
rect 9964 2080 10004 2120
rect 9868 1912 9908 1952
rect 10060 1744 10100 1784
rect 9484 1408 9524 1448
rect 9772 1408 9812 1448
rect 9388 988 9428 1028
rect 6604 736 6644 776
rect 5356 64 5396 104
rect 5644 64 5684 104
rect 6508 64 6548 104
rect 9676 1072 9716 1112
rect 9676 820 9716 860
rect 11116 6196 11156 6236
rect 11596 5692 11636 5732
rect 11500 5104 11540 5144
rect 11404 5020 11444 5060
rect 11308 4936 11348 4976
rect 11404 4852 11444 4892
rect 11404 3424 11444 3464
rect 11116 2752 11156 2792
rect 10636 2668 10676 2708
rect 11404 3004 11444 3044
rect 11212 2668 11252 2708
rect 11404 2584 11444 2624
rect 10540 2164 10580 2204
rect 10252 2080 10292 2120
rect 10348 1660 10388 1700
rect 10252 1156 10292 1196
rect 10636 1828 10676 1868
rect 10540 1660 10580 1700
rect 10444 1240 10484 1280
rect 10156 820 10196 860
rect 10252 568 10292 608
rect 10732 1072 10772 1112
rect 11116 1492 11156 1532
rect 10924 1408 10964 1448
rect 10924 1240 10964 1280
rect 10828 988 10868 1028
rect 11692 4936 11732 4976
rect 11596 3172 11636 3212
rect 11884 6700 11924 6740
rect 12652 8464 12692 8504
rect 12556 8296 12596 8336
rect 12364 7372 12404 7412
rect 12268 6448 12308 6488
rect 12172 6280 12212 6320
rect 12748 6028 12788 6068
rect 11884 5020 11924 5060
rect 12556 5356 12596 5396
rect 12268 5272 12308 5312
rect 12460 5272 12500 5312
rect 12076 4936 12116 4976
rect 11884 4432 11924 4472
rect 11788 3004 11828 3044
rect 11980 2752 12020 2792
rect 11788 2668 11828 2708
rect 11308 1744 11348 1784
rect 11692 1744 11732 1784
rect 11596 1072 11636 1112
rect 11020 904 11060 944
rect 10924 736 10964 776
rect 11404 988 11444 1028
rect 11788 1492 11828 1532
rect 11404 64 11444 104
rect 12076 2080 12116 2120
rect 11980 1240 12020 1280
rect 12268 4432 12308 4472
rect 12268 3928 12308 3968
rect 12556 4936 12596 4976
rect 12364 3760 12404 3800
rect 12268 3676 12308 3716
rect 12460 3676 12500 3716
rect 12460 3340 12500 3380
rect 12268 2668 12308 2708
rect 12460 2584 12500 2624
rect 12652 3340 12692 3380
rect 12940 8800 12980 8840
rect 13036 8632 13076 8672
rect 13228 8548 13268 8588
rect 12940 8296 12980 8336
rect 13132 8296 13172 8336
rect 13420 9640 13460 9680
rect 14284 9472 14324 9512
rect 14092 9136 14132 9176
rect 13708 8884 13748 8924
rect 13612 8716 13652 8756
rect 13516 8632 13556 8672
rect 13612 8464 13652 8504
rect 13420 8128 13460 8168
rect 13516 7288 13556 7328
rect 13900 8632 13940 8672
rect 13804 7960 13844 8000
rect 14188 8800 14228 8840
rect 14092 8464 14132 8504
rect 13996 8380 14036 8420
rect 13900 7876 13940 7916
rect 13708 7120 13748 7160
rect 16780 10648 16820 10688
rect 14764 9472 14804 9512
rect 14284 8128 14324 8168
rect 14284 7960 14324 8000
rect 13996 7372 14036 7412
rect 14188 7540 14228 7580
rect 14476 8632 14516 8672
rect 14380 7792 14420 7832
rect 14572 8464 14612 8504
rect 14476 7540 14516 7580
rect 14380 7372 14420 7412
rect 13132 6700 13172 6740
rect 13132 6532 13172 6572
rect 13036 6280 13076 6320
rect 13324 6196 13364 6236
rect 12940 5776 12980 5816
rect 12844 4264 12884 4304
rect 13228 5776 13268 5816
rect 13132 5356 13172 5396
rect 13804 6700 13844 6740
rect 13708 6112 13748 6152
rect 13420 5188 13460 5228
rect 13228 4768 13268 4808
rect 13132 3928 13172 3968
rect 13036 3676 13076 3716
rect 12940 3256 12980 3296
rect 12940 2836 12980 2876
rect 13036 2584 13076 2624
rect 12844 2416 12884 2456
rect 12748 2332 12788 2372
rect 12844 2248 12884 2288
rect 13036 2248 13076 2288
rect 12172 1576 12212 1616
rect 12172 1240 12212 1280
rect 12364 1240 12404 1280
rect 12748 1996 12788 2036
rect 12940 1912 12980 1952
rect 12652 1828 12692 1868
rect 12748 1324 12788 1364
rect 12556 568 12596 608
rect 13228 2836 13268 2876
rect 13708 5692 13748 5732
rect 13612 4852 13652 4892
rect 13612 4600 13652 4640
rect 14476 7120 14516 7160
rect 14476 6196 14516 6236
rect 13996 4936 14036 4976
rect 14284 4936 14324 4976
rect 13900 4096 13940 4136
rect 13900 3928 13940 3968
rect 13708 2584 13748 2624
rect 13612 2416 13652 2456
rect 13420 2332 13460 2372
rect 13420 1576 13460 1616
rect 13420 1408 13460 1448
rect 13324 1324 13364 1364
rect 13228 1240 13268 1280
rect 12844 1072 12884 1112
rect 13900 2752 13940 2792
rect 13900 2584 13940 2624
rect 13804 2080 13844 2120
rect 14284 4600 14324 4640
rect 14380 4180 14420 4220
rect 15436 8632 15476 8672
rect 15052 8548 15092 8588
rect 15340 8128 15380 8168
rect 16012 9472 16052 9512
rect 17452 9472 17492 9512
rect 17644 9472 17684 9512
rect 16396 9388 16436 9428
rect 16204 9220 16244 9260
rect 16588 9220 16628 9260
rect 16300 8800 16340 8840
rect 16204 8632 16244 8672
rect 16108 8548 16148 8588
rect 14668 7288 14708 7328
rect 14956 7288 14996 7328
rect 15436 7960 15476 8000
rect 16012 7876 16052 7916
rect 15052 6700 15092 6740
rect 15340 6532 15380 6572
rect 14956 6280 14996 6320
rect 16108 7372 16148 7412
rect 15724 7036 15764 7076
rect 15628 6952 15668 6992
rect 15436 6196 15476 6236
rect 14668 5272 14708 5312
rect 14860 4936 14900 4976
rect 15724 6616 15764 6656
rect 15724 6196 15764 6236
rect 15628 4768 15668 4808
rect 14860 4348 14900 4388
rect 14572 4264 14612 4304
rect 16204 6952 16244 6992
rect 16108 6868 16148 6908
rect 19372 9472 19412 9512
rect 19756 9472 19796 9512
rect 18124 9304 18164 9344
rect 19372 9136 19412 9176
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 17932 8800 17972 8840
rect 18124 8800 18164 8840
rect 17356 7960 17396 8000
rect 16684 7204 16724 7244
rect 16396 6616 16436 6656
rect 16108 6448 16148 6488
rect 16204 5608 16244 5648
rect 14284 3760 14324 3800
rect 14188 3592 14228 3632
rect 14188 3424 14228 3464
rect 14188 3088 14228 3128
rect 14668 3928 14708 3968
rect 14860 3508 14900 3548
rect 14668 3256 14708 3296
rect 14572 3088 14612 3128
rect 14476 2500 14516 2540
rect 14284 2164 14324 2204
rect 14092 1912 14132 1952
rect 13804 1576 13844 1616
rect 13708 1072 13748 1112
rect 13324 736 13364 776
rect 13516 820 13556 860
rect 13420 232 13460 272
rect 13996 1744 14036 1784
rect 13900 820 13940 860
rect 13804 736 13844 776
rect 13900 652 13940 692
rect 13708 64 13748 104
rect 14092 400 14132 440
rect 14572 2416 14612 2456
rect 15052 2584 15092 2624
rect 14956 2248 14996 2288
rect 15916 3928 15956 3968
rect 16108 3760 16148 3800
rect 16012 3424 16052 3464
rect 15820 3340 15860 3380
rect 15532 2668 15572 2708
rect 15244 2584 15284 2624
rect 15244 2332 15284 2372
rect 14956 1744 14996 1784
rect 15148 1744 15188 1784
rect 14668 1408 14708 1448
rect 15052 1408 15092 1448
rect 14860 1240 14900 1280
rect 14668 1072 14708 1112
rect 15148 1156 15188 1196
rect 14476 736 14516 776
rect 15052 820 15092 860
rect 14860 148 14900 188
rect 15148 568 15188 608
rect 15820 2500 15860 2540
rect 15436 1240 15476 1280
rect 15820 1828 15860 1868
rect 15436 1072 15476 1112
rect 15628 1156 15668 1196
rect 15532 988 15572 1028
rect 15628 736 15668 776
rect 16108 1408 16148 1448
rect 16684 4936 16724 4976
rect 16300 2836 16340 2876
rect 17164 5440 17204 5480
rect 17068 5104 17108 5144
rect 16780 2416 16820 2456
rect 16588 2164 16628 2204
rect 16492 1996 16532 2036
rect 16396 1912 16436 1952
rect 16300 1072 16340 1112
rect 16012 568 16052 608
rect 15724 484 15764 524
rect 16204 736 16244 776
rect 16012 232 16052 272
rect 16492 1324 16532 1364
rect 16396 316 16436 356
rect 16492 148 16532 188
rect 16780 2080 16820 2120
rect 16780 820 16820 860
rect 16876 652 16916 692
rect 18028 8632 18068 8672
rect 18508 8548 18548 8588
rect 17644 8212 17684 8252
rect 17452 7036 17492 7076
rect 17356 5608 17396 5648
rect 17548 6448 17588 6488
rect 17548 6280 17588 6320
rect 18412 8464 18452 8504
rect 18220 8380 18260 8420
rect 17740 7120 17780 7160
rect 18028 6952 18068 6992
rect 17932 6280 17972 6320
rect 17260 3676 17300 3716
rect 17164 2500 17204 2540
rect 17548 4936 17588 4976
rect 17644 4684 17684 4724
rect 17644 4096 17684 4136
rect 17644 3424 17684 3464
rect 17644 2752 17684 2792
rect 17068 2164 17108 2204
rect 17356 2248 17396 2288
rect 18316 8128 18356 8168
rect 18220 6616 18260 6656
rect 18124 6448 18164 6488
rect 18316 6280 18356 6320
rect 18508 7876 18548 7916
rect 18124 4971 18164 4976
rect 18124 4936 18164 4971
rect 18028 4852 18068 4892
rect 17932 4012 17972 4052
rect 17836 3592 17876 3632
rect 17740 2584 17780 2624
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 19756 8716 19796 8756
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 21484 9640 21524 9680
rect 21004 9556 21044 9596
rect 20044 8716 20084 8756
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 19756 7960 19796 8000
rect 19660 7876 19700 7916
rect 19372 7456 19412 7496
rect 18796 7288 18836 7328
rect 18988 7120 19028 7160
rect 19180 6784 19220 6824
rect 18796 6448 18836 6488
rect 18604 6280 18644 6320
rect 18604 5776 18644 5816
rect 18412 5608 18452 5648
rect 18508 5524 18548 5564
rect 18412 4936 18452 4976
rect 18316 4852 18356 4892
rect 18412 4684 18452 4724
rect 18028 2332 18068 2372
rect 18316 3004 18356 3044
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 20524 8128 20564 8168
rect 20812 8044 20852 8084
rect 20428 7876 20468 7916
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 20236 6616 20276 6656
rect 19852 6532 19892 6572
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 18892 3676 18932 3716
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 19660 4936 19700 4976
rect 20620 7120 20660 7160
rect 20716 5356 20756 5396
rect 20620 5272 20660 5312
rect 20620 5104 20660 5144
rect 21004 7540 21044 7580
rect 21004 7120 21044 7160
rect 21004 6616 21044 6656
rect 23692 10396 23732 10436
rect 22636 9556 22676 9596
rect 24460 9472 24500 9512
rect 23212 9388 23252 9428
rect 21484 8968 21524 9008
rect 21292 8800 21332 8840
rect 21292 8632 21332 8672
rect 22732 8800 22772 8840
rect 22540 8716 22580 8756
rect 22060 7540 22100 7580
rect 21484 7120 21524 7160
rect 21388 6868 21428 6908
rect 21004 6364 21044 6404
rect 21292 6364 21332 6404
rect 21100 6280 21140 6320
rect 21772 5944 21812 5984
rect 21100 5440 21140 5480
rect 21196 5272 21236 5312
rect 22540 7540 22580 7580
rect 22444 7456 22484 7496
rect 23020 8800 23060 8840
rect 22636 7456 22676 7496
rect 22444 6616 22484 6656
rect 22252 5860 22292 5900
rect 22348 5692 22388 5732
rect 22252 5440 22292 5480
rect 21772 5272 21812 5312
rect 20908 5020 20948 5060
rect 21388 5020 21428 5060
rect 21676 5020 21716 5060
rect 20236 4852 20276 4892
rect 20524 4852 20564 4892
rect 21004 4852 21044 4892
rect 21292 4852 21332 4892
rect 21100 4768 21140 4808
rect 20620 4264 20660 4304
rect 20044 4096 20084 4136
rect 20620 4012 20660 4052
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 18316 2584 18356 2624
rect 18412 2500 18452 2540
rect 18124 2248 18164 2288
rect 17644 1912 17684 1952
rect 18028 1492 18068 1532
rect 18124 1072 18164 1112
rect 17932 652 17972 692
rect 18220 736 18260 776
rect 18412 1996 18452 2036
rect 18412 1492 18452 1532
rect 18604 2584 18644 2624
rect 18604 1744 18644 1784
rect 19180 2584 19220 2624
rect 18604 904 18644 944
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 19372 3172 19412 3212
rect 19468 3004 19508 3044
rect 19372 2500 19412 2540
rect 20812 3928 20852 3968
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 20524 3676 20564 3716
rect 21100 3928 21140 3968
rect 21196 3760 21236 3800
rect 22060 4936 22100 4976
rect 23212 6868 23252 6908
rect 23116 6448 23156 6488
rect 23212 5692 23252 5732
rect 22540 5020 22580 5060
rect 21676 4684 21716 4724
rect 22444 4684 22484 4724
rect 22156 4432 22196 4472
rect 21868 4096 21908 4136
rect 22348 4012 22388 4052
rect 19660 3004 19700 3044
rect 20236 3004 20276 3044
rect 19660 2752 19700 2792
rect 19948 2500 19988 2540
rect 20140 2500 20180 2540
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 19564 2080 19604 2120
rect 19468 1912 19508 1952
rect 19372 1492 19412 1532
rect 19852 1996 19892 2036
rect 19564 1492 19604 1532
rect 20524 1240 20564 1280
rect 19660 1156 19700 1196
rect 19276 904 19316 944
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 20620 1156 20660 1196
rect 20236 568 20276 608
rect 20044 484 20084 524
rect 19852 232 19892 272
rect 20716 1072 20756 1112
rect 20908 988 20948 1028
rect 21292 3592 21332 3632
rect 21292 2752 21332 2792
rect 21100 1660 21140 1700
rect 21484 1324 21524 1364
rect 21388 568 21428 608
rect 21868 3844 21908 3884
rect 21772 2752 21812 2792
rect 22060 2836 22100 2876
rect 22348 3844 22388 3884
rect 22252 3760 22292 3800
rect 21868 2332 21908 2372
rect 21964 2248 22004 2288
rect 21868 2164 21908 2204
rect 21964 1744 22004 1784
rect 21868 1660 21908 1700
rect 21772 1072 21812 1112
rect 21772 904 21812 944
rect 21964 1072 22004 1112
rect 22156 1324 22196 1364
rect 22444 3592 22484 3632
rect 22444 2668 22484 2708
rect 22828 4264 22868 4304
rect 22732 3760 22772 3800
rect 23596 8380 23636 8420
rect 24076 8296 24116 8336
rect 23500 8212 23540 8252
rect 25996 10564 26036 10604
rect 27148 10480 27188 10520
rect 28300 9808 28340 9848
rect 27916 9724 27956 9764
rect 26284 9556 26324 9596
rect 25036 9472 25076 9512
rect 24748 8464 24788 8504
rect 25036 9052 25076 9092
rect 23500 7792 23540 7832
rect 24844 7960 24884 8000
rect 25900 8968 25940 9008
rect 25228 8632 25268 8672
rect 25612 8632 25652 8672
rect 25612 8464 25652 8504
rect 25516 8296 25556 8336
rect 24364 7540 24404 7580
rect 24652 7540 24692 7580
rect 23692 6700 23732 6740
rect 23884 6532 23924 6572
rect 23596 6280 23636 6320
rect 23308 4768 23348 4808
rect 23212 4516 23252 4556
rect 23116 4348 23156 4388
rect 23020 3424 23060 3464
rect 22444 2080 22484 2120
rect 22060 820 22100 860
rect 22252 820 22292 860
rect 22636 1324 22676 1364
rect 22636 484 22676 524
rect 23020 3004 23060 3044
rect 23116 2752 23156 2792
rect 23116 1828 23156 1868
rect 23116 1660 23156 1700
rect 23020 1240 23060 1280
rect 23500 3760 23540 3800
rect 24844 7204 24884 7244
rect 25228 7204 25268 7244
rect 24940 7036 24980 7076
rect 25708 8380 25748 8420
rect 25804 7204 25844 7244
rect 24940 6616 24980 6656
rect 24364 6532 24404 6572
rect 24460 5608 24500 5648
rect 23980 3424 24020 3464
rect 24940 5440 24980 5480
rect 24844 5104 24884 5144
rect 24556 4936 24596 4976
rect 25132 6364 25172 6404
rect 24460 4432 24500 4472
rect 24076 3004 24116 3044
rect 23692 2668 23732 2708
rect 24076 2668 24116 2708
rect 23308 1996 23348 2036
rect 23308 1324 23348 1364
rect 23212 1156 23252 1196
rect 24268 3760 24308 3800
rect 24556 3760 24596 3800
rect 24460 3088 24500 3128
rect 24268 2668 24308 2708
rect 23692 1660 23732 1700
rect 23884 1828 23924 1868
rect 24364 1576 24404 1616
rect 23596 1072 23636 1112
rect 23692 484 23732 524
rect 24172 1072 24212 1112
rect 24268 904 24308 944
rect 24076 820 24116 860
rect 24460 64 24500 104
rect 25228 6280 25268 6320
rect 24748 4096 24788 4136
rect 25516 6952 25556 6992
rect 25420 5776 25460 5816
rect 25324 3760 25364 3800
rect 24748 1912 24788 1952
rect 24844 1576 24884 1616
rect 25036 3004 25076 3044
rect 24940 1324 24980 1364
rect 24940 736 24980 776
rect 24844 316 24884 356
rect 25132 2164 25172 2204
rect 25324 3172 25364 3212
rect 25228 2080 25268 2120
rect 25228 1912 25268 1952
rect 25324 1828 25364 1868
rect 26188 8548 26228 8588
rect 26188 8296 26228 8336
rect 26668 9472 26708 9512
rect 29260 9640 29300 9680
rect 29452 9640 29492 9680
rect 27916 9052 27956 9092
rect 27340 8716 27380 8756
rect 26476 8380 26516 8420
rect 26284 8044 26324 8084
rect 26380 7204 26420 7244
rect 25804 6784 25844 6824
rect 25612 6700 25652 6740
rect 25516 3760 25556 3800
rect 25900 6616 25940 6656
rect 26188 6532 26228 6572
rect 26860 7036 26900 7076
rect 26860 6448 26900 6488
rect 27628 8380 27668 8420
rect 27916 8380 27956 8420
rect 27052 7540 27092 7580
rect 27148 7204 27188 7244
rect 27532 7036 27572 7076
rect 29548 9556 29588 9596
rect 29260 9304 29300 9344
rect 29740 8716 29780 8756
rect 28780 8632 28820 8672
rect 28588 8044 28628 8084
rect 29356 8044 29396 8084
rect 28492 7876 28532 7916
rect 28780 7876 28820 7916
rect 28972 7792 29012 7832
rect 28204 7204 28244 7244
rect 28780 7204 28820 7244
rect 27820 6952 27860 6992
rect 27436 6868 27476 6908
rect 27148 6784 27188 6824
rect 27436 6616 27476 6656
rect 26956 6280 26996 6320
rect 27148 6196 27188 6236
rect 26092 5692 26132 5732
rect 26476 5692 26516 5732
rect 26188 4936 26228 4976
rect 25804 4432 25844 4472
rect 25708 4348 25748 4388
rect 26188 4432 26228 4472
rect 25708 4012 25748 4052
rect 26092 4012 26132 4052
rect 25708 3760 25748 3800
rect 25612 3592 25652 3632
rect 25612 3256 25652 3296
rect 26092 3592 26132 3632
rect 25516 2752 25556 2792
rect 25708 2752 25748 2792
rect 26956 4852 26996 4892
rect 26572 4180 26612 4220
rect 26380 4012 26420 4052
rect 26668 4012 26708 4052
rect 25996 2584 26036 2624
rect 25996 2080 26036 2120
rect 26572 3424 26612 3464
rect 26476 2752 26516 2792
rect 26380 2332 26420 2372
rect 26284 2164 26324 2204
rect 26092 1912 26132 1952
rect 26380 1912 26420 1952
rect 26188 1408 26228 1448
rect 25996 1156 26036 1196
rect 25612 1072 25652 1112
rect 25516 652 25556 692
rect 25708 988 25748 1028
rect 25804 652 25844 692
rect 26860 4096 26900 4136
rect 26668 1744 26708 1784
rect 27052 4684 27092 4724
rect 27052 4348 27092 4388
rect 27340 4096 27380 4136
rect 27628 5860 27668 5900
rect 27628 5608 27668 5648
rect 27148 3844 27188 3884
rect 27436 3760 27476 3800
rect 27628 3760 27668 3800
rect 27244 3172 27284 3212
rect 26956 1912 26996 1952
rect 26860 1156 26900 1196
rect 26572 652 26612 692
rect 26572 400 26612 440
rect 26764 64 26804 104
rect 27052 820 27092 860
rect 27052 652 27092 692
rect 27628 3508 27668 3548
rect 27724 3256 27764 3296
rect 27436 1912 27476 1952
rect 27340 1828 27380 1868
rect 27340 1660 27380 1700
rect 27244 1240 27284 1280
rect 27148 316 27188 356
rect 28012 6028 28052 6068
rect 28108 5776 28148 5816
rect 29164 6364 29204 6404
rect 28204 5356 28244 5396
rect 29452 6196 29492 6236
rect 29452 5860 29492 5900
rect 29644 5776 29684 5816
rect 28780 5356 28820 5396
rect 28300 3256 28340 3296
rect 28300 3088 28340 3128
rect 28300 2584 28340 2624
rect 28012 2500 28052 2540
rect 27628 2248 27668 2288
rect 27532 1240 27572 1280
rect 27436 1072 27476 1112
rect 27532 316 27572 356
rect 27916 2416 27956 2456
rect 28588 4516 28628 4556
rect 28780 2836 28820 2876
rect 28012 2332 28052 2372
rect 27820 1660 27860 1700
rect 27916 1156 27956 1196
rect 28204 904 28244 944
rect 28108 232 28148 272
rect 28396 1828 28436 1868
rect 29164 5020 29204 5060
rect 29356 5020 29396 5060
rect 29260 4012 29300 4052
rect 29068 3760 29108 3800
rect 28684 1072 28724 1112
rect 30508 8884 30548 8924
rect 30220 8632 30260 8672
rect 30220 8044 30260 8084
rect 30220 7876 30260 7916
rect 29932 7792 29972 7832
rect 30028 7708 30068 7748
rect 30412 7708 30452 7748
rect 30412 7456 30452 7496
rect 30412 7204 30452 7244
rect 29932 6868 29972 6908
rect 29836 6784 29876 6824
rect 29932 6700 29972 6740
rect 30028 6616 30068 6656
rect 29836 5272 29876 5312
rect 29932 5020 29972 5060
rect 29548 3844 29588 3884
rect 29452 3592 29492 3632
rect 29164 2500 29204 2540
rect 29068 1660 29108 1700
rect 29548 3004 29588 3044
rect 29548 2080 29588 2120
rect 29452 1828 29492 1868
rect 29260 1660 29300 1700
rect 28492 652 28532 692
rect 28684 148 28724 188
rect 29164 1072 29204 1112
rect 29068 904 29108 944
rect 29548 1492 29588 1532
rect 29452 1324 29492 1364
rect 29932 3760 29972 3800
rect 29932 3592 29972 3632
rect 30700 8884 30740 8924
rect 30892 8800 30932 8840
rect 31084 8128 31124 8168
rect 31564 8128 31604 8168
rect 30700 7540 30740 7580
rect 30604 7456 30644 7496
rect 31564 7960 31604 8000
rect 32236 10648 32276 10688
rect 32332 10396 32372 10436
rect 31852 8716 31892 8756
rect 31852 8044 31892 8084
rect 31756 7876 31796 7916
rect 30316 7036 30356 7076
rect 30412 6448 30452 6488
rect 30412 5692 30452 5732
rect 30508 5356 30548 5396
rect 30220 4768 30260 4808
rect 30124 3844 30164 3884
rect 30028 3424 30068 3464
rect 30412 3424 30452 3464
rect 31084 7120 31124 7160
rect 32140 7708 32180 7748
rect 32044 7540 32084 7580
rect 31756 7204 31796 7244
rect 30700 6448 30740 6488
rect 30796 6364 30836 6404
rect 31564 6112 31604 6152
rect 31180 5272 31220 5312
rect 31372 5440 31412 5480
rect 31276 5104 31316 5144
rect 30700 4348 30740 4388
rect 30220 2836 30260 2876
rect 29932 2584 29972 2624
rect 29836 1912 29876 1952
rect 30028 2164 30068 2204
rect 30412 2500 30452 2540
rect 30316 2248 30356 2288
rect 30220 1240 30260 1280
rect 29932 1156 29972 1196
rect 29836 1072 29876 1112
rect 29932 400 29972 440
rect 30316 568 30356 608
rect 31276 4768 31316 4808
rect 31276 4348 31316 4388
rect 31084 4180 31124 4220
rect 30892 3172 30932 3212
rect 30796 2836 30836 2876
rect 30508 2080 30548 2120
rect 30700 1828 30740 1868
rect 30892 1408 30932 1448
rect 30796 1156 30836 1196
rect 30700 1072 30740 1112
rect 31468 4348 31508 4388
rect 31948 6952 31988 6992
rect 31852 6868 31892 6908
rect 31756 6448 31796 6488
rect 31948 6532 31988 6572
rect 31948 6364 31988 6404
rect 31852 6028 31892 6068
rect 31948 5944 31988 5984
rect 31564 3592 31604 3632
rect 31276 3004 31316 3044
rect 31180 2920 31220 2960
rect 31564 2920 31604 2960
rect 31372 2836 31412 2876
rect 31180 2668 31220 2708
rect 31276 2584 31316 2624
rect 31084 2416 31124 2456
rect 31564 2500 31604 2540
rect 31756 5524 31796 5564
rect 31660 2080 31700 2120
rect 31468 1996 31508 2036
rect 31852 4180 31892 4220
rect 32140 7204 32180 7244
rect 32908 9472 32948 9512
rect 32428 8800 32468 8840
rect 32812 8632 32852 8672
rect 32428 8044 32468 8084
rect 32812 7876 32852 7916
rect 32716 7708 32756 7748
rect 32524 6448 32564 6488
rect 32140 6028 32180 6068
rect 32140 5104 32180 5144
rect 32428 5020 32468 5060
rect 32524 4852 32564 4892
rect 32332 4684 32372 4724
rect 31852 3928 31892 3968
rect 31852 3592 31892 3632
rect 31276 1324 31316 1364
rect 31372 1240 31412 1280
rect 31756 1660 31796 1700
rect 31660 1492 31700 1532
rect 31660 736 31700 776
rect 31756 652 31796 692
rect 31948 2836 31988 2876
rect 31948 1828 31988 1868
rect 31948 1072 31988 1112
rect 32812 7540 32852 7580
rect 33196 7456 33236 7496
rect 32908 7120 32948 7160
rect 33100 6280 33140 6320
rect 33004 6196 33044 6236
rect 32716 5524 32756 5564
rect 32812 5020 32852 5060
rect 32716 4684 32756 4724
rect 33004 5020 33044 5060
rect 32908 4264 32948 4304
rect 32812 4012 32852 4052
rect 32332 3844 32372 3884
rect 32332 2080 32372 2120
rect 32140 1828 32180 1868
rect 32140 1492 32180 1532
rect 32620 3760 32660 3800
rect 32428 1408 32468 1448
rect 32044 988 32084 1028
rect 32332 736 32372 776
rect 31852 148 31892 188
rect 32140 148 32180 188
rect 32524 988 32564 1028
rect 32428 400 32468 440
rect 33004 3424 33044 3464
rect 32812 2668 32852 2708
rect 32812 1912 32852 1952
rect 33004 1660 33044 1700
rect 32908 1324 32948 1364
rect 33004 988 33044 1028
rect 33292 7120 33332 7160
rect 33292 6364 33332 6404
rect 33196 5188 33236 5228
rect 34060 9892 34100 9932
rect 34540 9808 34580 9848
rect 33772 9220 33812 9260
rect 34348 9220 34388 9260
rect 33676 7960 33716 8000
rect 33928 9052 33968 9092
rect 34010 9052 34050 9092
rect 34092 9052 34132 9092
rect 34174 9052 34214 9092
rect 34256 9052 34296 9092
rect 34540 8884 34580 8924
rect 33964 8548 34004 8588
rect 34444 8548 34484 8588
rect 34444 8044 34484 8084
rect 33928 7540 33968 7580
rect 34010 7540 34050 7580
rect 34092 7540 34132 7580
rect 34174 7540 34214 7580
rect 34256 7540 34296 7580
rect 33772 6952 33812 6992
rect 33484 6784 33524 6824
rect 33580 6196 33620 6236
rect 33388 5860 33428 5900
rect 33388 5692 33428 5732
rect 33484 5356 33524 5396
rect 33388 5272 33428 5312
rect 33484 5020 33524 5060
rect 33292 4684 33332 4724
rect 33484 4180 33524 4220
rect 33388 4096 33428 4136
rect 33292 1408 33332 1448
rect 34348 7204 34388 7244
rect 34732 7708 34772 7748
rect 34444 7036 34484 7076
rect 34348 6952 34388 6992
rect 34444 6868 34484 6908
rect 34252 6700 34292 6740
rect 34540 6616 34580 6656
rect 34060 6532 34100 6572
rect 33928 6028 33968 6068
rect 34010 6028 34050 6068
rect 34092 6028 34132 6068
rect 34174 6028 34214 6068
rect 34256 6028 34296 6068
rect 34252 5860 34292 5900
rect 34252 5524 34292 5564
rect 33676 4684 33716 4724
rect 34060 4684 34100 4724
rect 34348 5356 34388 5396
rect 34444 5272 34484 5312
rect 34732 5608 34772 5648
rect 34732 5356 34772 5396
rect 35168 9808 35208 9848
rect 35250 9808 35290 9848
rect 35332 9808 35372 9848
rect 35414 9808 35454 9848
rect 35496 9808 35536 9848
rect 34924 9304 34964 9344
rect 35884 9220 35924 9260
rect 35168 8296 35208 8336
rect 35250 8296 35290 8336
rect 35332 8296 35372 8336
rect 35414 8296 35454 8336
rect 35496 8296 35536 8336
rect 35116 7960 35156 8000
rect 35596 7960 35636 8000
rect 35500 7708 35540 7748
rect 35692 7204 35732 7244
rect 35596 7036 35636 7076
rect 35020 6952 35060 6992
rect 35168 6784 35208 6824
rect 35250 6784 35290 6824
rect 35332 6784 35372 6824
rect 35414 6784 35454 6824
rect 35496 6784 35536 6824
rect 34924 6448 34964 6488
rect 35500 6448 35540 6488
rect 35980 7120 36020 7160
rect 35788 6952 35828 6992
rect 35020 5524 35060 5564
rect 35168 5272 35208 5312
rect 35250 5272 35290 5312
rect 35332 5272 35372 5312
rect 35414 5272 35454 5312
rect 35496 5272 35536 5312
rect 34444 4852 34484 4892
rect 35308 5020 35348 5060
rect 33928 4516 33968 4556
rect 34010 4516 34050 4556
rect 34092 4516 34132 4556
rect 34174 4516 34214 4556
rect 34256 4516 34296 4556
rect 34060 4012 34100 4052
rect 34252 3928 34292 3968
rect 33868 3592 33908 3632
rect 34252 3508 34292 3548
rect 33676 3256 33716 3296
rect 33580 3172 33620 3212
rect 33580 1912 33620 1952
rect 33928 3004 33968 3044
rect 34010 3004 34050 3044
rect 34092 3004 34132 3044
rect 34174 3004 34214 3044
rect 34256 3004 34296 3044
rect 33772 2416 33812 2456
rect 34252 2248 34292 2288
rect 33964 2164 34004 2204
rect 34444 4012 34484 4052
rect 34444 3592 34484 3632
rect 34444 2500 34484 2540
rect 34444 2080 34484 2120
rect 34252 1660 34292 1700
rect 33928 1492 33968 1532
rect 34010 1492 34050 1532
rect 34092 1492 34132 1532
rect 34174 1492 34214 1532
rect 34256 1492 34296 1532
rect 33676 1324 33716 1364
rect 33772 1240 33812 1280
rect 34348 1240 34388 1280
rect 33580 1072 33620 1112
rect 33964 1072 34004 1112
rect 35020 4684 35060 4724
rect 34636 3592 34676 3632
rect 34636 2248 34676 2288
rect 35500 3928 35540 3968
rect 35168 3760 35208 3800
rect 35250 3760 35290 3800
rect 35332 3760 35372 3800
rect 35414 3760 35454 3800
rect 35496 3760 35536 3800
rect 35692 5440 35732 5480
rect 35884 6868 35924 6908
rect 36556 10564 36596 10604
rect 36940 10480 36980 10520
rect 37324 9640 37364 9680
rect 40972 10480 41012 10520
rect 40684 10144 40724 10184
rect 39340 9892 39380 9932
rect 38668 9640 38708 9680
rect 39724 9640 39764 9680
rect 40876 9724 40916 9764
rect 36364 9388 36404 9428
rect 36364 9220 36404 9260
rect 37132 9052 37172 9092
rect 36652 8716 36692 8756
rect 36556 8380 36596 8420
rect 36364 8128 36404 8168
rect 36268 7960 36308 8000
rect 36172 6784 36212 6824
rect 36076 6616 36116 6656
rect 36172 6532 36212 6572
rect 35884 5608 35924 5648
rect 35692 4180 35732 4220
rect 35692 3928 35732 3968
rect 35692 3760 35732 3800
rect 35020 3592 35060 3632
rect 34828 3508 34868 3548
rect 34924 2332 34964 2372
rect 35168 2248 35208 2288
rect 35250 2248 35290 2288
rect 35332 2248 35372 2288
rect 35414 2248 35454 2288
rect 35496 2248 35536 2288
rect 36364 7876 36404 7916
rect 36460 7204 36500 7244
rect 36364 7036 36404 7076
rect 36364 6616 36404 6656
rect 36460 6532 36500 6572
rect 36748 8380 36788 8420
rect 36748 8128 36788 8168
rect 36652 6700 36692 6740
rect 36940 8044 36980 8084
rect 36940 7708 36980 7748
rect 36844 7204 36884 7244
rect 36652 5860 36692 5900
rect 36652 5692 36692 5732
rect 36364 5440 36404 5480
rect 36748 4852 36788 4892
rect 36940 6868 36980 6908
rect 37420 8044 37460 8084
rect 38188 9388 38228 9428
rect 37708 9304 37748 9344
rect 38380 8632 38420 8672
rect 37804 7624 37844 7664
rect 37708 7288 37748 7328
rect 37516 7204 37556 7244
rect 37132 6700 37172 6740
rect 37708 6868 37748 6908
rect 37324 6784 37364 6824
rect 38092 7960 38132 8000
rect 37996 6364 38036 6404
rect 37612 6028 37652 6068
rect 37036 5440 37076 5480
rect 36940 5020 36980 5060
rect 37804 5692 37844 5732
rect 37996 5608 38036 5648
rect 37612 5524 37652 5564
rect 37612 5104 37652 5144
rect 37516 5020 37556 5060
rect 37228 4936 37268 4976
rect 37132 4852 37172 4892
rect 37612 4852 37652 4892
rect 37804 4852 37844 4892
rect 36076 3760 36116 3800
rect 35884 3424 35924 3464
rect 36076 3424 36116 3464
rect 36076 2836 36116 2876
rect 37036 4180 37076 4220
rect 36172 2752 36212 2792
rect 36556 2668 36596 2708
rect 36460 1996 36500 2036
rect 34732 1828 34772 1868
rect 34828 1660 34868 1700
rect 36556 1828 36596 1868
rect 35212 1324 35252 1364
rect 34636 1240 34676 1280
rect 35596 1240 35636 1280
rect 34636 1072 34676 1112
rect 35212 1072 35252 1112
rect 35596 1072 35636 1112
rect 36556 1156 36596 1196
rect 36268 904 36308 944
rect 35168 736 35208 776
rect 35250 736 35290 776
rect 35332 736 35372 776
rect 35414 736 35454 776
rect 35496 736 35536 776
rect 36940 3172 36980 3212
rect 37036 2584 37076 2624
rect 37516 3340 37556 3380
rect 37420 2836 37460 2876
rect 37516 2752 37556 2792
rect 37804 4012 37844 4052
rect 37708 3340 37748 3380
rect 37996 4096 38036 4136
rect 37708 2668 37748 2708
rect 37804 2584 37844 2624
rect 37324 2164 37364 2204
rect 37132 2080 37172 2120
rect 37324 1996 37364 2036
rect 36844 1912 36884 1952
rect 37228 1912 37268 1952
rect 36748 1156 36788 1196
rect 36748 988 36788 1028
rect 37804 2248 37844 2288
rect 38380 7120 38420 7160
rect 38956 8548 38996 8588
rect 38764 8380 38804 8420
rect 38572 7792 38612 7832
rect 39148 8632 39188 8672
rect 39052 8380 39092 8420
rect 39148 7708 39188 7748
rect 38956 7540 38996 7580
rect 38668 7120 38708 7160
rect 39052 7204 39092 7244
rect 39244 7204 39284 7244
rect 39148 7120 39188 7160
rect 39148 6868 39188 6908
rect 39340 7120 39380 7160
rect 38476 6112 38516 6152
rect 38380 6028 38420 6068
rect 38572 5860 38612 5900
rect 38380 4768 38420 4808
rect 38860 5104 38900 5144
rect 38764 5020 38804 5060
rect 38572 4684 38612 4724
rect 38284 3256 38324 3296
rect 37996 2836 38036 2876
rect 38380 2584 38420 2624
rect 37900 1912 37940 1952
rect 38380 2416 38420 2456
rect 38572 2668 38612 2708
rect 38476 2248 38516 2288
rect 38476 2080 38516 2120
rect 38572 1324 38612 1364
rect 39052 5020 39092 5060
rect 38956 4684 38996 4724
rect 39244 4516 39284 4556
rect 39628 8464 39668 8504
rect 39820 7960 39860 8000
rect 39820 7120 39860 7160
rect 39532 5944 39572 5984
rect 39820 5776 39860 5816
rect 39628 4516 39668 4556
rect 39148 2500 39188 2540
rect 39628 3508 39668 3548
rect 39916 5440 39956 5480
rect 40492 9388 40532 9428
rect 40780 8884 40820 8924
rect 40396 8632 40436 8672
rect 40396 7540 40436 7580
rect 40108 6616 40148 6656
rect 40684 7372 40724 7412
rect 40492 6952 40532 6992
rect 40588 6616 40628 6656
rect 40876 8716 40916 8756
rect 41068 9808 41108 9848
rect 41260 9556 41300 9596
rect 41452 9472 41492 9512
rect 41356 9136 41396 9176
rect 41164 8968 41204 9008
rect 41068 8128 41108 8168
rect 41260 8716 41300 8756
rect 41164 7708 41204 7748
rect 40972 7372 41012 7412
rect 40876 7036 40916 7076
rect 40876 6532 40916 6572
rect 41068 6784 41108 6824
rect 41068 6448 41108 6488
rect 40972 5944 41012 5984
rect 40780 5860 40820 5900
rect 40204 5776 40244 5816
rect 41068 5776 41108 5816
rect 40012 4348 40052 4388
rect 39820 3928 39860 3968
rect 39916 3844 39956 3884
rect 39340 2752 39380 2792
rect 39244 1996 39284 2036
rect 39052 1744 39092 1784
rect 39244 1744 39284 1784
rect 38380 1240 38420 1280
rect 38860 1072 38900 1112
rect 39532 2584 39572 2624
rect 39724 2668 39764 2708
rect 40108 3508 40148 3548
rect 39916 3172 39956 3212
rect 39820 2416 39860 2456
rect 39820 1912 39860 1952
rect 39916 1408 39956 1448
rect 39628 1324 39668 1364
rect 40492 5524 40532 5564
rect 40684 5440 40724 5480
rect 40876 5356 40916 5396
rect 41068 5104 41108 5144
rect 40876 4852 40916 4892
rect 40492 4768 40532 4808
rect 40684 4768 40724 4808
rect 41260 7456 41300 7496
rect 41260 6868 41300 6908
rect 41260 6364 41300 6404
rect 41260 5692 41300 5732
rect 41452 8464 41492 8504
rect 41452 7876 41492 7916
rect 41644 7792 41684 7832
rect 41452 7120 41492 7160
rect 41452 6196 41492 6236
rect 41452 5860 41492 5900
rect 41260 4600 41300 4640
rect 40876 4432 40916 4472
rect 41068 4432 41108 4472
rect 40396 4348 40436 4388
rect 40300 4264 40340 4304
rect 40492 4180 40532 4220
rect 41452 4096 41492 4136
rect 41068 3760 41108 3800
rect 41260 3676 41300 3716
rect 40684 3424 40724 3464
rect 40876 3340 40916 3380
rect 40204 2752 40244 2792
rect 40300 2416 40340 2456
rect 40108 1828 40148 1868
rect 40108 1324 40148 1364
rect 40012 1072 40052 1112
rect 39436 904 39476 944
rect 36844 820 36884 860
rect 36652 652 36692 692
rect 34540 484 34580 524
rect 33964 400 34004 440
rect 40780 3172 40820 3212
rect 41452 3172 41492 3212
rect 40588 2584 40628 2624
rect 40684 1660 40724 1700
rect 40588 1072 40628 1112
rect 41644 2752 41684 2792
rect 41452 2668 41492 2708
rect 40876 2500 40916 2540
rect 41260 2416 41300 2456
rect 41644 2080 41684 2120
rect 41068 1660 41108 1700
rect 40972 1240 41012 1280
rect 41452 1324 41492 1364
rect 40876 1156 40916 1196
rect 41260 820 41300 860
rect 40780 736 40820 776
rect 40396 400 40436 440
rect 40300 64 40340 104
rect 41452 64 41492 104
<< metal3 >>
rect 16771 10648 16780 10688
rect 16820 10648 32236 10688
rect 32276 10648 32285 10688
rect 25987 10564 25996 10604
rect 26036 10564 36556 10604
rect 36596 10564 36605 10604
rect 0 10520 80 10540
rect 42928 10520 43008 10540
rect 0 10480 12844 10520
rect 12884 10480 12893 10520
rect 27139 10480 27148 10520
rect 27188 10480 36940 10520
rect 36980 10480 36989 10520
rect 40963 10480 40972 10520
rect 41012 10480 43008 10520
rect 0 10460 80 10480
rect 42928 10460 43008 10480
rect 23683 10396 23692 10436
rect 23732 10396 32332 10436
rect 32372 10396 32381 10436
rect 0 10184 80 10204
rect 451 10184 509 10185
rect 42928 10184 43008 10204
rect 0 10144 460 10184
rect 500 10144 509 10184
rect 1411 10144 1420 10184
rect 1460 10144 8716 10184
rect 8756 10144 8765 10184
rect 40675 10144 40684 10184
rect 40724 10144 43008 10184
rect 0 10124 80 10144
rect 451 10143 509 10144
rect 42928 10124 43008 10144
rect 5635 10060 5644 10100
rect 5684 10060 11020 10100
rect 11060 10060 11069 10100
rect 34051 9892 34060 9932
rect 34100 9892 39340 9932
rect 39380 9892 39389 9932
rect 0 9848 80 9868
rect 42928 9848 43008 9868
rect 0 9808 2540 9848
rect 4919 9808 4928 9848
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 5296 9808 5305 9848
rect 20039 9808 20048 9848
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20416 9808 20425 9848
rect 28291 9808 28300 9848
rect 28340 9808 34540 9848
rect 34580 9808 34589 9848
rect 35159 9808 35168 9848
rect 35208 9808 35250 9848
rect 35290 9808 35332 9848
rect 35372 9808 35414 9848
rect 35454 9808 35496 9848
rect 35536 9808 35545 9848
rect 41059 9808 41068 9848
rect 41108 9808 43008 9848
rect 0 9788 80 9808
rect 2500 9764 2540 9808
rect 42928 9788 43008 9808
rect 2500 9724 9004 9764
rect 9044 9724 11500 9764
rect 11540 9724 11549 9764
rect 27907 9724 27916 9764
rect 27956 9724 40876 9764
rect 40916 9724 40925 9764
rect 2179 9640 2188 9680
rect 2228 9640 4492 9680
rect 4532 9640 4541 9680
rect 8611 9640 8620 9680
rect 8660 9640 13420 9680
rect 13460 9640 13469 9680
rect 21475 9640 21484 9680
rect 21524 9640 29260 9680
rect 29300 9640 29309 9680
rect 29443 9640 29452 9680
rect 29492 9640 37324 9680
rect 37364 9640 37373 9680
rect 38659 9640 38668 9680
rect 38708 9640 39724 9680
rect 39764 9640 39773 9680
rect 1699 9556 1708 9596
rect 1748 9556 2476 9596
rect 2516 9556 3820 9596
rect 3860 9556 3869 9596
rect 19372 9556 21004 9596
rect 21044 9556 22636 9596
rect 22676 9556 22685 9596
rect 26275 9556 26284 9596
rect 26324 9556 29548 9596
rect 29588 9556 41260 9596
rect 41300 9556 41309 9596
rect 0 9512 80 9532
rect 14755 9512 14813 9513
rect 19372 9512 19412 9556
rect 19747 9512 19805 9513
rect 32899 9512 32957 9513
rect 42928 9512 43008 9532
rect 0 9472 1420 9512
rect 1460 9472 1469 9512
rect 1603 9472 1612 9512
rect 1652 9472 2956 9512
rect 2996 9472 3005 9512
rect 3235 9472 3244 9512
rect 3284 9472 3628 9512
rect 3668 9472 5452 9512
rect 5492 9472 5501 9512
rect 7651 9472 7660 9512
rect 7700 9472 8716 9512
rect 8756 9472 8765 9512
rect 10723 9472 10732 9512
rect 10772 9472 11116 9512
rect 11156 9472 12748 9512
rect 12788 9472 14284 9512
rect 14324 9472 14333 9512
rect 14670 9472 14764 9512
rect 14804 9472 14813 9512
rect 16003 9472 16012 9512
rect 16052 9472 17452 9512
rect 17492 9472 17644 9512
rect 17684 9472 19372 9512
rect 19412 9472 19421 9512
rect 19662 9472 19756 9512
rect 19796 9472 19805 9512
rect 24451 9472 24460 9512
rect 24500 9472 25036 9512
rect 25076 9472 26668 9512
rect 26708 9472 26717 9512
rect 32814 9472 32908 9512
rect 32948 9472 32957 9512
rect 41443 9472 41452 9512
rect 41492 9472 43008 9512
rect 0 9452 80 9472
rect 14755 9471 14813 9472
rect 19747 9471 19805 9472
rect 32899 9471 32957 9472
rect 32908 9428 32948 9471
rect 42928 9452 43008 9472
rect 40483 9428 40541 9429
rect 4771 9388 4780 9428
rect 4820 9388 5068 9428
rect 5108 9388 5117 9428
rect 6691 9388 6700 9428
rect 6740 9388 16396 9428
rect 16436 9388 23212 9428
rect 23252 9388 32948 9428
rect 36355 9388 36364 9428
rect 36404 9388 38188 9428
rect 38228 9388 38237 9428
rect 40398 9388 40492 9428
rect 40532 9388 40541 9428
rect 40483 9387 40541 9388
rect 5251 9304 5260 9344
rect 5300 9304 7180 9344
rect 7220 9304 8332 9344
rect 8372 9304 8381 9344
rect 9859 9304 9868 9344
rect 9908 9304 18124 9344
rect 18164 9304 18173 9344
rect 29251 9304 29260 9344
rect 29300 9304 34924 9344
rect 34964 9304 37708 9344
rect 37748 9304 37757 9344
rect 4771 9220 4780 9260
rect 4820 9220 5356 9260
rect 5396 9220 5405 9260
rect 16195 9220 16204 9260
rect 16244 9220 16588 9260
rect 16628 9220 16637 9260
rect 33763 9220 33772 9260
rect 33812 9220 34348 9260
rect 34388 9220 34397 9260
rect 35875 9220 35884 9260
rect 35924 9220 36364 9260
rect 36404 9220 36413 9260
rect 0 9176 80 9196
rect 42928 9176 43008 9196
rect 0 9136 1228 9176
rect 1268 9136 1277 9176
rect 4195 9136 4204 9176
rect 4244 9136 8428 9176
rect 8468 9136 11116 9176
rect 11156 9136 14092 9176
rect 14132 9136 14141 9176
rect 19363 9136 19372 9176
rect 19412 9136 20180 9176
rect 41347 9136 41356 9176
rect 41396 9136 43008 9176
rect 0 9116 80 9136
rect 20140 9092 20180 9136
rect 42928 9116 43008 9136
rect 37123 9092 37181 9093
rect 3679 9052 3688 9092
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 4056 9052 4065 9092
rect 5443 9052 5452 9092
rect 5492 9052 7084 9092
rect 7124 9052 7372 9092
rect 7412 9052 8812 9092
rect 8852 9052 10732 9092
rect 10772 9052 10781 9092
rect 18799 9052 18808 9092
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 19176 9052 19185 9092
rect 20140 9052 25036 9092
rect 25076 9052 27916 9092
rect 27956 9052 27965 9092
rect 33919 9052 33928 9092
rect 33968 9052 34010 9092
rect 34050 9052 34092 9092
rect 34132 9052 34174 9092
rect 34214 9052 34256 9092
rect 34296 9052 34305 9092
rect 37038 9052 37132 9092
rect 37172 9052 37181 9092
rect 37123 9051 37181 9052
rect 1324 8968 5836 9008
rect 5876 8968 21484 9008
rect 21524 8968 21533 9008
rect 25891 8968 25900 9008
rect 25940 8968 41164 9008
rect 41204 8968 41213 9008
rect 1324 8924 1364 8968
rect 1132 8884 1364 8924
rect 1411 8884 1420 8924
rect 1460 8884 2540 8924
rect 7459 8884 7468 8924
rect 7508 8884 13708 8924
rect 13748 8884 13757 8924
rect 14284 8884 30508 8924
rect 30548 8884 30557 8924
rect 30691 8884 30700 8924
rect 30740 8884 34540 8924
rect 34580 8884 34589 8924
rect 40771 8884 40780 8924
rect 40820 8884 41600 8924
rect 0 8840 80 8860
rect 1132 8840 1172 8884
rect 2500 8841 2540 8884
rect 2467 8840 2540 8841
rect 4003 8840 4061 8841
rect 0 8800 1172 8840
rect 2460 8800 2476 8840
rect 2516 8800 2540 8840
rect 3918 8800 4012 8840
rect 4052 8800 4061 8840
rect 0 8780 80 8800
rect 2467 8799 2525 8800
rect 4003 8799 4061 8800
rect 4195 8840 4253 8841
rect 4195 8800 4204 8840
rect 4244 8800 4338 8840
rect 8800 8800 9716 8840
rect 10339 8800 10348 8840
rect 10388 8800 12748 8840
rect 12788 8800 12797 8840
rect 12931 8800 12940 8840
rect 12980 8800 14188 8840
rect 14228 8800 14237 8840
rect 4195 8799 4253 8800
rect 8131 8756 8189 8757
rect 8800 8756 8840 8800
rect 9571 8756 9629 8757
rect 1219 8716 1228 8756
rect 1268 8716 2540 8756
rect 1315 8672 1373 8673
rect 2371 8672 2429 8673
rect 1230 8632 1324 8672
rect 1364 8632 1373 8672
rect 2286 8632 2380 8672
rect 2420 8632 2429 8672
rect 2500 8672 2540 8716
rect 8131 8716 8140 8756
rect 8180 8716 8840 8756
rect 9475 8716 9484 8756
rect 9524 8716 9580 8756
rect 9620 8716 9629 8756
rect 9676 8756 9716 8800
rect 14284 8756 14324 8884
rect 41560 8840 41600 8884
rect 42928 8840 43008 8860
rect 16291 8800 16300 8840
rect 16340 8800 17932 8840
rect 17972 8800 17981 8840
rect 18115 8800 18124 8840
rect 18164 8800 21292 8840
rect 21332 8800 21341 8840
rect 22723 8800 22732 8840
rect 22772 8800 23020 8840
rect 23060 8800 23069 8840
rect 30883 8800 30892 8840
rect 30932 8800 32428 8840
rect 32468 8800 32477 8840
rect 41560 8800 43008 8840
rect 42928 8780 43008 8800
rect 41251 8756 41309 8757
rect 9676 8716 11020 8756
rect 11060 8716 11069 8756
rect 11500 8716 12076 8756
rect 12116 8716 12460 8756
rect 12500 8716 12509 8756
rect 12643 8716 12652 8756
rect 12692 8716 13612 8756
rect 13652 8716 14324 8756
rect 19747 8716 19756 8756
rect 19796 8716 20044 8756
rect 20084 8716 22540 8756
rect 22580 8716 22589 8756
rect 25228 8716 27340 8756
rect 27380 8716 27389 8756
rect 29731 8716 29740 8756
rect 29780 8716 31852 8756
rect 31892 8716 36652 8756
rect 36692 8716 36701 8756
rect 37780 8716 40876 8756
rect 40916 8716 40925 8756
rect 41166 8716 41260 8756
rect 41300 8716 41309 8756
rect 8131 8715 8189 8716
rect 9571 8715 9629 8716
rect 6115 8672 6173 8673
rect 7747 8672 7805 8673
rect 9763 8672 9821 8673
rect 11500 8672 11540 8716
rect 16195 8672 16253 8673
rect 21283 8672 21341 8673
rect 25228 8672 25268 8716
rect 33667 8672 33725 8673
rect 37780 8672 37820 8716
rect 41251 8715 41309 8716
rect 38371 8672 38429 8673
rect 2500 8632 6124 8672
rect 6164 8632 6173 8672
rect 6691 8632 6700 8672
rect 6740 8632 6749 8672
rect 7662 8632 7756 8672
rect 7796 8632 7805 8672
rect 9571 8632 9580 8672
rect 9620 8632 9629 8672
rect 9763 8632 9772 8672
rect 9812 8632 9906 8672
rect 10060 8632 10444 8672
rect 10484 8632 11540 8672
rect 11587 8632 11596 8672
rect 11636 8632 11884 8672
rect 11924 8632 11933 8672
rect 13027 8632 13036 8672
rect 13076 8632 13516 8672
rect 13556 8632 13900 8672
rect 13940 8632 13949 8672
rect 14467 8632 14476 8672
rect 14516 8632 15436 8672
rect 15476 8632 15485 8672
rect 16110 8632 16204 8672
rect 16244 8632 16253 8672
rect 18019 8632 18028 8672
rect 18068 8632 18077 8672
rect 21198 8632 21292 8672
rect 21332 8632 21341 8672
rect 1315 8631 1373 8632
rect 2371 8631 2429 8632
rect 6115 8631 6173 8632
rect 6700 8588 6740 8632
rect 7747 8631 7805 8632
rect 9580 8588 9620 8632
rect 9763 8631 9821 8632
rect 10060 8588 10100 8632
rect 16195 8631 16253 8632
rect 1036 8548 6740 8588
rect 8803 8548 8812 8588
rect 8852 8548 9004 8588
rect 9044 8548 9053 8588
rect 9580 8548 10100 8588
rect 10147 8548 10156 8588
rect 10196 8548 10540 8588
rect 10580 8548 10589 8588
rect 11011 8548 11020 8588
rect 11060 8548 13172 8588
rect 13219 8548 13228 8588
rect 13268 8548 15052 8588
rect 15092 8548 16108 8588
rect 16148 8548 16157 8588
rect 0 8504 80 8524
rect 1036 8504 1076 8548
rect 0 8464 1076 8504
rect 2851 8464 2860 8504
rect 2900 8464 4972 8504
rect 5012 8464 5021 8504
rect 5155 8464 5164 8504
rect 5204 8464 6700 8504
rect 6740 8464 6749 8504
rect 6979 8464 6988 8504
rect 7028 8464 7372 8504
rect 7412 8464 7421 8504
rect 8611 8464 8620 8504
rect 8660 8464 10636 8504
rect 10676 8464 12652 8504
rect 12692 8464 12701 8504
rect 0 8444 80 8464
rect 4387 8420 4445 8421
rect 13132 8420 13172 8548
rect 13612 8504 13652 8548
rect 13603 8464 13612 8504
rect 13652 8464 13661 8504
rect 14083 8464 14092 8504
rect 14132 8464 14572 8504
rect 14612 8464 14621 8504
rect 2755 8380 2764 8420
rect 2804 8380 3148 8420
rect 3188 8380 3197 8420
rect 3619 8380 3628 8420
rect 3668 8380 4396 8420
rect 4436 8380 7276 8420
rect 7316 8380 7325 8420
rect 9763 8380 9772 8420
rect 9812 8380 10060 8420
rect 10100 8380 10109 8420
rect 13132 8380 13996 8420
rect 14036 8380 14045 8420
rect 4387 8379 4445 8380
rect 4195 8336 4253 8337
rect 18028 8336 18068 8632
rect 21283 8631 21341 8632
rect 22732 8632 25228 8672
rect 25268 8632 25277 8672
rect 25603 8632 25612 8672
rect 25652 8632 25661 8672
rect 28771 8632 28780 8672
rect 28820 8632 30220 8672
rect 30260 8632 32812 8672
rect 32852 8632 32861 8672
rect 33667 8632 33676 8672
rect 33716 8632 37820 8672
rect 38286 8632 38380 8672
rect 38420 8632 39148 8672
rect 39188 8632 39197 8672
rect 40387 8632 40396 8672
rect 40436 8632 40445 8672
rect 22732 8588 22772 8632
rect 25612 8588 25652 8632
rect 33667 8631 33725 8632
rect 38371 8631 38429 8632
rect 40396 8588 40436 8632
rect 18499 8548 18508 8588
rect 18548 8548 22772 8588
rect 22828 8548 25652 8588
rect 26179 8548 26188 8588
rect 26228 8548 33964 8588
rect 34004 8548 34013 8588
rect 34435 8548 34444 8588
rect 34484 8548 38956 8588
rect 38996 8548 40436 8588
rect 22828 8504 22868 8548
rect 33964 8504 34004 8548
rect 42928 8504 43008 8524
rect 18403 8464 18412 8504
rect 18452 8464 22868 8504
rect 24739 8464 24748 8504
rect 24788 8464 25612 8504
rect 25652 8464 25661 8504
rect 33964 8464 39628 8504
rect 39668 8464 39677 8504
rect 41443 8464 41452 8504
rect 41492 8464 43008 8504
rect 42928 8444 43008 8464
rect 18211 8380 18220 8420
rect 18260 8380 23596 8420
rect 23636 8380 25708 8420
rect 25748 8380 26476 8420
rect 26516 8380 27628 8420
rect 27668 8380 27916 8420
rect 27956 8380 27965 8420
rect 36547 8380 36556 8420
rect 36596 8380 36748 8420
rect 36788 8380 36797 8420
rect 38755 8380 38764 8420
rect 38804 8380 39052 8420
rect 39092 8380 39101 8420
rect 4099 8296 4108 8336
rect 4148 8296 4204 8336
rect 4244 8296 4253 8336
rect 4919 8296 4928 8336
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 5296 8296 5305 8336
rect 8800 8296 9868 8336
rect 9908 8296 9917 8336
rect 10060 8296 10348 8336
rect 10388 8296 10397 8336
rect 11587 8296 11596 8336
rect 11636 8296 12556 8336
rect 12596 8296 12940 8336
rect 12980 8296 13132 8336
rect 13172 8296 18068 8336
rect 20039 8296 20048 8336
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20416 8296 20425 8336
rect 24067 8296 24076 8336
rect 24116 8296 25516 8336
rect 25556 8296 26188 8336
rect 26228 8296 26237 8336
rect 35159 8296 35168 8336
rect 35208 8296 35250 8336
rect 35290 8296 35332 8336
rect 35372 8296 35414 8336
rect 35454 8296 35496 8336
rect 35536 8296 35545 8336
rect 4195 8295 4253 8296
rect 8800 8252 8840 8296
rect 10060 8252 10100 8296
rect 2500 8212 8840 8252
rect 10051 8212 10060 8252
rect 10100 8212 10109 8252
rect 17635 8212 17644 8252
rect 17684 8212 23500 8252
rect 23540 8212 23549 8252
rect 0 8168 80 8188
rect 2500 8168 2540 8212
rect 42928 8168 43008 8188
rect 0 8128 2540 8168
rect 3043 8128 3052 8168
rect 3092 8128 3340 8168
rect 3380 8128 4684 8168
rect 4724 8128 4733 8168
rect 8131 8128 8140 8168
rect 8180 8128 8189 8168
rect 8899 8128 8908 8168
rect 8948 8128 9484 8168
rect 9524 8128 9533 8168
rect 9667 8128 9676 8168
rect 9716 8128 10156 8168
rect 10196 8128 10205 8168
rect 13411 8128 13420 8168
rect 13460 8128 14284 8168
rect 14324 8128 15340 8168
rect 15380 8128 15389 8168
rect 18307 8128 18316 8168
rect 18356 8128 20524 8168
rect 20564 8128 20573 8168
rect 31075 8128 31084 8168
rect 31124 8128 31564 8168
rect 31604 8128 31613 8168
rect 36355 8128 36364 8168
rect 36404 8128 36748 8168
rect 36788 8128 36797 8168
rect 41059 8128 41068 8168
rect 41108 8128 43008 8168
rect 0 8108 80 8128
rect 8140 8084 8180 8128
rect 42928 8108 43008 8128
rect 8140 8044 9388 8084
rect 9428 8044 9437 8084
rect 9484 8044 10636 8084
rect 10676 8044 20812 8084
rect 20852 8044 26284 8084
rect 26324 8044 26333 8084
rect 28579 8044 28588 8084
rect 28628 8044 29356 8084
rect 29396 8044 29405 8084
rect 30211 8044 30220 8084
rect 30260 8044 31852 8084
rect 31892 8044 32428 8084
rect 32468 8044 34444 8084
rect 34484 8044 34493 8084
rect 36931 8044 36940 8084
rect 36980 8044 37420 8084
rect 37460 8044 37469 8084
rect 4483 8000 4541 8001
rect 8707 8000 8765 8001
rect 9484 8000 9524 8044
rect 12067 8000 12125 8001
rect 2755 7960 2764 8000
rect 2804 7960 3244 8000
rect 3284 7960 3293 8000
rect 4398 7960 4492 8000
rect 4532 7960 4541 8000
rect 7651 7960 7660 8000
rect 7700 7960 8524 8000
rect 8564 7960 8573 8000
rect 8707 7960 8716 8000
rect 8756 7960 9524 8000
rect 9955 7960 9964 8000
rect 10004 7960 11404 8000
rect 11444 7960 11453 8000
rect 11982 7960 12076 8000
rect 12116 7960 12125 8000
rect 4483 7959 4541 7960
rect 8707 7959 8765 7960
rect 12067 7959 12125 7960
rect 13699 8000 13757 8001
rect 33667 8000 33725 8001
rect 13699 7960 13708 8000
rect 13748 7960 13804 8000
rect 13844 7960 13853 8000
rect 14275 7960 14284 8000
rect 14324 7960 15436 8000
rect 15476 7960 15485 8000
rect 17347 7960 17356 8000
rect 17396 7960 19756 8000
rect 19796 7960 19805 8000
rect 24835 7960 24844 8000
rect 24884 7960 31564 8000
rect 31604 7960 31613 8000
rect 33582 7960 33676 8000
rect 33716 7960 33725 8000
rect 35107 7960 35116 8000
rect 35156 7960 35596 8000
rect 35636 7960 36268 8000
rect 36308 7960 36317 8000
rect 36364 7960 38092 8000
rect 38132 7960 39820 8000
rect 39860 7960 39869 8000
rect 13699 7959 13757 7960
rect 33667 7959 33725 7960
rect 18499 7916 18557 7917
rect 36364 7916 36404 7960
rect 36547 7916 36605 7917
rect 2179 7876 2188 7916
rect 2228 7876 3052 7916
rect 3092 7876 3101 7916
rect 4579 7876 4588 7916
rect 4628 7876 5260 7916
rect 5300 7876 8620 7916
rect 8660 7876 8669 7916
rect 13891 7876 13900 7916
rect 13940 7876 16012 7916
rect 16052 7876 16061 7916
rect 18414 7876 18508 7916
rect 18548 7876 18557 7916
rect 19651 7876 19660 7916
rect 19700 7876 20428 7916
rect 20468 7876 20477 7916
rect 28483 7876 28492 7916
rect 28532 7876 28780 7916
rect 28820 7876 30220 7916
rect 30260 7876 30269 7916
rect 31747 7876 31756 7916
rect 31796 7876 31805 7916
rect 32803 7876 32812 7916
rect 32852 7876 36364 7916
rect 36404 7876 36413 7916
rect 36547 7876 36556 7916
rect 36596 7876 41452 7916
rect 41492 7876 41501 7916
rect 18499 7875 18557 7876
rect 0 7832 80 7852
rect 1219 7832 1277 7833
rect 4675 7832 4733 7833
rect 8131 7832 8189 7833
rect 23491 7832 23549 7833
rect 31756 7832 31796 7876
rect 36547 7875 36605 7876
rect 42928 7832 43008 7852
rect 0 7792 1228 7832
rect 1268 7792 1277 7832
rect 4195 7792 4204 7832
rect 4244 7792 4684 7832
rect 4724 7792 5356 7832
rect 5396 7792 8140 7832
rect 8180 7792 8189 7832
rect 9667 7792 9676 7832
rect 9716 7792 14380 7832
rect 14420 7792 14429 7832
rect 23406 7792 23500 7832
rect 23540 7792 28972 7832
rect 29012 7792 29932 7832
rect 29972 7792 29981 7832
rect 31756 7792 38572 7832
rect 38612 7792 38621 7832
rect 41635 7792 41644 7832
rect 41684 7792 43008 7832
rect 0 7772 80 7792
rect 1219 7791 1277 7792
rect 4675 7791 4733 7792
rect 8131 7791 8189 7792
rect 23491 7791 23549 7792
rect 42928 7772 43008 7792
rect 11779 7748 11837 7749
rect 16099 7748 16157 7749
rect 9676 7708 11596 7748
rect 11636 7708 11645 7748
rect 11694 7708 11788 7748
rect 11828 7708 16108 7748
rect 16148 7708 16157 7748
rect 30019 7708 30028 7748
rect 30068 7708 30412 7748
rect 30452 7708 30461 7748
rect 32131 7708 32140 7748
rect 32180 7708 32660 7748
rect 32707 7708 32716 7748
rect 32756 7708 34732 7748
rect 34772 7708 34781 7748
rect 35491 7708 35500 7748
rect 35540 7708 36940 7748
rect 36980 7708 36989 7748
rect 39139 7708 39148 7748
rect 39188 7708 41164 7748
rect 41204 7708 41213 7748
rect 9676 7664 9716 7708
rect 11779 7707 11837 7708
rect 16099 7707 16157 7708
rect 10147 7664 10205 7665
rect 32620 7664 32660 7708
rect 1603 7624 1612 7664
rect 1652 7624 4780 7664
rect 4820 7624 4829 7664
rect 6403 7624 6412 7664
rect 6452 7624 9620 7664
rect 9667 7624 9676 7664
rect 9716 7624 9725 7664
rect 9772 7624 10156 7664
rect 10196 7624 32180 7664
rect 32620 7624 37804 7664
rect 37844 7624 37853 7664
rect 1795 7580 1853 7581
rect 9580 7580 9620 7624
rect 9772 7580 9812 7624
rect 10147 7623 10205 7624
rect 25795 7580 25853 7581
rect 32140 7580 32180 7624
rect 1710 7540 1804 7580
rect 1844 7540 1853 7580
rect 3679 7540 3688 7580
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 4056 7540 4065 7580
rect 6787 7540 6796 7580
rect 6836 7540 7756 7580
rect 7796 7540 7805 7580
rect 9580 7540 9812 7580
rect 10243 7540 10252 7580
rect 10292 7540 11596 7580
rect 11636 7540 11645 7580
rect 14179 7540 14188 7580
rect 14228 7540 14476 7580
rect 14516 7540 14525 7580
rect 18799 7540 18808 7580
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 19176 7540 19185 7580
rect 20995 7540 21004 7580
rect 21044 7540 22060 7580
rect 22100 7540 22109 7580
rect 22531 7540 22540 7580
rect 22580 7540 24364 7580
rect 24404 7540 24652 7580
rect 24692 7540 24701 7580
rect 25795 7540 25804 7580
rect 25844 7540 27052 7580
rect 27092 7540 27101 7580
rect 30691 7540 30700 7580
rect 30740 7540 32044 7580
rect 32084 7540 32093 7580
rect 32140 7540 32812 7580
rect 32852 7540 32861 7580
rect 33919 7540 33928 7580
rect 33968 7540 34010 7580
rect 34050 7540 34092 7580
rect 34132 7540 34174 7580
rect 34214 7540 34256 7580
rect 34296 7540 34305 7580
rect 38947 7540 38956 7580
rect 38996 7540 40396 7580
rect 40436 7540 40445 7580
rect 1795 7539 1853 7540
rect 25795 7539 25853 7540
rect 0 7496 80 7516
rect 42928 7496 43008 7516
rect 0 7456 10924 7496
rect 10964 7456 10973 7496
rect 11491 7456 11500 7496
rect 11540 7456 19372 7496
rect 19412 7456 19421 7496
rect 22435 7456 22444 7496
rect 22484 7456 22636 7496
rect 22676 7456 22685 7496
rect 30403 7456 30412 7496
rect 30452 7456 30604 7496
rect 30644 7456 33196 7496
rect 33236 7456 33245 7496
rect 41251 7456 41260 7496
rect 41300 7456 43008 7496
rect 0 7436 80 7456
rect 42928 7436 43008 7456
rect 1987 7372 1996 7412
rect 2036 7372 3532 7412
rect 3572 7372 3581 7412
rect 7843 7372 7852 7412
rect 7892 7372 9004 7412
rect 9044 7372 9053 7412
rect 11875 7372 11884 7412
rect 11924 7372 12364 7412
rect 12404 7372 13652 7412
rect 13987 7372 13996 7412
rect 14036 7372 14380 7412
rect 14420 7372 14429 7412
rect 16099 7372 16108 7412
rect 16148 7372 20180 7412
rect 40675 7372 40684 7412
rect 40724 7372 40972 7412
rect 41012 7372 41021 7412
rect 13612 7328 13652 7372
rect 20140 7328 20180 7372
rect 2947 7288 2956 7328
rect 2996 7288 4204 7328
rect 4244 7288 4972 7328
rect 5012 7288 5021 7328
rect 7267 7288 7276 7328
rect 7316 7288 8044 7328
rect 8084 7288 8093 7328
rect 8611 7288 8620 7328
rect 8660 7288 13516 7328
rect 13556 7288 13565 7328
rect 13612 7288 14668 7328
rect 14708 7288 14956 7328
rect 14996 7288 18796 7328
rect 18836 7288 18845 7328
rect 20140 7288 37708 7328
rect 37748 7288 37757 7328
rect 3235 7204 3244 7244
rect 3284 7204 4492 7244
rect 4532 7204 4541 7244
rect 11491 7204 11500 7244
rect 11540 7204 16684 7244
rect 16724 7204 16733 7244
rect 24835 7204 24844 7244
rect 24884 7204 25228 7244
rect 25268 7204 25277 7244
rect 25795 7204 25804 7244
rect 25844 7204 26380 7244
rect 26420 7204 27148 7244
rect 27188 7204 28204 7244
rect 28244 7204 28780 7244
rect 28820 7204 28829 7244
rect 28960 7204 30412 7244
rect 30452 7204 30461 7244
rect 31747 7204 31756 7244
rect 31796 7204 32140 7244
rect 32180 7204 32189 7244
rect 34339 7204 34348 7244
rect 34388 7204 35692 7244
rect 35732 7204 36460 7244
rect 36500 7204 36509 7244
rect 36835 7204 36844 7244
rect 36884 7204 37516 7244
rect 37556 7204 37565 7244
rect 37780 7204 39052 7244
rect 39092 7204 39244 7244
rect 39284 7204 39293 7244
rect 0 7160 80 7180
rect 4387 7160 4445 7161
rect 14467 7160 14525 7161
rect 17731 7160 17789 7161
rect 21379 7160 21437 7161
rect 28960 7160 29000 7204
rect 0 7120 1420 7160
rect 1460 7120 2476 7160
rect 2516 7120 2525 7160
rect 3907 7120 3916 7160
rect 3956 7120 4396 7160
rect 4436 7120 4445 7160
rect 9571 7120 9580 7160
rect 9620 7120 13708 7160
rect 13748 7120 13757 7160
rect 14382 7120 14476 7160
rect 14516 7120 14525 7160
rect 17646 7120 17740 7160
rect 17780 7120 17789 7160
rect 18979 7120 18988 7160
rect 19028 7120 20620 7160
rect 20660 7120 21004 7160
rect 21044 7120 21053 7160
rect 21360 7120 21388 7160
rect 21428 7120 21484 7160
rect 21524 7120 29000 7160
rect 30019 7160 30077 7161
rect 32899 7160 32957 7161
rect 37780 7160 37820 7204
rect 42928 7160 43008 7180
rect 30019 7120 30028 7160
rect 30068 7120 31084 7160
rect 31124 7120 31133 7160
rect 32814 7120 32908 7160
rect 32948 7120 33292 7160
rect 33332 7120 33341 7160
rect 35971 7120 35980 7160
rect 36020 7120 37820 7160
rect 38371 7120 38380 7160
rect 38420 7120 38668 7160
rect 38708 7120 38717 7160
rect 39139 7120 39148 7160
rect 39188 7120 39340 7160
rect 39380 7120 39820 7160
rect 39860 7120 39869 7160
rect 41443 7120 41452 7160
rect 41492 7120 43008 7160
rect 0 7100 80 7120
rect 4387 7119 4445 7120
rect 14467 7119 14525 7120
rect 17731 7119 17789 7120
rect 21379 7119 21437 7120
rect 30019 7119 30077 7120
rect 32899 7119 32957 7120
rect 1507 7076 1565 7077
rect 4579 7076 4637 7077
rect 11875 7076 11933 7077
rect 17740 7076 17780 7119
rect 42928 7100 43008 7120
rect 27523 7076 27581 7077
rect 36547 7076 36605 7077
rect 1422 7036 1516 7076
rect 1556 7036 1565 7076
rect 4494 7036 4588 7076
rect 4628 7036 4637 7076
rect 4771 7036 4780 7076
rect 4820 7036 7564 7076
rect 7604 7036 11500 7076
rect 11540 7036 11549 7076
rect 11790 7036 11884 7076
rect 11924 7036 11933 7076
rect 15715 7036 15724 7076
rect 15764 7036 17452 7076
rect 17492 7036 17501 7076
rect 17740 7036 24940 7076
rect 24980 7036 24989 7076
rect 26851 7036 26860 7076
rect 26900 7036 27532 7076
rect 27572 7036 27581 7076
rect 30307 7036 30316 7076
rect 30356 7036 34444 7076
rect 34484 7036 34493 7076
rect 35587 7036 35596 7076
rect 35636 7036 36364 7076
rect 36404 7036 36413 7076
rect 36547 7036 36556 7076
rect 36596 7036 40876 7076
rect 40916 7036 40925 7076
rect 1507 7035 1565 7036
rect 4579 7035 4637 7036
rect 11875 7035 11933 7036
rect 27523 7035 27581 7036
rect 36547 7035 36605 7036
rect 13795 6992 13853 6993
rect 2500 6952 3340 6992
rect 3380 6952 4972 6992
rect 5012 6952 5021 6992
rect 6019 6952 6028 6992
rect 6068 6952 7180 6992
rect 7220 6952 7229 6992
rect 10915 6952 10924 6992
rect 10964 6952 11308 6992
rect 11348 6952 13804 6992
rect 13844 6952 13853 6992
rect 15619 6952 15628 6992
rect 15668 6952 16204 6992
rect 16244 6952 18028 6992
rect 18068 6952 18077 6992
rect 19180 6952 25516 6992
rect 25556 6952 25565 6992
rect 27811 6952 27820 6992
rect 27860 6952 31948 6992
rect 31988 6952 31997 6992
rect 33763 6952 33772 6992
rect 33812 6952 34348 6992
rect 34388 6952 34397 6992
rect 35011 6952 35020 6992
rect 35060 6952 35788 6992
rect 35828 6952 35837 6992
rect 2500 6908 2540 6952
rect 13795 6951 13853 6952
rect 1315 6868 1324 6908
rect 1364 6868 2540 6908
rect 3811 6868 3820 6908
rect 3860 6868 4684 6908
rect 4724 6868 8428 6908
rect 8468 6868 9676 6908
rect 9716 6868 9725 6908
rect 11875 6868 11884 6908
rect 11924 6868 16108 6908
rect 16148 6868 16157 6908
rect 0 6824 80 6844
rect 1795 6824 1853 6825
rect 3820 6824 3860 6868
rect 19180 6824 19220 6952
rect 21379 6868 21388 6908
rect 21428 6868 23212 6908
rect 23252 6868 27436 6908
rect 27476 6868 27485 6908
rect 29923 6868 29932 6908
rect 29972 6868 31852 6908
rect 31892 6868 31901 6908
rect 34435 6868 34444 6908
rect 34484 6868 35884 6908
rect 35924 6868 36940 6908
rect 36980 6868 36989 6908
rect 27148 6824 27188 6868
rect 37324 6824 37364 7036
rect 40387 6992 40445 6993
rect 40387 6952 40396 6992
rect 40436 6952 40492 6992
rect 40532 6952 40541 6992
rect 40387 6951 40445 6952
rect 37699 6868 37708 6908
rect 37748 6868 39148 6908
rect 39188 6868 41260 6908
rect 41300 6868 41309 6908
rect 42928 6824 43008 6844
rect 0 6784 1804 6824
rect 1844 6784 1853 6824
rect 1987 6784 1996 6824
rect 2036 6784 3860 6824
rect 4919 6784 4928 6824
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 5296 6784 5305 6824
rect 9091 6784 9100 6824
rect 9140 6784 9580 6824
rect 9620 6784 9629 6824
rect 11779 6784 11788 6824
rect 11828 6784 19180 6824
rect 19220 6784 19229 6824
rect 20039 6784 20048 6824
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20416 6784 20425 6824
rect 23596 6784 25804 6824
rect 25844 6784 25853 6824
rect 27139 6784 27148 6824
rect 27188 6784 27197 6824
rect 28960 6784 29836 6824
rect 29876 6784 33484 6824
rect 33524 6784 33533 6824
rect 35159 6784 35168 6824
rect 35208 6784 35250 6824
rect 35290 6784 35332 6824
rect 35372 6784 35414 6824
rect 35454 6784 35496 6824
rect 35536 6784 35545 6824
rect 36163 6784 36172 6824
rect 36212 6784 36252 6824
rect 37315 6784 37324 6824
rect 37364 6784 37373 6824
rect 41059 6784 41068 6824
rect 41108 6784 43008 6824
rect 0 6764 80 6784
rect 1795 6783 1853 6784
rect 23596 6740 23636 6784
rect 28960 6740 29000 6784
rect 36172 6740 36212 6784
rect 42928 6764 43008 6784
rect 2467 6700 2476 6740
rect 2516 6700 11884 6740
rect 11924 6700 11933 6740
rect 13123 6700 13132 6740
rect 13172 6700 13804 6740
rect 13844 6700 15052 6740
rect 15092 6700 23636 6740
rect 23683 6700 23692 6740
rect 23732 6700 25612 6740
rect 25652 6700 29000 6740
rect 29923 6700 29932 6740
rect 29972 6700 34252 6740
rect 34292 6700 34301 6740
rect 35980 6700 36652 6740
rect 36692 6700 37132 6740
rect 37172 6700 37181 6740
rect 20236 6656 20276 6700
rect 1507 6616 1516 6656
rect 1556 6616 2284 6656
rect 2324 6616 2860 6656
rect 2900 6616 3148 6656
rect 3188 6616 6508 6656
rect 6548 6616 6557 6656
rect 6988 6616 8140 6656
rect 8180 6616 8716 6656
rect 8756 6616 8765 6656
rect 9283 6616 9292 6656
rect 9332 6616 9341 6656
rect 13132 6616 15724 6656
rect 15764 6616 15773 6656
rect 16387 6616 16396 6656
rect 16436 6616 18220 6656
rect 18260 6616 18269 6656
rect 20227 6616 20236 6656
rect 20276 6616 20285 6656
rect 20995 6616 21004 6656
rect 21044 6616 22444 6656
rect 22484 6616 22493 6656
rect 24931 6616 24940 6656
rect 24980 6616 25900 6656
rect 25940 6616 25949 6656
rect 26188 6616 27436 6656
rect 27476 6616 29000 6656
rect 30019 6616 30028 6656
rect 30068 6616 34540 6656
rect 34580 6616 34589 6656
rect 6988 6572 7028 6616
rect 3427 6532 3436 6572
rect 3476 6532 3485 6572
rect 5731 6532 5740 6572
rect 5780 6532 6988 6572
rect 7028 6532 7037 6572
rect 7651 6532 7660 6572
rect 7700 6532 7709 6572
rect 0 6488 80 6508
rect 1699 6488 1757 6489
rect 0 6448 1708 6488
rect 1748 6448 1757 6488
rect 0 6428 80 6448
rect 1699 6447 1757 6448
rect 3436 6404 3476 6532
rect 4003 6488 4061 6489
rect 7660 6488 7700 6532
rect 8131 6488 8189 6489
rect 3907 6448 3916 6488
rect 3956 6448 4012 6488
rect 4052 6448 4061 6488
rect 4195 6448 4204 6488
rect 4244 6448 4588 6488
rect 4628 6448 5164 6488
rect 5204 6448 5213 6488
rect 5827 6448 5836 6488
rect 5876 6448 6700 6488
rect 6740 6448 7700 6488
rect 8046 6448 8140 6488
rect 8180 6448 8189 6488
rect 4003 6447 4061 6448
rect 5164 6404 5204 6448
rect 8131 6447 8189 6448
rect 3436 6364 4436 6404
rect 5164 6364 6124 6404
rect 6164 6364 6173 6404
rect 6403 6364 6412 6404
rect 6452 6364 6796 6404
rect 6836 6364 7276 6404
rect 7316 6364 8620 6404
rect 8660 6364 8669 6404
rect 1795 6320 1853 6321
rect 4396 6320 4436 6364
rect 9292 6320 9332 6616
rect 13132 6572 13172 6616
rect 17731 6572 17789 6573
rect 26188 6572 26228 6616
rect 28960 6572 29000 6616
rect 35980 6572 36020 6700
rect 36067 6616 36076 6656
rect 36116 6616 36364 6656
rect 36404 6616 36413 6656
rect 40099 6616 40108 6656
rect 40148 6616 40588 6656
rect 40628 6616 40637 6656
rect 13123 6532 13132 6572
rect 13172 6532 13181 6572
rect 15331 6532 15340 6572
rect 15380 6532 17740 6572
rect 17780 6532 17789 6572
rect 19843 6532 19852 6572
rect 19892 6532 23884 6572
rect 23924 6532 23933 6572
rect 24355 6532 24364 6572
rect 24404 6532 26188 6572
rect 26228 6532 26237 6572
rect 28960 6532 29204 6572
rect 31939 6532 31948 6572
rect 31988 6532 34060 6572
rect 34100 6532 36020 6572
rect 36163 6532 36172 6572
rect 36212 6532 36460 6572
rect 36500 6532 36509 6572
rect 36556 6532 40876 6572
rect 40916 6532 40925 6572
rect 17731 6531 17789 6532
rect 16099 6488 16157 6489
rect 23107 6488 23165 6489
rect 11491 6448 11500 6488
rect 11540 6448 12268 6488
rect 12308 6448 12317 6488
rect 16014 6448 16108 6488
rect 16148 6448 16157 6488
rect 17539 6448 17548 6488
rect 17588 6448 18124 6488
rect 18164 6448 18173 6488
rect 18787 6448 18796 6488
rect 18836 6448 21332 6488
rect 23022 6448 23116 6488
rect 23156 6448 26860 6488
rect 26900 6448 26909 6488
rect 16099 6447 16157 6448
rect 21292 6404 21332 6448
rect 23107 6447 23165 6448
rect 29164 6404 29204 6532
rect 30403 6488 30461 6489
rect 30691 6488 30749 6489
rect 35491 6488 35549 6489
rect 30318 6448 30412 6488
rect 30452 6448 30461 6488
rect 30606 6448 30700 6488
rect 30740 6448 30749 6488
rect 31747 6448 31756 6488
rect 31796 6448 32524 6488
rect 32564 6448 34924 6488
rect 34964 6448 34973 6488
rect 35406 6448 35500 6488
rect 35540 6448 35549 6488
rect 30403 6447 30461 6448
rect 30691 6447 30749 6448
rect 35491 6447 35549 6448
rect 33283 6404 33341 6405
rect 10819 6364 10828 6404
rect 10868 6364 11308 6404
rect 11348 6364 21004 6404
rect 21044 6364 21053 6404
rect 21283 6364 21292 6404
rect 21332 6364 25132 6404
rect 25172 6364 25181 6404
rect 29155 6364 29164 6404
rect 29204 6364 30796 6404
rect 30836 6364 31948 6404
rect 31988 6364 31997 6404
rect 33198 6364 33292 6404
rect 33332 6364 33341 6404
rect 33283 6363 33341 6364
rect 34723 6404 34781 6405
rect 36556 6404 36596 6532
rect 42928 6488 43008 6508
rect 41059 6448 41068 6488
rect 41108 6448 43008 6488
rect 42928 6428 43008 6448
rect 41251 6404 41309 6405
rect 34723 6364 34732 6404
rect 34772 6364 36596 6404
rect 37780 6364 37996 6404
rect 38036 6364 38045 6404
rect 41166 6364 41260 6404
rect 41300 6364 41309 6404
rect 34723 6363 34781 6364
rect 14947 6320 15005 6321
rect 37780 6320 37820 6364
rect 41251 6363 41309 6364
rect 1710 6280 1804 6320
rect 1844 6280 1853 6320
rect 3235 6280 3244 6320
rect 3284 6280 4300 6320
rect 4340 6280 4349 6320
rect 4396 6280 4820 6320
rect 4867 6280 4876 6320
rect 4916 6280 6028 6320
rect 6068 6280 6077 6320
rect 6499 6280 6508 6320
rect 6548 6280 7084 6320
rect 7124 6280 8812 6320
rect 8852 6280 9332 6320
rect 12163 6280 12172 6320
rect 12212 6280 13036 6320
rect 13076 6280 13085 6320
rect 14862 6280 14956 6320
rect 14996 6280 15005 6320
rect 17539 6280 17548 6320
rect 17588 6280 17932 6320
rect 17972 6280 17981 6320
rect 18307 6280 18316 6320
rect 18356 6280 18604 6320
rect 18644 6280 18653 6320
rect 21091 6280 21100 6320
rect 21140 6280 23596 6320
rect 23636 6280 23645 6320
rect 25219 6280 25228 6320
rect 25268 6280 26956 6320
rect 26996 6280 27005 6320
rect 33091 6280 33100 6320
rect 33140 6280 37820 6320
rect 1795 6279 1853 6280
rect 4780 6236 4820 6280
rect 14947 6279 15005 6280
rect 22627 6236 22685 6237
rect 1315 6196 1324 6236
rect 1364 6196 4396 6236
rect 4436 6196 4445 6236
rect 4780 6196 7220 6236
rect 7267 6196 7276 6236
rect 7316 6196 7660 6236
rect 7700 6196 8524 6236
rect 8564 6196 8573 6236
rect 8620 6196 11116 6236
rect 11156 6196 11165 6236
rect 13315 6196 13324 6236
rect 13364 6196 14476 6236
rect 14516 6196 14525 6236
rect 15427 6196 15436 6236
rect 15476 6196 15724 6236
rect 15764 6196 20180 6236
rect 0 6152 80 6172
rect 1507 6152 1565 6153
rect 7180 6152 7220 6196
rect 8620 6152 8660 6196
rect 0 6112 1516 6152
rect 1556 6112 1565 6152
rect 2275 6112 2284 6152
rect 2324 6112 6604 6152
rect 6644 6112 6892 6152
rect 6932 6112 6941 6152
rect 7180 6112 8660 6152
rect 8707 6112 8716 6152
rect 8756 6112 13708 6152
rect 13748 6112 13757 6152
rect 0 6092 80 6112
rect 1507 6111 1565 6112
rect 20140 6068 20180 6196
rect 22627 6196 22636 6236
rect 22676 6196 27148 6236
rect 27188 6196 27197 6236
rect 29443 6196 29452 6236
rect 29492 6196 33004 6236
rect 33044 6196 33580 6236
rect 33620 6196 33629 6236
rect 41443 6196 41452 6236
rect 41492 6196 41600 6236
rect 22627 6195 22685 6196
rect 41560 6152 41600 6196
rect 42928 6152 43008 6172
rect 31555 6112 31564 6152
rect 31604 6112 38476 6152
rect 38516 6112 38525 6152
rect 41560 6112 43008 6152
rect 42928 6092 43008 6112
rect 3679 6028 3688 6068
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 4056 6028 4065 6068
rect 7363 6028 7372 6068
rect 7412 6028 12748 6068
rect 12788 6028 12797 6068
rect 18799 6028 18808 6068
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 19176 6028 19185 6068
rect 20140 6028 28012 6068
rect 28052 6028 28061 6068
rect 31843 6028 31852 6068
rect 31892 6028 32140 6068
rect 32180 6028 32189 6068
rect 33919 6028 33928 6068
rect 33968 6028 34010 6068
rect 34050 6028 34092 6068
rect 34132 6028 34174 6068
rect 34214 6028 34256 6068
rect 34296 6028 34305 6068
rect 37603 6028 37612 6068
rect 37652 6028 38380 6068
rect 38420 6028 38429 6068
rect 21763 5984 21821 5985
rect 3139 5944 3148 5984
rect 3188 5944 3340 5984
rect 3380 5944 3389 5984
rect 8995 5944 9004 5984
rect 9044 5944 9292 5984
rect 9332 5944 9341 5984
rect 21678 5944 21772 5984
rect 21812 5944 29000 5984
rect 31939 5944 31948 5984
rect 31988 5944 39532 5984
rect 39572 5944 39581 5984
rect 39628 5944 40972 5984
rect 41012 5944 41021 5984
rect 21763 5943 21821 5944
rect 28960 5900 29000 5944
rect 6595 5860 6604 5900
rect 6644 5860 7468 5900
rect 7508 5860 7517 5900
rect 20140 5860 22252 5900
rect 22292 5860 22301 5900
rect 27619 5860 27628 5900
rect 27668 5860 28244 5900
rect 28960 5860 29452 5900
rect 29492 5860 29501 5900
rect 33379 5860 33388 5900
rect 33428 5860 34252 5900
rect 34292 5860 34301 5900
rect 36643 5860 36652 5900
rect 36692 5860 38572 5900
rect 38612 5860 38621 5900
rect 0 5816 80 5836
rect 2371 5816 2429 5817
rect 20140 5816 20180 5860
rect 28204 5816 28244 5860
rect 39628 5816 39668 5944
rect 40771 5860 40780 5900
rect 40820 5860 41452 5900
rect 41492 5860 41501 5900
rect 42928 5816 43008 5836
rect 0 5776 2380 5816
rect 2420 5776 2429 5816
rect 3331 5776 3340 5816
rect 3380 5776 4684 5816
rect 4724 5776 4733 5816
rect 5443 5776 5452 5816
rect 5492 5776 6316 5816
rect 6356 5776 7180 5816
rect 7220 5776 7229 5816
rect 9100 5776 9196 5816
rect 9236 5776 9245 5816
rect 12931 5776 12940 5816
rect 12980 5776 13228 5816
rect 13268 5776 13277 5816
rect 18595 5776 18604 5816
rect 18644 5776 20180 5816
rect 22252 5776 25420 5816
rect 25460 5776 28108 5816
rect 28148 5776 28157 5816
rect 28204 5776 29644 5816
rect 29684 5776 39668 5816
rect 39811 5776 39820 5816
rect 39860 5776 40204 5816
rect 40244 5776 40253 5816
rect 41059 5776 41068 5816
rect 41108 5776 43008 5816
rect 0 5756 80 5776
rect 2371 5775 2429 5776
rect 2563 5692 2572 5732
rect 2612 5692 2956 5732
rect 2996 5692 3005 5732
rect 8227 5692 8236 5732
rect 8276 5692 8428 5732
rect 8468 5692 8477 5732
rect 9100 5648 9140 5776
rect 22252 5732 22292 5776
rect 11587 5692 11596 5732
rect 11636 5692 13708 5732
rect 13748 5692 22292 5732
rect 22339 5692 22348 5732
rect 22388 5692 23212 5732
rect 23252 5692 23261 5732
rect 26083 5692 26092 5732
rect 26132 5692 26476 5732
rect 26516 5692 26525 5732
rect 16195 5648 16253 5649
rect 18403 5648 18461 5649
rect 1315 5608 1324 5648
rect 1364 5608 1373 5648
rect 1507 5608 1516 5648
rect 1556 5608 3724 5648
rect 3764 5608 3773 5648
rect 3907 5608 3916 5648
rect 3956 5608 6892 5648
rect 6932 5608 6941 5648
rect 8707 5608 8716 5648
rect 8756 5608 9100 5648
rect 9140 5608 9149 5648
rect 16110 5608 16204 5648
rect 16244 5608 16253 5648
rect 17347 5608 17356 5648
rect 17396 5608 18412 5648
rect 18452 5608 18461 5648
rect 1324 5564 1364 5608
rect 16195 5607 16253 5608
rect 18403 5607 18461 5608
rect 22819 5648 22877 5649
rect 27619 5648 27677 5649
rect 22819 5608 22828 5648
rect 22868 5608 24460 5648
rect 24500 5608 24509 5648
rect 27534 5608 27628 5648
rect 27668 5608 27677 5648
rect 28108 5648 28148 5776
rect 42928 5756 43008 5776
rect 29740 5692 30412 5732
rect 30452 5692 30461 5732
rect 33379 5692 33388 5732
rect 33428 5692 36652 5732
rect 36692 5692 36701 5732
rect 37795 5692 37804 5732
rect 37844 5692 41260 5732
rect 41300 5692 41309 5732
rect 29740 5648 29780 5692
rect 34723 5648 34781 5649
rect 28108 5608 29780 5648
rect 34638 5608 34732 5648
rect 34772 5608 34781 5648
rect 22819 5607 22877 5608
rect 27619 5607 27677 5608
rect 34723 5607 34781 5608
rect 35299 5648 35357 5649
rect 35299 5608 35308 5648
rect 35348 5608 35884 5648
rect 35924 5608 37996 5648
rect 38036 5608 38045 5648
rect 35299 5607 35357 5608
rect 14659 5564 14717 5565
rect 1324 5524 2036 5564
rect 3523 5524 3532 5564
rect 3572 5524 3581 5564
rect 4003 5524 4012 5564
rect 4052 5524 5356 5564
rect 5396 5524 5405 5564
rect 9964 5524 12596 5564
rect 0 5480 80 5500
rect 0 5440 1900 5480
rect 1940 5440 1949 5480
rect 0 5420 80 5440
rect 1996 5396 2036 5524
rect 3532 5480 3572 5524
rect 4291 5480 4349 5481
rect 3532 5440 4300 5480
rect 4340 5440 4349 5480
rect 4675 5440 4684 5480
rect 4724 5440 6508 5480
rect 6548 5440 6557 5480
rect 8323 5440 8332 5480
rect 8372 5440 9580 5480
rect 9620 5440 9629 5480
rect 4291 5439 4349 5440
rect 4483 5396 4541 5397
rect 9964 5396 10004 5524
rect 10243 5440 10252 5480
rect 10292 5440 10636 5480
rect 10676 5440 10685 5480
rect 12556 5396 12596 5524
rect 14659 5524 14668 5564
rect 14708 5524 18508 5564
rect 18548 5524 31700 5564
rect 31747 5524 31756 5564
rect 31796 5524 32716 5564
rect 32756 5524 32765 5564
rect 34243 5524 34252 5564
rect 34292 5524 35020 5564
rect 35060 5524 35069 5564
rect 35692 5524 37612 5564
rect 37652 5524 37661 5564
rect 37780 5524 40492 5564
rect 40532 5524 40541 5564
rect 14659 5523 14717 5524
rect 31660 5480 31700 5524
rect 35692 5480 35732 5524
rect 36355 5480 36413 5481
rect 37027 5480 37085 5481
rect 37780 5480 37820 5524
rect 17155 5440 17164 5480
rect 17204 5440 21100 5480
rect 21140 5440 21149 5480
rect 22243 5440 22252 5480
rect 22292 5440 24940 5480
rect 24980 5440 31372 5480
rect 31412 5440 31421 5480
rect 31660 5440 35692 5480
rect 35732 5440 35741 5480
rect 36270 5440 36364 5480
rect 36404 5440 36413 5480
rect 36942 5440 37036 5480
rect 37076 5440 37085 5480
rect 36355 5439 36413 5440
rect 37027 5439 37085 5440
rect 37132 5440 37820 5480
rect 37891 5480 37949 5481
rect 42928 5480 43008 5500
rect 37891 5440 37900 5480
rect 37940 5440 39916 5480
rect 39956 5440 39965 5480
rect 40675 5440 40684 5480
rect 40724 5440 43008 5480
rect 1996 5356 3532 5396
rect 3572 5356 3581 5396
rect 3628 5356 4492 5396
rect 4532 5356 10004 5396
rect 11320 5356 12500 5396
rect 12547 5356 12556 5396
rect 12596 5356 12605 5396
rect 13123 5356 13132 5396
rect 13172 5356 20716 5396
rect 20756 5356 20765 5396
rect 28195 5356 28204 5396
rect 28244 5356 28780 5396
rect 28820 5356 28829 5396
rect 30499 5356 30508 5396
rect 30548 5356 33484 5396
rect 33524 5356 33533 5396
rect 34339 5356 34348 5396
rect 34388 5356 34732 5396
rect 34772 5356 34781 5396
rect 3628 5312 3668 5356
rect 4483 5355 4541 5356
rect 11320 5312 11360 5356
rect 12259 5312 12317 5313
rect 12460 5312 12500 5356
rect 13132 5312 13172 5356
rect 21667 5312 21725 5313
rect 34531 5312 34589 5313
rect 2500 5272 3668 5312
rect 4919 5272 4928 5312
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 5296 5272 5305 5312
rect 6499 5272 6508 5312
rect 6548 5272 6796 5312
rect 6836 5272 6845 5312
rect 8428 5272 11360 5312
rect 12174 5272 12268 5312
rect 12308 5272 12317 5312
rect 12365 5272 12460 5312
rect 12500 5272 13172 5312
rect 14659 5272 14668 5312
rect 14708 5272 18452 5312
rect 20039 5272 20048 5312
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20416 5272 20425 5312
rect 20611 5272 20620 5312
rect 20660 5272 21196 5312
rect 21236 5272 21245 5312
rect 21648 5272 21676 5312
rect 21716 5272 21772 5312
rect 21812 5272 29836 5312
rect 29876 5272 31180 5312
rect 31220 5272 31229 5312
rect 33100 5272 33388 5312
rect 33428 5272 33437 5312
rect 34435 5272 34444 5312
rect 34484 5272 34540 5312
rect 34580 5272 34589 5312
rect 35159 5272 35168 5312
rect 35208 5272 35250 5312
rect 35290 5272 35332 5312
rect 35372 5272 35414 5312
rect 35454 5272 35496 5312
rect 35536 5272 35545 5312
rect 0 5144 80 5164
rect 2500 5144 2540 5272
rect 4291 5228 4349 5229
rect 8428 5228 8468 5272
rect 12259 5271 12317 5272
rect 14668 5228 14708 5272
rect 4291 5188 4300 5228
rect 4340 5188 7852 5228
rect 7892 5188 8428 5228
rect 8468 5188 8477 5228
rect 9475 5188 9484 5228
rect 9524 5188 13420 5228
rect 13460 5188 14708 5228
rect 18412 5228 18452 5272
rect 21667 5271 21725 5272
rect 33100 5228 33140 5272
rect 34531 5271 34589 5272
rect 37132 5228 37172 5440
rect 37891 5439 37949 5440
rect 42928 5420 43008 5440
rect 37780 5356 40876 5396
rect 40916 5356 40925 5396
rect 37780 5228 37820 5356
rect 18412 5188 33140 5228
rect 33187 5188 33196 5228
rect 33236 5188 37172 5228
rect 37228 5188 37820 5228
rect 4291 5187 4349 5188
rect 6691 5144 6749 5145
rect 26563 5144 26621 5145
rect 37228 5144 37268 5188
rect 42928 5144 43008 5164
rect 0 5104 2540 5144
rect 3427 5104 3436 5144
rect 3476 5104 5452 5144
rect 5492 5104 5501 5144
rect 6691 5104 6700 5144
rect 6740 5104 7276 5144
rect 7316 5104 7325 5144
rect 8899 5104 8908 5144
rect 8948 5104 9140 5144
rect 11491 5104 11500 5144
rect 11540 5104 14324 5144
rect 17059 5104 17068 5144
rect 17108 5104 20620 5144
rect 20660 5104 20669 5144
rect 20812 5104 24844 5144
rect 24884 5104 24893 5144
rect 26563 5104 26572 5144
rect 26612 5104 31276 5144
rect 31316 5104 31325 5144
rect 32131 5104 32140 5144
rect 32180 5104 37268 5144
rect 37603 5104 37612 5144
rect 37652 5104 38860 5144
rect 38900 5104 38909 5144
rect 41059 5104 41068 5144
rect 41108 5104 43008 5144
rect 0 5084 80 5104
rect 6691 5103 6749 5104
rect 9100 5060 9140 5104
rect 9571 5060 9629 5061
rect 11875 5060 11933 5061
rect 3811 5020 3820 5060
rect 3860 5020 4012 5060
rect 4052 5020 4061 5060
rect 4876 5020 7660 5060
rect 7700 5020 7709 5060
rect 8515 5020 8524 5060
rect 8564 5020 9004 5060
rect 9044 5020 9053 5060
rect 9100 5020 9388 5060
rect 9428 5020 9437 5060
rect 9571 5020 9580 5060
rect 9620 5020 11404 5060
rect 11444 5020 11453 5060
rect 11790 5020 11884 5060
rect 11924 5020 11933 5060
rect 14284 5060 14324 5104
rect 20812 5060 20852 5104
rect 24844 5060 24884 5104
rect 26563 5103 26621 5104
rect 42928 5084 43008 5104
rect 14284 5020 20852 5060
rect 20899 5020 20908 5060
rect 20948 5020 21388 5060
rect 21428 5020 21437 5060
rect 21667 5020 21676 5060
rect 21716 5020 22540 5060
rect 22580 5020 22589 5060
rect 24844 5020 29164 5060
rect 29204 5020 29356 5060
rect 29396 5020 29932 5060
rect 29972 5020 29981 5060
rect 32419 5020 32428 5060
rect 32468 5020 32812 5060
rect 32852 5020 33004 5060
rect 33044 5020 33053 5060
rect 33475 5020 33484 5060
rect 33524 5020 35308 5060
rect 35348 5020 35357 5060
rect 36931 5020 36940 5060
rect 36980 5020 37516 5060
rect 37556 5020 37565 5060
rect 37612 5020 38764 5060
rect 38804 5020 39052 5060
rect 39092 5020 39101 5060
rect 1315 4976 1373 4977
rect 4483 4976 4541 4977
rect 4876 4976 4916 5020
rect 9571 5019 9629 5020
rect 11875 5019 11933 5020
rect 5059 4976 5117 4977
rect 6595 4976 6653 4977
rect 12547 4976 12605 4977
rect 14851 4976 14909 4977
rect 22051 4976 22109 4977
rect 24547 4976 24605 4977
rect 26851 4976 26909 4977
rect 1230 4936 1324 4976
rect 1364 4936 1373 4976
rect 2851 4936 2860 4976
rect 2900 4936 3244 4976
rect 3284 4936 3293 4976
rect 4099 4936 4108 4976
rect 4148 4936 4492 4976
rect 4532 4936 4588 4976
rect 4628 4936 4637 4976
rect 4867 4936 4876 4976
rect 4916 4936 4925 4976
rect 4974 4936 5068 4976
rect 5108 4936 5117 4976
rect 5539 4936 5548 4976
rect 5588 4936 6604 4976
rect 6644 4936 6653 4976
rect 7267 4936 7276 4976
rect 7316 4936 8620 4976
rect 8660 4936 8669 4976
rect 10339 4936 10348 4976
rect 10388 4936 11308 4976
rect 11348 4936 11692 4976
rect 11732 4936 11741 4976
rect 12067 4936 12076 4976
rect 12116 4936 12125 4976
rect 12462 4936 12556 4976
rect 12596 4936 12605 4976
rect 13987 4936 13996 4976
rect 14036 4936 14284 4976
rect 14324 4936 14333 4976
rect 14766 4936 14860 4976
rect 14900 4936 14909 4976
rect 16675 4936 16684 4976
rect 16724 4936 16733 4976
rect 17539 4936 17548 4976
rect 17588 4936 18124 4976
rect 18164 4936 18173 4976
rect 18220 4936 18412 4976
rect 18452 4936 18461 4976
rect 19651 4936 19660 4976
rect 19700 4936 21044 4976
rect 21966 4936 22060 4976
rect 22100 4936 22109 4976
rect 24462 4936 24556 4976
rect 24596 4936 26188 4976
rect 26228 4936 26237 4976
rect 26851 4936 26860 4976
rect 26900 4936 37228 4976
rect 37268 4936 37277 4976
rect 1315 4935 1373 4936
rect 4483 4935 4541 4936
rect 5059 4935 5117 4936
rect 6595 4935 6653 4936
rect 12076 4892 12116 4936
rect 12547 4935 12605 4936
rect 14851 4935 14909 4936
rect 16684 4892 16724 4936
rect 18220 4892 18260 4936
rect 21004 4892 21044 4936
rect 22051 4935 22109 4936
rect 24547 4935 24605 4936
rect 26851 4935 26909 4936
rect 26947 4892 27005 4893
rect 31555 4892 31613 4893
rect 37612 4892 37652 5020
rect 2500 4852 6452 4892
rect 6787 4852 6796 4892
rect 6836 4852 7564 4892
rect 7604 4852 10540 4892
rect 10580 4852 10589 4892
rect 11395 4852 11404 4892
rect 11444 4852 12116 4892
rect 13603 4852 13612 4892
rect 13652 4852 16724 4892
rect 18019 4852 18028 4892
rect 18068 4852 18260 4892
rect 18307 4852 18316 4892
rect 18356 4852 20236 4892
rect 20276 4852 20285 4892
rect 20515 4852 20524 4892
rect 20564 4852 20573 4892
rect 20995 4852 21004 4892
rect 21044 4852 21053 4892
rect 21283 4852 21292 4892
rect 21332 4852 23348 4892
rect 26862 4852 26956 4892
rect 26996 4852 27005 4892
rect 0 4808 80 4828
rect 2500 4808 2540 4852
rect 6412 4808 6452 4852
rect 12076 4808 12116 4852
rect 20524 4808 20564 4852
rect 23308 4808 23348 4852
rect 26947 4851 27005 4852
rect 30220 4852 31564 4892
rect 31604 4852 32524 4892
rect 32564 4852 34444 4892
rect 34484 4852 34493 4892
rect 36739 4852 36748 4892
rect 36788 4852 37132 4892
rect 37172 4852 37612 4892
rect 37652 4852 37661 4892
rect 37795 4852 37804 4892
rect 37844 4852 40876 4892
rect 40916 4852 40925 4892
rect 30220 4808 30260 4852
rect 31555 4851 31613 4852
rect 42928 4808 43008 4828
rect 0 4768 2540 4808
rect 2755 4768 2764 4808
rect 2804 4768 4972 4808
rect 5012 4768 5021 4808
rect 6412 4768 10156 4808
rect 10196 4768 10924 4808
rect 10964 4768 10973 4808
rect 12076 4768 13228 4808
rect 13268 4768 15628 4808
rect 15668 4768 15677 4808
rect 20524 4768 21100 4808
rect 21140 4768 21149 4808
rect 23299 4768 23308 4808
rect 23348 4768 30220 4808
rect 30260 4768 30269 4808
rect 31267 4768 31276 4808
rect 31316 4768 38380 4808
rect 38420 4768 40492 4808
rect 40532 4768 40541 4808
rect 40675 4768 40684 4808
rect 40724 4768 43008 4808
rect 0 4748 80 4768
rect 2764 4724 2804 4768
rect 6595 4724 6653 4725
rect 6787 4724 6845 4725
rect 1315 4684 1324 4724
rect 1364 4684 2804 4724
rect 3907 4684 3916 4724
rect 3956 4684 4300 4724
rect 4340 4684 4349 4724
rect 4771 4684 4780 4724
rect 4820 4684 6412 4724
rect 6452 4684 6461 4724
rect 6595 4684 6604 4724
rect 6644 4684 6738 4724
rect 6787 4684 6796 4724
rect 6836 4684 9772 4724
rect 9812 4684 9821 4724
rect 17635 4684 17644 4724
rect 17684 4684 18412 4724
rect 18452 4684 21676 4724
rect 21716 4684 21725 4724
rect 22435 4684 22444 4724
rect 22484 4684 27052 4724
rect 27092 4684 27101 4724
rect 6595 4683 6653 4684
rect 6787 4683 6845 4684
rect 31276 4640 31316 4768
rect 42928 4748 43008 4768
rect 32323 4684 32332 4724
rect 32372 4684 32716 4724
rect 32756 4684 32765 4724
rect 33283 4684 33292 4724
rect 33332 4684 33676 4724
rect 33716 4684 33725 4724
rect 34051 4684 34060 4724
rect 34100 4684 35020 4724
rect 35060 4684 35069 4724
rect 38563 4684 38572 4724
rect 38612 4684 38956 4724
rect 38996 4684 39005 4724
rect 5059 4600 5068 4640
rect 5108 4600 5356 4640
rect 5396 4600 9388 4640
rect 9428 4600 13612 4640
rect 13652 4600 14284 4640
rect 14324 4600 14333 4640
rect 15724 4600 31316 4640
rect 32707 4640 32765 4641
rect 32707 4600 32716 4640
rect 32756 4600 41260 4640
rect 41300 4600 41309 4640
rect 15724 4556 15764 4600
rect 32707 4599 32765 4600
rect 3679 4516 3688 4556
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 4056 4516 4065 4556
rect 10915 4516 10924 4556
rect 10964 4516 15764 4556
rect 18799 4516 18808 4556
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 19176 4516 19185 4556
rect 23203 4516 23212 4556
rect 23252 4516 28588 4556
rect 28628 4516 28637 4556
rect 33919 4516 33928 4556
rect 33968 4516 34010 4556
rect 34050 4516 34092 4556
rect 34132 4516 34174 4556
rect 34214 4516 34256 4556
rect 34296 4516 34305 4556
rect 39235 4516 39244 4556
rect 39284 4516 39628 4556
rect 39668 4516 39677 4556
rect 0 4472 80 4492
rect 355 4472 413 4473
rect 6691 4472 6749 4473
rect 22147 4472 22205 4473
rect 42928 4472 43008 4492
rect 0 4432 364 4472
rect 404 4432 413 4472
rect 1699 4432 1708 4472
rect 1748 4432 2956 4472
rect 2996 4432 3005 4472
rect 6606 4432 6700 4472
rect 6740 4432 6749 4472
rect 8611 4432 8620 4472
rect 8660 4432 11360 4472
rect 11875 4432 11884 4472
rect 11924 4432 12268 4472
rect 12308 4432 12317 4472
rect 22062 4432 22156 4472
rect 22196 4432 22205 4472
rect 24451 4432 24460 4472
rect 24500 4432 25804 4472
rect 25844 4432 25853 4472
rect 26179 4432 26188 4472
rect 26228 4432 40876 4472
rect 40916 4432 40925 4472
rect 41059 4432 41068 4472
rect 41108 4432 43008 4472
rect 0 4412 80 4432
rect 355 4431 413 4432
rect 6691 4431 6749 4432
rect 11320 4388 11360 4432
rect 22147 4431 22205 4432
rect 42928 4412 43008 4432
rect 12547 4388 12605 4389
rect 4195 4348 4204 4388
rect 4244 4348 7372 4388
rect 7412 4348 7421 4388
rect 8995 4348 9004 4388
rect 9044 4348 10060 4388
rect 10100 4348 10109 4388
rect 11320 4348 12556 4388
rect 12596 4348 12605 4388
rect 14851 4348 14860 4388
rect 14900 4348 23116 4388
rect 23156 4348 23165 4388
rect 25699 4348 25708 4388
rect 25748 4348 26804 4388
rect 27043 4348 27052 4388
rect 27092 4348 30700 4388
rect 30740 4348 30749 4388
rect 31267 4348 31276 4388
rect 31316 4348 31468 4388
rect 31508 4348 40012 4388
rect 40052 4348 40396 4388
rect 40436 4348 40445 4388
rect 12547 4347 12605 4348
rect 4099 4304 4157 4305
rect 13315 4304 13373 4305
rect 14563 4304 14621 4305
rect 26764 4304 26804 4348
rect 40291 4304 40349 4305
rect 3715 4264 3724 4304
rect 3764 4264 4108 4304
rect 4148 4264 7180 4304
rect 7220 4264 7229 4304
rect 9187 4264 9196 4304
rect 9236 4264 12844 4304
rect 12884 4264 13324 4304
rect 13364 4264 13373 4304
rect 14478 4264 14572 4304
rect 14612 4264 14621 4304
rect 20611 4264 20620 4304
rect 20660 4264 22828 4304
rect 22868 4264 26708 4304
rect 26764 4264 32908 4304
rect 32948 4264 32957 4304
rect 40206 4264 40300 4304
rect 40340 4264 40349 4304
rect 4099 4263 4157 4264
rect 13315 4263 13373 4264
rect 14563 4263 14621 4264
rect 4675 4220 4733 4221
rect 12259 4220 12317 4221
rect 26668 4220 26708 4264
rect 40291 4263 40349 4264
rect 2947 4180 2956 4220
rect 2996 4180 3244 4220
rect 3284 4180 4492 4220
rect 4532 4180 4541 4220
rect 4675 4180 4684 4220
rect 4724 4180 4818 4220
rect 5347 4180 5356 4220
rect 5396 4180 6124 4220
rect 6164 4180 6173 4220
rect 10060 4180 12268 4220
rect 12308 4180 12317 4220
rect 14371 4180 14380 4220
rect 14420 4180 26572 4220
rect 26612 4180 26621 4220
rect 26668 4180 29000 4220
rect 31075 4180 31084 4220
rect 31124 4180 31852 4220
rect 31892 4180 31901 4220
rect 33475 4180 33484 4220
rect 33524 4180 35692 4220
rect 35732 4180 35741 4220
rect 37027 4180 37036 4220
rect 37076 4180 40492 4220
rect 40532 4180 40541 4220
rect 4675 4179 4733 4180
rect 0 4136 80 4156
rect 5059 4136 5117 4137
rect 0 4096 5068 4136
rect 5108 4096 5117 4136
rect 5251 4096 5260 4136
rect 5300 4096 5548 4136
rect 5588 4096 5597 4136
rect 5827 4096 5836 4136
rect 5876 4096 9964 4136
rect 10004 4096 10013 4136
rect 0 4076 80 4096
rect 5059 4095 5117 4096
rect 4387 4052 4445 4053
rect 7363 4052 7421 4053
rect 10060 4052 10100 4180
rect 12259 4179 12317 4180
rect 10243 4136 10301 4137
rect 20035 4136 20093 4137
rect 28960 4136 29000 4180
rect 42928 4136 43008 4156
rect 10243 4096 10252 4136
rect 10292 4096 10828 4136
rect 10868 4096 10877 4136
rect 11320 4096 13900 4136
rect 13940 4096 17644 4136
rect 17684 4096 17693 4136
rect 17740 4096 20044 4136
rect 20084 4096 20093 4136
rect 21859 4096 21868 4136
rect 21908 4096 24748 4136
rect 24788 4096 24797 4136
rect 26851 4096 26860 4136
rect 26900 4096 27340 4136
rect 27380 4096 27389 4136
rect 28960 4096 33388 4136
rect 33428 4096 37996 4136
rect 38036 4096 38045 4136
rect 41443 4096 41452 4136
rect 41492 4096 43008 4136
rect 10243 4095 10301 4096
rect 2500 4012 4396 4052
rect 4436 4012 4445 4052
rect 4675 4012 4684 4052
rect 4724 4012 6316 4052
rect 6356 4012 7180 4052
rect 7220 4012 7229 4052
rect 7363 4012 7372 4052
rect 7412 4012 8620 4052
rect 8660 4012 10100 4052
rect 2500 3968 2540 4012
rect 4387 4011 4445 4012
rect 7363 4011 7421 4012
rect 11320 3968 11360 4096
rect 11875 4052 11933 4053
rect 17740 4052 17780 4096
rect 20035 4095 20093 4096
rect 42928 4076 43008 4096
rect 37795 4052 37853 4053
rect 11875 4012 11884 4052
rect 11924 4012 17780 4052
rect 17923 4012 17932 4052
rect 17972 4012 20620 4052
rect 20660 4012 20669 4052
rect 22339 4012 22348 4052
rect 22388 4012 25708 4052
rect 25748 4012 25757 4052
rect 26083 4012 26092 4052
rect 26132 4012 26380 4052
rect 26420 4012 26429 4052
rect 26659 4012 26668 4052
rect 26708 4012 29260 4052
rect 29300 4012 29309 4052
rect 31660 4012 32812 4052
rect 32852 4012 32861 4052
rect 34051 4012 34060 4052
rect 34100 4012 34444 4052
rect 34484 4012 34493 4052
rect 37710 4012 37804 4052
rect 37844 4012 37853 4052
rect 11875 4011 11933 4012
rect 1795 3928 1804 3968
rect 1844 3928 2540 3968
rect 3523 3928 3532 3968
rect 3572 3928 5932 3968
rect 5972 3928 5981 3968
rect 6595 3928 6604 3968
rect 6644 3928 7372 3968
rect 7412 3928 8524 3968
rect 8564 3928 11360 3968
rect 7363 3884 7421 3885
rect 2500 3844 4492 3884
rect 4532 3844 4541 3884
rect 4588 3844 7372 3884
rect 7412 3844 7421 3884
rect 7555 3844 7564 3884
rect 7604 3844 9580 3884
rect 9620 3844 9629 3884
rect 0 3800 80 3820
rect 2500 3800 2540 3844
rect 4387 3800 4445 3801
rect 4588 3800 4628 3844
rect 7363 3843 7421 3844
rect 7651 3800 7709 3801
rect 12076 3800 12116 4012
rect 22147 3968 22205 3969
rect 31660 3968 31700 4012
rect 37795 4011 37853 4012
rect 31843 3968 31901 3969
rect 34243 3968 34301 3969
rect 12259 3928 12268 3968
rect 12308 3928 13132 3968
rect 13172 3928 13181 3968
rect 13891 3928 13900 3968
rect 13940 3928 14668 3968
rect 14708 3928 14717 3968
rect 15907 3928 15916 3968
rect 15956 3928 20812 3968
rect 20852 3928 20861 3968
rect 21091 3928 21100 3968
rect 21140 3928 22004 3968
rect 12163 3884 12221 3885
rect 12547 3884 12605 3885
rect 21964 3884 22004 3928
rect 22147 3928 22156 3968
rect 22196 3928 31700 3968
rect 31758 3928 31852 3968
rect 31892 3928 31901 3968
rect 34158 3928 34252 3968
rect 34292 3928 34301 3968
rect 22147 3927 22205 3928
rect 31843 3927 31901 3928
rect 34243 3927 34301 3928
rect 34348 3928 35500 3968
rect 35540 3928 35549 3968
rect 35683 3928 35692 3968
rect 35732 3928 39820 3968
rect 39860 3928 39869 3968
rect 12163 3844 12172 3884
rect 12212 3844 12556 3884
rect 12596 3844 21868 3884
rect 21908 3844 21917 3884
rect 21964 3844 22348 3884
rect 22388 3844 22397 3884
rect 27139 3844 27148 3884
rect 27188 3844 27668 3884
rect 29539 3844 29548 3884
rect 29588 3844 30124 3884
rect 30164 3844 32332 3884
rect 32372 3844 32381 3884
rect 12163 3843 12221 3844
rect 12547 3843 12605 3844
rect 27628 3800 27668 3844
rect 34348 3800 34388 3928
rect 34435 3884 34493 3885
rect 34435 3844 34444 3884
rect 34484 3844 39916 3884
rect 39956 3844 39965 3884
rect 34435 3843 34493 3844
rect 42928 3800 43008 3820
rect 0 3760 2540 3800
rect 2851 3760 2860 3800
rect 2900 3760 3244 3800
rect 3284 3760 3293 3800
rect 4387 3760 4396 3800
rect 4436 3760 4628 3800
rect 4919 3760 4928 3800
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 5296 3760 5305 3800
rect 5539 3760 5548 3800
rect 5588 3760 6028 3800
rect 6068 3760 6077 3800
rect 7566 3760 7660 3800
rect 7700 3760 7709 3800
rect 8995 3760 9004 3800
rect 9044 3760 12116 3800
rect 12355 3760 12364 3800
rect 12404 3760 14284 3800
rect 14324 3760 14333 3800
rect 16099 3760 16108 3800
rect 16148 3760 16157 3800
rect 20039 3760 20048 3800
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20416 3760 20425 3800
rect 21187 3760 21196 3800
rect 21236 3760 22252 3800
rect 22292 3760 22301 3800
rect 22723 3760 22732 3800
rect 22772 3760 23500 3800
rect 23540 3760 23549 3800
rect 24259 3760 24268 3800
rect 24308 3760 24556 3800
rect 24596 3760 24605 3800
rect 25315 3760 25324 3800
rect 25364 3760 25516 3800
rect 25556 3760 25565 3800
rect 25699 3760 25708 3800
rect 25748 3760 27436 3800
rect 27476 3760 27485 3800
rect 27619 3760 27628 3800
rect 27668 3760 27677 3800
rect 29059 3760 29068 3800
rect 29108 3760 29932 3800
rect 29972 3760 29981 3800
rect 32611 3760 32620 3800
rect 32660 3760 34388 3800
rect 35159 3760 35168 3800
rect 35208 3760 35250 3800
rect 35290 3760 35332 3800
rect 35372 3760 35414 3800
rect 35454 3760 35496 3800
rect 35536 3760 35545 3800
rect 35683 3760 35692 3800
rect 35732 3760 36076 3800
rect 36116 3760 36125 3800
rect 41059 3760 41068 3800
rect 41108 3760 43008 3800
rect 0 3740 80 3760
rect 4387 3759 4445 3760
rect 7651 3759 7709 3760
rect 1411 3716 1469 3717
rect 12451 3716 12509 3717
rect 16108 3716 16148 3760
rect 42928 3740 43008 3760
rect 20515 3716 20573 3717
rect 1326 3676 1420 3716
rect 1460 3676 1469 3716
rect 1603 3676 1612 3716
rect 1652 3676 2540 3716
rect 2659 3676 2668 3716
rect 2708 3676 4684 3716
rect 4724 3676 5740 3716
rect 5780 3676 6412 3716
rect 6452 3676 6796 3716
rect 6836 3676 8908 3716
rect 8948 3676 8957 3716
rect 10627 3676 10636 3716
rect 10676 3676 12268 3716
rect 12308 3676 12317 3716
rect 12451 3676 12460 3716
rect 12500 3676 12594 3716
rect 13027 3676 13036 3716
rect 13076 3676 17260 3716
rect 17300 3676 18892 3716
rect 18932 3676 20180 3716
rect 20430 3676 20524 3716
rect 20564 3676 41260 3716
rect 41300 3676 41309 3716
rect 1411 3675 1469 3676
rect 2500 3632 2540 3676
rect 12451 3675 12509 3676
rect 12460 3632 12500 3675
rect 20140 3632 20180 3676
rect 20515 3675 20573 3676
rect 2500 3592 12500 3632
rect 14179 3592 14188 3632
rect 14228 3592 17836 3632
rect 17876 3592 17885 3632
rect 20140 3592 21292 3632
rect 21332 3592 21341 3632
rect 22435 3592 22444 3632
rect 22484 3592 25612 3632
rect 25652 3592 26092 3632
rect 26132 3592 26141 3632
rect 29443 3592 29452 3632
rect 29492 3592 29932 3632
rect 29972 3592 29981 3632
rect 31555 3592 31564 3632
rect 31604 3592 31852 3632
rect 31892 3592 31901 3632
rect 33859 3592 33868 3632
rect 33908 3592 34444 3632
rect 34484 3592 34493 3632
rect 34627 3592 34636 3632
rect 34676 3592 35020 3632
rect 35060 3592 35069 3632
rect 30019 3548 30077 3549
rect 2659 3508 2668 3548
rect 2708 3508 2860 3548
rect 2900 3508 2909 3548
rect 7939 3508 7948 3548
rect 7988 3508 9292 3548
rect 9332 3508 9341 3548
rect 14851 3508 14860 3548
rect 14900 3508 27628 3548
rect 27668 3508 27677 3548
rect 29164 3508 30028 3548
rect 30068 3508 30077 3548
rect 0 3464 80 3484
rect 1411 3464 1469 3465
rect 16003 3464 16061 3465
rect 17635 3464 17693 3465
rect 29164 3464 29204 3508
rect 30019 3507 30077 3508
rect 31555 3548 31613 3549
rect 40867 3548 40925 3549
rect 31555 3508 31564 3548
rect 31604 3508 34252 3548
rect 34292 3508 34828 3548
rect 34868 3508 35300 3548
rect 31555 3507 31613 3508
rect 32995 3464 33053 3465
rect 0 3424 1420 3464
rect 1460 3424 1469 3464
rect 1891 3424 1900 3464
rect 1940 3424 3820 3464
rect 3860 3424 3869 3464
rect 4003 3424 4012 3464
rect 4052 3424 9236 3464
rect 11395 3424 11404 3464
rect 11444 3424 14188 3464
rect 14228 3424 14237 3464
rect 15918 3424 16012 3464
rect 16052 3424 16061 3464
rect 17550 3424 17644 3464
rect 17684 3424 17693 3464
rect 23011 3424 23020 3464
rect 23060 3424 23980 3464
rect 24020 3424 26572 3464
rect 26612 3424 29204 3464
rect 30019 3424 30028 3464
rect 30068 3424 30412 3464
rect 30452 3424 30461 3464
rect 32910 3424 33004 3464
rect 33044 3424 33053 3464
rect 35260 3464 35300 3508
rect 36076 3508 39628 3548
rect 39668 3508 39677 3548
rect 40099 3508 40108 3548
rect 40148 3508 40876 3548
rect 40916 3508 40925 3548
rect 36076 3465 36116 3508
rect 40867 3507 40925 3508
rect 36067 3464 36125 3465
rect 42928 3464 43008 3484
rect 35260 3424 35884 3464
rect 35924 3424 35933 3464
rect 35982 3424 36076 3464
rect 36116 3424 36125 3464
rect 40675 3424 40684 3464
rect 40724 3424 43008 3464
rect 0 3404 80 3424
rect 1411 3423 1469 3424
rect 6979 3380 7037 3381
rect 3427 3340 3436 3380
rect 3476 3340 5068 3380
rect 5108 3340 5117 3380
rect 6979 3340 6988 3380
rect 7028 3340 7084 3380
rect 7124 3340 7133 3380
rect 6979 3339 7037 3340
rect 9196 3296 9236 3424
rect 16003 3423 16061 3424
rect 17635 3423 17693 3424
rect 32995 3423 33053 3424
rect 36067 3423 36125 3424
rect 42928 3404 43008 3424
rect 12451 3340 12460 3380
rect 12500 3340 12652 3380
rect 12692 3340 12701 3380
rect 15811 3340 15820 3380
rect 15860 3340 37516 3380
rect 37556 3340 37565 3380
rect 37699 3340 37708 3380
rect 37748 3340 40876 3380
rect 40916 3340 40925 3380
rect 1507 3256 1516 3296
rect 1556 3256 1804 3296
rect 1844 3256 1853 3296
rect 2755 3256 2764 3296
rect 2804 3256 3532 3296
rect 3572 3256 3581 3296
rect 5635 3256 5644 3296
rect 5684 3256 7276 3296
rect 7316 3256 7325 3296
rect 8611 3256 8620 3296
rect 8660 3256 9100 3296
rect 9140 3256 9149 3296
rect 9196 3256 12940 3296
rect 12980 3256 12989 3296
rect 14659 3256 14668 3296
rect 14708 3256 25612 3296
rect 25652 3256 27724 3296
rect 27764 3256 28300 3296
rect 28340 3256 28349 3296
rect 33667 3256 33676 3296
rect 33716 3256 38284 3296
rect 38324 3256 38333 3296
rect 9763 3212 9821 3213
rect 36931 3212 36989 3213
rect 3139 3172 3148 3212
rect 3188 3172 3724 3212
rect 3764 3172 3773 3212
rect 5923 3172 5932 3212
rect 5972 3172 7468 3212
rect 7508 3172 8428 3212
rect 8468 3172 8477 3212
rect 9763 3172 9772 3212
rect 9812 3172 11596 3212
rect 11636 3172 19372 3212
rect 19412 3172 19421 3212
rect 25315 3172 25324 3212
rect 25364 3172 27244 3212
rect 27284 3172 27293 3212
rect 30883 3172 30892 3212
rect 30932 3172 33580 3212
rect 33620 3172 33629 3212
rect 36846 3172 36940 3212
rect 36980 3172 36989 3212
rect 39907 3172 39916 3212
rect 39956 3172 40780 3212
rect 40820 3172 40829 3212
rect 41443 3172 41452 3212
rect 41492 3172 41600 3212
rect 9763 3171 9821 3172
rect 36931 3171 36989 3172
rect 0 3128 80 3148
rect 14467 3128 14525 3129
rect 41560 3128 41600 3172
rect 42928 3128 43008 3148
rect 0 3088 1612 3128
rect 1652 3088 1661 3128
rect 5827 3088 5836 3128
rect 5876 3088 6220 3128
rect 6260 3088 7948 3128
rect 7988 3088 7997 3128
rect 8044 3088 14188 3128
rect 14228 3088 14237 3128
rect 14467 3088 14476 3128
rect 14516 3088 14572 3128
rect 14612 3088 14621 3128
rect 24451 3088 24460 3128
rect 24500 3088 28300 3128
rect 28340 3088 28349 3128
rect 41560 3088 43008 3128
rect 0 3068 80 3088
rect 8044 3044 8084 3088
rect 14467 3087 14525 3088
rect 42928 3068 43008 3088
rect 29539 3044 29597 3045
rect 3679 3004 3688 3044
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 4056 3004 4065 3044
rect 7075 3004 7084 3044
rect 7124 3004 8084 3044
rect 10051 3004 10060 3044
rect 10100 3004 11404 3044
rect 11444 3004 11453 3044
rect 11779 3004 11788 3044
rect 11828 3004 18316 3044
rect 18356 3004 18365 3044
rect 18799 3004 18808 3044
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 19176 3004 19185 3044
rect 19459 3004 19468 3044
rect 19508 3004 19660 3044
rect 19700 3004 19709 3044
rect 20227 3004 20236 3044
rect 20276 3004 23020 3044
rect 23060 3004 23069 3044
rect 24067 3004 24076 3044
rect 24116 3004 25036 3044
rect 25076 3004 25085 3044
rect 29454 3004 29548 3044
rect 29588 3004 31276 3044
rect 31316 3004 31325 3044
rect 33919 3004 33928 3044
rect 33968 3004 34010 3044
rect 34050 3004 34092 3044
rect 34132 3004 34174 3044
rect 34214 3004 34256 3044
rect 34296 3004 34305 3044
rect 29539 3003 29597 3004
rect 31555 2960 31613 2961
rect 1603 2920 1612 2960
rect 1652 2920 2956 2960
rect 2996 2920 3005 2960
rect 4483 2920 4492 2960
rect 4532 2920 31180 2960
rect 31220 2920 31229 2960
rect 31470 2920 31564 2960
rect 31604 2920 31613 2960
rect 31555 2919 31613 2920
rect 1315 2876 1373 2877
rect 1795 2876 1853 2877
rect 12547 2876 12605 2877
rect 36067 2876 36125 2877
rect 1228 2836 1324 2876
rect 1364 2836 1373 2876
rect 1710 2836 1804 2876
rect 1844 2836 1853 2876
rect 0 2792 80 2812
rect 1228 2792 1268 2836
rect 1315 2835 1373 2836
rect 1795 2835 1853 2836
rect 2500 2836 12556 2876
rect 12596 2836 12605 2876
rect 12931 2836 12940 2876
rect 12980 2836 13228 2876
rect 13268 2836 13277 2876
rect 16291 2836 16300 2876
rect 16340 2836 22060 2876
rect 22100 2836 28780 2876
rect 28820 2836 28829 2876
rect 30211 2836 30220 2876
rect 30260 2836 30796 2876
rect 30836 2836 30845 2876
rect 31363 2836 31372 2876
rect 31412 2836 31948 2876
rect 31988 2836 31997 2876
rect 35982 2836 36076 2876
rect 36116 2836 36125 2876
rect 37411 2836 37420 2876
rect 37460 2836 37996 2876
rect 38036 2836 38045 2876
rect 2500 2792 2540 2836
rect 12547 2835 12605 2836
rect 36067 2835 36125 2836
rect 14467 2792 14525 2793
rect 19459 2792 19517 2793
rect 42928 2792 43008 2812
rect 0 2752 1268 2792
rect 1315 2752 1324 2792
rect 1364 2752 2540 2792
rect 3139 2752 3148 2792
rect 3188 2752 7084 2792
rect 7124 2752 7133 2792
rect 11107 2752 11116 2792
rect 11156 2752 11360 2792
rect 11971 2752 11980 2792
rect 12020 2752 13900 2792
rect 13940 2752 13949 2792
rect 14467 2752 14476 2792
rect 14516 2752 17644 2792
rect 17684 2752 19468 2792
rect 19508 2752 19517 2792
rect 19651 2752 19660 2792
rect 19700 2752 21292 2792
rect 21332 2752 21772 2792
rect 21812 2752 21821 2792
rect 23107 2752 23116 2792
rect 23156 2752 24308 2792
rect 25507 2752 25516 2792
rect 25556 2752 25708 2792
rect 25748 2752 25757 2792
rect 26467 2752 26476 2792
rect 26516 2752 36172 2792
rect 36212 2752 36221 2792
rect 37507 2752 37516 2792
rect 37556 2752 39340 2792
rect 39380 2752 40204 2792
rect 40244 2752 40253 2792
rect 41635 2752 41644 2792
rect 41684 2752 43008 2792
rect 0 2732 80 2752
rect 11320 2708 11360 2752
rect 14467 2751 14525 2752
rect 19459 2751 19517 2752
rect 24268 2709 24308 2752
rect 42928 2732 43008 2752
rect 24259 2708 24317 2709
rect 41443 2708 41501 2709
rect 3235 2668 3244 2708
rect 3284 2668 4972 2708
rect 5012 2668 5021 2708
rect 8419 2668 8428 2708
rect 8468 2668 9236 2708
rect 9667 2668 9676 2708
rect 9716 2668 10636 2708
rect 10676 2668 11212 2708
rect 11252 2668 11261 2708
rect 11320 2668 11788 2708
rect 11828 2668 11837 2708
rect 12259 2668 12268 2708
rect 12308 2668 15532 2708
rect 15572 2668 15581 2708
rect 18604 2668 22444 2708
rect 22484 2668 22493 2708
rect 23683 2668 23692 2708
rect 23732 2668 24076 2708
rect 24116 2668 24125 2708
rect 24259 2668 24268 2708
rect 24308 2668 24402 2708
rect 31171 2668 31180 2708
rect 31220 2668 32812 2708
rect 32852 2668 36556 2708
rect 36596 2668 37708 2708
rect 37748 2668 37757 2708
rect 38563 2668 38572 2708
rect 38612 2668 39724 2708
rect 39764 2668 39773 2708
rect 41358 2668 41452 2708
rect 41492 2668 41501 2708
rect 8803 2624 8861 2625
rect 9196 2624 9236 2668
rect 12451 2624 12509 2625
rect 15235 2624 15293 2625
rect 18604 2624 18644 2668
rect 24259 2667 24317 2668
rect 41443 2667 41501 2668
rect 19459 2624 19517 2625
rect 1315 2584 1324 2624
rect 1364 2584 5260 2624
rect 5300 2584 5309 2624
rect 8718 2584 8812 2624
rect 8852 2584 8861 2624
rect 9187 2584 9196 2624
rect 9236 2584 10060 2624
rect 10100 2584 10109 2624
rect 11395 2584 11404 2624
rect 11444 2584 12308 2624
rect 12366 2584 12460 2624
rect 12500 2584 12509 2624
rect 8803 2583 8861 2584
rect 3331 2540 3389 2541
rect 7171 2540 7229 2541
rect 12268 2540 12308 2584
rect 12451 2583 12509 2584
rect 12556 2584 13036 2624
rect 13076 2584 13708 2624
rect 13748 2584 13757 2624
rect 13891 2584 13900 2624
rect 13940 2584 15052 2624
rect 15092 2584 15101 2624
rect 15150 2584 15244 2624
rect 15284 2584 15293 2624
rect 17731 2584 17740 2624
rect 17780 2584 18260 2624
rect 18307 2584 18316 2624
rect 18356 2584 18604 2624
rect 18644 2584 18653 2624
rect 19171 2584 19180 2624
rect 19220 2584 19412 2624
rect 12556 2540 12596 2584
rect 15235 2583 15293 2584
rect 14467 2540 14525 2541
rect 17155 2540 17213 2541
rect 3246 2500 3340 2540
rect 3380 2500 3389 2540
rect 6948 2500 6988 2540
rect 7028 2500 7037 2540
rect 7171 2500 7180 2540
rect 7220 2500 7314 2540
rect 12268 2500 12596 2540
rect 14382 2500 14476 2540
rect 14516 2500 14525 2540
rect 15811 2500 15820 2540
rect 15860 2500 15869 2540
rect 17070 2500 17164 2540
rect 17204 2500 17213 2540
rect 18220 2540 18260 2584
rect 19372 2540 19412 2584
rect 19459 2584 19468 2624
rect 19508 2584 25996 2624
rect 26036 2584 26045 2624
rect 28291 2584 28300 2624
rect 28340 2584 29932 2624
rect 29972 2584 29981 2624
rect 31267 2584 31276 2624
rect 31316 2584 37036 2624
rect 37076 2584 37085 2624
rect 37795 2584 37804 2624
rect 37844 2584 38380 2624
rect 38420 2584 38429 2624
rect 39523 2584 39532 2624
rect 39572 2584 40588 2624
rect 40628 2584 40637 2624
rect 19459 2583 19517 2584
rect 19939 2540 19997 2541
rect 18220 2500 18412 2540
rect 18452 2500 18461 2540
rect 19332 2500 19372 2540
rect 19412 2500 19421 2540
rect 19854 2500 19948 2540
rect 19988 2500 19997 2540
rect 20131 2500 20140 2540
rect 20180 2500 20220 2540
rect 28003 2500 28012 2540
rect 28052 2500 29164 2540
rect 29204 2500 29213 2540
rect 30403 2500 30412 2540
rect 30452 2500 31564 2540
rect 31604 2500 31613 2540
rect 34404 2500 34444 2540
rect 34484 2500 34493 2540
rect 37780 2500 38420 2540
rect 39139 2500 39148 2540
rect 39188 2500 40876 2540
rect 40916 2500 40925 2540
rect 3331 2499 3389 2500
rect 0 2456 80 2476
rect 1795 2456 1853 2457
rect 0 2416 1804 2456
rect 1844 2416 1853 2456
rect 6988 2456 7028 2500
rect 7171 2499 7229 2500
rect 14467 2499 14525 2500
rect 12835 2456 12893 2457
rect 6988 2416 9388 2456
rect 9428 2416 9437 2456
rect 12750 2416 12844 2456
rect 12884 2416 12893 2456
rect 13603 2416 13612 2456
rect 13652 2416 14572 2456
rect 14612 2416 14621 2456
rect 0 2396 80 2416
rect 1795 2415 1853 2416
rect 12835 2415 12893 2416
rect 14563 2372 14621 2373
rect 15820 2372 15860 2500
rect 17155 2499 17213 2500
rect 19372 2456 19412 2500
rect 19939 2499 19997 2500
rect 20140 2456 20180 2500
rect 34444 2456 34484 2500
rect 16771 2416 16780 2456
rect 16820 2416 18164 2456
rect 19372 2416 20180 2456
rect 27907 2416 27916 2456
rect 27956 2416 31084 2456
rect 31124 2416 31133 2456
rect 33763 2416 33772 2456
rect 33812 2416 34484 2456
rect 18124 2372 18164 2416
rect 28963 2372 29021 2373
rect 37780 2372 37820 2500
rect 38380 2456 38420 2500
rect 42928 2456 43008 2476
rect 38371 2416 38380 2456
rect 38420 2416 38429 2456
rect 39811 2416 39820 2456
rect 39860 2416 40300 2456
rect 40340 2416 40349 2456
rect 41251 2416 41260 2456
rect 41300 2416 43008 2456
rect 42928 2396 43008 2416
rect 4291 2332 4300 2372
rect 4340 2332 9772 2372
rect 9812 2332 9821 2372
rect 12739 2332 12748 2372
rect 12788 2332 12980 2372
rect 13411 2332 13420 2372
rect 13460 2332 14572 2372
rect 14612 2332 14621 2372
rect 15235 2332 15244 2372
rect 15284 2332 15860 2372
rect 15916 2332 18028 2372
rect 18068 2332 18077 2372
rect 18124 2332 21868 2372
rect 21908 2332 21917 2372
rect 26371 2332 26380 2372
rect 26420 2332 28012 2372
rect 28052 2332 28061 2372
rect 28963 2332 28972 2372
rect 29012 2332 34924 2372
rect 34964 2332 37820 2372
rect 10531 2288 10589 2289
rect 1411 2248 1420 2288
rect 1460 2248 2188 2288
rect 2228 2248 2237 2288
rect 3235 2248 3244 2288
rect 3284 2248 3293 2288
rect 4919 2248 4928 2288
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 5296 2248 5305 2288
rect 5731 2248 5740 2288
rect 5780 2248 6892 2288
rect 6932 2248 10540 2288
rect 10580 2248 10589 2288
rect 3244 2204 3284 2248
rect 10531 2247 10589 2248
rect 11320 2248 12844 2288
rect 12884 2248 12893 2288
rect 11320 2204 11360 2248
rect 1507 2164 1516 2204
rect 1556 2164 2540 2204
rect 3244 2164 10540 2204
rect 10580 2164 11360 2204
rect 0 2120 80 2140
rect 2500 2120 2540 2164
rect 4483 2120 4541 2121
rect 12940 2120 12980 2332
rect 14563 2331 14621 2332
rect 13027 2248 13036 2288
rect 13076 2248 14956 2288
rect 14996 2248 15005 2288
rect 15916 2204 15956 2332
rect 28963 2331 29021 2332
rect 22723 2288 22781 2289
rect 17347 2248 17356 2288
rect 17396 2248 18124 2288
rect 18164 2248 18173 2288
rect 20039 2248 20048 2288
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20416 2248 20425 2288
rect 21772 2248 21964 2288
rect 22004 2248 22013 2288
rect 22723 2248 22732 2288
rect 22772 2248 27628 2288
rect 27668 2248 30316 2288
rect 30356 2248 30365 2288
rect 34243 2248 34252 2288
rect 34292 2248 34636 2288
rect 34676 2248 34685 2288
rect 35159 2248 35168 2288
rect 35208 2248 35250 2288
rect 35290 2248 35332 2288
rect 35372 2248 35414 2288
rect 35454 2248 35496 2288
rect 35536 2248 35545 2288
rect 37795 2248 37804 2288
rect 37844 2248 38476 2288
rect 38516 2248 38525 2288
rect 21772 2204 21812 2248
rect 22723 2247 22781 2248
rect 30019 2204 30077 2205
rect 14275 2164 14284 2204
rect 14324 2164 15956 2204
rect 16579 2164 16588 2204
rect 16628 2164 17068 2204
rect 17108 2164 21812 2204
rect 21859 2164 21868 2204
rect 21908 2164 25132 2204
rect 25172 2164 26284 2204
rect 26324 2164 26333 2204
rect 29934 2164 30028 2204
rect 30068 2164 30077 2204
rect 33955 2164 33964 2204
rect 34004 2164 37324 2204
rect 37364 2164 37373 2204
rect 30019 2163 30077 2164
rect 19555 2120 19613 2121
rect 36067 2120 36125 2121
rect 42928 2120 43008 2140
rect 0 2080 212 2120
rect 2500 2080 4492 2120
rect 4532 2080 7564 2120
rect 7604 2080 7613 2120
rect 9955 2080 9964 2120
rect 10004 2080 10252 2120
rect 10292 2080 10301 2120
rect 12067 2080 12076 2120
rect 12116 2080 12980 2120
rect 13795 2080 13804 2120
rect 13844 2080 16780 2120
rect 16820 2080 16829 2120
rect 19470 2080 19564 2120
rect 19604 2080 19613 2120
rect 0 2060 80 2080
rect 172 1952 212 2080
rect 4483 2079 4541 2080
rect 9571 2036 9629 2037
rect 12940 2036 12980 2080
rect 19555 2079 19613 2080
rect 19660 2080 22444 2120
rect 22484 2080 22493 2120
rect 25219 2080 25228 2120
rect 25268 2080 25996 2120
rect 26036 2080 26045 2120
rect 29539 2080 29548 2120
rect 29588 2080 30508 2120
rect 30548 2080 30557 2120
rect 31276 2080 31660 2120
rect 31700 2080 32332 2120
rect 32372 2080 34444 2120
rect 34484 2080 34493 2120
rect 36067 2080 36076 2120
rect 36116 2080 37076 2120
rect 37123 2080 37132 2120
rect 37172 2080 38476 2120
rect 38516 2080 38525 2120
rect 41635 2080 41644 2120
rect 41684 2080 43008 2120
rect 19660 2036 19700 2080
rect 31276 2036 31316 2080
rect 36067 2079 36125 2080
rect 31459 2036 31517 2037
rect 37036 2036 37076 2080
rect 42928 2060 43008 2080
rect 37795 2036 37853 2037
rect 4867 1996 4876 2036
rect 4916 1996 7852 2036
rect 7892 1996 7901 2036
rect 9486 1996 9580 2036
rect 9620 1996 9629 2036
rect 12739 1996 12748 2036
rect 12788 1996 12797 2036
rect 12940 1996 16492 2036
rect 16532 1996 16541 2036
rect 18403 1996 18412 2036
rect 18452 1996 19700 2036
rect 19843 1996 19852 2036
rect 19892 1996 23308 2036
rect 23348 1996 23357 2036
rect 24748 1996 31316 2036
rect 31374 1996 31468 2036
rect 31508 1996 31517 2036
rect 9571 1995 9629 1996
rect 1795 1952 1853 1953
rect 12748 1952 12788 1996
rect 16387 1952 16445 1953
rect 24748 1952 24788 1996
rect 31459 1995 31517 1996
rect 31756 1996 36460 2036
rect 36500 1996 36509 2036
rect 37036 1996 37324 2036
rect 37364 1996 37373 2036
rect 37795 1996 37804 2036
rect 37844 1996 39244 2036
rect 39284 1996 39293 2036
rect 26755 1952 26813 1953
rect 31756 1952 31796 1996
rect 37795 1995 37853 1996
rect 36835 1952 36893 1953
rect 172 1912 1804 1952
rect 1844 1912 1853 1952
rect 5251 1912 5260 1952
rect 5300 1912 5836 1952
rect 5876 1912 5885 1952
rect 9859 1912 9868 1952
rect 9908 1912 12788 1952
rect 12931 1912 12940 1952
rect 12980 1912 14092 1952
rect 14132 1912 14141 1952
rect 16302 1912 16396 1952
rect 16436 1912 16445 1952
rect 17635 1912 17644 1952
rect 17684 1912 19468 1952
rect 19508 1912 19517 1952
rect 20140 1912 24748 1952
rect 24788 1912 24797 1952
rect 25219 1912 25228 1952
rect 25268 1912 26092 1952
rect 26132 1912 26141 1952
rect 26371 1912 26380 1952
rect 26420 1912 26764 1952
rect 26804 1912 26813 1952
rect 26947 1912 26956 1952
rect 26996 1912 27436 1952
rect 27476 1912 27485 1952
rect 29827 1912 29836 1952
rect 29876 1912 31796 1952
rect 32803 1912 32812 1952
rect 32852 1912 33580 1952
rect 33620 1912 33629 1952
rect 36750 1912 36844 1952
rect 36884 1912 36893 1952
rect 37219 1912 37228 1952
rect 37268 1912 37900 1952
rect 37940 1912 39820 1952
rect 39860 1912 39869 1952
rect 1795 1911 1853 1912
rect 16387 1911 16445 1912
rect 6979 1868 7037 1869
rect 6211 1828 6220 1868
rect 6260 1828 6988 1868
rect 7028 1828 8428 1868
rect 8468 1828 10636 1868
rect 10676 1828 10685 1868
rect 12643 1828 12652 1868
rect 12692 1828 15820 1868
rect 15860 1828 15869 1868
rect 6979 1827 7037 1828
rect 0 1784 80 1804
rect 0 1744 1172 1784
rect 1411 1744 1420 1784
rect 1460 1744 2284 1784
rect 2324 1744 2333 1784
rect 5347 1744 5356 1784
rect 5396 1744 7180 1784
rect 7220 1744 7229 1784
rect 10051 1744 10060 1784
rect 10100 1744 11308 1784
rect 11348 1744 11357 1784
rect 11683 1744 11692 1784
rect 11732 1744 13996 1784
rect 14036 1744 14045 1784
rect 14947 1744 14956 1784
rect 14996 1744 15148 1784
rect 15188 1744 18604 1784
rect 18644 1744 18653 1784
rect 0 1724 80 1744
rect 1132 1700 1172 1744
rect 10531 1700 10589 1701
rect 20140 1700 20180 1912
rect 26755 1911 26813 1912
rect 36835 1911 36893 1912
rect 25315 1868 25373 1869
rect 28867 1868 28925 1869
rect 23107 1828 23116 1868
rect 23156 1828 23884 1868
rect 23924 1828 23933 1868
rect 25230 1828 25324 1868
rect 25364 1828 25373 1868
rect 27331 1828 27340 1868
rect 27380 1828 28396 1868
rect 28436 1828 28445 1868
rect 28867 1828 28876 1868
rect 28916 1828 29452 1868
rect 29492 1828 29501 1868
rect 30691 1828 30700 1868
rect 30740 1828 31948 1868
rect 31988 1828 31997 1868
rect 32131 1828 32140 1868
rect 32180 1828 34732 1868
rect 34772 1828 34781 1868
rect 36547 1828 36556 1868
rect 36596 1828 40108 1868
rect 40148 1828 40157 1868
rect 25315 1827 25373 1828
rect 28867 1827 28925 1828
rect 42928 1784 43008 1804
rect 21955 1744 21964 1784
rect 22004 1744 26668 1784
rect 26708 1744 26717 1784
rect 26764 1744 39052 1784
rect 39092 1744 39244 1784
rect 39284 1744 39293 1784
rect 41068 1744 43008 1784
rect 26179 1700 26237 1701
rect 26764 1700 26804 1744
rect 28291 1700 28349 1701
rect 32803 1700 32861 1701
rect 40675 1700 40733 1701
rect 41068 1700 41108 1744
rect 42928 1724 43008 1744
rect 1132 1660 1804 1700
rect 1844 1660 1853 1700
rect 4099 1660 4108 1700
rect 4148 1660 4492 1700
rect 4532 1660 4541 1700
rect 5635 1660 5644 1700
rect 5684 1660 6508 1700
rect 6548 1660 7948 1700
rect 7988 1660 10348 1700
rect 10388 1660 10397 1700
rect 10531 1660 10540 1700
rect 10580 1660 10674 1700
rect 14860 1660 20180 1700
rect 21091 1660 21100 1700
rect 21140 1660 21868 1700
rect 21908 1660 21917 1700
rect 23107 1660 23116 1700
rect 23156 1660 23692 1700
rect 23732 1660 23741 1700
rect 26179 1660 26188 1700
rect 26228 1660 26804 1700
rect 27331 1660 27340 1700
rect 27380 1660 27820 1700
rect 27860 1660 27869 1700
rect 28291 1660 28300 1700
rect 28340 1660 29068 1700
rect 29108 1660 29117 1700
rect 29251 1660 29260 1700
rect 29300 1660 31756 1700
rect 31796 1660 31805 1700
rect 32803 1660 32812 1700
rect 32852 1660 33004 1700
rect 33044 1660 33053 1700
rect 34243 1660 34252 1700
rect 34292 1660 34828 1700
rect 34868 1660 34877 1700
rect 40590 1660 40684 1700
rect 40724 1660 40733 1700
rect 41059 1660 41068 1700
rect 41108 1660 41117 1700
rect 10531 1659 10589 1660
rect 14860 1616 14900 1660
rect 26179 1659 26237 1660
rect 28291 1659 28349 1660
rect 32803 1659 32861 1660
rect 34252 1616 34292 1660
rect 40675 1659 40733 1660
rect 5155 1576 5164 1616
rect 5204 1576 12172 1616
rect 12212 1576 13420 1616
rect 13460 1576 13469 1616
rect 13795 1576 13804 1616
rect 13844 1576 14900 1616
rect 14956 1576 24364 1616
rect 24404 1576 24413 1616
rect 24835 1576 24844 1616
rect 24884 1576 34292 1616
rect 4291 1532 4349 1533
rect 14563 1532 14621 1533
rect 14956 1532 14996 1576
rect 1603 1492 1612 1532
rect 1652 1492 1900 1532
rect 1940 1492 1949 1532
rect 3679 1492 3688 1532
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 4056 1492 4065 1532
rect 4206 1492 4300 1532
rect 4340 1492 4349 1532
rect 5539 1492 5548 1532
rect 5588 1492 8332 1532
rect 8372 1492 11116 1532
rect 11156 1492 11165 1532
rect 11779 1492 11788 1532
rect 11828 1492 14572 1532
rect 14612 1492 14996 1532
rect 18019 1492 18028 1532
rect 18068 1492 18412 1532
rect 18452 1492 18461 1532
rect 18799 1492 18808 1532
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 19176 1492 19185 1532
rect 19363 1492 19372 1532
rect 19412 1492 19564 1532
rect 19604 1492 19613 1532
rect 23920 1492 29548 1532
rect 29588 1492 29597 1532
rect 31651 1492 31660 1532
rect 31700 1492 32140 1532
rect 32180 1492 32189 1532
rect 33919 1492 33928 1532
rect 33968 1492 34010 1532
rect 34050 1492 34092 1532
rect 34132 1492 34174 1532
rect 34214 1492 34256 1532
rect 34296 1492 34305 1532
rect 4291 1491 4349 1492
rect 14563 1491 14621 1492
rect 0 1448 80 1468
rect 16291 1448 16349 1449
rect 23920 1448 23960 1492
rect 40867 1448 40925 1449
rect 42928 1448 43008 1468
rect 0 1408 3340 1448
rect 3380 1408 3389 1448
rect 5827 1408 5836 1448
rect 5876 1408 6644 1448
rect 9475 1408 9484 1448
rect 9524 1408 9772 1448
rect 9812 1408 10924 1448
rect 10964 1408 10973 1448
rect 13411 1408 13420 1448
rect 13460 1408 14668 1448
rect 14708 1408 15052 1448
rect 15092 1408 15101 1448
rect 16099 1408 16108 1448
rect 16148 1408 16157 1448
rect 16291 1408 16300 1448
rect 16340 1408 23960 1448
rect 26179 1408 26188 1448
rect 26228 1408 30892 1448
rect 30932 1408 30941 1448
rect 32419 1408 32428 1448
rect 32468 1408 32477 1448
rect 33283 1408 33292 1448
rect 33332 1408 39916 1448
rect 39956 1408 39965 1448
rect 40867 1408 40876 1448
rect 40916 1408 43008 1448
rect 0 1388 80 1408
rect 6604 1364 6644 1408
rect 10243 1364 10301 1365
rect 6604 1324 10252 1364
rect 10292 1324 10301 1364
rect 12739 1324 12748 1364
rect 12788 1324 13324 1364
rect 13364 1324 13373 1364
rect 10243 1323 10301 1324
rect 12163 1280 12221 1281
rect 16108 1280 16148 1408
rect 16291 1407 16349 1408
rect 29251 1364 29309 1365
rect 16483 1324 16492 1364
rect 16532 1324 21484 1364
rect 21524 1324 21533 1364
rect 22147 1324 22156 1364
rect 22196 1324 22205 1364
rect 22627 1324 22636 1364
rect 22676 1324 23156 1364
rect 23299 1324 23308 1364
rect 23348 1324 24940 1364
rect 24980 1324 24989 1364
rect 26668 1324 29260 1364
rect 29300 1324 29309 1364
rect 29443 1324 29452 1364
rect 29492 1324 31276 1364
rect 31316 1324 31325 1364
rect 22156 1280 22196 1324
rect 23116 1280 23156 1324
rect 26668 1280 26708 1324
rect 29251 1323 29309 1324
rect 1315 1240 1324 1280
rect 1364 1240 3724 1280
rect 3764 1240 3773 1280
rect 3820 1240 4684 1280
rect 4724 1240 5068 1280
rect 5108 1240 5117 1280
rect 7747 1240 7756 1280
rect 7796 1240 10444 1280
rect 10484 1240 10493 1280
rect 10915 1240 10924 1280
rect 10964 1240 11980 1280
rect 12020 1240 12029 1280
rect 12078 1240 12172 1280
rect 12212 1240 12221 1280
rect 12355 1240 12364 1280
rect 12404 1240 13228 1280
rect 13268 1240 13277 1280
rect 14851 1240 14860 1280
rect 14900 1240 15436 1280
rect 15476 1240 15485 1280
rect 16108 1240 20524 1280
rect 20564 1240 20573 1280
rect 22156 1240 23020 1280
rect 23060 1240 23069 1280
rect 23116 1240 26708 1280
rect 26755 1280 26813 1281
rect 28963 1280 29021 1281
rect 31363 1280 31421 1281
rect 26755 1240 26764 1280
rect 26804 1240 26813 1280
rect 27235 1240 27244 1280
rect 27284 1240 27532 1280
rect 27572 1240 27581 1280
rect 28963 1240 28972 1280
rect 29012 1240 30220 1280
rect 30260 1240 30269 1280
rect 31278 1240 31372 1280
rect 31412 1240 31421 1280
rect 3820 1196 3860 1240
rect 12163 1239 12221 1240
rect 26755 1239 26813 1240
rect 28963 1239 29021 1240
rect 31363 1239 31421 1240
rect 4579 1196 4637 1197
rect 10147 1196 10205 1197
rect 14947 1196 15005 1197
rect 20611 1196 20669 1197
rect 26563 1196 26621 1197
rect 1219 1156 1228 1196
rect 1268 1156 3860 1196
rect 4012 1156 4588 1196
rect 4628 1156 4637 1196
rect 5443 1156 5452 1196
rect 5492 1156 7988 1196
rect 8899 1156 8908 1196
rect 8948 1156 9812 1196
rect 0 1112 80 1132
rect 3619 1112 3677 1113
rect 4012 1112 4052 1156
rect 4579 1155 4637 1156
rect 7948 1113 7988 1156
rect 0 1072 3436 1112
rect 3476 1072 3628 1112
rect 3668 1072 3677 1112
rect 3811 1072 3820 1112
rect 3860 1072 4052 1112
rect 4099 1112 4157 1113
rect 7939 1112 7997 1113
rect 9772 1112 9812 1156
rect 10147 1156 10156 1196
rect 10196 1156 10252 1196
rect 10292 1156 10301 1196
rect 14947 1156 14956 1196
rect 14996 1156 15148 1196
rect 15188 1156 15197 1196
rect 15619 1156 15628 1196
rect 15668 1156 19660 1196
rect 19700 1156 19709 1196
rect 20526 1156 20620 1196
rect 20660 1156 20669 1196
rect 10147 1155 10205 1156
rect 14947 1155 15005 1156
rect 20611 1155 20669 1156
rect 20812 1156 23212 1196
rect 23252 1156 23261 1196
rect 25987 1156 25996 1196
rect 26036 1156 26572 1196
rect 26612 1156 26621 1196
rect 11587 1112 11645 1113
rect 18115 1112 18173 1113
rect 20707 1112 20765 1113
rect 4099 1072 4108 1112
rect 4148 1072 4396 1112
rect 4436 1072 4445 1112
rect 5155 1072 5164 1112
rect 5204 1072 5932 1112
rect 5972 1072 5981 1112
rect 6883 1072 6892 1112
rect 6932 1072 7372 1112
rect 7412 1072 7421 1112
rect 7854 1072 7948 1112
rect 7988 1072 7997 1112
rect 8611 1072 8620 1112
rect 8660 1072 9676 1112
rect 9716 1072 9725 1112
rect 9772 1072 10732 1112
rect 10772 1072 10781 1112
rect 11502 1072 11596 1112
rect 11636 1072 11645 1112
rect 12835 1072 12844 1112
rect 12884 1072 13708 1112
rect 13748 1072 14668 1112
rect 14708 1072 14717 1112
rect 15427 1072 15436 1112
rect 15476 1072 16300 1112
rect 16340 1072 16349 1112
rect 18030 1072 18124 1112
rect 18164 1072 18173 1112
rect 20622 1072 20716 1112
rect 20756 1072 20765 1112
rect 0 1052 80 1072
rect 3619 1071 3677 1072
rect 4099 1071 4157 1072
rect 5932 944 5972 1072
rect 7939 1071 7997 1072
rect 11587 1071 11645 1072
rect 18115 1071 18173 1072
rect 20707 1071 20765 1072
rect 20812 1028 20852 1156
rect 26563 1155 26621 1156
rect 26659 1112 26717 1113
rect 21763 1072 21772 1112
rect 21812 1072 21964 1112
rect 22004 1072 23596 1112
rect 23636 1072 24172 1112
rect 24212 1072 25172 1112
rect 25603 1072 25612 1112
rect 25652 1072 26668 1112
rect 26708 1072 26717 1112
rect 26764 1112 26804 1239
rect 32428 1196 32468 1408
rect 40867 1407 40925 1408
rect 42928 1388 43008 1408
rect 32899 1324 32908 1364
rect 32948 1324 33676 1364
rect 33716 1324 33725 1364
rect 35203 1324 35212 1364
rect 35252 1324 38572 1364
rect 38612 1324 38621 1364
rect 39619 1324 39628 1364
rect 39668 1324 40108 1364
rect 40148 1324 41452 1364
rect 41492 1324 41501 1364
rect 33763 1240 33772 1280
rect 33812 1240 34348 1280
rect 34388 1240 34397 1280
rect 34627 1240 34636 1280
rect 34676 1240 35596 1280
rect 35636 1240 35645 1280
rect 38371 1240 38380 1280
rect 38420 1240 40972 1280
rect 41012 1240 41021 1280
rect 26851 1156 26860 1196
rect 26900 1156 27916 1196
rect 27956 1156 27965 1196
rect 28492 1156 29932 1196
rect 29972 1156 29981 1196
rect 30787 1156 30796 1196
rect 30836 1156 32468 1196
rect 32524 1156 36556 1196
rect 36596 1156 36605 1196
rect 36739 1156 36748 1196
rect 36788 1156 40876 1196
rect 40916 1156 40925 1196
rect 28492 1112 28532 1156
rect 28675 1112 28733 1113
rect 32524 1112 32564 1156
rect 33571 1112 33629 1113
rect 35203 1112 35261 1113
rect 42928 1112 43008 1132
rect 26764 1072 27436 1112
rect 27476 1072 28532 1112
rect 28590 1072 28684 1112
rect 28724 1072 29108 1112
rect 29155 1072 29164 1112
rect 29204 1072 29836 1112
rect 29876 1072 30700 1112
rect 30740 1072 30749 1112
rect 31939 1072 31948 1112
rect 31988 1072 32564 1112
rect 33486 1072 33580 1112
rect 33620 1072 33629 1112
rect 33955 1072 33964 1112
rect 34004 1072 34636 1112
rect 34676 1072 34685 1112
rect 35118 1072 35212 1112
rect 35252 1072 35261 1112
rect 35587 1072 35596 1112
rect 35636 1072 38860 1112
rect 38900 1072 40012 1112
rect 40052 1072 40061 1112
rect 40579 1072 40588 1112
rect 40628 1072 43008 1112
rect 25027 1028 25085 1029
rect 9379 988 9388 1028
rect 9428 988 10828 1028
rect 10868 988 10877 1028
rect 11395 988 11404 1028
rect 11444 988 15532 1028
rect 15572 988 15581 1028
rect 16396 988 20852 1028
rect 20899 988 20908 1028
rect 20948 988 25036 1028
rect 25076 988 25085 1028
rect 25132 1028 25172 1072
rect 26659 1071 26717 1072
rect 28675 1071 28733 1072
rect 28963 1028 29021 1029
rect 25132 988 25708 1028
rect 25748 988 28972 1028
rect 29012 988 29021 1028
rect 29068 1028 29108 1072
rect 31948 1028 31988 1072
rect 33571 1071 33629 1072
rect 35203 1071 35261 1072
rect 42928 1052 43008 1072
rect 29068 988 31988 1028
rect 32035 988 32044 1028
rect 32084 988 32524 1028
rect 32564 988 32573 1028
rect 32995 988 33004 1028
rect 33044 988 36748 1028
rect 36788 988 36797 1028
rect 16291 944 16349 945
rect 2083 904 2092 944
rect 2132 904 3532 944
rect 3572 904 3581 944
rect 5932 904 11020 944
rect 11060 904 16300 944
rect 16340 904 16349 944
rect 16291 903 16349 904
rect 16396 860 16436 988
rect 25027 987 25085 988
rect 28963 987 29021 988
rect 24067 944 24125 945
rect 18595 904 18604 944
rect 18644 904 19276 944
rect 19316 904 19325 944
rect 21763 904 21772 944
rect 21812 904 24076 944
rect 24116 904 24125 944
rect 24259 904 24268 944
rect 24308 904 28204 944
rect 28244 904 28253 944
rect 29059 904 29068 944
rect 29108 904 36268 944
rect 36308 904 36317 944
rect 36844 904 39436 944
rect 39476 904 39485 944
rect 24067 903 24125 904
rect 22243 860 22301 861
rect 26467 860 26525 861
rect 27043 860 27101 861
rect 36844 860 36884 904
rect 1603 820 1612 860
rect 1652 820 3244 860
rect 3284 820 4492 860
rect 4532 820 6644 860
rect 9667 820 9676 860
rect 9716 820 10156 860
rect 10196 820 10205 860
rect 13507 820 13516 860
rect 13556 820 13900 860
rect 13940 820 13949 860
rect 15043 820 15052 860
rect 15092 820 16436 860
rect 16771 820 16780 860
rect 16820 820 22060 860
rect 22100 820 22109 860
rect 22158 820 22252 860
rect 22292 820 22301 860
rect 24067 820 24076 860
rect 24116 820 26476 860
rect 26516 820 26525 860
rect 26958 820 27052 860
rect 27092 820 36844 860
rect 36884 820 36893 860
rect 37780 820 41260 860
rect 41300 820 41309 860
rect 0 776 80 796
rect 6604 776 6644 820
rect 22243 819 22301 820
rect 26467 819 26525 820
rect 27043 819 27101 820
rect 14659 776 14717 777
rect 15619 776 15677 777
rect 34531 776 34589 777
rect 0 736 2540 776
rect 4919 736 4928 776
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 5296 736 5305 776
rect 6595 736 6604 776
rect 6644 736 10924 776
rect 10964 736 10973 776
rect 13315 736 13324 776
rect 13364 736 13804 776
rect 13844 736 13853 776
rect 14467 736 14476 776
rect 14516 736 14668 776
rect 14708 736 14717 776
rect 15534 736 15628 776
rect 15668 736 15677 776
rect 16195 736 16204 776
rect 16244 736 18220 776
rect 18260 736 18269 776
rect 20039 736 20048 776
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20416 736 20425 776
rect 24931 736 24940 776
rect 24980 736 31660 776
rect 31700 736 31709 776
rect 32323 736 32332 776
rect 32372 736 34540 776
rect 34580 736 34589 776
rect 35159 736 35168 776
rect 35208 736 35250 776
rect 35290 736 35332 776
rect 35372 736 35414 776
rect 35454 736 35496 776
rect 35536 736 35545 776
rect 0 716 80 736
rect 2500 692 2540 736
rect 14659 735 14717 736
rect 15619 735 15677 736
rect 34531 735 34589 736
rect 25315 692 25373 693
rect 2500 652 5452 692
rect 5492 652 5501 692
rect 13891 652 13900 692
rect 13940 652 16876 692
rect 16916 652 16925 692
rect 17923 652 17932 692
rect 17972 652 25324 692
rect 25364 652 25373 692
rect 25315 651 25373 652
rect 25507 692 25565 693
rect 25795 692 25853 693
rect 25507 652 25516 692
rect 25556 652 25650 692
rect 25795 652 25804 692
rect 25844 652 25938 692
rect 26563 652 26572 692
rect 26612 652 27052 692
rect 27092 652 27101 692
rect 28483 652 28492 692
rect 28532 652 29000 692
rect 31747 652 31756 692
rect 31796 652 36652 692
rect 36692 652 36701 692
rect 25507 651 25565 652
rect 25795 651 25853 652
rect 1795 608 1853 609
rect 10243 608 10301 609
rect 27619 608 27677 609
rect 1710 568 1804 608
rect 1844 568 1853 608
rect 10158 568 10252 608
rect 10292 568 10301 608
rect 12547 568 12556 608
rect 12596 568 15148 608
rect 15188 568 15197 608
rect 16003 568 16012 608
rect 16052 568 20236 608
rect 20276 568 20285 608
rect 21379 568 21388 608
rect 21428 568 27628 608
rect 27668 568 27677 608
rect 1795 567 1853 568
rect 10243 567 10301 568
rect 27619 567 27677 568
rect 20227 524 20285 525
rect 27523 524 27581 525
rect 15715 484 15724 524
rect 15764 484 20044 524
rect 20084 484 20093 524
rect 20227 484 20236 524
rect 20276 484 22636 524
rect 22676 484 22685 524
rect 23683 484 23692 524
rect 23732 484 27532 524
rect 27572 484 27581 524
rect 28960 524 29000 652
rect 37780 608 37820 820
rect 42928 776 43008 796
rect 40771 736 40780 776
rect 40820 736 43008 776
rect 42928 716 43008 736
rect 30307 568 30316 608
rect 30356 568 37820 608
rect 28960 484 34540 524
rect 34580 484 34589 524
rect 20227 483 20285 484
rect 27523 483 27581 484
rect 0 440 80 460
rect 8803 440 8861 441
rect 17539 440 17597 441
rect 26851 440 26909 441
rect 42928 440 43008 460
rect 0 400 8812 440
rect 8852 400 8861 440
rect 14083 400 14092 440
rect 14132 400 17548 440
rect 17588 400 17597 440
rect 26563 400 26572 440
rect 26612 400 26860 440
rect 26900 400 26909 440
rect 29923 400 29932 440
rect 29972 400 32428 440
rect 32468 400 33964 440
rect 34004 400 34013 440
rect 40387 400 40396 440
rect 40436 400 43008 440
rect 0 380 80 400
rect 8803 399 8861 400
rect 17539 399 17597 400
rect 26851 399 26909 400
rect 42928 380 43008 400
rect 12835 356 12893 357
rect 12835 316 12844 356
rect 12884 316 16340 356
rect 16387 316 16396 356
rect 16436 316 24844 356
rect 24884 316 24893 356
rect 27139 316 27148 356
rect 27188 316 27532 356
rect 27572 316 27581 356
rect 12835 315 12893 316
rect 13411 272 13469 273
rect 16003 272 16061 273
rect 13326 232 13420 272
rect 13460 232 14996 272
rect 15918 232 16012 272
rect 16052 232 16061 272
rect 16300 272 16340 316
rect 28099 272 28157 273
rect 16300 232 19852 272
rect 19892 232 19901 272
rect 28014 232 28108 272
rect 28148 232 28157 272
rect 13411 231 13469 232
rect 14851 188 14909 189
rect 14766 148 14860 188
rect 14900 148 14909 188
rect 14956 188 14996 232
rect 16003 231 16061 232
rect 28099 231 28157 232
rect 28675 188 28733 189
rect 14956 148 16492 188
rect 16532 148 16541 188
rect 28590 148 28684 188
rect 28724 148 28733 188
rect 31843 148 31852 188
rect 31892 148 32140 188
rect 32180 148 32189 188
rect 14851 147 14909 148
rect 28675 147 28733 148
rect 0 104 80 124
rect 22147 104 22205 105
rect 24451 104 24509 105
rect 42928 104 43008 124
rect 0 64 5356 104
rect 5396 64 5405 104
rect 5635 64 5644 104
rect 5684 64 6508 104
rect 6548 64 11404 104
rect 11444 64 11453 104
rect 13699 64 13708 104
rect 13748 64 22156 104
rect 22196 64 22205 104
rect 24366 64 24460 104
rect 24500 64 24509 104
rect 26755 64 26764 104
rect 26804 64 40300 104
rect 40340 64 40349 104
rect 41443 64 41452 104
rect 41492 64 43008 104
rect 0 44 80 64
rect 22147 63 22205 64
rect 24451 63 24509 64
rect 42928 44 43008 64
<< via3 >>
rect 460 10144 500 10184
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 35168 9808 35208 9848
rect 35250 9808 35290 9848
rect 35332 9808 35372 9848
rect 35414 9808 35454 9848
rect 35496 9808 35536 9848
rect 14764 9472 14804 9512
rect 19756 9472 19796 9512
rect 32908 9472 32948 9512
rect 40492 9388 40532 9428
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 33928 9052 33968 9092
rect 34010 9052 34050 9092
rect 34092 9052 34132 9092
rect 34174 9052 34214 9092
rect 34256 9052 34296 9092
rect 37132 9052 37172 9092
rect 2476 8800 2516 8840
rect 4012 8800 4052 8840
rect 4204 8800 4244 8840
rect 1324 8632 1364 8672
rect 2380 8632 2420 8672
rect 8140 8716 8180 8756
rect 9580 8716 9620 8756
rect 41260 8716 41300 8756
rect 6124 8632 6164 8672
rect 7756 8632 7796 8672
rect 9772 8632 9812 8672
rect 16204 8632 16244 8672
rect 21292 8632 21332 8672
rect 4396 8380 4436 8420
rect 33676 8632 33716 8672
rect 38380 8632 38420 8672
rect 4204 8296 4244 8336
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 35168 8296 35208 8336
rect 35250 8296 35290 8336
rect 35332 8296 35372 8336
rect 35414 8296 35454 8336
rect 35496 8296 35536 8336
rect 4492 7960 4532 8000
rect 8716 7960 8756 8000
rect 12076 7960 12116 8000
rect 13708 7960 13748 8000
rect 33676 7960 33716 8000
rect 18508 7876 18548 7916
rect 36556 7876 36596 7916
rect 1228 7792 1268 7832
rect 4684 7792 4724 7832
rect 8140 7792 8180 7832
rect 23500 7792 23540 7832
rect 11788 7708 11828 7748
rect 16108 7708 16148 7748
rect 10156 7624 10196 7664
rect 1804 7540 1844 7580
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 25804 7540 25844 7580
rect 33928 7540 33968 7580
rect 34010 7540 34050 7580
rect 34092 7540 34132 7580
rect 34174 7540 34214 7580
rect 34256 7540 34296 7580
rect 4396 7120 4436 7160
rect 14476 7120 14516 7160
rect 17740 7120 17780 7160
rect 21388 7120 21428 7160
rect 30028 7120 30068 7160
rect 32908 7120 32948 7160
rect 1516 7036 1556 7076
rect 4588 7036 4628 7076
rect 11884 7036 11924 7076
rect 27532 7036 27572 7076
rect 36556 7036 36596 7076
rect 13804 6952 13844 6992
rect 40396 6952 40436 6992
rect 1804 6784 1844 6824
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 35168 6784 35208 6824
rect 35250 6784 35290 6824
rect 35332 6784 35372 6824
rect 35414 6784 35454 6824
rect 35496 6784 35536 6824
rect 1708 6448 1748 6488
rect 4012 6448 4052 6488
rect 8140 6448 8180 6488
rect 17740 6532 17780 6572
rect 16108 6448 16148 6488
rect 23116 6448 23156 6488
rect 30412 6448 30452 6488
rect 30700 6448 30740 6488
rect 35500 6448 35540 6488
rect 33292 6364 33332 6404
rect 34732 6364 34772 6404
rect 41260 6364 41300 6404
rect 1804 6280 1844 6320
rect 14956 6280 14996 6320
rect 1516 6112 1556 6152
rect 22636 6196 22676 6236
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 33928 6028 33968 6068
rect 34010 6028 34050 6068
rect 34092 6028 34132 6068
rect 34174 6028 34214 6068
rect 34256 6028 34296 6068
rect 21772 5944 21812 5984
rect 2380 5776 2420 5816
rect 16204 5608 16244 5648
rect 18412 5608 18452 5648
rect 22828 5608 22868 5648
rect 27628 5608 27668 5648
rect 34732 5608 34772 5648
rect 35308 5608 35348 5648
rect 4300 5440 4340 5480
rect 14668 5524 14708 5564
rect 36364 5440 36404 5480
rect 37036 5440 37076 5480
rect 37900 5440 37940 5480
rect 4492 5356 4532 5396
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 12268 5272 12308 5312
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 21676 5272 21716 5312
rect 34540 5272 34580 5312
rect 35168 5272 35208 5312
rect 35250 5272 35290 5312
rect 35332 5272 35372 5312
rect 35414 5272 35454 5312
rect 35496 5272 35536 5312
rect 4300 5188 4340 5228
rect 6700 5104 6740 5144
rect 26572 5104 26612 5144
rect 9580 5020 9620 5060
rect 11884 5020 11924 5060
rect 1324 4936 1364 4976
rect 4492 4936 4532 4976
rect 5068 4936 5108 4976
rect 6604 4936 6644 4976
rect 12556 4936 12596 4976
rect 14860 4936 14900 4976
rect 22060 4936 22100 4976
rect 24556 4936 24596 4976
rect 26860 4936 26900 4976
rect 26956 4852 26996 4892
rect 31564 4852 31604 4892
rect 6604 4684 6644 4724
rect 6796 4684 6836 4724
rect 32716 4600 32756 4640
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 33928 4516 33968 4556
rect 34010 4516 34050 4556
rect 34092 4516 34132 4556
rect 34174 4516 34214 4556
rect 34256 4516 34296 4556
rect 364 4432 404 4472
rect 6700 4432 6740 4472
rect 22156 4432 22196 4472
rect 12556 4348 12596 4388
rect 4108 4264 4148 4304
rect 13324 4264 13364 4304
rect 14572 4264 14612 4304
rect 40300 4264 40340 4304
rect 4684 4180 4724 4220
rect 12268 4180 12308 4220
rect 5068 4096 5108 4136
rect 10252 4096 10292 4136
rect 20044 4096 20084 4136
rect 4396 4012 4436 4052
rect 7372 4012 7412 4052
rect 11884 4012 11924 4052
rect 37804 4012 37844 4052
rect 7372 3844 7412 3884
rect 22156 3928 22196 3968
rect 31852 3928 31892 3968
rect 34252 3928 34292 3968
rect 12172 3844 12212 3884
rect 12556 3844 12596 3884
rect 34444 3844 34484 3884
rect 4396 3760 4436 3800
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 7660 3760 7700 3800
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 35168 3760 35208 3800
rect 35250 3760 35290 3800
rect 35332 3760 35372 3800
rect 35414 3760 35454 3800
rect 35496 3760 35536 3800
rect 1420 3676 1460 3716
rect 12460 3676 12500 3716
rect 20524 3676 20564 3716
rect 30028 3508 30068 3548
rect 31564 3508 31604 3548
rect 1420 3424 1460 3464
rect 16012 3424 16052 3464
rect 17644 3424 17684 3464
rect 33004 3424 33044 3464
rect 40876 3508 40916 3548
rect 36076 3424 36116 3464
rect 6988 3340 7028 3380
rect 9772 3172 9812 3212
rect 36940 3172 36980 3212
rect 14476 3088 14516 3128
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 29548 3004 29588 3044
rect 33928 3004 33968 3044
rect 34010 3004 34050 3044
rect 34092 3004 34132 3044
rect 34174 3004 34214 3044
rect 34256 3004 34296 3044
rect 31564 2920 31604 2960
rect 1324 2836 1364 2876
rect 1804 2836 1844 2876
rect 12556 2836 12596 2876
rect 36076 2836 36116 2876
rect 14476 2752 14516 2792
rect 19468 2752 19508 2792
rect 24268 2668 24308 2708
rect 41452 2668 41492 2708
rect 8812 2584 8852 2624
rect 12460 2584 12500 2624
rect 15244 2584 15284 2624
rect 3340 2500 3380 2540
rect 7180 2500 7220 2540
rect 14476 2500 14516 2540
rect 17164 2500 17204 2540
rect 19468 2584 19508 2624
rect 19948 2500 19988 2540
rect 1804 2416 1844 2456
rect 12844 2416 12884 2456
rect 14572 2332 14612 2372
rect 28972 2332 29012 2372
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 10540 2248 10580 2288
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 22732 2248 22772 2288
rect 35168 2248 35208 2288
rect 35250 2248 35290 2288
rect 35332 2248 35372 2288
rect 35414 2248 35454 2288
rect 35496 2248 35536 2288
rect 30028 2164 30068 2204
rect 4492 2080 4532 2120
rect 19564 2080 19604 2120
rect 36076 2080 36116 2120
rect 9580 1996 9620 2036
rect 31468 1996 31508 2036
rect 37804 1996 37844 2036
rect 1804 1912 1844 1952
rect 16396 1912 16436 1952
rect 26764 1912 26804 1952
rect 36844 1912 36884 1952
rect 6988 1828 7028 1868
rect 25324 1828 25364 1868
rect 28876 1828 28916 1868
rect 10540 1660 10580 1700
rect 26188 1660 26228 1700
rect 28300 1660 28340 1700
rect 32812 1660 32852 1700
rect 40684 1660 40724 1700
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 4300 1492 4340 1532
rect 14572 1492 14612 1532
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 33928 1492 33968 1532
rect 34010 1492 34050 1532
rect 34092 1492 34132 1532
rect 34174 1492 34214 1532
rect 34256 1492 34296 1532
rect 16300 1408 16340 1448
rect 40876 1408 40916 1448
rect 10252 1324 10292 1364
rect 29260 1324 29300 1364
rect 12172 1240 12212 1280
rect 26764 1240 26804 1280
rect 28972 1240 29012 1280
rect 31372 1240 31412 1280
rect 4588 1156 4628 1196
rect 3628 1072 3668 1112
rect 10156 1156 10196 1196
rect 14956 1156 14996 1196
rect 20620 1156 20660 1196
rect 26572 1156 26612 1196
rect 4108 1072 4148 1112
rect 7948 1072 7988 1112
rect 11596 1072 11636 1112
rect 18124 1072 18164 1112
rect 20716 1072 20756 1112
rect 26668 1072 26708 1112
rect 28684 1072 28724 1112
rect 33580 1072 33620 1112
rect 35212 1072 35252 1112
rect 25036 988 25076 1028
rect 28972 988 29012 1028
rect 16300 904 16340 944
rect 24076 904 24116 944
rect 22252 820 22292 860
rect 26476 820 26516 860
rect 27052 820 27092 860
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 14668 736 14708 776
rect 15628 736 15668 776
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 34540 736 34580 776
rect 35168 736 35208 776
rect 35250 736 35290 776
rect 35332 736 35372 776
rect 35414 736 35454 776
rect 35496 736 35536 776
rect 25324 652 25364 692
rect 25516 652 25556 692
rect 25804 652 25844 692
rect 1804 568 1844 608
rect 10252 568 10292 608
rect 27628 568 27668 608
rect 20236 484 20276 524
rect 27532 484 27572 524
rect 8812 400 8852 440
rect 17548 400 17588 440
rect 26860 400 26900 440
rect 12844 316 12884 356
rect 13420 232 13460 272
rect 16012 232 16052 272
rect 28108 232 28148 272
rect 14860 148 14900 188
rect 28684 148 28724 188
rect 22156 64 22196 104
rect 24460 64 24500 104
<< metal4 >>
rect 460 10184 500 10193
rect 460 8009 500 10144
rect 4928 9848 5296 9857
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 4928 9799 5296 9808
rect 20048 9848 20416 9857
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20048 9799 20416 9808
rect 35168 9848 35536 9857
rect 35208 9808 35250 9848
rect 35290 9808 35332 9848
rect 35372 9808 35414 9848
rect 35454 9808 35496 9848
rect 35168 9799 35536 9808
rect 14764 9512 14804 9521
rect 3688 9092 4056 9101
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 3688 9043 4056 9052
rect 2476 8840 2516 8849
rect 1323 8756 1365 8765
rect 1323 8716 1324 8756
rect 1364 8716 1365 8756
rect 1323 8707 1365 8716
rect 1803 8756 1845 8765
rect 1803 8716 1804 8756
rect 1844 8716 1845 8756
rect 1803 8707 1845 8716
rect 1324 8672 1364 8707
rect 1324 8621 1364 8632
rect 459 8000 501 8009
rect 459 7960 460 8000
rect 500 7960 501 8000
rect 459 7951 501 7960
rect 1227 7832 1269 7841
rect 1227 7792 1228 7832
rect 1268 7792 1269 7832
rect 1227 7783 1269 7792
rect 1228 7698 1268 7783
rect 1804 7580 1844 8707
rect 2379 8672 2421 8681
rect 2379 8632 2380 8672
rect 2420 8632 2421 8672
rect 2379 8623 2421 8632
rect 1804 7531 1844 7540
rect 1515 7160 1557 7169
rect 1515 7120 1516 7160
rect 1556 7120 1557 7160
rect 1515 7111 1557 7120
rect 1516 7076 1556 7111
rect 1516 6152 1556 7036
rect 1803 7076 1845 7085
rect 1803 7036 1804 7076
rect 1844 7036 1845 7076
rect 1803 7027 1845 7036
rect 1804 6824 1844 7027
rect 1707 6488 1749 6497
rect 1707 6448 1708 6488
rect 1748 6448 1749 6488
rect 1707 6439 1749 6448
rect 1708 6354 1748 6439
rect 1804 6320 1844 6784
rect 1804 6271 1844 6280
rect 1516 6103 1556 6112
rect 2380 5816 2420 8623
rect 2476 8513 2516 8800
rect 4012 8840 4052 8849
rect 2475 8504 2517 8513
rect 2475 8464 2476 8504
rect 2516 8464 2517 8504
rect 2475 8455 2517 8464
rect 4012 8177 4052 8800
rect 4204 8840 4244 8849
rect 4204 8336 4244 8800
rect 14764 8765 14804 9472
rect 19756 9512 19796 9521
rect 18808 9092 19176 9101
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 18808 9043 19176 9052
rect 8140 8756 8180 8765
rect 6124 8672 6164 8683
rect 6124 8597 6164 8632
rect 7756 8672 7796 8681
rect 6123 8588 6165 8597
rect 6123 8548 6124 8588
rect 6164 8548 6165 8588
rect 6123 8539 6165 8548
rect 7756 8513 7796 8632
rect 7755 8504 7797 8513
rect 7755 8464 7756 8504
rect 7796 8464 7797 8504
rect 7755 8455 7797 8464
rect 4204 8287 4244 8296
rect 4396 8420 4436 8429
rect 4011 8168 4053 8177
rect 4011 8128 4012 8168
rect 4052 8128 4053 8168
rect 4011 8119 4053 8128
rect 3688 7580 4056 7589
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 3688 7531 4056 7540
rect 4396 7160 4436 8380
rect 4928 8336 5296 8345
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 4928 8287 5296 8296
rect 6795 8168 6837 8177
rect 6795 8128 6796 8168
rect 6836 8128 6837 8168
rect 6795 8119 6837 8128
rect 4012 6488 4052 6497
rect 4012 6236 4052 6448
rect 4012 6196 4148 6236
rect 3688 6068 4056 6077
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 3688 6019 4056 6028
rect 2380 5767 2420 5776
rect 1324 4976 1364 4985
rect 1324 4817 1364 4936
rect 1323 4808 1365 4817
rect 1323 4768 1324 4808
rect 1364 4768 1365 4808
rect 1323 4759 1365 4768
rect 364 4472 404 4481
rect 364 3977 404 4432
rect 363 3968 405 3977
rect 363 3928 364 3968
rect 404 3928 405 3968
rect 363 3919 405 3928
rect 1324 2876 1364 4759
rect 3688 4556 4056 4565
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 3688 4507 4056 4516
rect 4108 4304 4148 6196
rect 1803 4220 1845 4229
rect 1803 4180 1804 4220
rect 1844 4180 1845 4220
rect 1803 4171 1845 4180
rect 1324 2827 1364 2836
rect 1420 3716 1460 3725
rect 1420 3464 1460 3676
rect 1420 2801 1460 3424
rect 1804 2876 1844 4171
rect 3688 3044 4056 3053
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 3688 2995 4056 3004
rect 1419 2792 1461 2801
rect 1419 2752 1420 2792
rect 1460 2752 1461 2792
rect 1419 2743 1461 2752
rect 1804 2456 1844 2836
rect 3339 2708 3381 2717
rect 3339 2668 3340 2708
rect 3380 2668 3381 2708
rect 3339 2659 3381 2668
rect 3340 2540 3380 2659
rect 3340 2491 3380 2500
rect 1804 2407 1844 2416
rect 1803 1952 1845 1961
rect 1803 1912 1804 1952
rect 1844 1912 1845 1952
rect 1803 1903 1845 1912
rect 1804 1818 1844 1903
rect 3688 1532 4056 1541
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 3688 1483 4056 1492
rect 3628 1112 3668 1123
rect 3628 1037 3668 1072
rect 4108 1112 4148 4264
rect 4300 5480 4340 5489
rect 4300 5228 4340 5440
rect 4300 1532 4340 5188
rect 4396 4052 4436 7120
rect 4492 8000 4532 8009
rect 4492 5396 4532 7960
rect 4684 7832 4724 7841
rect 4492 5347 4532 5356
rect 4588 7076 4628 7085
rect 4396 3800 4436 4012
rect 4396 3751 4436 3760
rect 4492 4976 4532 4985
rect 4492 2120 4532 4936
rect 4492 2071 4532 2080
rect 4300 1483 4340 1492
rect 4588 1196 4628 7036
rect 4684 4220 4724 7792
rect 4928 6824 5296 6833
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 4928 6775 5296 6784
rect 4928 5312 5296 5321
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 4928 5263 5296 5272
rect 6700 5144 6740 5153
rect 5067 4976 5109 4985
rect 5067 4936 5068 4976
rect 5108 4936 5109 4976
rect 5067 4927 5109 4936
rect 6604 4976 6644 4985
rect 4684 4171 4724 4180
rect 5068 4136 5108 4927
rect 6604 4724 6644 4936
rect 6604 4675 6644 4684
rect 6700 4472 6740 5104
rect 6796 4724 6836 8119
rect 8140 7832 8180 8716
rect 9580 8756 9620 8765
rect 8715 8504 8757 8513
rect 8715 8464 8716 8504
rect 8756 8464 8757 8504
rect 8715 8455 8757 8464
rect 8716 8000 8756 8455
rect 8716 7951 8756 7960
rect 8140 6488 8180 7792
rect 8140 6439 8180 6448
rect 9580 5060 9620 8716
rect 14763 8756 14805 8765
rect 14763 8716 14764 8756
rect 14804 8716 14805 8756
rect 14763 8707 14805 8716
rect 9580 5011 9620 5020
rect 9772 8672 9812 8681
rect 7659 4892 7701 4901
rect 7659 4852 7660 4892
rect 7700 4852 7701 4892
rect 7659 4843 7701 4852
rect 6796 4675 6836 4684
rect 6700 4423 6740 4432
rect 5068 4087 5108 4096
rect 7372 4052 7412 4061
rect 7372 3884 7412 4012
rect 7660 3977 7700 4843
rect 7659 3968 7701 3977
rect 7659 3928 7660 3968
rect 7700 3928 7701 3968
rect 7659 3919 7701 3928
rect 7372 3835 7412 3844
rect 4928 3800 5296 3809
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 4928 3751 5296 3760
rect 7660 3800 7700 3919
rect 7660 3751 7700 3760
rect 6988 3380 7028 3389
rect 4928 2288 5296 2297
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 4928 2239 5296 2248
rect 6988 1868 7028 3340
rect 9772 3212 9812 8632
rect 14764 8177 14804 8707
rect 16203 8672 16245 8681
rect 16203 8632 16204 8672
rect 16244 8632 16245 8672
rect 16203 8623 16245 8632
rect 14763 8168 14805 8177
rect 14763 8128 14764 8168
rect 14804 8128 14805 8168
rect 14763 8119 14805 8128
rect 16204 8009 16244 8623
rect 19756 8597 19796 9472
rect 32908 9512 32948 9521
rect 32908 8765 32948 9472
rect 40492 9428 40532 9437
rect 33928 9092 34296 9101
rect 33968 9052 34010 9092
rect 34050 9052 34092 9092
rect 34132 9052 34174 9092
rect 34214 9052 34256 9092
rect 33928 9043 34296 9052
rect 37132 9092 37172 9101
rect 32907 8756 32949 8765
rect 32907 8716 32908 8756
rect 32948 8716 32949 8756
rect 32907 8707 32949 8716
rect 21292 8672 21332 8683
rect 21292 8597 21332 8632
rect 33676 8672 33716 8712
rect 33676 8597 33716 8632
rect 19755 8588 19797 8597
rect 19755 8548 19756 8588
rect 19796 8548 19797 8588
rect 19755 8539 19797 8548
rect 21291 8588 21333 8597
rect 21291 8548 21292 8588
rect 21332 8548 21333 8588
rect 21291 8539 21333 8548
rect 33675 8588 33717 8597
rect 33675 8548 33676 8588
rect 33716 8548 33717 8588
rect 33675 8539 33717 8548
rect 20048 8336 20416 8345
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20048 8287 20416 8296
rect 21387 8168 21429 8177
rect 21387 8128 21388 8168
rect 21428 8128 21429 8168
rect 21387 8119 21429 8128
rect 12075 8000 12117 8009
rect 12075 7960 12076 8000
rect 12116 7960 12117 8000
rect 12075 7951 12117 7960
rect 13708 8000 13748 8009
rect 12076 7866 12116 7951
rect 11787 7748 11829 7757
rect 11787 7708 11788 7748
rect 11828 7708 11829 7748
rect 11787 7699 11829 7708
rect 9772 3163 9812 3172
rect 10156 7664 10196 7673
rect 8812 2624 8852 2633
rect 7179 2540 7221 2549
rect 7179 2500 7180 2540
rect 7220 2500 7221 2540
rect 7179 2491 7221 2500
rect 7180 2406 7220 2491
rect 6988 1819 7028 1828
rect 8812 1205 8852 2584
rect 9579 2036 9621 2045
rect 9579 1996 9580 2036
rect 9620 1996 9621 2036
rect 9579 1987 9621 1996
rect 9580 1902 9620 1987
rect 4588 1147 4628 1156
rect 8811 1196 8853 1205
rect 8811 1156 8812 1196
rect 8852 1156 8853 1196
rect 8811 1147 8853 1156
rect 10156 1196 10196 7624
rect 11788 7614 11828 7699
rect 11883 7160 11925 7169
rect 11883 7120 11884 7160
rect 11924 7120 11925 7160
rect 11883 7111 11925 7120
rect 11884 7076 11924 7111
rect 11884 7025 11924 7036
rect 13708 6581 13748 7960
rect 16203 8000 16245 8009
rect 16203 7960 16204 8000
rect 16244 7960 16245 8000
rect 16203 7951 16245 7960
rect 18508 7916 18548 7925
rect 16108 7748 16148 7757
rect 14476 7160 14516 7171
rect 14476 7085 14516 7120
rect 14475 7076 14517 7085
rect 14475 7036 14476 7076
rect 14516 7036 14517 7076
rect 14475 7027 14517 7036
rect 13803 6992 13845 7001
rect 13803 6952 13804 6992
rect 13844 6952 13845 6992
rect 13803 6943 13845 6952
rect 13804 6858 13844 6943
rect 13707 6572 13749 6581
rect 13707 6532 13708 6572
rect 13748 6532 13749 6572
rect 13707 6523 13749 6532
rect 16108 6488 16148 7708
rect 17740 7160 17780 7169
rect 17740 7001 17780 7120
rect 18508 7085 18548 7876
rect 18808 7580 19176 7589
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 18808 7531 19176 7540
rect 21388 7160 21428 8119
rect 23499 8000 23541 8009
rect 23499 7960 23500 8000
rect 23540 7960 23541 8000
rect 23499 7951 23541 7960
rect 33676 8000 33716 8539
rect 35168 8336 35536 8345
rect 35208 8296 35250 8336
rect 35290 8296 35332 8336
rect 35372 8296 35414 8336
rect 35454 8296 35496 8336
rect 35168 8287 35536 8296
rect 33676 7951 33716 7960
rect 23500 7832 23540 7951
rect 23500 7783 23540 7792
rect 36556 7916 36596 7925
rect 31371 7748 31413 7757
rect 31371 7708 31372 7748
rect 31412 7708 31413 7748
rect 31371 7699 31413 7708
rect 22635 7580 22677 7589
rect 22635 7540 22636 7580
rect 22676 7540 22677 7580
rect 22635 7531 22677 7540
rect 25804 7580 25844 7589
rect 22636 7169 22676 7531
rect 21388 7111 21428 7120
rect 22635 7160 22677 7169
rect 22635 7120 22636 7160
rect 22676 7120 22677 7160
rect 22635 7111 22677 7120
rect 18507 7076 18549 7085
rect 18507 7036 18508 7076
rect 18548 7036 18549 7076
rect 18507 7027 18549 7036
rect 17739 6992 17781 7001
rect 17739 6952 17740 6992
rect 17780 6952 17781 6992
rect 17739 6943 17781 6952
rect 20048 6824 20416 6833
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20048 6775 20416 6784
rect 16108 6413 16148 6448
rect 17740 6572 17780 6581
rect 16107 6404 16149 6413
rect 16107 6364 16108 6404
rect 16148 6364 16149 6404
rect 16107 6355 16149 6364
rect 14956 6320 14996 6329
rect 14668 5564 14708 5573
rect 12268 5312 12308 5321
rect 11884 5060 11924 5069
rect 10251 4808 10293 4817
rect 10251 4768 10252 4808
rect 10292 4768 10293 4808
rect 10251 4759 10293 4768
rect 10252 4136 10292 4759
rect 10252 3473 10292 4096
rect 11884 4052 11924 5020
rect 12268 4220 12308 5272
rect 13323 5060 13365 5069
rect 13323 5020 13324 5060
rect 13364 5020 13365 5060
rect 13323 5011 13365 5020
rect 12556 4976 12596 4985
rect 12556 4733 12596 4936
rect 12555 4724 12597 4733
rect 12555 4684 12556 4724
rect 12596 4684 12597 4724
rect 12555 4675 12597 4684
rect 12268 4171 12308 4180
rect 12556 4388 12596 4397
rect 11884 4003 11924 4012
rect 12172 3884 12212 3893
rect 10251 3464 10293 3473
rect 10251 3424 10252 3464
rect 10292 3424 10293 3464
rect 10251 3415 10293 3424
rect 10540 2288 10580 2297
rect 10540 1877 10580 2248
rect 10539 1868 10581 1877
rect 10539 1828 10540 1868
rect 10580 1828 10581 1868
rect 10539 1819 10581 1828
rect 10540 1700 10580 1819
rect 10540 1651 10580 1660
rect 10252 1364 10292 1404
rect 10252 1289 10292 1324
rect 10251 1280 10293 1289
rect 10251 1240 10252 1280
rect 10292 1240 10293 1280
rect 10251 1231 10293 1240
rect 12172 1280 12212 3844
rect 12556 3884 12596 4348
rect 13324 4304 13364 5011
rect 13324 4255 13364 4264
rect 14572 4304 14612 4313
rect 12556 3835 12596 3844
rect 12460 3716 12500 3725
rect 12460 3557 12500 3676
rect 12459 3548 12501 3557
rect 12459 3508 12460 3548
rect 12500 3508 12501 3548
rect 12459 3499 12501 3508
rect 14476 3128 14516 3137
rect 12555 2876 12597 2885
rect 12555 2836 12556 2876
rect 12596 2836 12597 2876
rect 12555 2827 12597 2836
rect 12556 2742 12596 2827
rect 14476 2792 14516 3088
rect 12460 2717 12500 2719
rect 12459 2708 12501 2717
rect 12459 2668 12460 2708
rect 12500 2668 12501 2708
rect 12459 2659 12501 2668
rect 12172 1231 12212 1240
rect 12460 2624 12500 2659
rect 10156 1147 10196 1156
rect 4108 1063 4148 1072
rect 7948 1112 7988 1121
rect 3627 1028 3669 1037
rect 3627 988 3628 1028
rect 3668 988 3669 1028
rect 3627 979 3669 988
rect 7948 953 7988 1072
rect 7947 944 7989 953
rect 7947 904 7948 944
rect 7988 904 7989 944
rect 7947 895 7989 904
rect 4928 776 5296 785
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 4928 727 5296 736
rect 1803 608 1845 617
rect 1803 568 1804 608
rect 1844 568 1845 608
rect 1803 559 1845 568
rect 1804 474 1844 559
rect 8812 440 8852 1147
rect 10252 608 10292 1231
rect 11596 1112 11636 1123
rect 12460 1121 12500 2584
rect 14476 2540 14516 2752
rect 14476 2491 14516 2500
rect 12844 2456 12884 2465
rect 11596 1037 11636 1072
rect 12459 1112 12501 1121
rect 12459 1072 12460 1112
rect 12500 1072 12501 1112
rect 12459 1063 12501 1072
rect 11595 1028 11637 1037
rect 11595 988 11596 1028
rect 11636 988 11637 1028
rect 11595 979 11637 988
rect 10252 559 10292 568
rect 8812 391 8852 400
rect 12844 356 12884 2416
rect 14572 2372 14612 4264
rect 14572 1532 14612 2332
rect 14572 1483 14612 1492
rect 14668 776 14708 5524
rect 14859 4976 14901 4985
rect 14859 4936 14860 4976
rect 14900 4936 14901 4976
rect 14859 4927 14901 4936
rect 14860 4842 14900 4927
rect 14956 1196 14996 6280
rect 17740 6245 17780 6532
rect 23116 6488 23156 6499
rect 23116 6413 23156 6448
rect 23115 6404 23157 6413
rect 23115 6364 23116 6404
rect 23156 6364 23157 6404
rect 23115 6355 23157 6364
rect 17739 6236 17781 6245
rect 17739 6196 17740 6236
rect 17780 6196 17781 6236
rect 17739 6187 17781 6196
rect 22635 6236 22677 6245
rect 22635 6196 22636 6236
rect 22676 6196 22677 6236
rect 22635 6187 22677 6196
rect 22636 6102 22676 6187
rect 18808 6068 19176 6077
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 18808 6019 19176 6028
rect 21772 5984 21812 5993
rect 16204 5648 16244 5657
rect 16204 4901 16244 5608
rect 18411 5648 18453 5657
rect 18411 5608 18412 5648
rect 18452 5608 18453 5648
rect 18411 5599 18453 5608
rect 18412 5514 18452 5599
rect 20048 5312 20416 5321
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20048 5263 20416 5272
rect 21676 5312 21716 5321
rect 17547 5144 17589 5153
rect 17547 5104 17548 5144
rect 17588 5104 17589 5144
rect 17547 5095 17589 5104
rect 16203 4892 16245 4901
rect 16203 4852 16204 4892
rect 16244 4852 16245 4892
rect 16203 4843 16245 4852
rect 17163 4892 17205 4901
rect 17163 4852 17164 4892
rect 17204 4852 17205 4892
rect 17163 4843 17205 4852
rect 16011 3464 16053 3473
rect 16011 3424 16012 3464
rect 16052 3424 16053 3464
rect 16011 3415 16053 3424
rect 16012 3330 16052 3415
rect 15243 2876 15285 2885
rect 15243 2836 15244 2876
rect 15284 2836 15285 2876
rect 15243 2827 15285 2836
rect 15244 2624 15284 2827
rect 15244 2575 15284 2584
rect 17164 2540 17204 4843
rect 17451 3296 17493 3305
rect 17451 3256 17452 3296
rect 17492 3256 17493 3296
rect 17451 3247 17493 3256
rect 17164 2491 17204 2500
rect 15627 2372 15669 2381
rect 15627 2332 15628 2372
rect 15668 2332 15669 2372
rect 15627 2323 15669 2332
rect 14956 1147 14996 1156
rect 14668 727 14708 736
rect 15628 776 15668 2323
rect 17452 1961 17492 3247
rect 16396 1952 16436 1961
rect 16396 1793 16436 1912
rect 17451 1952 17493 1961
rect 17451 1912 17452 1952
rect 17492 1912 17493 1952
rect 17451 1903 17493 1912
rect 16395 1784 16437 1793
rect 16395 1744 16396 1784
rect 16436 1744 16437 1784
rect 16395 1735 16437 1744
rect 16300 1448 16340 1457
rect 16300 944 16340 1408
rect 16300 895 16340 904
rect 15628 727 15668 736
rect 13419 608 13461 617
rect 13419 568 13420 608
rect 13460 568 13461 608
rect 13419 559 13461 568
rect 12844 307 12884 316
rect 13420 272 13460 559
rect 16011 524 16053 533
rect 16011 484 16012 524
rect 16052 484 16053 524
rect 16011 475 16053 484
rect 13420 223 13460 232
rect 16012 272 16052 475
rect 17548 440 17588 5095
rect 21676 4901 21716 5272
rect 21772 5153 21812 5944
rect 25323 5732 25365 5741
rect 25323 5692 25324 5732
rect 25364 5692 25365 5732
rect 25323 5683 25365 5692
rect 22828 5648 22868 5657
rect 21771 5144 21813 5153
rect 21771 5104 21772 5144
rect 21812 5104 21813 5144
rect 21771 5095 21813 5104
rect 22059 5060 22101 5069
rect 22059 5020 22060 5060
rect 22100 5020 22101 5060
rect 22059 5011 22101 5020
rect 22060 4976 22100 5011
rect 22060 4925 22100 4936
rect 21675 4892 21717 4901
rect 21675 4852 21676 4892
rect 21716 4852 21717 4892
rect 21675 4843 21717 4852
rect 18808 4556 19176 4565
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 18808 4507 19176 4516
rect 22156 4472 22196 4481
rect 20619 4304 20661 4313
rect 20619 4264 20620 4304
rect 20660 4264 20661 4304
rect 20619 4255 20661 4264
rect 20043 4136 20085 4145
rect 20043 4096 20044 4136
rect 20084 4096 20085 4136
rect 20043 4087 20085 4096
rect 20044 4002 20084 4087
rect 20048 3800 20416 3809
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20048 3751 20416 3760
rect 20524 3716 20564 3725
rect 20524 3557 20564 3676
rect 17643 3548 17685 3557
rect 17643 3508 17644 3548
rect 17684 3508 17685 3548
rect 17643 3499 17685 3508
rect 20523 3548 20565 3557
rect 20523 3508 20524 3548
rect 20564 3508 20565 3548
rect 20523 3499 20565 3508
rect 17644 3464 17684 3499
rect 17644 3413 17684 3424
rect 18808 3044 19176 3053
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 18808 2995 19176 3004
rect 19468 2792 19508 2801
rect 19468 2624 19508 2752
rect 19468 2575 19508 2584
rect 19948 2549 19988 2634
rect 19947 2540 19989 2549
rect 19947 2500 19948 2540
rect 19988 2500 19989 2540
rect 19947 2491 19989 2500
rect 20048 2288 20416 2297
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20048 2239 20416 2248
rect 19563 2120 19605 2129
rect 19563 2080 19564 2120
rect 19604 2080 19605 2120
rect 19563 2071 19605 2080
rect 19564 1986 19604 2071
rect 18808 1532 19176 1541
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 18808 1483 19176 1492
rect 20620 1196 20660 4255
rect 22156 3968 22196 4432
rect 20620 1147 20660 1156
rect 20715 1196 20757 1205
rect 20715 1156 20716 1196
rect 20756 1156 20757 1196
rect 20715 1147 20757 1156
rect 18123 1112 18165 1121
rect 18123 1072 18124 1112
rect 18164 1072 18165 1112
rect 18123 1063 18165 1072
rect 20716 1112 20756 1147
rect 18124 978 18164 1063
rect 20716 1061 20756 1072
rect 20048 776 20416 785
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20048 727 20416 736
rect 20139 524 20181 533
rect 20236 524 20276 533
rect 20139 484 20140 524
rect 20180 484 20236 524
rect 20139 475 20181 484
rect 20236 475 20276 484
rect 20140 456 20180 475
rect 17548 391 17588 400
rect 16012 223 16052 232
rect 14859 188 14901 197
rect 14859 148 14860 188
rect 14900 148 14901 188
rect 14859 139 14901 148
rect 14860 54 14900 139
rect 22156 104 22196 3928
rect 22251 3464 22293 3473
rect 22251 3424 22252 3464
rect 22292 3424 22293 3464
rect 22251 3415 22293 3424
rect 22252 2717 22292 3415
rect 22251 2708 22293 2717
rect 22251 2668 22252 2708
rect 22292 2668 22293 2708
rect 22251 2659 22293 2668
rect 22252 860 22292 2659
rect 22731 2624 22773 2633
rect 22731 2584 22732 2624
rect 22772 2584 22773 2624
rect 22731 2575 22773 2584
rect 22732 2288 22772 2575
rect 22828 2465 22868 5608
rect 24075 5480 24117 5489
rect 24075 5440 24076 5480
rect 24116 5440 24117 5480
rect 24075 5431 24117 5440
rect 22827 2456 22869 2465
rect 22827 2416 22828 2456
rect 22868 2416 22869 2456
rect 22827 2407 22869 2416
rect 22732 2239 22772 2248
rect 24076 944 24116 5431
rect 24555 4976 24597 4985
rect 24555 4936 24556 4976
rect 24596 4936 24597 4976
rect 24555 4927 24597 4936
rect 24556 4842 24596 4927
rect 25035 3800 25077 3809
rect 25035 3760 25036 3800
rect 25076 3760 25077 3800
rect 25035 3751 25077 3760
rect 24268 2708 24308 2719
rect 24268 2633 24308 2668
rect 24267 2624 24309 2633
rect 24267 2584 24268 2624
rect 24308 2584 24309 2624
rect 24267 2575 24309 2584
rect 25036 1028 25076 3751
rect 25036 979 25076 988
rect 25324 1868 25364 5683
rect 24076 895 24116 904
rect 22252 811 22292 820
rect 25324 692 25364 1828
rect 25515 1028 25557 1037
rect 25515 988 25516 1028
rect 25556 988 25557 1028
rect 25515 979 25557 988
rect 25516 785 25556 979
rect 25515 776 25557 785
rect 25515 736 25516 776
rect 25556 736 25557 776
rect 25515 727 25557 736
rect 25324 643 25364 652
rect 25516 692 25556 727
rect 25516 642 25556 652
rect 25804 692 25844 7540
rect 27531 7244 27573 7253
rect 27531 7204 27532 7244
rect 27572 7204 27573 7244
rect 27531 7195 27573 7204
rect 27532 7076 27572 7195
rect 27532 7027 27572 7036
rect 30028 7160 30068 7169
rect 26955 6488 26997 6497
rect 26955 6448 26956 6488
rect 26996 6448 26997 6488
rect 26955 6439 26997 6448
rect 26572 5144 26612 5153
rect 25804 643 25844 652
rect 26188 1700 26228 1709
rect 24460 113 24500 198
rect 26188 197 26228 1660
rect 26475 1700 26517 1709
rect 26475 1660 26476 1700
rect 26516 1660 26517 1700
rect 26475 1651 26517 1660
rect 26476 860 26516 1651
rect 26572 1196 26612 5104
rect 26667 5144 26709 5153
rect 26667 5104 26668 5144
rect 26708 5104 26709 5144
rect 26667 5095 26709 5104
rect 26572 1147 26612 1156
rect 26668 1112 26708 5095
rect 26860 4976 26900 4985
rect 26764 1952 26804 1961
rect 26764 1280 26804 1912
rect 26764 1231 26804 1240
rect 26668 1063 26708 1072
rect 26476 811 26516 820
rect 26860 440 26900 4936
rect 26956 4892 26996 6439
rect 27628 5648 27668 5657
rect 27628 5069 27668 5608
rect 27627 5060 27669 5069
rect 27627 5020 27628 5060
rect 27668 5020 27669 5060
rect 27627 5011 27669 5020
rect 26956 4145 26996 4852
rect 28971 4220 29013 4229
rect 28971 4180 28972 4220
rect 29012 4180 29013 4220
rect 28971 4171 29013 4180
rect 26955 4136 26997 4145
rect 26955 4096 26956 4136
rect 26996 4096 26997 4136
rect 26955 4087 26997 4096
rect 27627 3968 27669 3977
rect 27627 3928 27628 3968
rect 27668 3928 27669 3968
rect 27627 3919 27669 3928
rect 27531 3212 27573 3221
rect 27531 3172 27532 3212
rect 27572 3172 27573 3212
rect 27531 3163 27573 3172
rect 27051 860 27093 869
rect 27051 820 27052 860
rect 27092 820 27093 860
rect 27051 811 27093 820
rect 27052 726 27092 811
rect 27532 524 27572 3163
rect 27628 608 27668 3919
rect 28972 2372 29012 4171
rect 30028 3548 30068 7120
rect 30411 6656 30453 6665
rect 30411 6616 30412 6656
rect 30452 6616 30453 6656
rect 30411 6607 30453 6616
rect 30412 6497 30452 6607
rect 30699 6572 30741 6581
rect 30699 6532 30700 6572
rect 30740 6532 30741 6572
rect 30699 6523 30741 6532
rect 30411 6488 30453 6497
rect 30411 6448 30412 6488
rect 30452 6448 30453 6488
rect 30411 6439 30453 6448
rect 30700 6488 30740 6523
rect 30412 6354 30452 6439
rect 30700 6437 30740 6448
rect 29548 3044 29588 3053
rect 29548 2801 29588 3004
rect 29547 2792 29589 2801
rect 29547 2752 29548 2792
rect 29588 2752 29589 2792
rect 29547 2743 29589 2752
rect 28972 2323 29012 2332
rect 30028 2204 30068 3508
rect 30028 2155 30068 2164
rect 28875 1868 28917 1877
rect 28875 1828 28876 1868
rect 28916 1828 28917 1868
rect 28875 1819 28917 1828
rect 28876 1734 28916 1819
rect 28300 1700 28340 1709
rect 28300 1289 28340 1660
rect 29259 1364 29301 1373
rect 29259 1324 29260 1364
rect 29300 1324 29301 1364
rect 29259 1315 29301 1324
rect 28299 1280 28341 1289
rect 28299 1240 28300 1280
rect 28340 1240 28341 1280
rect 28299 1231 28341 1240
rect 28972 1280 29012 1289
rect 28683 1196 28725 1205
rect 28683 1156 28684 1196
rect 28724 1156 28725 1196
rect 28683 1147 28725 1156
rect 28684 1112 28724 1147
rect 28684 1061 28724 1072
rect 28972 1028 29012 1240
rect 29260 1230 29300 1315
rect 31372 1280 31412 7699
rect 32907 7580 32949 7589
rect 32907 7540 32908 7580
rect 32948 7540 32949 7580
rect 32907 7531 32949 7540
rect 33928 7580 34296 7589
rect 33968 7540 34010 7580
rect 34050 7540 34092 7580
rect 34132 7540 34174 7580
rect 34214 7540 34256 7580
rect 33928 7531 34296 7540
rect 32908 7160 32948 7531
rect 36556 7253 36596 7876
rect 37132 7757 37172 9052
rect 38379 8672 38421 8681
rect 38379 8632 38380 8672
rect 38420 8632 38421 8672
rect 38379 8623 38421 8632
rect 38380 8538 38420 8623
rect 37131 7748 37173 7757
rect 37131 7708 37132 7748
rect 37172 7708 37173 7748
rect 37131 7699 37173 7708
rect 36555 7244 36597 7253
rect 36555 7204 36556 7244
rect 36596 7204 36597 7244
rect 36555 7195 36597 7204
rect 32908 7111 32948 7120
rect 36556 7076 36596 7087
rect 36556 7001 36596 7036
rect 36555 6992 36597 7001
rect 36555 6952 36556 6992
rect 36596 6952 36597 6992
rect 36555 6943 36597 6952
rect 40396 6992 40436 7001
rect 35168 6824 35536 6833
rect 35208 6784 35250 6824
rect 35290 6784 35332 6824
rect 35372 6784 35414 6824
rect 35454 6784 35496 6824
rect 35168 6775 35536 6784
rect 34731 6572 34773 6581
rect 34731 6532 34732 6572
rect 34772 6532 34773 6572
rect 34731 6523 34773 6532
rect 33291 6404 33333 6413
rect 33291 6364 33292 6404
rect 33332 6364 33333 6404
rect 33291 6355 33333 6364
rect 34732 6404 34772 6523
rect 33292 6270 33332 6355
rect 33928 6068 34296 6077
rect 33968 6028 34010 6068
rect 34050 6028 34092 6068
rect 34132 6028 34174 6068
rect 34214 6028 34256 6068
rect 33928 6019 34296 6028
rect 34732 5648 34772 6364
rect 35500 6488 35540 6497
rect 35500 5741 35540 6448
rect 35499 5732 35541 5741
rect 35499 5692 35500 5732
rect 35540 5692 35541 5732
rect 35499 5683 35541 5692
rect 34732 5599 34772 5608
rect 35308 5648 35348 5659
rect 35308 5573 35348 5608
rect 35307 5564 35349 5573
rect 35307 5524 35308 5564
rect 35348 5524 35349 5564
rect 35307 5515 35349 5524
rect 36363 5480 36405 5489
rect 36363 5440 36364 5480
rect 36404 5440 36405 5480
rect 36363 5431 36405 5440
rect 37036 5480 37076 5489
rect 36364 5346 36404 5431
rect 34540 5312 34580 5321
rect 31564 4892 31604 4901
rect 31564 3548 31604 4852
rect 33003 4724 33045 4733
rect 33003 4684 33004 4724
rect 33044 4684 33045 4724
rect 33003 4675 33045 4684
rect 32716 4640 32756 4649
rect 31852 3968 31892 3977
rect 31852 3809 31892 3928
rect 31851 3800 31893 3809
rect 31851 3760 31852 3800
rect 31892 3760 31893 3800
rect 31851 3751 31893 3760
rect 31564 2960 31604 3508
rect 31564 2911 31604 2920
rect 32716 2633 32756 4600
rect 33004 4061 33044 4675
rect 33928 4556 34296 4565
rect 33968 4516 34010 4556
rect 34050 4516 34092 4556
rect 34132 4516 34174 4556
rect 34214 4516 34256 4556
rect 33928 4507 34296 4516
rect 33003 4052 33045 4061
rect 33003 4012 33004 4052
rect 33044 4012 33045 4052
rect 33003 4003 33045 4012
rect 33004 3464 33044 4003
rect 34251 3968 34293 3977
rect 34251 3928 34252 3968
rect 34292 3928 34293 3968
rect 34251 3919 34293 3928
rect 34252 3834 34292 3919
rect 34444 3884 34484 3893
rect 33004 3415 33044 3424
rect 33928 3044 34296 3053
rect 33968 3004 34010 3044
rect 34050 3004 34092 3044
rect 34132 3004 34174 3044
rect 34214 3004 34256 3044
rect 33928 2995 34296 3004
rect 32715 2624 32757 2633
rect 32715 2584 32716 2624
rect 32756 2584 32757 2624
rect 32715 2575 32757 2584
rect 31467 2036 31509 2045
rect 31467 1996 31468 2036
rect 31508 1996 31509 2036
rect 31467 1987 31509 1996
rect 31468 1902 31508 1987
rect 32715 1784 32757 1793
rect 32715 1744 32716 1784
rect 32756 1744 32852 1784
rect 32715 1735 32757 1744
rect 32812 1700 32852 1744
rect 32812 1651 32852 1660
rect 33928 1532 34296 1541
rect 33968 1492 34010 1532
rect 34050 1492 34092 1532
rect 34132 1492 34174 1532
rect 34214 1492 34256 1532
rect 33928 1483 34296 1492
rect 31372 1231 31412 1240
rect 34444 1121 34484 3844
rect 33579 1112 33621 1121
rect 33579 1072 33580 1112
rect 33620 1072 33621 1112
rect 33579 1063 33621 1072
rect 34443 1112 34485 1121
rect 34443 1072 34444 1112
rect 34484 1072 34485 1112
rect 34443 1063 34485 1072
rect 28972 979 29012 988
rect 33580 978 33620 1063
rect 34540 776 34580 5272
rect 35168 5312 35536 5321
rect 35208 5272 35250 5312
rect 35290 5272 35332 5312
rect 35372 5272 35414 5312
rect 35454 5272 35496 5312
rect 35168 5263 35536 5272
rect 37036 5153 37076 5440
rect 37900 5480 37940 5489
rect 37035 5144 37077 5153
rect 37035 5104 37036 5144
rect 37076 5104 37077 5144
rect 37035 5095 37077 5104
rect 37803 4052 37845 4061
rect 37803 4012 37804 4052
rect 37844 4012 37845 4052
rect 37803 4003 37845 4012
rect 37804 3918 37844 4003
rect 35168 3800 35536 3809
rect 35208 3760 35250 3800
rect 35290 3760 35332 3800
rect 35372 3760 35414 3800
rect 35454 3760 35496 3800
rect 35168 3751 35536 3760
rect 36076 3464 36116 3473
rect 36076 3305 36116 3424
rect 36075 3296 36117 3305
rect 36075 3256 36076 3296
rect 36116 3256 36117 3296
rect 36075 3247 36117 3256
rect 36939 3212 36981 3221
rect 36939 3172 36940 3212
rect 36980 3172 36981 3212
rect 36939 3163 36981 3172
rect 36940 3078 36980 3163
rect 36076 2876 36116 2885
rect 35168 2288 35536 2297
rect 35208 2248 35250 2288
rect 35290 2248 35332 2288
rect 35372 2248 35414 2288
rect 35454 2248 35496 2288
rect 35168 2239 35536 2248
rect 36076 2129 36116 2836
rect 36075 2120 36117 2129
rect 36075 2080 36076 2120
rect 36116 2080 36117 2120
rect 36075 2071 36117 2080
rect 36076 1985 36116 2071
rect 37804 2036 37844 2045
rect 36844 1952 36884 1961
rect 36844 1373 36884 1912
rect 36843 1364 36885 1373
rect 36843 1324 36844 1364
rect 36884 1324 36885 1364
rect 36843 1315 36885 1324
rect 35212 1112 35252 1123
rect 35212 1037 35252 1072
rect 35211 1028 35253 1037
rect 35211 988 35212 1028
rect 35252 988 35253 1028
rect 35211 979 35253 988
rect 34540 727 34580 736
rect 35168 776 35536 785
rect 35208 736 35250 776
rect 35290 736 35332 776
rect 35372 736 35414 776
rect 35454 736 35496 776
rect 35168 727 35536 736
rect 27628 559 27668 568
rect 27532 475 27572 484
rect 26860 391 26900 400
rect 28107 272 28149 281
rect 28107 232 28108 272
rect 28148 232 28149 272
rect 28107 223 28149 232
rect 26187 188 26229 197
rect 26187 148 26188 188
rect 26228 148 26229 188
rect 26187 139 26229 148
rect 28108 138 28148 223
rect 28683 188 28725 197
rect 28683 148 28684 188
rect 28724 148 28725 188
rect 28683 139 28725 148
rect 22156 55 22196 64
rect 24459 104 24501 113
rect 24459 64 24460 104
rect 24500 64 24501 104
rect 24459 55 24501 64
rect 28684 54 28724 139
rect 37804 113 37844 1996
rect 37900 281 37940 5440
rect 40299 4304 40341 4313
rect 40299 4264 40300 4304
rect 40340 4264 40341 4304
rect 40299 4255 40341 4264
rect 40300 4170 40340 4255
rect 37899 272 37941 281
rect 37899 232 37900 272
rect 37940 232 37941 272
rect 37899 223 37941 232
rect 40396 197 40436 6952
rect 40492 6665 40532 9388
rect 41259 8756 41301 8765
rect 41259 8716 41260 8756
rect 41300 8716 41301 8756
rect 41259 8707 41301 8716
rect 41260 8622 41300 8707
rect 40491 6656 40533 6665
rect 40491 6616 40492 6656
rect 40532 6616 40533 6656
rect 40491 6607 40533 6616
rect 41260 6413 41300 6498
rect 41259 6404 41301 6413
rect 41259 6364 41260 6404
rect 41300 6364 41301 6404
rect 41259 6355 41301 6364
rect 40876 3548 40916 3557
rect 40683 1700 40725 1709
rect 40683 1660 40684 1700
rect 40724 1660 40725 1700
rect 40683 1651 40725 1660
rect 40684 1566 40724 1651
rect 40876 1448 40916 3508
rect 41451 2708 41493 2717
rect 41451 2668 41452 2708
rect 41492 2668 41493 2708
rect 41451 2659 41493 2668
rect 41452 2574 41492 2659
rect 40876 1399 40916 1408
rect 40395 188 40437 197
rect 40395 148 40396 188
rect 40436 148 40437 188
rect 40395 139 40437 148
rect 37803 104 37845 113
rect 37803 64 37804 104
rect 37844 64 37845 104
rect 37803 55 37845 64
<< via4 >>
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 35168 9808 35208 9848
rect 35250 9808 35290 9848
rect 35332 9808 35372 9848
rect 35414 9808 35454 9848
rect 35496 9808 35536 9848
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 1324 8716 1364 8756
rect 1804 8716 1844 8756
rect 460 7960 500 8000
rect 1228 7792 1268 7832
rect 2380 8632 2420 8672
rect 1516 7120 1556 7160
rect 1804 7036 1844 7076
rect 1708 6448 1748 6488
rect 2476 8464 2516 8504
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 6124 8548 6164 8588
rect 7756 8464 7796 8504
rect 4012 8128 4052 8168
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 6796 8128 6836 8168
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 1324 4768 1364 4808
rect 364 3928 404 3968
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 1804 4180 1844 4220
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 1420 2752 1460 2792
rect 3340 2668 3380 2708
rect 1804 1912 1844 1952
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 5068 4936 5108 4976
rect 8716 8464 8756 8504
rect 14764 8716 14804 8756
rect 7660 4852 7700 4892
rect 7660 3928 7700 3968
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 16204 8632 16244 8672
rect 14764 8128 14804 8168
rect 33928 9052 33968 9092
rect 34010 9052 34050 9092
rect 34092 9052 34132 9092
rect 34174 9052 34214 9092
rect 34256 9052 34296 9092
rect 32908 8716 32948 8756
rect 19756 8548 19796 8588
rect 21292 8548 21332 8588
rect 33676 8548 33716 8588
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 21388 8128 21428 8168
rect 12076 7960 12116 8000
rect 11788 7708 11828 7748
rect 7180 2500 7220 2540
rect 9580 1996 9620 2036
rect 8812 1156 8852 1196
rect 11884 7120 11924 7160
rect 16204 7960 16244 8000
rect 14476 7036 14516 7076
rect 13804 6952 13844 6992
rect 13708 6532 13748 6572
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 23500 7960 23540 8000
rect 35168 8296 35208 8336
rect 35250 8296 35290 8336
rect 35332 8296 35372 8336
rect 35414 8296 35454 8336
rect 35496 8296 35536 8336
rect 31372 7708 31412 7748
rect 22636 7540 22676 7580
rect 22636 7120 22676 7160
rect 18508 7036 18548 7076
rect 17740 6952 17780 6992
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 16108 6364 16148 6404
rect 10252 4768 10292 4808
rect 13324 5020 13364 5060
rect 12556 4684 12596 4724
rect 10252 3424 10292 3464
rect 10540 1828 10580 1868
rect 10252 1240 10292 1280
rect 12460 3508 12500 3548
rect 12556 2836 12596 2876
rect 12460 2668 12500 2708
rect 3628 988 3668 1028
rect 7948 904 7988 944
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 1804 568 1844 608
rect 12460 1072 12500 1112
rect 11596 988 11636 1028
rect 14860 4936 14900 4976
rect 23116 6364 23156 6404
rect 17740 6196 17780 6236
rect 22636 6196 22676 6236
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 18412 5608 18452 5648
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 17548 5104 17588 5144
rect 16204 4852 16244 4892
rect 17164 4852 17204 4892
rect 16012 3424 16052 3464
rect 15244 2836 15284 2876
rect 17452 3256 17492 3296
rect 15628 2332 15668 2372
rect 17452 1912 17492 1952
rect 16396 1744 16436 1784
rect 13420 568 13460 608
rect 16012 484 16052 524
rect 25324 5692 25364 5732
rect 21772 5104 21812 5144
rect 22060 5020 22100 5060
rect 21676 4852 21716 4892
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 20620 4264 20660 4304
rect 20044 4096 20084 4136
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 17644 3508 17684 3548
rect 20524 3508 20564 3548
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 19948 2500 19988 2540
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 19564 2080 19604 2120
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 20716 1156 20756 1196
rect 18124 1072 18164 1112
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 20140 484 20180 524
rect 14860 148 14900 188
rect 22252 3424 22292 3464
rect 22252 2668 22292 2708
rect 22732 2584 22772 2624
rect 24076 5440 24116 5480
rect 22828 2416 22868 2456
rect 24556 4936 24596 4976
rect 25036 3760 25076 3800
rect 24268 2584 24308 2624
rect 25516 988 25556 1028
rect 25516 736 25556 776
rect 27532 7204 27572 7244
rect 26956 6448 26996 6488
rect 26476 1660 26516 1700
rect 26668 5104 26708 5144
rect 27628 5020 27668 5060
rect 28972 4180 29012 4220
rect 26956 4096 26996 4136
rect 27628 3928 27668 3968
rect 27532 3172 27572 3212
rect 27052 820 27092 860
rect 30412 6616 30452 6656
rect 30700 6532 30740 6572
rect 30412 6448 30452 6488
rect 29548 2752 29588 2792
rect 28876 1828 28916 1868
rect 29260 1324 29300 1364
rect 28300 1240 28340 1280
rect 28684 1156 28724 1196
rect 32908 7540 32948 7580
rect 33928 7540 33968 7580
rect 34010 7540 34050 7580
rect 34092 7540 34132 7580
rect 34174 7540 34214 7580
rect 34256 7540 34296 7580
rect 38380 8632 38420 8672
rect 37132 7708 37172 7748
rect 36556 7204 36596 7244
rect 36556 6952 36596 6992
rect 35168 6784 35208 6824
rect 35250 6784 35290 6824
rect 35332 6784 35372 6824
rect 35414 6784 35454 6824
rect 35496 6784 35536 6824
rect 34732 6532 34772 6572
rect 33292 6364 33332 6404
rect 33928 6028 33968 6068
rect 34010 6028 34050 6068
rect 34092 6028 34132 6068
rect 34174 6028 34214 6068
rect 34256 6028 34296 6068
rect 35500 5692 35540 5732
rect 35308 5524 35348 5564
rect 36364 5440 36404 5480
rect 33004 4684 33044 4724
rect 31852 3760 31892 3800
rect 33928 4516 33968 4556
rect 34010 4516 34050 4556
rect 34092 4516 34132 4556
rect 34174 4516 34214 4556
rect 34256 4516 34296 4556
rect 33004 4012 33044 4052
rect 34252 3928 34292 3968
rect 33928 3004 33968 3044
rect 34010 3004 34050 3044
rect 34092 3004 34132 3044
rect 34174 3004 34214 3044
rect 34256 3004 34296 3044
rect 32716 2584 32756 2624
rect 31468 1996 31508 2036
rect 32716 1744 32756 1784
rect 33928 1492 33968 1532
rect 34010 1492 34050 1532
rect 34092 1492 34132 1532
rect 34174 1492 34214 1532
rect 34256 1492 34296 1532
rect 33580 1072 33620 1112
rect 34444 1072 34484 1112
rect 35168 5272 35208 5312
rect 35250 5272 35290 5312
rect 35332 5272 35372 5312
rect 35414 5272 35454 5312
rect 35496 5272 35536 5312
rect 37036 5104 37076 5144
rect 37804 4012 37844 4052
rect 35168 3760 35208 3800
rect 35250 3760 35290 3800
rect 35332 3760 35372 3800
rect 35414 3760 35454 3800
rect 35496 3760 35536 3800
rect 36076 3256 36116 3296
rect 36940 3172 36980 3212
rect 35168 2248 35208 2288
rect 35250 2248 35290 2288
rect 35332 2248 35372 2288
rect 35414 2248 35454 2288
rect 35496 2248 35536 2288
rect 36076 2080 36116 2120
rect 36844 1324 36884 1364
rect 35212 988 35252 1028
rect 35168 736 35208 776
rect 35250 736 35290 776
rect 35332 736 35372 776
rect 35414 736 35454 776
rect 35496 736 35536 776
rect 28108 232 28148 272
rect 26188 148 26228 188
rect 28684 148 28724 188
rect 24460 64 24500 104
rect 40300 4264 40340 4304
rect 37900 232 37940 272
rect 41260 8716 41300 8756
rect 40492 6616 40532 6656
rect 41260 6364 41300 6404
rect 40684 1660 40724 1700
rect 41452 2668 41492 2708
rect 40396 148 40436 188
rect 37804 64 37844 104
<< metal5 >>
rect 4919 9871 5305 9890
rect 4919 9848 4985 9871
rect 5071 9848 5153 9871
rect 5239 9848 5305 9871
rect 4919 9808 4928 9848
rect 4968 9808 4985 9848
rect 5071 9808 5092 9848
rect 5132 9808 5153 9848
rect 5239 9808 5256 9848
rect 5296 9808 5305 9848
rect 4919 9785 4985 9808
rect 5071 9785 5153 9808
rect 5239 9785 5305 9808
rect 4919 9766 5305 9785
rect 20039 9871 20425 9890
rect 20039 9848 20105 9871
rect 20191 9848 20273 9871
rect 20359 9848 20425 9871
rect 20039 9808 20048 9848
rect 20088 9808 20105 9848
rect 20191 9808 20212 9848
rect 20252 9808 20273 9848
rect 20359 9808 20376 9848
rect 20416 9808 20425 9848
rect 20039 9785 20105 9808
rect 20191 9785 20273 9808
rect 20359 9785 20425 9808
rect 20039 9766 20425 9785
rect 35159 9871 35545 9890
rect 35159 9848 35225 9871
rect 35311 9848 35393 9871
rect 35479 9848 35545 9871
rect 35159 9808 35168 9848
rect 35208 9808 35225 9848
rect 35311 9808 35332 9848
rect 35372 9808 35393 9848
rect 35479 9808 35496 9848
rect 35536 9808 35545 9848
rect 35159 9785 35225 9808
rect 35311 9785 35393 9808
rect 35479 9785 35545 9808
rect 35159 9766 35545 9785
rect 3679 9115 4065 9134
rect 3679 9092 3745 9115
rect 3831 9092 3913 9115
rect 3999 9092 4065 9115
rect 3679 9052 3688 9092
rect 3728 9052 3745 9092
rect 3831 9052 3852 9092
rect 3892 9052 3913 9092
rect 3999 9052 4016 9092
rect 4056 9052 4065 9092
rect 3679 9029 3745 9052
rect 3831 9029 3913 9052
rect 3999 9029 4065 9052
rect 3679 9010 4065 9029
rect 18799 9115 19185 9134
rect 18799 9092 18865 9115
rect 18951 9092 19033 9115
rect 19119 9092 19185 9115
rect 18799 9052 18808 9092
rect 18848 9052 18865 9092
rect 18951 9052 18972 9092
rect 19012 9052 19033 9092
rect 19119 9052 19136 9092
rect 19176 9052 19185 9092
rect 18799 9029 18865 9052
rect 18951 9029 19033 9052
rect 19119 9029 19185 9052
rect 18799 9010 19185 9029
rect 33919 9115 34305 9134
rect 33919 9092 33985 9115
rect 34071 9092 34153 9115
rect 34239 9092 34305 9115
rect 33919 9052 33928 9092
rect 33968 9052 33985 9092
rect 34071 9052 34092 9092
rect 34132 9052 34153 9092
rect 34239 9052 34256 9092
rect 34296 9052 34305 9092
rect 33919 9029 33985 9052
rect 34071 9029 34153 9052
rect 34239 9029 34305 9052
rect 33919 9010 34305 9029
rect 1315 8716 1324 8756
rect 1364 8716 1804 8756
rect 1844 8716 14764 8756
rect 14804 8716 14813 8756
rect 32899 8716 32908 8756
rect 32948 8716 41260 8756
rect 41300 8716 41309 8756
rect 2371 8632 2380 8672
rect 2420 8632 16204 8672
rect 16244 8632 16253 8672
rect 20140 8632 38380 8672
rect 38420 8632 38429 8672
rect 20140 8588 20180 8632
rect 6115 8548 6124 8588
rect 6164 8548 19756 8588
rect 19796 8548 20180 8588
rect 21283 8548 21292 8588
rect 21332 8548 33676 8588
rect 33716 8548 33725 8588
rect 2467 8464 2476 8504
rect 2516 8464 7756 8504
rect 7796 8464 8716 8504
rect 8756 8464 8765 8504
rect 4919 8359 5305 8378
rect 4919 8336 4985 8359
rect 5071 8336 5153 8359
rect 5239 8336 5305 8359
rect 4919 8296 4928 8336
rect 4968 8296 4985 8336
rect 5071 8296 5092 8336
rect 5132 8296 5153 8336
rect 5239 8296 5256 8336
rect 5296 8296 5305 8336
rect 4919 8273 4985 8296
rect 5071 8273 5153 8296
rect 5239 8273 5305 8296
rect 4919 8254 5305 8273
rect 20039 8359 20425 8378
rect 20039 8336 20105 8359
rect 20191 8336 20273 8359
rect 20359 8336 20425 8359
rect 20039 8296 20048 8336
rect 20088 8296 20105 8336
rect 20191 8296 20212 8336
rect 20252 8296 20273 8336
rect 20359 8296 20376 8336
rect 20416 8296 20425 8336
rect 20039 8273 20105 8296
rect 20191 8273 20273 8296
rect 20359 8273 20425 8296
rect 20039 8254 20425 8273
rect 35159 8359 35545 8378
rect 35159 8336 35225 8359
rect 35311 8336 35393 8359
rect 35479 8336 35545 8359
rect 35159 8296 35168 8336
rect 35208 8296 35225 8336
rect 35311 8296 35332 8336
rect 35372 8296 35393 8336
rect 35479 8296 35496 8336
rect 35536 8296 35545 8336
rect 35159 8273 35225 8296
rect 35311 8273 35393 8296
rect 35479 8273 35545 8296
rect 35159 8254 35545 8273
rect 4003 8128 4012 8168
rect 4052 8128 6796 8168
rect 6836 8128 6845 8168
rect 14755 8128 14764 8168
rect 14804 8128 21388 8168
rect 21428 8128 21437 8168
rect 451 7960 460 8000
rect 500 7960 12076 8000
rect 12116 7960 12125 8000
rect 16195 7960 16204 8000
rect 16244 7960 23500 8000
rect 23540 7960 23549 8000
rect 1219 7792 1228 7832
rect 1268 7792 2540 7832
rect 2500 7748 2540 7792
rect 2500 7708 11788 7748
rect 11828 7708 11837 7748
rect 31363 7708 31372 7748
rect 31412 7708 37132 7748
rect 37172 7708 37181 7748
rect 3679 7603 4065 7622
rect 3679 7580 3745 7603
rect 3831 7580 3913 7603
rect 3999 7580 4065 7603
rect 3679 7540 3688 7580
rect 3728 7540 3745 7580
rect 3831 7540 3852 7580
rect 3892 7540 3913 7580
rect 3999 7540 4016 7580
rect 4056 7540 4065 7580
rect 3679 7517 3745 7540
rect 3831 7517 3913 7540
rect 3999 7517 4065 7540
rect 3679 7498 4065 7517
rect 18799 7603 19185 7622
rect 18799 7580 18865 7603
rect 18951 7580 19033 7603
rect 19119 7580 19185 7603
rect 33919 7603 34305 7622
rect 33919 7580 33985 7603
rect 34071 7580 34153 7603
rect 34239 7580 34305 7603
rect 18799 7540 18808 7580
rect 18848 7540 18865 7580
rect 18951 7540 18972 7580
rect 19012 7540 19033 7580
rect 19119 7540 19136 7580
rect 19176 7540 19185 7580
rect 22627 7540 22636 7580
rect 22676 7540 32908 7580
rect 32948 7540 32957 7580
rect 33919 7540 33928 7580
rect 33968 7540 33985 7580
rect 34071 7540 34092 7580
rect 34132 7540 34153 7580
rect 34239 7540 34256 7580
rect 34296 7540 34305 7580
rect 18799 7517 18865 7540
rect 18951 7517 19033 7540
rect 19119 7517 19185 7540
rect 18799 7498 19185 7517
rect 33919 7517 33985 7540
rect 34071 7517 34153 7540
rect 34239 7517 34305 7540
rect 33919 7498 34305 7517
rect 27523 7204 27532 7244
rect 27572 7204 36556 7244
rect 36596 7204 36605 7244
rect 1507 7120 1516 7160
rect 1556 7120 11884 7160
rect 11924 7120 22636 7160
rect 22676 7120 22685 7160
rect 1795 7036 1804 7076
rect 1844 7036 14476 7076
rect 14516 7036 18508 7076
rect 18548 7036 20180 7076
rect 20140 6992 20180 7036
rect 13795 6952 13804 6992
rect 13844 6952 17740 6992
rect 17780 6952 17789 6992
rect 20140 6952 36556 6992
rect 36596 6952 36605 6992
rect 4919 6847 5305 6866
rect 4919 6824 4985 6847
rect 5071 6824 5153 6847
rect 5239 6824 5305 6847
rect 4919 6784 4928 6824
rect 4968 6784 4985 6824
rect 5071 6784 5092 6824
rect 5132 6784 5153 6824
rect 5239 6784 5256 6824
rect 5296 6784 5305 6824
rect 4919 6761 4985 6784
rect 5071 6761 5153 6784
rect 5239 6761 5305 6784
rect 4919 6742 5305 6761
rect 20039 6847 20425 6866
rect 20039 6824 20105 6847
rect 20191 6824 20273 6847
rect 20359 6824 20425 6847
rect 20039 6784 20048 6824
rect 20088 6784 20105 6824
rect 20191 6784 20212 6824
rect 20252 6784 20273 6824
rect 20359 6784 20376 6824
rect 20416 6784 20425 6824
rect 20039 6761 20105 6784
rect 20191 6761 20273 6784
rect 20359 6761 20425 6784
rect 20039 6742 20425 6761
rect 35159 6847 35545 6866
rect 35159 6824 35225 6847
rect 35311 6824 35393 6847
rect 35479 6824 35545 6847
rect 35159 6784 35168 6824
rect 35208 6784 35225 6824
rect 35311 6784 35332 6824
rect 35372 6784 35393 6824
rect 35479 6784 35496 6824
rect 35536 6784 35545 6824
rect 35159 6761 35225 6784
rect 35311 6761 35393 6784
rect 35479 6761 35545 6784
rect 35159 6742 35545 6761
rect 30403 6616 30412 6656
rect 30452 6616 40492 6656
rect 40532 6616 40541 6656
rect 2500 6532 13708 6572
rect 13748 6532 30700 6572
rect 30740 6532 34732 6572
rect 34772 6532 34781 6572
rect 2500 6488 2540 6532
rect 1699 6448 1708 6488
rect 1748 6448 2540 6488
rect 26947 6448 26956 6488
rect 26996 6448 30412 6488
rect 30452 6448 30461 6488
rect 16099 6364 16108 6404
rect 16148 6364 23116 6404
rect 23156 6364 23165 6404
rect 33283 6364 33292 6404
rect 33332 6364 41260 6404
rect 41300 6364 41309 6404
rect 17731 6196 17740 6236
rect 17780 6196 22636 6236
rect 22676 6196 22685 6236
rect 3679 6091 4065 6110
rect 3679 6068 3745 6091
rect 3831 6068 3913 6091
rect 3999 6068 4065 6091
rect 3679 6028 3688 6068
rect 3728 6028 3745 6068
rect 3831 6028 3852 6068
rect 3892 6028 3913 6068
rect 3999 6028 4016 6068
rect 4056 6028 4065 6068
rect 3679 6005 3745 6028
rect 3831 6005 3913 6028
rect 3999 6005 4065 6028
rect 3679 5986 4065 6005
rect 18799 6091 19185 6110
rect 18799 6068 18865 6091
rect 18951 6068 19033 6091
rect 19119 6068 19185 6091
rect 18799 6028 18808 6068
rect 18848 6028 18865 6068
rect 18951 6028 18972 6068
rect 19012 6028 19033 6068
rect 19119 6028 19136 6068
rect 19176 6028 19185 6068
rect 18799 6005 18865 6028
rect 18951 6005 19033 6028
rect 19119 6005 19185 6028
rect 18799 5986 19185 6005
rect 33919 6091 34305 6110
rect 33919 6068 33985 6091
rect 34071 6068 34153 6091
rect 34239 6068 34305 6091
rect 33919 6028 33928 6068
rect 33968 6028 33985 6068
rect 34071 6028 34092 6068
rect 34132 6028 34153 6068
rect 34239 6028 34256 6068
rect 34296 6028 34305 6068
rect 33919 6005 33985 6028
rect 34071 6005 34153 6028
rect 34239 6005 34305 6028
rect 33919 5986 34305 6005
rect 25315 5692 25324 5732
rect 25364 5692 35500 5732
rect 35540 5692 35549 5732
rect 18403 5608 18412 5648
rect 18452 5608 20180 5648
rect 20140 5564 20180 5608
rect 20140 5524 35308 5564
rect 35348 5524 35357 5564
rect 24067 5440 24076 5480
rect 24116 5440 36364 5480
rect 36404 5440 36413 5480
rect 4919 5335 5305 5354
rect 4919 5312 4985 5335
rect 5071 5312 5153 5335
rect 5239 5312 5305 5335
rect 4919 5272 4928 5312
rect 4968 5272 4985 5312
rect 5071 5272 5092 5312
rect 5132 5272 5153 5312
rect 5239 5272 5256 5312
rect 5296 5272 5305 5312
rect 4919 5249 4985 5272
rect 5071 5249 5153 5272
rect 5239 5249 5305 5272
rect 4919 5230 5305 5249
rect 20039 5335 20425 5354
rect 20039 5312 20105 5335
rect 20191 5312 20273 5335
rect 20359 5312 20425 5335
rect 20039 5272 20048 5312
rect 20088 5272 20105 5312
rect 20191 5272 20212 5312
rect 20252 5272 20273 5312
rect 20359 5272 20376 5312
rect 20416 5272 20425 5312
rect 20039 5249 20105 5272
rect 20191 5249 20273 5272
rect 20359 5249 20425 5272
rect 20039 5230 20425 5249
rect 35159 5335 35545 5354
rect 35159 5312 35225 5335
rect 35311 5312 35393 5335
rect 35479 5312 35545 5335
rect 35159 5272 35168 5312
rect 35208 5272 35225 5312
rect 35311 5272 35332 5312
rect 35372 5272 35393 5312
rect 35479 5272 35496 5312
rect 35536 5272 35545 5312
rect 35159 5249 35225 5272
rect 35311 5249 35393 5272
rect 35479 5249 35545 5272
rect 35159 5230 35545 5249
rect 17539 5104 17548 5144
rect 17588 5104 21772 5144
rect 21812 5104 21821 5144
rect 26659 5104 26668 5144
rect 26708 5104 37036 5144
rect 37076 5104 37085 5144
rect 13315 5020 13324 5060
rect 13364 5020 22060 5060
rect 22100 5020 27628 5060
rect 27668 5020 27677 5060
rect 5059 4936 5068 4976
rect 5108 4936 14860 4976
rect 14900 4936 14909 4976
rect 16268 4936 24556 4976
rect 24596 4936 24605 4976
rect 16268 4892 16308 4936
rect 7651 4852 7660 4892
rect 7700 4852 16204 4892
rect 16244 4852 16308 4892
rect 17155 4852 17164 4892
rect 17204 4852 21676 4892
rect 21716 4852 21725 4892
rect 1315 4768 1324 4808
rect 1364 4768 10252 4808
rect 10292 4768 10301 4808
rect 12547 4684 12556 4724
rect 12596 4684 33004 4724
rect 33044 4684 33053 4724
rect 3679 4579 4065 4598
rect 3679 4556 3745 4579
rect 3831 4556 3913 4579
rect 3999 4556 4065 4579
rect 3679 4516 3688 4556
rect 3728 4516 3745 4556
rect 3831 4516 3852 4556
rect 3892 4516 3913 4556
rect 3999 4516 4016 4556
rect 4056 4516 4065 4556
rect 3679 4493 3745 4516
rect 3831 4493 3913 4516
rect 3999 4493 4065 4516
rect 3679 4474 4065 4493
rect 18799 4579 19185 4598
rect 18799 4556 18865 4579
rect 18951 4556 19033 4579
rect 19119 4556 19185 4579
rect 18799 4516 18808 4556
rect 18848 4516 18865 4556
rect 18951 4516 18972 4556
rect 19012 4516 19033 4556
rect 19119 4516 19136 4556
rect 19176 4516 19185 4556
rect 18799 4493 18865 4516
rect 18951 4493 19033 4516
rect 19119 4493 19185 4516
rect 18799 4474 19185 4493
rect 33919 4579 34305 4598
rect 33919 4556 33985 4579
rect 34071 4556 34153 4579
rect 34239 4556 34305 4579
rect 33919 4516 33928 4556
rect 33968 4516 33985 4556
rect 34071 4516 34092 4556
rect 34132 4516 34153 4556
rect 34239 4516 34256 4556
rect 34296 4516 34305 4556
rect 33919 4493 33985 4516
rect 34071 4493 34153 4516
rect 34239 4493 34305 4516
rect 33919 4474 34305 4493
rect 20611 4264 20620 4304
rect 20660 4264 40300 4304
rect 40340 4264 40349 4304
rect 1795 4180 1804 4220
rect 1844 4180 28972 4220
rect 29012 4180 29021 4220
rect 20035 4096 20044 4136
rect 20084 4096 26956 4136
rect 26996 4096 27005 4136
rect 32995 4012 33004 4052
rect 33044 4012 37804 4052
rect 37844 4012 37853 4052
rect 355 3928 364 3968
rect 404 3928 7660 3968
rect 7700 3928 7709 3968
rect 27619 3928 27628 3968
rect 27668 3928 34252 3968
rect 34292 3928 34301 3968
rect 4919 3823 5305 3842
rect 4919 3800 4985 3823
rect 5071 3800 5153 3823
rect 5239 3800 5305 3823
rect 4919 3760 4928 3800
rect 4968 3760 4985 3800
rect 5071 3760 5092 3800
rect 5132 3760 5153 3800
rect 5239 3760 5256 3800
rect 5296 3760 5305 3800
rect 4919 3737 4985 3760
rect 5071 3737 5153 3760
rect 5239 3737 5305 3760
rect 4919 3718 5305 3737
rect 20039 3823 20425 3842
rect 20039 3800 20105 3823
rect 20191 3800 20273 3823
rect 20359 3800 20425 3823
rect 35159 3823 35545 3842
rect 35159 3800 35225 3823
rect 35311 3800 35393 3823
rect 35479 3800 35545 3823
rect 20039 3760 20048 3800
rect 20088 3760 20105 3800
rect 20191 3760 20212 3800
rect 20252 3760 20273 3800
rect 20359 3760 20376 3800
rect 20416 3760 20425 3800
rect 25027 3760 25036 3800
rect 25076 3760 31852 3800
rect 31892 3760 31901 3800
rect 35159 3760 35168 3800
rect 35208 3760 35225 3800
rect 35311 3760 35332 3800
rect 35372 3760 35393 3800
rect 35479 3760 35496 3800
rect 35536 3760 35545 3800
rect 20039 3737 20105 3760
rect 20191 3737 20273 3760
rect 20359 3737 20425 3760
rect 20039 3718 20425 3737
rect 35159 3737 35225 3760
rect 35311 3737 35393 3760
rect 35479 3737 35545 3760
rect 35159 3718 35545 3737
rect 12451 3508 12460 3548
rect 12500 3508 17644 3548
rect 17684 3508 20524 3548
rect 20564 3508 20573 3548
rect 10243 3424 10252 3464
rect 10292 3424 16012 3464
rect 16052 3424 22252 3464
rect 22292 3424 22301 3464
rect 17443 3256 17452 3296
rect 17492 3256 36076 3296
rect 36116 3256 36125 3296
rect 27523 3172 27532 3212
rect 27572 3172 36940 3212
rect 36980 3172 36989 3212
rect 3679 3067 4065 3086
rect 3679 3044 3745 3067
rect 3831 3044 3913 3067
rect 3999 3044 4065 3067
rect 3679 3004 3688 3044
rect 3728 3004 3745 3044
rect 3831 3004 3852 3044
rect 3892 3004 3913 3044
rect 3999 3004 4016 3044
rect 4056 3004 4065 3044
rect 3679 2981 3745 3004
rect 3831 2981 3913 3004
rect 3999 2981 4065 3004
rect 3679 2962 4065 2981
rect 18799 3067 19185 3086
rect 18799 3044 18865 3067
rect 18951 3044 19033 3067
rect 19119 3044 19185 3067
rect 18799 3004 18808 3044
rect 18848 3004 18865 3044
rect 18951 3004 18972 3044
rect 19012 3004 19033 3044
rect 19119 3004 19136 3044
rect 19176 3004 19185 3044
rect 18799 2981 18865 3004
rect 18951 2981 19033 3004
rect 19119 2981 19185 3004
rect 18799 2962 19185 2981
rect 33919 3067 34305 3086
rect 33919 3044 33985 3067
rect 34071 3044 34153 3067
rect 34239 3044 34305 3067
rect 33919 3004 33928 3044
rect 33968 3004 33985 3044
rect 34071 3004 34092 3044
rect 34132 3004 34153 3044
rect 34239 3004 34256 3044
rect 34296 3004 34305 3044
rect 33919 2981 33985 3004
rect 34071 2981 34153 3004
rect 34239 2981 34305 3004
rect 33919 2962 34305 2981
rect 12547 2836 12556 2876
rect 12596 2836 15244 2876
rect 15284 2836 15293 2876
rect 1411 2752 1420 2792
rect 1460 2752 29548 2792
rect 29588 2752 29597 2792
rect 3331 2668 3340 2708
rect 3380 2668 12460 2708
rect 12500 2668 12509 2708
rect 22243 2668 22252 2708
rect 22292 2668 41452 2708
rect 41492 2668 41501 2708
rect 19460 2584 19956 2624
rect 7171 2500 7180 2540
rect 7220 2500 8840 2540
rect 8800 2456 8840 2500
rect 19460 2456 19500 2584
rect 19916 2540 19956 2584
rect 20140 2584 22732 2624
rect 22772 2584 22781 2624
rect 24259 2584 24268 2624
rect 24308 2584 32716 2624
rect 32756 2584 32765 2624
rect 20140 2540 20180 2584
rect 19916 2500 19948 2540
rect 19988 2500 20180 2540
rect 8800 2416 19500 2456
rect 19916 2416 22828 2456
rect 22868 2416 22877 2456
rect 19916 2372 19956 2416
rect 15619 2332 15628 2372
rect 15668 2332 19956 2372
rect 4919 2311 5305 2330
rect 4919 2288 4985 2311
rect 5071 2288 5153 2311
rect 5239 2288 5305 2311
rect 4919 2248 4928 2288
rect 4968 2248 4985 2288
rect 5071 2248 5092 2288
rect 5132 2248 5153 2288
rect 5239 2248 5256 2288
rect 5296 2248 5305 2288
rect 4919 2225 4985 2248
rect 5071 2225 5153 2248
rect 5239 2225 5305 2248
rect 4919 2206 5305 2225
rect 20039 2311 20425 2330
rect 20039 2288 20105 2311
rect 20191 2288 20273 2311
rect 20359 2288 20425 2311
rect 20039 2248 20048 2288
rect 20088 2248 20105 2288
rect 20191 2248 20212 2288
rect 20252 2248 20273 2288
rect 20359 2248 20376 2288
rect 20416 2248 20425 2288
rect 20039 2225 20105 2248
rect 20191 2225 20273 2248
rect 20359 2225 20425 2248
rect 20039 2206 20425 2225
rect 35159 2311 35545 2330
rect 35159 2288 35225 2311
rect 35311 2288 35393 2311
rect 35479 2288 35545 2311
rect 35159 2248 35168 2288
rect 35208 2248 35225 2288
rect 35311 2248 35332 2288
rect 35372 2248 35393 2288
rect 35479 2248 35496 2288
rect 35536 2248 35545 2288
rect 35159 2225 35225 2248
rect 35311 2225 35393 2248
rect 35479 2225 35545 2248
rect 35159 2206 35545 2225
rect 19555 2080 19564 2120
rect 19604 2080 36076 2120
rect 36116 2080 36125 2120
rect 9571 1996 9580 2036
rect 9620 1996 31468 2036
rect 31508 1996 31517 2036
rect 1795 1912 1804 1952
rect 1844 1912 17452 1952
rect 17492 1912 17501 1952
rect 10531 1828 10540 1868
rect 10580 1828 28876 1868
rect 28916 1828 28925 1868
rect 16387 1744 16396 1784
rect 16436 1744 32716 1784
rect 32756 1744 32765 1784
rect 26467 1660 26476 1700
rect 26516 1660 40684 1700
rect 40724 1660 40733 1700
rect 3679 1555 4065 1574
rect 3679 1532 3745 1555
rect 3831 1532 3913 1555
rect 3999 1532 4065 1555
rect 3679 1492 3688 1532
rect 3728 1492 3745 1532
rect 3831 1492 3852 1532
rect 3892 1492 3913 1532
rect 3999 1492 4016 1532
rect 4056 1492 4065 1532
rect 3679 1469 3745 1492
rect 3831 1469 3913 1492
rect 3999 1469 4065 1492
rect 3679 1450 4065 1469
rect 18799 1555 19185 1574
rect 18799 1532 18865 1555
rect 18951 1532 19033 1555
rect 19119 1532 19185 1555
rect 18799 1492 18808 1532
rect 18848 1492 18865 1532
rect 18951 1492 18972 1532
rect 19012 1492 19033 1532
rect 19119 1492 19136 1532
rect 19176 1492 19185 1532
rect 18799 1469 18865 1492
rect 18951 1469 19033 1492
rect 19119 1469 19185 1492
rect 18799 1450 19185 1469
rect 33919 1555 34305 1574
rect 33919 1532 33985 1555
rect 34071 1532 34153 1555
rect 34239 1532 34305 1555
rect 33919 1492 33928 1532
rect 33968 1492 33985 1532
rect 34071 1492 34092 1532
rect 34132 1492 34153 1532
rect 34239 1492 34256 1532
rect 34296 1492 34305 1532
rect 33919 1469 33985 1492
rect 34071 1469 34153 1492
rect 34239 1469 34305 1492
rect 33919 1450 34305 1469
rect 29251 1324 29260 1364
rect 29300 1324 36844 1364
rect 36884 1324 36893 1364
rect 10243 1240 10252 1280
rect 10292 1240 28300 1280
rect 28340 1240 28349 1280
rect 8803 1156 8812 1196
rect 8852 1156 20716 1196
rect 20756 1156 28684 1196
rect 28724 1156 28733 1196
rect 12451 1072 12460 1112
rect 12500 1072 18124 1112
rect 18164 1072 33580 1112
rect 33620 1072 34444 1112
rect 34484 1072 34493 1112
rect 3619 988 3628 1028
rect 3668 988 11596 1028
rect 11636 988 25428 1028
rect 25507 988 25516 1028
rect 25556 988 35212 1028
rect 35252 988 35261 1028
rect 7939 904 7948 944
rect 7988 904 24516 944
rect 4919 799 5305 818
rect 4919 776 4985 799
rect 5071 776 5153 799
rect 5239 776 5305 799
rect 4919 736 4928 776
rect 4968 736 4985 776
rect 5071 736 5092 776
rect 5132 736 5153 776
rect 5239 736 5256 776
rect 5296 736 5305 776
rect 4919 713 4985 736
rect 5071 713 5153 736
rect 5239 713 5305 736
rect 4919 694 5305 713
rect 20039 799 20425 818
rect 20039 776 20105 799
rect 20191 776 20273 799
rect 20359 776 20425 799
rect 20039 736 20048 776
rect 20088 736 20105 776
rect 20191 736 20212 776
rect 20252 736 20273 776
rect 20359 736 20376 776
rect 20416 736 20425 776
rect 24476 776 24516 904
rect 25388 860 25428 988
rect 25388 820 27052 860
rect 27092 820 27101 860
rect 35159 799 35545 818
rect 35159 776 35225 799
rect 35311 776 35393 799
rect 35479 776 35545 799
rect 24476 736 25516 776
rect 25556 736 25565 776
rect 35159 736 35168 776
rect 35208 736 35225 776
rect 35311 736 35332 776
rect 35372 736 35393 776
rect 35479 736 35496 776
rect 35536 736 35545 776
rect 20039 713 20105 736
rect 20191 713 20273 736
rect 20359 713 20425 736
rect 20039 694 20425 713
rect 35159 713 35225 736
rect 35311 713 35393 736
rect 35479 713 35545 736
rect 35159 694 35545 713
rect 1795 568 1804 608
rect 1844 568 13420 608
rect 13460 568 13469 608
rect 16003 484 16012 524
rect 16052 484 20140 524
rect 20180 484 20189 524
rect 28099 232 28108 272
rect 28148 232 37900 272
rect 37940 232 37949 272
rect 14851 148 14860 188
rect 14900 148 26188 188
rect 26228 148 26237 188
rect 28675 148 28684 188
rect 28724 148 40396 188
rect 40436 148 40445 188
rect 24451 64 24460 104
rect 24500 64 37804 104
rect 37844 64 37853 104
<< via5 >>
rect 4985 9848 5071 9871
rect 5153 9848 5239 9871
rect 4985 9808 5010 9848
rect 5010 9808 5050 9848
rect 5050 9808 5071 9848
rect 5153 9808 5174 9848
rect 5174 9808 5214 9848
rect 5214 9808 5239 9848
rect 4985 9785 5071 9808
rect 5153 9785 5239 9808
rect 20105 9848 20191 9871
rect 20273 9848 20359 9871
rect 20105 9808 20130 9848
rect 20130 9808 20170 9848
rect 20170 9808 20191 9848
rect 20273 9808 20294 9848
rect 20294 9808 20334 9848
rect 20334 9808 20359 9848
rect 20105 9785 20191 9808
rect 20273 9785 20359 9808
rect 35225 9848 35311 9871
rect 35393 9848 35479 9871
rect 35225 9808 35250 9848
rect 35250 9808 35290 9848
rect 35290 9808 35311 9848
rect 35393 9808 35414 9848
rect 35414 9808 35454 9848
rect 35454 9808 35479 9848
rect 35225 9785 35311 9808
rect 35393 9785 35479 9808
rect 3745 9092 3831 9115
rect 3913 9092 3999 9115
rect 3745 9052 3770 9092
rect 3770 9052 3810 9092
rect 3810 9052 3831 9092
rect 3913 9052 3934 9092
rect 3934 9052 3974 9092
rect 3974 9052 3999 9092
rect 3745 9029 3831 9052
rect 3913 9029 3999 9052
rect 18865 9092 18951 9115
rect 19033 9092 19119 9115
rect 18865 9052 18890 9092
rect 18890 9052 18930 9092
rect 18930 9052 18951 9092
rect 19033 9052 19054 9092
rect 19054 9052 19094 9092
rect 19094 9052 19119 9092
rect 18865 9029 18951 9052
rect 19033 9029 19119 9052
rect 33985 9092 34071 9115
rect 34153 9092 34239 9115
rect 33985 9052 34010 9092
rect 34010 9052 34050 9092
rect 34050 9052 34071 9092
rect 34153 9052 34174 9092
rect 34174 9052 34214 9092
rect 34214 9052 34239 9092
rect 33985 9029 34071 9052
rect 34153 9029 34239 9052
rect 4985 8336 5071 8359
rect 5153 8336 5239 8359
rect 4985 8296 5010 8336
rect 5010 8296 5050 8336
rect 5050 8296 5071 8336
rect 5153 8296 5174 8336
rect 5174 8296 5214 8336
rect 5214 8296 5239 8336
rect 4985 8273 5071 8296
rect 5153 8273 5239 8296
rect 20105 8336 20191 8359
rect 20273 8336 20359 8359
rect 20105 8296 20130 8336
rect 20130 8296 20170 8336
rect 20170 8296 20191 8336
rect 20273 8296 20294 8336
rect 20294 8296 20334 8336
rect 20334 8296 20359 8336
rect 20105 8273 20191 8296
rect 20273 8273 20359 8296
rect 35225 8336 35311 8359
rect 35393 8336 35479 8359
rect 35225 8296 35250 8336
rect 35250 8296 35290 8336
rect 35290 8296 35311 8336
rect 35393 8296 35414 8336
rect 35414 8296 35454 8336
rect 35454 8296 35479 8336
rect 35225 8273 35311 8296
rect 35393 8273 35479 8296
rect 3745 7580 3831 7603
rect 3913 7580 3999 7603
rect 3745 7540 3770 7580
rect 3770 7540 3810 7580
rect 3810 7540 3831 7580
rect 3913 7540 3934 7580
rect 3934 7540 3974 7580
rect 3974 7540 3999 7580
rect 3745 7517 3831 7540
rect 3913 7517 3999 7540
rect 18865 7580 18951 7603
rect 19033 7580 19119 7603
rect 33985 7580 34071 7603
rect 34153 7580 34239 7603
rect 18865 7540 18890 7580
rect 18890 7540 18930 7580
rect 18930 7540 18951 7580
rect 19033 7540 19054 7580
rect 19054 7540 19094 7580
rect 19094 7540 19119 7580
rect 33985 7540 34010 7580
rect 34010 7540 34050 7580
rect 34050 7540 34071 7580
rect 34153 7540 34174 7580
rect 34174 7540 34214 7580
rect 34214 7540 34239 7580
rect 18865 7517 18951 7540
rect 19033 7517 19119 7540
rect 33985 7517 34071 7540
rect 34153 7517 34239 7540
rect 4985 6824 5071 6847
rect 5153 6824 5239 6847
rect 4985 6784 5010 6824
rect 5010 6784 5050 6824
rect 5050 6784 5071 6824
rect 5153 6784 5174 6824
rect 5174 6784 5214 6824
rect 5214 6784 5239 6824
rect 4985 6761 5071 6784
rect 5153 6761 5239 6784
rect 20105 6824 20191 6847
rect 20273 6824 20359 6847
rect 20105 6784 20130 6824
rect 20130 6784 20170 6824
rect 20170 6784 20191 6824
rect 20273 6784 20294 6824
rect 20294 6784 20334 6824
rect 20334 6784 20359 6824
rect 20105 6761 20191 6784
rect 20273 6761 20359 6784
rect 35225 6824 35311 6847
rect 35393 6824 35479 6847
rect 35225 6784 35250 6824
rect 35250 6784 35290 6824
rect 35290 6784 35311 6824
rect 35393 6784 35414 6824
rect 35414 6784 35454 6824
rect 35454 6784 35479 6824
rect 35225 6761 35311 6784
rect 35393 6761 35479 6784
rect 3745 6068 3831 6091
rect 3913 6068 3999 6091
rect 3745 6028 3770 6068
rect 3770 6028 3810 6068
rect 3810 6028 3831 6068
rect 3913 6028 3934 6068
rect 3934 6028 3974 6068
rect 3974 6028 3999 6068
rect 3745 6005 3831 6028
rect 3913 6005 3999 6028
rect 18865 6068 18951 6091
rect 19033 6068 19119 6091
rect 18865 6028 18890 6068
rect 18890 6028 18930 6068
rect 18930 6028 18951 6068
rect 19033 6028 19054 6068
rect 19054 6028 19094 6068
rect 19094 6028 19119 6068
rect 18865 6005 18951 6028
rect 19033 6005 19119 6028
rect 33985 6068 34071 6091
rect 34153 6068 34239 6091
rect 33985 6028 34010 6068
rect 34010 6028 34050 6068
rect 34050 6028 34071 6068
rect 34153 6028 34174 6068
rect 34174 6028 34214 6068
rect 34214 6028 34239 6068
rect 33985 6005 34071 6028
rect 34153 6005 34239 6028
rect 4985 5312 5071 5335
rect 5153 5312 5239 5335
rect 4985 5272 5010 5312
rect 5010 5272 5050 5312
rect 5050 5272 5071 5312
rect 5153 5272 5174 5312
rect 5174 5272 5214 5312
rect 5214 5272 5239 5312
rect 4985 5249 5071 5272
rect 5153 5249 5239 5272
rect 20105 5312 20191 5335
rect 20273 5312 20359 5335
rect 20105 5272 20130 5312
rect 20130 5272 20170 5312
rect 20170 5272 20191 5312
rect 20273 5272 20294 5312
rect 20294 5272 20334 5312
rect 20334 5272 20359 5312
rect 20105 5249 20191 5272
rect 20273 5249 20359 5272
rect 35225 5312 35311 5335
rect 35393 5312 35479 5335
rect 35225 5272 35250 5312
rect 35250 5272 35290 5312
rect 35290 5272 35311 5312
rect 35393 5272 35414 5312
rect 35414 5272 35454 5312
rect 35454 5272 35479 5312
rect 35225 5249 35311 5272
rect 35393 5249 35479 5272
rect 3745 4556 3831 4579
rect 3913 4556 3999 4579
rect 3745 4516 3770 4556
rect 3770 4516 3810 4556
rect 3810 4516 3831 4556
rect 3913 4516 3934 4556
rect 3934 4516 3974 4556
rect 3974 4516 3999 4556
rect 3745 4493 3831 4516
rect 3913 4493 3999 4516
rect 18865 4556 18951 4579
rect 19033 4556 19119 4579
rect 18865 4516 18890 4556
rect 18890 4516 18930 4556
rect 18930 4516 18951 4556
rect 19033 4516 19054 4556
rect 19054 4516 19094 4556
rect 19094 4516 19119 4556
rect 18865 4493 18951 4516
rect 19033 4493 19119 4516
rect 33985 4556 34071 4579
rect 34153 4556 34239 4579
rect 33985 4516 34010 4556
rect 34010 4516 34050 4556
rect 34050 4516 34071 4556
rect 34153 4516 34174 4556
rect 34174 4516 34214 4556
rect 34214 4516 34239 4556
rect 33985 4493 34071 4516
rect 34153 4493 34239 4516
rect 4985 3800 5071 3823
rect 5153 3800 5239 3823
rect 4985 3760 5010 3800
rect 5010 3760 5050 3800
rect 5050 3760 5071 3800
rect 5153 3760 5174 3800
rect 5174 3760 5214 3800
rect 5214 3760 5239 3800
rect 4985 3737 5071 3760
rect 5153 3737 5239 3760
rect 20105 3800 20191 3823
rect 20273 3800 20359 3823
rect 35225 3800 35311 3823
rect 35393 3800 35479 3823
rect 20105 3760 20130 3800
rect 20130 3760 20170 3800
rect 20170 3760 20191 3800
rect 20273 3760 20294 3800
rect 20294 3760 20334 3800
rect 20334 3760 20359 3800
rect 35225 3760 35250 3800
rect 35250 3760 35290 3800
rect 35290 3760 35311 3800
rect 35393 3760 35414 3800
rect 35414 3760 35454 3800
rect 35454 3760 35479 3800
rect 20105 3737 20191 3760
rect 20273 3737 20359 3760
rect 35225 3737 35311 3760
rect 35393 3737 35479 3760
rect 3745 3044 3831 3067
rect 3913 3044 3999 3067
rect 3745 3004 3770 3044
rect 3770 3004 3810 3044
rect 3810 3004 3831 3044
rect 3913 3004 3934 3044
rect 3934 3004 3974 3044
rect 3974 3004 3999 3044
rect 3745 2981 3831 3004
rect 3913 2981 3999 3004
rect 18865 3044 18951 3067
rect 19033 3044 19119 3067
rect 18865 3004 18890 3044
rect 18890 3004 18930 3044
rect 18930 3004 18951 3044
rect 19033 3004 19054 3044
rect 19054 3004 19094 3044
rect 19094 3004 19119 3044
rect 18865 2981 18951 3004
rect 19033 2981 19119 3004
rect 33985 3044 34071 3067
rect 34153 3044 34239 3067
rect 33985 3004 34010 3044
rect 34010 3004 34050 3044
rect 34050 3004 34071 3044
rect 34153 3004 34174 3044
rect 34174 3004 34214 3044
rect 34214 3004 34239 3044
rect 33985 2981 34071 3004
rect 34153 2981 34239 3004
rect 4985 2288 5071 2311
rect 5153 2288 5239 2311
rect 4985 2248 5010 2288
rect 5010 2248 5050 2288
rect 5050 2248 5071 2288
rect 5153 2248 5174 2288
rect 5174 2248 5214 2288
rect 5214 2248 5239 2288
rect 4985 2225 5071 2248
rect 5153 2225 5239 2248
rect 20105 2288 20191 2311
rect 20273 2288 20359 2311
rect 20105 2248 20130 2288
rect 20130 2248 20170 2288
rect 20170 2248 20191 2288
rect 20273 2248 20294 2288
rect 20294 2248 20334 2288
rect 20334 2248 20359 2288
rect 20105 2225 20191 2248
rect 20273 2225 20359 2248
rect 35225 2288 35311 2311
rect 35393 2288 35479 2311
rect 35225 2248 35250 2288
rect 35250 2248 35290 2288
rect 35290 2248 35311 2288
rect 35393 2248 35414 2288
rect 35414 2248 35454 2288
rect 35454 2248 35479 2288
rect 35225 2225 35311 2248
rect 35393 2225 35479 2248
rect 3745 1532 3831 1555
rect 3913 1532 3999 1555
rect 3745 1492 3770 1532
rect 3770 1492 3810 1532
rect 3810 1492 3831 1532
rect 3913 1492 3934 1532
rect 3934 1492 3974 1532
rect 3974 1492 3999 1532
rect 3745 1469 3831 1492
rect 3913 1469 3999 1492
rect 18865 1532 18951 1555
rect 19033 1532 19119 1555
rect 18865 1492 18890 1532
rect 18890 1492 18930 1532
rect 18930 1492 18951 1532
rect 19033 1492 19054 1532
rect 19054 1492 19094 1532
rect 19094 1492 19119 1532
rect 18865 1469 18951 1492
rect 19033 1469 19119 1492
rect 33985 1532 34071 1555
rect 34153 1532 34239 1555
rect 33985 1492 34010 1532
rect 34010 1492 34050 1532
rect 34050 1492 34071 1532
rect 34153 1492 34174 1532
rect 34174 1492 34214 1532
rect 34214 1492 34239 1532
rect 33985 1469 34071 1492
rect 34153 1469 34239 1492
rect 4985 776 5071 799
rect 5153 776 5239 799
rect 4985 736 5010 776
rect 5010 736 5050 776
rect 5050 736 5071 776
rect 5153 736 5174 776
rect 5174 736 5214 776
rect 5214 736 5239 776
rect 4985 713 5071 736
rect 5153 713 5239 736
rect 20105 776 20191 799
rect 20273 776 20359 799
rect 20105 736 20130 776
rect 20130 736 20170 776
rect 20170 736 20191 776
rect 20273 736 20294 776
rect 20294 736 20334 776
rect 20334 736 20359 776
rect 35225 776 35311 799
rect 35393 776 35479 799
rect 35225 736 35250 776
rect 35250 736 35290 776
rect 35290 736 35311 776
rect 35393 736 35414 776
rect 35414 736 35454 776
rect 35454 736 35479 776
rect 20105 713 20191 736
rect 20273 713 20359 736
rect 35225 713 35311 736
rect 35393 713 35479 736
<< metal6 >>
rect 3652 9115 4092 10752
rect 3652 9029 3745 9115
rect 3831 9029 3913 9115
rect 3999 9029 4092 9115
rect 3652 7603 4092 9029
rect 3652 7517 3745 7603
rect 3831 7517 3913 7603
rect 3999 7517 4092 7603
rect 3652 6091 4092 7517
rect 3652 6005 3745 6091
rect 3831 6005 3913 6091
rect 3999 6005 4092 6091
rect 3652 4579 4092 6005
rect 3652 4493 3745 4579
rect 3831 4493 3913 4579
rect 3999 4493 4092 4579
rect 3652 3067 4092 4493
rect 3652 2981 3745 3067
rect 3831 2981 3913 3067
rect 3999 2981 4092 3067
rect 3652 1555 4092 2981
rect 3652 1469 3745 1555
rect 3831 1469 3913 1555
rect 3999 1469 4092 1555
rect 3652 0 4092 1469
rect 4892 9871 5332 10752
rect 4892 9785 4985 9871
rect 5071 9785 5153 9871
rect 5239 9785 5332 9871
rect 4892 8359 5332 9785
rect 4892 8273 4985 8359
rect 5071 8273 5153 8359
rect 5239 8273 5332 8359
rect 4892 6847 5332 8273
rect 4892 6761 4985 6847
rect 5071 6761 5153 6847
rect 5239 6761 5332 6847
rect 4892 5335 5332 6761
rect 4892 5249 4985 5335
rect 5071 5249 5153 5335
rect 5239 5249 5332 5335
rect 4892 3823 5332 5249
rect 4892 3737 4985 3823
rect 5071 3737 5153 3823
rect 5239 3737 5332 3823
rect 4892 2311 5332 3737
rect 4892 2225 4985 2311
rect 5071 2225 5153 2311
rect 5239 2225 5332 2311
rect 4892 799 5332 2225
rect 4892 713 4985 799
rect 5071 713 5153 799
rect 5239 713 5332 799
rect 4892 0 5332 713
rect 18772 9115 19212 10752
rect 18772 9029 18865 9115
rect 18951 9029 19033 9115
rect 19119 9029 19212 9115
rect 18772 7603 19212 9029
rect 18772 7517 18865 7603
rect 18951 7517 19033 7603
rect 19119 7517 19212 7603
rect 18772 6091 19212 7517
rect 18772 6005 18865 6091
rect 18951 6005 19033 6091
rect 19119 6005 19212 6091
rect 18772 4579 19212 6005
rect 18772 4493 18865 4579
rect 18951 4493 19033 4579
rect 19119 4493 19212 4579
rect 18772 3067 19212 4493
rect 18772 2981 18865 3067
rect 18951 2981 19033 3067
rect 19119 2981 19212 3067
rect 18772 1555 19212 2981
rect 18772 1469 18865 1555
rect 18951 1469 19033 1555
rect 19119 1469 19212 1555
rect 18772 0 19212 1469
rect 20012 9871 20452 10752
rect 20012 9785 20105 9871
rect 20191 9785 20273 9871
rect 20359 9785 20452 9871
rect 20012 8359 20452 9785
rect 20012 8273 20105 8359
rect 20191 8273 20273 8359
rect 20359 8273 20452 8359
rect 20012 6847 20452 8273
rect 20012 6761 20105 6847
rect 20191 6761 20273 6847
rect 20359 6761 20452 6847
rect 20012 5335 20452 6761
rect 20012 5249 20105 5335
rect 20191 5249 20273 5335
rect 20359 5249 20452 5335
rect 20012 3823 20452 5249
rect 20012 3737 20105 3823
rect 20191 3737 20273 3823
rect 20359 3737 20452 3823
rect 20012 2311 20452 3737
rect 20012 2225 20105 2311
rect 20191 2225 20273 2311
rect 20359 2225 20452 2311
rect 20012 799 20452 2225
rect 20012 713 20105 799
rect 20191 713 20273 799
rect 20359 713 20452 799
rect 20012 0 20452 713
rect 33892 9115 34332 10752
rect 33892 9029 33985 9115
rect 34071 9029 34153 9115
rect 34239 9029 34332 9115
rect 33892 7603 34332 9029
rect 33892 7517 33985 7603
rect 34071 7517 34153 7603
rect 34239 7517 34332 7603
rect 33892 6091 34332 7517
rect 33892 6005 33985 6091
rect 34071 6005 34153 6091
rect 34239 6005 34332 6091
rect 33892 4579 34332 6005
rect 33892 4493 33985 4579
rect 34071 4493 34153 4579
rect 34239 4493 34332 4579
rect 33892 3067 34332 4493
rect 33892 2981 33985 3067
rect 34071 2981 34153 3067
rect 34239 2981 34332 3067
rect 33892 1555 34332 2981
rect 33892 1469 33985 1555
rect 34071 1469 34153 1555
rect 34239 1469 34332 1555
rect 33892 0 34332 1469
rect 35132 9871 35572 10752
rect 35132 9785 35225 9871
rect 35311 9785 35393 9871
rect 35479 9785 35572 9871
rect 35132 8359 35572 9785
rect 35132 8273 35225 8359
rect 35311 8273 35393 8359
rect 35479 8273 35572 8359
rect 35132 6847 35572 8273
rect 35132 6761 35225 6847
rect 35311 6761 35393 6847
rect 35479 6761 35572 6847
rect 35132 5335 35572 6761
rect 35132 5249 35225 5335
rect 35311 5249 35393 5335
rect 35479 5249 35572 5335
rect 35132 3823 35572 5249
rect 35132 3737 35225 3823
rect 35311 3737 35393 3823
rect 35479 3737 35572 3823
rect 35132 2311 35572 3737
rect 35132 2225 35225 2311
rect 35311 2225 35393 2311
rect 35479 2225 35572 2311
rect 35132 799 35572 2225
rect 35132 713 35225 799
rect 35311 713 35393 799
rect 35479 713 35572 799
rect 35132 0 35572 713
use sg13g2_inv_1  _083_
timestamp 1676382929
transform -1 0 7104 0 -1 9828
box -48 -56 336 834
use sg13g2_inv_1  _084_
timestamp 1676382929
transform -1 0 1440 0 1 6804
box -48 -56 336 834
use sg13g2_inv_1  _085_
timestamp 1676382929
transform 1 0 4896 0 -1 9828
box -48 -56 336 834
use sg13g2_inv_1  _086_
timestamp 1676382929
transform 1 0 10464 0 1 5292
box -48 -56 336 834
use sg13g2_mux4_1  _087_
timestamp 1677257233
transform 1 0 32160 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _088_
timestamp 1677257233
transform 1 0 16416 0 -1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _089_
timestamp 1677257233
transform 1 0 30240 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _090_
timestamp 1677257233
transform 1 0 17376 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _091_
timestamp 1677257233
transform 1 0 35136 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _092_
timestamp 1677257233
transform 1 0 13728 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _093_
timestamp 1677257233
transform 1 0 10656 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _094_
timestamp 1677257233
transform 1 0 9504 0 1 756
box -48 -56 2064 834
use sg13g2_mux4_1  _095_
timestamp 1677257233
transform 1 0 10560 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _096_
timestamp 1677257233
transform 1 0 10368 0 1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _097_
timestamp 1677257233
transform -1 0 4992 0 1 3780
box -48 -56 2064 834
use sg13g2_o21ai_1  _098_
timestamp 1685175443
transform -1 0 1728 0 1 2268
box -48 -56 538 834
use sg13g2_nor2_1  _099_
timestamp 1676627187
transform -1 0 4992 0 1 5292
box -48 -56 432 834
use sg13g2_nand2_1  _100_
timestamp 1676557249
transform 1 0 3264 0 1 5292
box -48 -56 432 834
use sg13g2_nand3_1  _101_
timestamp 1683988354
transform -1 0 5472 0 1 2268
box -48 -56 528 834
use sg13g2_o21ai_1  _102_
timestamp 1685175443
transform 1 0 3168 0 -1 3780
box -48 -56 538 834
use sg13g2_mux4_1  _103_
timestamp 1677257233
transform -1 0 4896 0 1 8316
box -48 -56 2064 834
use sg13g2_o21ai_1  _104_
timestamp 1685175443
transform -1 0 1728 0 -1 2268
box -48 -56 538 834
use sg13g2_nor2_1  _105_
timestamp 1676627187
transform -1 0 3456 0 1 6804
box -48 -56 432 834
use sg13g2_nand2_1  _106_
timestamp 1676557249
transform 1 0 4416 0 1 6804
box -48 -56 432 834
use sg13g2_nand3_1  _107_
timestamp 1683988354
transform -1 0 3936 0 1 756
box -48 -56 528 834
use sg13g2_o21ai_1  _108_
timestamp 1685175443
transform -1 0 1824 0 -1 9828
box -48 -56 538 834
use sg13g2_nand2b_1  _109_
timestamp 1676567195
transform 1 0 12384 0 1 8316
box -48 -56 528 834
use sg13g2_mux4_1  _110_
timestamp 1677257233
transform 1 0 10368 0 1 8316
box -48 -56 2064 834
use sg13g2_o21ai_1  _111_
timestamp 1685175443
transform 1 0 9408 0 1 8316
box -48 -56 538 834
use sg13g2_o21ai_1  _112_
timestamp 1685175443
transform -1 0 10272 0 -1 8316
box -48 -56 538 834
use sg13g2_nand2b_1  _113_
timestamp 1676567195
transform 1 0 9888 0 1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _114_
timestamp 1685175443
transform 1 0 11328 0 -1 6804
box -48 -56 538 834
use sg13g2_nand2b_1  _115_
timestamp 1676567195
transform -1 0 13344 0 1 8316
box -48 -56 528 834
use sg13g2_mux4_1  _116_
timestamp 1677257233
transform 1 0 13344 0 1 8316
box -48 -56 2064 834
use sg13g2_o21ai_1  _117_
timestamp 1685175443
transform -1 0 16320 0 -1 8316
box -48 -56 538 834
use sg13g2_o21ai_1  _118_
timestamp 1685175443
transform 1 0 13920 0 1 6804
box -48 -56 538 834
use sg13g2_nand2b_1  _119_
timestamp 1676567195
transform 1 0 15360 0 -1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _120_
timestamp 1685175443
transform 1 0 15360 0 1 8316
box -48 -56 538 834
use sg13g2_nand2_1  _121_
timestamp 1676557249
transform 1 0 9408 0 1 6804
box -48 -56 432 834
use sg13g2_nand2b_1  _122_
timestamp 1676567195
transform 1 0 7104 0 -1 9828
box -48 -56 528 834
use sg13g2_a21oi_1  _123_
timestamp 1683973020
transform 1 0 13440 0 1 6804
box -48 -56 528 834
use sg13g2_nor2b_1  _124_
timestamp 1685181386
transform -1 0 9408 0 1 6804
box -54 -56 528 834
use sg13g2_o21ai_1  _125_
timestamp 1685175443
transform 1 0 4512 0 -1 5292
box -48 -56 538 834
use sg13g2_o21ai_1  _126_
timestamp 1685175443
transform -1 0 8064 0 -1 9828
box -48 -56 538 834
use sg13g2_mux2_1  _127_
timestamp 1677247768
transform -1 0 9024 0 1 5292
box -48 -56 1008 834
use sg13g2_or2_1  _128_
timestamp 1684236171
transform -1 0 8544 0 -1 9828
box -48 -56 528 834
use sg13g2_a21oi_1  _129_
timestamp 1683973020
transform -1 0 6912 0 -1 6804
box -48 -56 528 834
use sg13g2_a221oi_1  _130_
timestamp 1685197497
transform 1 0 7584 0 -1 8316
box -48 -56 816 834
use sg13g2_o21ai_1  _131_
timestamp 1685175443
transform 1 0 8544 0 -1 9828
box -48 -56 538 834
use sg13g2_mux4_1  _132_
timestamp 1677257233
transform 1 0 6912 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _133_
timestamp 1677257233
transform 1 0 6912 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux2_1  _134_
timestamp 1677247768
transform 1 0 8352 0 -1 8316
box -48 -56 1008 834
use sg13g2_nand2b_1  _135_
timestamp 1676567195
transform 1 0 9024 0 -1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _136_
timestamp 1685175443
transform 1 0 9312 0 -1 8316
box -48 -56 538 834
use sg13g2_mux2_1  _137_
timestamp 1677247768
transform -1 0 4416 0 -1 6804
box -48 -56 1008 834
use sg13g2_mux2_1  _138_
timestamp 1677247768
transform -1 0 4416 0 -1 5292
box -48 -56 1008 834
use sg13g2_nand2b_1  _139_
timestamp 1676567195
transform -1 0 1632 0 -1 6804
box -48 -56 528 834
use sg13g2_a21oi_1  _140_
timestamp 1683973020
transform 1 0 2976 0 -1 5292
box -48 -56 528 834
use sg13g2_mux2_1  _141_
timestamp 1677247768
transform -1 0 4416 0 1 6804
box -48 -56 1008 834
use sg13g2_nand2b_1  _142_
timestamp 1676567195
transform 1 0 1824 0 -1 9828
box -48 -56 528 834
use sg13g2_mux2_1  _143_
timestamp 1677247768
transform -1 0 4608 0 1 5292
box -48 -56 1008 834
use sg13g2_a21oi_1  _144_
timestamp 1683973020
transform 1 0 1152 0 1 5292
box -48 -56 528 834
use sg13g2_a221oi_1  _145_
timestamp 1685197497
transform -1 0 4896 0 -1 9828
box -48 -56 816 834
use sg13g2_mux2_1  _146_
timestamp 1677247768
transform -1 0 6336 0 -1 6804
box -48 -56 1008 834
use sg13g2_mux2_1  _147_
timestamp 1677247768
transform 1 0 4416 0 -1 6804
box -48 -56 1008 834
use sg13g2_mux2_1  _148_
timestamp 1677247768
transform 1 0 4800 0 -1 8316
box -48 -56 1008 834
use sg13g2_mux2_1  _149_
timestamp 1677247768
transform 1 0 4992 0 1 5292
box -48 -56 1008 834
use sg13g2_mux4_1  _150_
timestamp 1677257233
transform 1 0 4800 0 1 6804
box -48 -56 2064 834
use sg13g2_a21o_1  _151_
timestamp 1677175127
transform -1 0 5760 0 1 8316
box -48 -56 720 834
use sg13g2_mux4_1  _152_
timestamp 1677257233
transform 1 0 6624 0 -1 5292
box -48 -56 2064 834
use sg13g2_mux2_1  _153_
timestamp 1677247768
transform 1 0 8160 0 1 3780
box -48 -56 1008 834
use sg13g2_nor2b_1  _154_
timestamp 1685181386
transform -1 0 5472 0 1 3780
box -54 -56 528 834
use sg13g2_o21ai_1  _155_
timestamp 1685175443
transform -1 0 7680 0 -1 2268
box -48 -56 538 834
use sg13g2_o21ai_1  _156_
timestamp 1685175443
transform 1 0 5472 0 1 3780
box -48 -56 538 834
use sg13g2_a21oi_1  _157_
timestamp 1683973020
transform 1 0 9984 0 1 5292
box -48 -56 528 834
use sg13g2_o21ai_1  _158_
timestamp 1685175443
transform 1 0 8928 0 -1 6804
box -48 -56 538 834
use sg13g2_mux4_1  _159_
timestamp 1677257233
transform 1 0 5952 0 1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _160_
timestamp 1677257233
transform 1 0 5952 0 1 3780
box -48 -56 2064 834
use sg13g2_mux2_1  _161_
timestamp 1677247768
transform 1 0 7776 0 -1 3780
box -48 -56 1008 834
use sg13g2_nand2b_1  _162_
timestamp 1676567195
transform 1 0 9024 0 1 5292
box -48 -56 528 834
use sg13g2_o21ai_1  _163_
timestamp 1685175443
transform -1 0 9984 0 1 5292
box -48 -56 538 834
use sg13g2_mux2_1  _164_
timestamp 1677247768
transform -1 0 4896 0 1 756
box -48 -56 1008 834
use sg13g2_or2_1  _165_
timestamp 1684236171
transform -1 0 13632 0 -1 2268
box -48 -56 528 834
use sg13g2_a21oi_1  _166_
timestamp 1683973020
transform -1 0 1728 0 1 756
box -48 -56 528 834
use sg13g2_a221oi_1  _167_
timestamp 1685197497
transform 1 0 3648 0 -1 3780
box -48 -56 816 834
use sg13g2_nor2b_1  _168_
timestamp 1685181386
transform -1 0 14976 0 1 2268
box -54 -56 528 834
use sg13g2_o21ai_1  _169_
timestamp 1685175443
transform 1 0 12000 0 -1 5292
box -48 -56 538 834
use sg13g2_nand2_1  _170_
timestamp 1676557249
transform 1 0 1152 0 -1 3780
box -48 -56 432 834
use sg13g2_nand2b_1  _171_
timestamp 1676567195
transform 1 0 14976 0 1 756
box -48 -56 528 834
use sg13g2_a21oi_1  _172_
timestamp 1683973020
transform 1 0 14976 0 1 2268
box -48 -56 528 834
use sg13g2_o21ai_1  _173_
timestamp 1685175443
transform -1 0 14496 0 1 2268
box -48 -56 538 834
use sg13g2_o21ai_1  _174_
timestamp 1685175443
transform -1 0 13152 0 -1 2268
box -48 -56 538 834
use sg13g2_mux4_1  _175_
timestamp 1677257233
transform 1 0 4992 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _176_
timestamp 1677257233
transform 1 0 4896 0 1 756
box -48 -56 2064 834
use sg13g2_mux2_1  _177_
timestamp 1677247768
transform 1 0 6912 0 1 756
box -48 -56 1008 834
use sg13g2_nand2b_1  _178_
timestamp 1676567195
transform -1 0 10656 0 -1 2268
box -48 -56 528 834
use sg13g2_o21ai_1  _179_
timestamp 1685175443
transform 1 0 9696 0 -1 2268
box -48 -56 538 834
use sg13g2_mux4_1  _180_
timestamp 1677257233
transform 1 0 7680 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _181_
timestamp 1677257233
transform 1 0 28800 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _182_
timestamp 1677257233
transform 1 0 27936 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _183_
timestamp 1677257233
transform 1 0 26688 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _184_
timestamp 1677257233
transform 1 0 38592 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _185_
timestamp 1677257233
transform 1 0 32256 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _186_
timestamp 1677257233
transform 1 0 26880 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _187_
timestamp 1677257233
transform 1 0 38400 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _188_
timestamp 1677257233
transform 1 0 13440 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _189_
timestamp 1677257233
transform 1 0 29856 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _190_
timestamp 1677257233
transform 1 0 12480 0 1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _191_
timestamp 1677257233
transform 1 0 24096 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _192_
timestamp 1677257233
transform 1 0 28032 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _193_
timestamp 1677257233
transform 1 0 12960 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _194_
timestamp 1677257233
transform 1 0 38592 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _195_
timestamp 1677257233
transform 1 0 32064 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _196_
timestamp 1677257233
transform 1 0 34176 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _197_
timestamp 1677257233
transform 1 0 26016 0 1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _198_
timestamp 1677257233
transform 1 0 29184 0 1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _199_
timestamp 1677257233
transform 1 0 24960 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _200_
timestamp 1677257233
transform 1 0 35712 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _201_
timestamp 1677257233
transform 1 0 22848 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _202_
timestamp 1677257233
transform 1 0 24192 0 1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _203_
timestamp 1677257233
transform 1 0 17952 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _204_
timestamp 1677257233
transform 1 0 32160 0 1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _205_
timestamp 1677257233
transform 1 0 22944 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _206_
timestamp 1677257233
transform 1 0 37344 0 1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _207_
timestamp 1677257233
transform 1 0 25344 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _208_
timestamp 1677257233
transform 1 0 37248 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _209_
timestamp 1677257233
transform 1 0 21792 0 1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _210_
timestamp 1677257233
transform 1 0 36576 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _211_
timestamp 1677257233
transform 1 0 17952 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _212_
timestamp 1677257233
transform 1 0 24096 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _213_
timestamp 1677257233
transform 1 0 21216 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _214_
timestamp 1677257233
transform 1 0 21600 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _215_
timestamp 1677257233
transform 1 0 20448 0 1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _216_
timestamp 1677257233
transform 1 0 21024 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _217_
timestamp 1677257233
transform 1 0 17760 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _218_
timestamp 1677257233
transform 1 0 17760 0 1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _219_
timestamp 1677257233
transform 1 0 14016 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _220_
timestamp 1677257233
transform 1 0 34272 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _221_
timestamp 1677257233
transform 1 0 16416 0 -1 8316
box -48 -56 2064 834
use sg13g2_dlhq_1  _222_
timestamp 1678805552
transform 1 0 10368 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _223_
timestamp 1678805552
transform 1 0 9504 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _224_
timestamp 1678805552
transform 1 0 8928 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _225_
timestamp 1678805552
transform 1 0 9120 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _226_
timestamp 1678805552
transform 1 0 7104 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _227_
timestamp 1678805552
transform 1 0 8736 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _228_
timestamp 1678805552
transform 1 0 7872 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _229_
timestamp 1678805552
transform 1 0 11520 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _230_
timestamp 1678805552
transform 1 0 12384 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _231_
timestamp 1678805552
transform 1 0 13344 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _232_
timestamp 1678805552
transform -1 0 36192 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _233_
timestamp 1678805552
transform 1 0 34848 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _234_
timestamp 1678805552
transform 1 0 15936 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _235_
timestamp 1678805552
transform 1 0 17568 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _236_
timestamp 1678805552
transform -1 0 31584 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _237_
timestamp 1678805552
transform -1 0 32928 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _238_
timestamp 1678805552
transform 1 0 14784 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _239_
timestamp 1678805552
transform 1 0 16128 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _240_
timestamp 1678805552
transform 1 0 31200 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _241_
timestamp 1678805552
transform 1 0 32928 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _242_
timestamp 1678805552
transform 1 0 14688 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _243_
timestamp 1678805552
transform 1 0 16128 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _244_
timestamp 1678805552
transform 1 0 33120 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _245_
timestamp 1678805552
transform 1 0 34656 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _246_
timestamp 1678805552
transform 1 0 14400 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _247_
timestamp 1678805552
transform 1 0 11808 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _248_
timestamp 1678805552
transform 1 0 17664 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _249_
timestamp 1678805552
transform 1 0 16032 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _250_
timestamp 1678805552
transform 1 0 18048 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _251_
timestamp 1678805552
transform 1 0 16320 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _252_
timestamp 1678805552
transform 1 0 21312 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _253_
timestamp 1678805552
transform 1 0 19680 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _254_
timestamp 1678805552
transform 1 0 20736 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _255_
timestamp 1678805552
transform 1 0 19296 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _256_
timestamp 1678805552
transform 1 0 19968 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _257_
timestamp 1678805552
transform 1 0 21984 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _258_
timestamp 1678805552
transform 1 0 19968 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _259_
timestamp 1678805552
transform 1 0 20640 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _260_
timestamp 1678805552
transform -1 0 25536 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _261_
timestamp 1678805552
transform -1 0 27168 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _262_
timestamp 1678805552
transform 1 0 18048 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _263_
timestamp 1678805552
transform 1 0 16320 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _264_
timestamp 1678805552
transform -1 0 39744 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _265_
timestamp 1678805552
transform -1 0 38592 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _266_
timestamp 1678805552
transform 1 0 22272 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _267_
timestamp 1678805552
transform 1 0 20448 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _268_
timestamp 1678805552
transform -1 0 40128 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _269_
timestamp 1678805552
transform 1 0 36480 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _270_
timestamp 1678805552
transform 1 0 24192 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _271_
timestamp 1678805552
transform 1 0 26112 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _272_
timestamp 1678805552
transform -1 0 38496 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _273_
timestamp 1678805552
transform 1 0 37728 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _274_
timestamp 1678805552
transform 1 0 21312 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _275_
timestamp 1678805552
transform 1 0 23424 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _276_
timestamp 1678805552
transform 1 0 32832 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _277_
timestamp 1678805552
transform 1 0 30624 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _278_
timestamp 1678805552
transform 1 0 18432 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _279_
timestamp 1678805552
transform 1 0 16032 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _280_
timestamp 1678805552
transform 1 0 24864 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _281_
timestamp 1678805552
transform 1 0 23040 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _282_
timestamp 1678805552
transform 1 0 21216 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _283_
timestamp 1678805552
transform 1 0 23136 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _284_
timestamp 1678805552
transform 1 0 34848 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _285_
timestamp 1678805552
transform -1 0 38496 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _286_
timestamp 1678805552
transform -1 0 26400 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _287_
timestamp 1678805552
transform -1 0 28032 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _288_
timestamp 1678805552
transform -1 0 30528 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _289_
timestamp 1678805552
transform 1 0 29568 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _290_
timestamp 1678805552
transform -1 0 27744 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _291_
timestamp 1678805552
transform -1 0 28800 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _292_
timestamp 1678805552
transform -1 0 35328 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _293_
timestamp 1678805552
transform -1 0 36960 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _294_
timestamp 1678805552
transform -1 0 33696 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _295_
timestamp 1678805552
transform 1 0 32928 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _296_
timestamp 1678805552
transform -1 0 40224 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _297_
timestamp 1678805552
transform -1 0 41376 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _298_
timestamp 1678805552
transform 1 0 10752 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _299_
timestamp 1678805552
transform 1 0 12384 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _300_
timestamp 1678805552
transform -1 0 29664 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _301_
timestamp 1678805552
transform -1 0 31296 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _302_
timestamp 1678805552
transform 1 0 23040 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _303_
timestamp 1678805552
transform 1 0 24480 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _304_
timestamp 1678805552
transform 1 0 10848 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _305_
timestamp 1678805552
transform 1 0 12480 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _306_
timestamp 1678805552
transform 1 0 30528 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _307_
timestamp 1678805552
transform 1 0 28896 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _308_
timestamp 1678805552
transform 1 0 11808 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _309_
timestamp 1678805552
transform 1 0 13728 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _310_
timestamp 1678805552
transform 1 0 37248 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _311_
timestamp 1678805552
transform 1 0 39072 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _312_
timestamp 1678805552
transform 1 0 25824 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _313_
timestamp 1678805552
transform 1 0 27456 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _314_
timestamp 1678805552
transform -1 0 33792 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _315_
timestamp 1678805552
transform 1 0 32832 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _316_
timestamp 1678805552
transform 1 0 37632 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _317_
timestamp 1678805552
transform 1 0 39072 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _318_
timestamp 1678805552
transform -1 0 29664 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _319_
timestamp 1678805552
transform 1 0 25056 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _320_
timestamp 1678805552
transform 1 0 26880 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _321_
timestamp 1678805552
transform 1 0 27552 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _322_
timestamp 1678805552
transform -1 0 30432 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _323_
timestamp 1678805552
transform -1 0 32064 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _324_
timestamp 1678805552
transform 1 0 5472 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _325_
timestamp 1678805552
transform 1 0 3360 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _326_
timestamp 1678805552
transform 1 0 3360 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _327_
timestamp 1678805552
transform 1 0 1728 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _328_
timestamp 1678805552
transform 1 0 1728 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _329_
timestamp 1678805552
transform 1 0 1728 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _330_
timestamp 1678805552
transform 1 0 1248 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _331_
timestamp 1678805552
transform 1 0 1536 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _332_
timestamp 1678805552
transform 1 0 1344 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _333_
timestamp 1678805552
transform 1 0 4416 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _334_
timestamp 1678805552
transform 1 0 4992 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _335_
timestamp 1678805552
transform -1 0 7776 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _336_
timestamp 1678805552
transform -1 0 10272 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _337_
timestamp 1678805552
transform -1 0 4608 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _338_
timestamp 1678805552
transform 1 0 1248 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _339_
timestamp 1678805552
transform 1 0 2304 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _340_
timestamp 1678805552
transform 1 0 1440 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _341_
timestamp 1678805552
transform 1 0 1632 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _342_
timestamp 1678805552
transform 1 0 1632 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _343_
timestamp 1678805552
transform 1 0 1344 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _344_
timestamp 1678805552
transform -1 0 11424 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _345_
timestamp 1678805552
transform -1 0 11904 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _346_
timestamp 1678805552
transform 1 0 9792 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _347_
timestamp 1678805552
transform -1 0 6816 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _348_
timestamp 1678805552
transform 1 0 5760 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _349_
timestamp 1678805552
transform 1 0 6048 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _350_
timestamp 1678805552
transform 1 0 7680 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _351_
timestamp 1678805552
transform 1 0 11424 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _352_
timestamp 1678805552
transform 1 0 12096 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _353_
timestamp 1678805552
transform 1 0 13056 0 -1 9828
box -50 -56 1692 834
use sg13g2_dfrbpq_1  _354_
timestamp 1746535128
transform -1 0 30144 0 1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _355_
timestamp 1746535128
transform -1 0 36480 0 -1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _356_
timestamp 1746535128
transform 1 0 31488 0 1 8316
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _357_
timestamp 1746535128
transform -1 0 36864 0 1 8316
box -48 -56 2640 834
use sg13g2_tiehi  _358_
timestamp 1680000651
transform -1 0 38112 0 -1 8316
box -48 -56 432 834
use sg13g2_tiehi  _359_
timestamp 1680000651
transform -1 0 37056 0 -1 6804
box -48 -56 432 834
use sg13g2_tiehi  _360_
timestamp 1680000651
transform -1 0 29856 0 1 6804
box -48 -56 432 834
use sg13g2_tiehi  _361_
timestamp 1680000651
transform -1 0 36672 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _362_
timestamp 1676381911
transform 1 0 41184 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _363_
timestamp 1676381911
transform 1 0 40032 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _364_
timestamp 1676381911
transform 1 0 39648 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _365_
timestamp 1676381911
transform 1 0 39264 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _366_
timestamp 1676381911
transform 1 0 39840 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _367_
timestamp 1676381911
transform 1 0 40800 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _368_
timestamp 1676381911
transform 1 0 41376 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _369_
timestamp 1676381911
transform 1 0 40992 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _370_
timestamp 1676381911
transform 1 0 41376 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _371_
timestamp 1676381911
transform 1 0 41184 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _372_
timestamp 1676381911
transform 1 0 40416 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _373_
timestamp 1676381911
transform 1 0 40800 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _374_
timestamp 1676381911
transform 1 0 41184 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _375_
timestamp 1676381911
transform 1 0 40800 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _376_
timestamp 1676381911
transform 1 0 40416 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _377_
timestamp 1676381911
transform 1 0 40800 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _378_
timestamp 1676381911
transform 1 0 40416 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _379_
timestamp 1676381911
transform 1 0 40800 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _380_
timestamp 1676381911
transform 1 0 41184 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _381_
timestamp 1676381911
transform 1 0 40800 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _382_
timestamp 1676381911
transform 1 0 40800 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _383_
timestamp 1676381911
transform 1 0 41184 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _384_
timestamp 1676381911
transform 1 0 40992 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _385_
timestamp 1676381911
transform 1 0 41376 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _386_
timestamp 1676381911
transform 1 0 40800 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _387_
timestamp 1676381911
transform 1 0 41184 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _388_
timestamp 1676381911
transform 1 0 41184 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _389_
timestamp 1676381911
transform 1 0 41184 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _390_
timestamp 1676381911
transform 1 0 41184 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _391_
timestamp 1676381911
transform 1 0 40800 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _392_
timestamp 1676381911
transform 1 0 40416 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _393_
timestamp 1676381911
transform 1 0 40608 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _394_
timestamp 1676381911
transform 1 0 15648 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _395_
timestamp 1676381911
transform -1 0 20352 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _396_
timestamp 1676381911
transform 1 0 19968 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _397_
timestamp 1676381911
transform 1 0 20832 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _398_
timestamp 1676381911
transform -1 0 22752 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _399_
timestamp 1676381911
transform -1 0 32640 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _400_
timestamp 1676381911
transform -1 0 31968 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _401_
timestamp 1676381911
transform -1 0 36864 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _402_
timestamp 1676381911
transform -1 0 37248 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _403_
timestamp 1676381911
transform -1 0 34848 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _404_
timestamp 1676381911
transform -1 0 37632 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _405_
timestamp 1676381911
transform -1 0 32640 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _406_
timestamp 1676381911
transform -1 0 38880 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _407_
timestamp 1676381911
transform -1 0 34560 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _408_
timestamp 1676381911
transform -1 0 39648 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _409_
timestamp 1676381911
transform -1 0 35520 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _410_
timestamp 1676381911
transform -1 0 38496 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _411_
timestamp 1676381911
transform -1 0 38112 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _412_
timestamp 1676381911
transform -1 0 40032 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _413_
timestamp 1676381911
transform -1 0 40416 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _414_
timestamp 1676381911
transform 1 0 15456 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _415_
timestamp 1676381911
transform 1 0 12576 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _416_
timestamp 1676381911
transform 1 0 15456 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _417_
timestamp 1676381911
transform 1 0 15744 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _418_
timestamp 1676381911
transform 1 0 15840 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _419_
timestamp 1676381911
transform -1 0 40608 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _420_
timestamp 1676381911
transform 1 0 19872 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _421_
timestamp 1676381911
transform -1 0 32160 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _422_
timestamp 1676381911
transform 1 0 20160 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _423_
timestamp 1676381911
transform -1 0 34560 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _424_
timestamp 1676381911
transform 1 0 20448 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _425_
timestamp 1676381911
transform -1 0 36672 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _426_
timestamp 1676381911
transform 1 0 20832 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _427_
timestamp 1676381911
transform 1 0 20928 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _428_
timestamp 1676381911
transform 1 0 20352 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _429_
timestamp 1676381911
transform -1 0 22944 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _430_
timestamp 1676381911
transform -1 0 23328 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _431_
timestamp 1676381911
transform 1 0 22656 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _432_
timestamp 1676381911
transform -1 0 24000 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _433_
timestamp 1676381911
transform -1 0 25344 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _434_
timestamp 1676381911
transform 1 0 23232 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _435_
timestamp 1676381911
transform -1 0 37248 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _436_
timestamp 1676381911
transform -1 0 24192 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _437_
timestamp 1676381911
transform -1 0 40992 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _438_
timestamp 1676381911
transform -1 0 28512 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _439_
timestamp 1676381911
transform -1 0 39744 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _440_
timestamp 1676381911
transform -1 0 25344 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _441_
timestamp 1676381911
transform -1 0 35136 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _442_
timestamp 1676381911
transform 1 0 23808 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _443_
timestamp 1676381911
transform -1 0 26592 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _444_
timestamp 1676381911
transform -1 0 25728 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _445_
timestamp 1676381911
transform -1 0 37344 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _446_
timestamp 1676381911
transform -1 0 27360 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _447_
timestamp 1676381911
transform -1 0 31584 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _448_
timestamp 1676381911
transform -1 0 31200 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _449_
timestamp 1676381911
transform -1 0 36576 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _450_
timestamp 1676381911
transform -1 0 37536 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _451_
timestamp 1676381911
transform -1 0 40608 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _452_
timestamp 1676381911
transform -1 0 27744 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _453_
timestamp 1676381911
transform -1 0 29568 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _454_
timestamp 1676381911
transform -1 0 28128 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _455_
timestamp 1676381911
transform 1 0 26496 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _456_
timestamp 1676381911
transform -1 0 32256 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _457_
timestamp 1676381911
transform 1 0 27072 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _458_
timestamp 1676381911
transform -1 0 40224 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _459_
timestamp 1676381911
transform -1 0 28896 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _460_
timestamp 1676381911
transform -1 0 35136 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _461_
timestamp 1676381911
transform -1 0 40800 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _462_
timestamp 1676381911
transform -1 0 29472 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _463_
timestamp 1676381911
transform -1 0 36576 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _464_
timestamp 1676381911
transform -1 0 32064 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _465_
timestamp 1676381911
transform -1 0 31584 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _466_
timestamp 1676381911
transform -1 0 32544 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_8  clkbuf_0_UserCLK
timestamp 1676451365
transform -1 0 32160 0 -1 9828
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_0_UserCLK_regs
timestamp 1676451365
transform -1 0 35712 0 1 6804
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_1_0__f_UserCLK_regs
timestamp 1676451365
transform -1 0 30912 0 -1 9828
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_1_0__f_UserCLK
timestamp 1676451365
transform -1 0 31392 0 1 8316
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_1_1__f_UserCLK_regs
timestamp 1676451365
transform 1 0 35616 0 -1 5292
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_regs_0_UserCLK
timestamp 1676451365
transform 1 0 36480 0 -1 8316
box -48 -56 1296 834
use sg13g2_fill_1  FILLER_0_0
timestamp 1677579658
transform 1 0 1152 0 1 756
box -48 -56 144 834
use sg13g2_fill_1  FILLER_0_23
timestamp 1677579658
transform 1 0 3360 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_125
timestamp 1677580104
transform 1 0 13152 0 1 756
box -48 -56 240 834
use sg13g2_decap_8  FILLER_0_153
timestamp 1679581782
transform 1 0 15840 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_160
timestamp 1679581782
transform 1 0 16512 0 1 756
box -48 -56 720 834
use sg13g2_decap_8  FILLER_0_167
timestamp 1679581782
transform 1 0 17184 0 1 756
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_174
timestamp 1677580104
transform 1 0 17856 0 1 756
box -48 -56 240 834
use sg13g2_decap_8  FILLER_0_193
timestamp 1679581782
transform 1 0 19680 0 1 756
box -48 -56 720 834
use sg13g2_fill_2  FILLER_0_200
timestamp 1677580104
transform 1 0 20352 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_202
timestamp 1677579658
transform 1 0 20544 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_411
timestamp 1677580104
transform 1 0 40608 0 1 756
box -48 -56 240 834
use sg13g2_fill_2  FILLER_0_421
timestamp 1677580104
transform 1 0 41568 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_423
timestamp 1677579658
transform 1 0 41760 0 1 756
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_0
timestamp 1677579658
transform 1 0 1152 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_61
timestamp 1677580104
transform 1 0 7008 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_130
timestamp 1677579658
transform 1 0 13632 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_156
timestamp 1677580104
transform 1 0 16128 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_8  FILLER_1_196
timestamp 1679581782
transform 1 0 19968 0 -1 2268
box -48 -56 720 834
use sg13g2_fill_2  FILLER_1_203
timestamp 1677580104
transform 1 0 20640 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_238
timestamp 1677579658
transform 1 0 24000 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_285
timestamp 1677580104
transform 1 0 28512 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_287
timestamp 1677579658
transform 1 0 28704 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_317
timestamp 1677579658
transform 1 0 31584 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_343
timestamp 1677579658
transform 1 0 34080 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_423
timestamp 1677579658
transform 1 0 41760 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_0
timestamp 1677579658
transform 1 0 1152 0 1 2268
box -48 -56 144 834
use sg13g2_decap_8  FILLER_2_157
timestamp 1679581782
transform 1 0 16224 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_164
timestamp 1679581782
transform 1 0 16896 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_171
timestamp 1679581782
transform 1 0 17568 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_178
timestamp 1679581782
transform 1 0 18240 0 1 2268
box -48 -56 720 834
use sg13g2_decap_8  FILLER_2_185
timestamp 1679581782
transform 1 0 18912 0 1 2268
box -48 -56 720 834
use sg13g2_decap_4  FILLER_2_192
timestamp 1679577901
transform 1 0 19584 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_213
timestamp 1677580104
transform 1 0 21600 0 1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_257
timestamp 1677580104
transform 1 0 25824 0 1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_348
timestamp 1677580104
transform 1 0 34560 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_350
timestamp 1677579658
transform 1 0 34752 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_423
timestamp 1677579658
transform 1 0 41760 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_51
timestamp 1677579658
transform 1 0 6048 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_79
timestamp 1677580104
transform 1 0 8736 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_3_144
timestamp 1679581782
transform 1 0 14976 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_151
timestamp 1677580104
transform 1 0 15648 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_153
timestamp 1677579658
transform 1 0 15840 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_3_188
timestamp 1679581782
transform 1 0 19200 0 -1 3780
box -48 -56 720 834
use sg13g2_fill_2  FILLER_3_199
timestamp 1677580104
transform 1 0 20256 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_4  FILLER_3_218
timestamp 1679577901
transform 1 0 22080 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_222
timestamp 1677580104
transform 1 0 22464 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_245
timestamp 1677580104
transform 1 0 24672 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_247
timestamp 1677579658
transform 1 0 24864 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_277
timestamp 1677580104
transform 1 0 27744 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_279
timestamp 1677579658
transform 1 0 27936 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_301
timestamp 1677580104
transform 1 0 30048 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_328
timestamp 1677580104
transform 1 0 32640 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_330
timestamp 1677579658
transform 1 0 32832 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_369
timestamp 1677580104
transform 1 0 36576 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_371
timestamp 1677579658
transform 1 0 36768 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_421
timestamp 1677580104
transform 1 0 41568 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_423
timestamp 1677579658
transform 1 0 41760 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_0
timestamp 1677580104
transform 1 0 1152 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_71
timestamp 1677580104
transform 1 0 7968 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_155
timestamp 1679581782
transform 1 0 16032 0 1 3780
box -48 -56 720 834
use sg13g2_decap_8  FILLER_4_162
timestamp 1679581782
transform 1 0 16704 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_190
timestamp 1679577901
transform 1 0 19392 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_194
timestamp 1677580104
transform 1 0 19776 0 1 3780
box -48 -56 240 834
use sg13g2_decap_4  FILLER_4_234
timestamp 1679577901
transform 1 0 23616 0 1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_238
timestamp 1677579658
transform 1 0 24000 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_277
timestamp 1677580104
transform 1 0 27744 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_317
timestamp 1677580104
transform 1 0 31584 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_348
timestamp 1677580104
transform 1 0 34560 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_379
timestamp 1677580104
transform 1 0 37536 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_402
timestamp 1677579658
transform 1 0 39744 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_411
timestamp 1677580104
transform 1 0 40608 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_421
timestamp 1677580104
transform 1 0 41568 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_423
timestamp 1677579658
transform 1 0 41760 0 1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_0
timestamp 1677579658
transform 1 0 1152 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_18
timestamp 1677579658
transform 1 0 2880 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_34
timestamp 1677579658
transform 1 0 4416 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_95
timestamp 1677579658
transform 1 0 10272 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_135
timestamp 1679581782
transform 1 0 14112 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_180
timestamp 1679581782
transform 1 0 18432 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_187
timestamp 1679581782
transform 1 0 19104 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_4  FILLER_5_194
timestamp 1679577901
transform 1 0 19776 0 -1 5292
box -48 -56 432 834
use sg13g2_decap_4  FILLER_5_202
timestamp 1679577901
transform 1 0 20544 0 -1 5292
box -48 -56 432 834
use sg13g2_decap_8  FILLER_5_210
timestamp 1679581782
transform 1 0 21312 0 -1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_5_234
timestamp 1679581782
transform 1 0 23616 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_241
timestamp 1677580104
transform 1 0 24288 0 -1 5292
box -48 -56 240 834
use sg13g2_decap_4  FILLER_5_260
timestamp 1679577901
transform 1 0 26112 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_5_289
timestamp 1677580104
transform 1 0 28896 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_291
timestamp 1677579658
transform 1 0 29088 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_330
timestamp 1677580104
transform 1 0 32832 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_332
timestamp 1677579658
transform 1 0 33024 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_358
timestamp 1677579658
transform 1 0 35520 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_406
timestamp 1677580104
transform 1 0 40128 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_408
timestamp 1677579658
transform 1 0 40320 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_421
timestamp 1677580104
transform 1 0 41568 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_423
timestamp 1677579658
transform 1 0 41760 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_71
timestamp 1677579658
transform 1 0 7968 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_100
timestamp 1677579658
transform 1 0 10752 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_139
timestamp 1679581782
transform 1 0 14496 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_146
timestamp 1679581782
transform 1 0 15168 0 1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_6_153
timestamp 1677580104
transform 1 0 15840 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_155
timestamp 1677579658
transform 1 0 16032 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_194
timestamp 1679581782
transform 1 0 19776 0 1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_222
timestamp 1677579658
transform 1 0 22464 0 1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_6_231
timestamp 1679577901
transform 1 0 23328 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_235
timestamp 1677579658
transform 1 0 23712 0 1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_6_265
timestamp 1679577901
transform 1 0 26592 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_269
timestamp 1677579658
transform 1 0 26976 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_274
timestamp 1677579658
transform 1 0 27456 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_321
timestamp 1677580104
transform 1 0 31968 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_348
timestamp 1677579658
transform 1 0 34560 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_370
timestamp 1677580104
transform 1 0 36672 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_372
timestamp 1677579658
transform 1 0 36864 0 1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_6_398
timestamp 1679577901
transform 1 0 39360 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_402
timestamp 1677579658
transform 1 0 39744 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_407
timestamp 1677580104
transform 1 0 40224 0 1 5292
box -48 -56 240 834
use sg13g2_fill_2  FILLER_6_421
timestamp 1677580104
transform 1 0 41568 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_423
timestamp 1677579658
transform 1 0 41760 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_22
timestamp 1677580104
transform 1 0 3264 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_54
timestamp 1677579658
transform 1 0 6336 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_86
timestamp 1677579658
transform 1 0 9408 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_104
timestamp 1677580104
transform 1 0 11136 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_149
timestamp 1677580104
transform 1 0 15456 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_172
timestamp 1677580104
transform 1 0 17664 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_174
timestamp 1677579658
transform 1 0 17856 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_200
timestamp 1679581782
transform 1 0 20352 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_245
timestamp 1677580104
transform 1 0 24672 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_4  FILLER_7_264
timestamp 1679577901
transform 1 0 26496 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_7_306
timestamp 1677579658
transform 1 0 30528 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_374
timestamp 1677580104
transform 1 0 37056 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_393
timestamp 1677580104
transform 1 0 38880 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_412
timestamp 1677579658
transform 1 0 40704 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_421
timestamp 1677580104
transform 1 0 41568 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_423
timestamp 1677579658
transform 1 0 41760 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_59
timestamp 1677579658
transform 1 0 6816 0 1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_107
timestamp 1679577901
transform 1 0 11424 0 1 6804
box -48 -56 432 834
use sg13g2_decap_4  FILLER_8_206
timestamp 1679577901
transform 1 0 20928 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_256
timestamp 1677579658
transform 1 0 25728 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_328
timestamp 1677580104
transform 1 0 32640 0 1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_385
timestamp 1677580104
transform 1 0 38112 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_387
timestamp 1677579658
transform 1 0 38304 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_421
timestamp 1677580104
transform 1 0 41568 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_423
timestamp 1677579658
transform 1 0 41760 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_0
timestamp 1677580104
transform 1 0 1152 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_36
timestamp 1677580104
transform 1 0 4608 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_65
timestamp 1677580104
transform 1 0 7392 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_112
timestamp 1677580104
transform 1 0 11904 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_158
timestamp 1677579658
transform 1 0 16320 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_197
timestamp 1677580104
transform 1 0 20064 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_199
timestamp 1677579658
transform 1 0 20256 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_225
timestamp 1679581782
transform 1 0 22752 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_287
timestamp 1677580104
transform 1 0 28704 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_340
timestamp 1677579658
transform 1 0 33792 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_389
timestamp 1677579658
transform 1 0 38496 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_423
timestamp 1677579658
transform 1 0 41760 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_0
timestamp 1677579658
transform 1 0 1152 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_39
timestamp 1677580104
transform 1 0 4896 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_48
timestamp 1677580104
transform 1 0 5760 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_50
timestamp 1677579658
transform 1 0 5952 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_85
timestamp 1677579658
transform 1 0 9312 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_153
timestamp 1677580104
transform 1 0 15840 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_155
timestamp 1677579658
transform 1 0 16032 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_194
timestamp 1677580104
transform 1 0 19776 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_200
timestamp 1677579658
transform 1 0 20352 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_247
timestamp 1677579658
transform 1 0 24864 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_273
timestamp 1677580104
transform 1 0 27360 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_315
timestamp 1677579658
transform 1 0 31392 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_343
timestamp 1677580104
transform 1 0 34080 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_393
timestamp 1677580104
transform 1 0 38880 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_412
timestamp 1677579658
transform 1 0 40704 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_421
timestamp 1677580104
transform 1 0 41568 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_423
timestamp 1677579658
transform 1 0 41760 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_0
timestamp 1677580104
transform 1 0 1152 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_29
timestamp 1677580104
transform 1 0 3936 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_87
timestamp 1677580104
transform 1 0 9504 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_89
timestamp 1677579658
transform 1 0 9696 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_175
timestamp 1677579658
transform 1 0 17952 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_227
timestamp 1677580104
transform 1 0 22944 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_327
timestamp 1677580104
transform 1 0 32544 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_329
timestamp 1677579658
transform 1 0 32736 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_421
timestamp 1677580104
transform 1 0 41568 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_423
timestamp 1677579658
transform 1 0 41760 0 -1 9828
box -48 -56 144 834
<< labels >>
flabel metal2 s 4088 10672 4168 10752 0 FreeSans 320 0 0 0 A_I_top
port 0 nsew signal output
flabel metal2 s 2936 10672 3016 10752 0 FreeSans 320 0 0 0 A_O_top
port 1 nsew signal input
flabel metal2 s 5240 10672 5320 10752 0 FreeSans 320 0 0 0 A_T_top
port 2 nsew signal output
flabel metal2 s 7544 10672 7624 10752 0 FreeSans 320 0 0 0 B_I_top
port 3 nsew signal output
flabel metal2 s 6392 10672 6472 10752 0 FreeSans 320 0 0 0 B_O_top
port 4 nsew signal input
flabel metal2 s 8696 10672 8776 10752 0 FreeSans 320 0 0 0 B_T_top
port 5 nsew signal output
flabel metal2 s 11000 10672 11080 10752 0 FreeSans 320 0 0 0 C_I_top
port 6 nsew signal output
flabel metal2 s 9848 10672 9928 10752 0 FreeSans 320 0 0 0 C_O_top
port 7 nsew signal input
flabel metal2 s 12152 10672 12232 10752 0 FreeSans 320 0 0 0 C_T_top
port 8 nsew signal output
flabel metal2 s 19448 0 19528 80 0 FreeSans 320 0 0 0 Ci
port 9 nsew signal input
flabel metal2 s 14456 10672 14536 10752 0 FreeSans 320 0 0 0 D_I_top
port 10 nsew signal output
flabel metal2 s 13304 10672 13384 10752 0 FreeSans 320 0 0 0 D_O_top
port 11 nsew signal input
flabel metal2 s 15608 10672 15688 10752 0 FreeSans 320 0 0 0 D_T_top
port 12 nsew signal output
flabel metal3 s 0 44 80 124 0 FreeSans 320 0 0 0 FrameData[0]
port 13 nsew signal input
flabel metal3 s 0 3404 80 3484 0 FreeSans 320 0 0 0 FrameData[10]
port 14 nsew signal input
flabel metal3 s 0 3740 80 3820 0 FreeSans 320 0 0 0 FrameData[11]
port 15 nsew signal input
flabel metal3 s 0 4076 80 4156 0 FreeSans 320 0 0 0 FrameData[12]
port 16 nsew signal input
flabel metal3 s 0 4412 80 4492 0 FreeSans 320 0 0 0 FrameData[13]
port 17 nsew signal input
flabel metal3 s 0 4748 80 4828 0 FreeSans 320 0 0 0 FrameData[14]
port 18 nsew signal input
flabel metal3 s 0 5084 80 5164 0 FreeSans 320 0 0 0 FrameData[15]
port 19 nsew signal input
flabel metal3 s 0 5420 80 5500 0 FreeSans 320 0 0 0 FrameData[16]
port 20 nsew signal input
flabel metal3 s 0 5756 80 5836 0 FreeSans 320 0 0 0 FrameData[17]
port 21 nsew signal input
flabel metal3 s 0 6092 80 6172 0 FreeSans 320 0 0 0 FrameData[18]
port 22 nsew signal input
flabel metal3 s 0 6428 80 6508 0 FreeSans 320 0 0 0 FrameData[19]
port 23 nsew signal input
flabel metal3 s 0 380 80 460 0 FreeSans 320 0 0 0 FrameData[1]
port 24 nsew signal input
flabel metal3 s 0 6764 80 6844 0 FreeSans 320 0 0 0 FrameData[20]
port 25 nsew signal input
flabel metal3 s 0 7100 80 7180 0 FreeSans 320 0 0 0 FrameData[21]
port 26 nsew signal input
flabel metal3 s 0 7436 80 7516 0 FreeSans 320 0 0 0 FrameData[22]
port 27 nsew signal input
flabel metal3 s 0 7772 80 7852 0 FreeSans 320 0 0 0 FrameData[23]
port 28 nsew signal input
flabel metal3 s 0 8108 80 8188 0 FreeSans 320 0 0 0 FrameData[24]
port 29 nsew signal input
flabel metal3 s 0 8444 80 8524 0 FreeSans 320 0 0 0 FrameData[25]
port 30 nsew signal input
flabel metal3 s 0 8780 80 8860 0 FreeSans 320 0 0 0 FrameData[26]
port 31 nsew signal input
flabel metal3 s 0 9116 80 9196 0 FreeSans 320 0 0 0 FrameData[27]
port 32 nsew signal input
flabel metal3 s 0 9452 80 9532 0 FreeSans 320 0 0 0 FrameData[28]
port 33 nsew signal input
flabel metal3 s 0 9788 80 9868 0 FreeSans 320 0 0 0 FrameData[29]
port 34 nsew signal input
flabel metal3 s 0 716 80 796 0 FreeSans 320 0 0 0 FrameData[2]
port 35 nsew signal input
flabel metal3 s 0 10124 80 10204 0 FreeSans 320 0 0 0 FrameData[30]
port 36 nsew signal input
flabel metal3 s 0 10460 80 10540 0 FreeSans 320 0 0 0 FrameData[31]
port 37 nsew signal input
flabel metal3 s 0 1052 80 1132 0 FreeSans 320 0 0 0 FrameData[3]
port 38 nsew signal input
flabel metal3 s 0 1388 80 1468 0 FreeSans 320 0 0 0 FrameData[4]
port 39 nsew signal input
flabel metal3 s 0 1724 80 1804 0 FreeSans 320 0 0 0 FrameData[5]
port 40 nsew signal input
flabel metal3 s 0 2060 80 2140 0 FreeSans 320 0 0 0 FrameData[6]
port 41 nsew signal input
flabel metal3 s 0 2396 80 2476 0 FreeSans 320 0 0 0 FrameData[7]
port 42 nsew signal input
flabel metal3 s 0 2732 80 2812 0 FreeSans 320 0 0 0 FrameData[8]
port 43 nsew signal input
flabel metal3 s 0 3068 80 3148 0 FreeSans 320 0 0 0 FrameData[9]
port 44 nsew signal input
flabel metal3 s 42928 44 43008 124 0 FreeSans 320 0 0 0 FrameData_O[0]
port 45 nsew signal output
flabel metal3 s 42928 3404 43008 3484 0 FreeSans 320 0 0 0 FrameData_O[10]
port 46 nsew signal output
flabel metal3 s 42928 3740 43008 3820 0 FreeSans 320 0 0 0 FrameData_O[11]
port 47 nsew signal output
flabel metal3 s 42928 4076 43008 4156 0 FreeSans 320 0 0 0 FrameData_O[12]
port 48 nsew signal output
flabel metal3 s 42928 4412 43008 4492 0 FreeSans 320 0 0 0 FrameData_O[13]
port 49 nsew signal output
flabel metal3 s 42928 4748 43008 4828 0 FreeSans 320 0 0 0 FrameData_O[14]
port 50 nsew signal output
flabel metal3 s 42928 5084 43008 5164 0 FreeSans 320 0 0 0 FrameData_O[15]
port 51 nsew signal output
flabel metal3 s 42928 5420 43008 5500 0 FreeSans 320 0 0 0 FrameData_O[16]
port 52 nsew signal output
flabel metal3 s 42928 5756 43008 5836 0 FreeSans 320 0 0 0 FrameData_O[17]
port 53 nsew signal output
flabel metal3 s 42928 6092 43008 6172 0 FreeSans 320 0 0 0 FrameData_O[18]
port 54 nsew signal output
flabel metal3 s 42928 6428 43008 6508 0 FreeSans 320 0 0 0 FrameData_O[19]
port 55 nsew signal output
flabel metal3 s 42928 380 43008 460 0 FreeSans 320 0 0 0 FrameData_O[1]
port 56 nsew signal output
flabel metal3 s 42928 6764 43008 6844 0 FreeSans 320 0 0 0 FrameData_O[20]
port 57 nsew signal output
flabel metal3 s 42928 7100 43008 7180 0 FreeSans 320 0 0 0 FrameData_O[21]
port 58 nsew signal output
flabel metal3 s 42928 7436 43008 7516 0 FreeSans 320 0 0 0 FrameData_O[22]
port 59 nsew signal output
flabel metal3 s 42928 7772 43008 7852 0 FreeSans 320 0 0 0 FrameData_O[23]
port 60 nsew signal output
flabel metal3 s 42928 8108 43008 8188 0 FreeSans 320 0 0 0 FrameData_O[24]
port 61 nsew signal output
flabel metal3 s 42928 8444 43008 8524 0 FreeSans 320 0 0 0 FrameData_O[25]
port 62 nsew signal output
flabel metal3 s 42928 8780 43008 8860 0 FreeSans 320 0 0 0 FrameData_O[26]
port 63 nsew signal output
flabel metal3 s 42928 9116 43008 9196 0 FreeSans 320 0 0 0 FrameData_O[27]
port 64 nsew signal output
flabel metal3 s 42928 9452 43008 9532 0 FreeSans 320 0 0 0 FrameData_O[28]
port 65 nsew signal output
flabel metal3 s 42928 9788 43008 9868 0 FreeSans 320 0 0 0 FrameData_O[29]
port 66 nsew signal output
flabel metal3 s 42928 716 43008 796 0 FreeSans 320 0 0 0 FrameData_O[2]
port 67 nsew signal output
flabel metal3 s 42928 10124 43008 10204 0 FreeSans 320 0 0 0 FrameData_O[30]
port 68 nsew signal output
flabel metal3 s 42928 10460 43008 10540 0 FreeSans 320 0 0 0 FrameData_O[31]
port 69 nsew signal output
flabel metal3 s 42928 1052 43008 1132 0 FreeSans 320 0 0 0 FrameData_O[3]
port 70 nsew signal output
flabel metal3 s 42928 1388 43008 1468 0 FreeSans 320 0 0 0 FrameData_O[4]
port 71 nsew signal output
flabel metal3 s 42928 1724 43008 1804 0 FreeSans 320 0 0 0 FrameData_O[5]
port 72 nsew signal output
flabel metal3 s 42928 2060 43008 2140 0 FreeSans 320 0 0 0 FrameData_O[6]
port 73 nsew signal output
flabel metal3 s 42928 2396 43008 2476 0 FreeSans 320 0 0 0 FrameData_O[7]
port 74 nsew signal output
flabel metal3 s 42928 2732 43008 2812 0 FreeSans 320 0 0 0 FrameData_O[8]
port 75 nsew signal output
flabel metal3 s 42928 3068 43008 3148 0 FreeSans 320 0 0 0 FrameData_O[9]
port 76 nsew signal output
flabel metal2 s 29816 0 29896 80 0 FreeSans 320 0 0 0 FrameStrobe[0]
port 77 nsew signal input
flabel metal2 s 31736 0 31816 80 0 FreeSans 320 0 0 0 FrameStrobe[10]
port 78 nsew signal input
flabel metal2 s 31928 0 32008 80 0 FreeSans 320 0 0 0 FrameStrobe[11]
port 79 nsew signal input
flabel metal2 s 32120 0 32200 80 0 FreeSans 320 0 0 0 FrameStrobe[12]
port 80 nsew signal input
flabel metal2 s 32312 0 32392 80 0 FreeSans 320 0 0 0 FrameStrobe[13]
port 81 nsew signal input
flabel metal2 s 32504 0 32584 80 0 FreeSans 320 0 0 0 FrameStrobe[14]
port 82 nsew signal input
flabel metal2 s 32696 0 32776 80 0 FreeSans 320 0 0 0 FrameStrobe[15]
port 83 nsew signal input
flabel metal2 s 32888 0 32968 80 0 FreeSans 320 0 0 0 FrameStrobe[16]
port 84 nsew signal input
flabel metal2 s 33080 0 33160 80 0 FreeSans 320 0 0 0 FrameStrobe[17]
port 85 nsew signal input
flabel metal2 s 33272 0 33352 80 0 FreeSans 320 0 0 0 FrameStrobe[18]
port 86 nsew signal input
flabel metal2 s 33464 0 33544 80 0 FreeSans 320 0 0 0 FrameStrobe[19]
port 87 nsew signal input
flabel metal2 s 30008 0 30088 80 0 FreeSans 320 0 0 0 FrameStrobe[1]
port 88 nsew signal input
flabel metal2 s 30200 0 30280 80 0 FreeSans 320 0 0 0 FrameStrobe[2]
port 89 nsew signal input
flabel metal2 s 30392 0 30472 80 0 FreeSans 320 0 0 0 FrameStrobe[3]
port 90 nsew signal input
flabel metal2 s 30584 0 30664 80 0 FreeSans 320 0 0 0 FrameStrobe[4]
port 91 nsew signal input
flabel metal2 s 30776 0 30856 80 0 FreeSans 320 0 0 0 FrameStrobe[5]
port 92 nsew signal input
flabel metal2 s 30968 0 31048 80 0 FreeSans 320 0 0 0 FrameStrobe[6]
port 93 nsew signal input
flabel metal2 s 31160 0 31240 80 0 FreeSans 320 0 0 0 FrameStrobe[7]
port 94 nsew signal input
flabel metal2 s 31352 0 31432 80 0 FreeSans 320 0 0 0 FrameStrobe[8]
port 95 nsew signal input
flabel metal2 s 31544 0 31624 80 0 FreeSans 320 0 0 0 FrameStrobe[9]
port 96 nsew signal input
flabel metal2 s 17912 10672 17992 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[0]
port 97 nsew signal output
flabel metal2 s 29432 10672 29512 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[10]
port 98 nsew signal output
flabel metal2 s 30584 10672 30664 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[11]
port 99 nsew signal output
flabel metal2 s 31736 10672 31816 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[12]
port 100 nsew signal output
flabel metal2 s 32888 10672 32968 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[13]
port 101 nsew signal output
flabel metal2 s 34040 10672 34120 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[14]
port 102 nsew signal output
flabel metal2 s 35192 10672 35272 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[15]
port 103 nsew signal output
flabel metal2 s 36344 10672 36424 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[16]
port 104 nsew signal output
flabel metal2 s 37496 10672 37576 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[17]
port 105 nsew signal output
flabel metal2 s 38648 10672 38728 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[18]
port 106 nsew signal output
flabel metal2 s 39800 10672 39880 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[19]
port 107 nsew signal output
flabel metal2 s 19064 10672 19144 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[1]
port 108 nsew signal output
flabel metal2 s 20216 10672 20296 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[2]
port 109 nsew signal output
flabel metal2 s 21368 10672 21448 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[3]
port 110 nsew signal output
flabel metal2 s 22520 10672 22600 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[4]
port 111 nsew signal output
flabel metal2 s 23672 10672 23752 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[5]
port 112 nsew signal output
flabel metal2 s 24824 10672 24904 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[6]
port 113 nsew signal output
flabel metal2 s 25976 10672 26056 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[7]
port 114 nsew signal output
flabel metal2 s 27128 10672 27208 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[8]
port 115 nsew signal output
flabel metal2 s 28280 10672 28360 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[9]
port 116 nsew signal output
flabel metal2 s 9464 0 9544 80 0 FreeSans 320 0 0 0 N1END[0]
port 117 nsew signal input
flabel metal2 s 9656 0 9736 80 0 FreeSans 320 0 0 0 N1END[1]
port 118 nsew signal input
flabel metal2 s 9848 0 9928 80 0 FreeSans 320 0 0 0 N1END[2]
port 119 nsew signal input
flabel metal2 s 10040 0 10120 80 0 FreeSans 320 0 0 0 N1END[3]
port 120 nsew signal input
flabel metal2 s 11768 0 11848 80 0 FreeSans 320 0 0 0 N2END[0]
port 121 nsew signal input
flabel metal2 s 11960 0 12040 80 0 FreeSans 320 0 0 0 N2END[1]
port 122 nsew signal input
flabel metal2 s 12152 0 12232 80 0 FreeSans 320 0 0 0 N2END[2]
port 123 nsew signal input
flabel metal2 s 12344 0 12424 80 0 FreeSans 320 0 0 0 N2END[3]
port 124 nsew signal input
flabel metal2 s 12536 0 12616 80 0 FreeSans 320 0 0 0 N2END[4]
port 125 nsew signal input
flabel metal2 s 12728 0 12808 80 0 FreeSans 320 0 0 0 N2END[5]
port 126 nsew signal input
flabel metal2 s 12920 0 13000 80 0 FreeSans 320 0 0 0 N2END[6]
port 127 nsew signal input
flabel metal2 s 13112 0 13192 80 0 FreeSans 320 0 0 0 N2END[7]
port 128 nsew signal input
flabel metal2 s 10232 0 10312 80 0 FreeSans 320 0 0 0 N2MID[0]
port 129 nsew signal input
flabel metal2 s 10424 0 10504 80 0 FreeSans 320 0 0 0 N2MID[1]
port 130 nsew signal input
flabel metal2 s 10616 0 10696 80 0 FreeSans 320 0 0 0 N2MID[2]
port 131 nsew signal input
flabel metal2 s 10808 0 10888 80 0 FreeSans 320 0 0 0 N2MID[3]
port 132 nsew signal input
flabel metal2 s 11000 0 11080 80 0 FreeSans 320 0 0 0 N2MID[4]
port 133 nsew signal input
flabel metal2 s 11192 0 11272 80 0 FreeSans 320 0 0 0 N2MID[5]
port 134 nsew signal input
flabel metal2 s 11384 0 11464 80 0 FreeSans 320 0 0 0 N2MID[6]
port 135 nsew signal input
flabel metal2 s 11576 0 11656 80 0 FreeSans 320 0 0 0 N2MID[7]
port 136 nsew signal input
flabel metal2 s 13304 0 13384 80 0 FreeSans 320 0 0 0 N4END[0]
port 137 nsew signal input
flabel metal2 s 15224 0 15304 80 0 FreeSans 320 0 0 0 N4END[10]
port 138 nsew signal input
flabel metal2 s 15416 0 15496 80 0 FreeSans 320 0 0 0 N4END[11]
port 139 nsew signal input
flabel metal2 s 15608 0 15688 80 0 FreeSans 320 0 0 0 N4END[12]
port 140 nsew signal input
flabel metal2 s 15800 0 15880 80 0 FreeSans 320 0 0 0 N4END[13]
port 141 nsew signal input
flabel metal2 s 15992 0 16072 80 0 FreeSans 320 0 0 0 N4END[14]
port 142 nsew signal input
flabel metal2 s 16184 0 16264 80 0 FreeSans 320 0 0 0 N4END[15]
port 143 nsew signal input
flabel metal2 s 13496 0 13576 80 0 FreeSans 320 0 0 0 N4END[1]
port 144 nsew signal input
flabel metal2 s 13688 0 13768 80 0 FreeSans 320 0 0 0 N4END[2]
port 145 nsew signal input
flabel metal2 s 13880 0 13960 80 0 FreeSans 320 0 0 0 N4END[3]
port 146 nsew signal input
flabel metal2 s 14072 0 14152 80 0 FreeSans 320 0 0 0 N4END[4]
port 147 nsew signal input
flabel metal2 s 14264 0 14344 80 0 FreeSans 320 0 0 0 N4END[5]
port 148 nsew signal input
flabel metal2 s 14456 0 14536 80 0 FreeSans 320 0 0 0 N4END[6]
port 149 nsew signal input
flabel metal2 s 14648 0 14728 80 0 FreeSans 320 0 0 0 N4END[7]
port 150 nsew signal input
flabel metal2 s 14840 0 14920 80 0 FreeSans 320 0 0 0 N4END[8]
port 151 nsew signal input
flabel metal2 s 15032 0 15112 80 0 FreeSans 320 0 0 0 N4END[9]
port 152 nsew signal input
flabel metal2 s 16376 0 16456 80 0 FreeSans 320 0 0 0 NN4END[0]
port 153 nsew signal input
flabel metal2 s 18296 0 18376 80 0 FreeSans 320 0 0 0 NN4END[10]
port 154 nsew signal input
flabel metal2 s 18488 0 18568 80 0 FreeSans 320 0 0 0 NN4END[11]
port 155 nsew signal input
flabel metal2 s 18680 0 18760 80 0 FreeSans 320 0 0 0 NN4END[12]
port 156 nsew signal input
flabel metal2 s 18872 0 18952 80 0 FreeSans 320 0 0 0 NN4END[13]
port 157 nsew signal input
flabel metal2 s 19064 0 19144 80 0 FreeSans 320 0 0 0 NN4END[14]
port 158 nsew signal input
flabel metal2 s 19256 0 19336 80 0 FreeSans 320 0 0 0 NN4END[15]
port 159 nsew signal input
flabel metal2 s 16568 0 16648 80 0 FreeSans 320 0 0 0 NN4END[1]
port 160 nsew signal input
flabel metal2 s 16760 0 16840 80 0 FreeSans 320 0 0 0 NN4END[2]
port 161 nsew signal input
flabel metal2 s 16952 0 17032 80 0 FreeSans 320 0 0 0 NN4END[3]
port 162 nsew signal input
flabel metal2 s 17144 0 17224 80 0 FreeSans 320 0 0 0 NN4END[4]
port 163 nsew signal input
flabel metal2 s 17336 0 17416 80 0 FreeSans 320 0 0 0 NN4END[5]
port 164 nsew signal input
flabel metal2 s 17528 0 17608 80 0 FreeSans 320 0 0 0 NN4END[6]
port 165 nsew signal input
flabel metal2 s 17720 0 17800 80 0 FreeSans 320 0 0 0 NN4END[7]
port 166 nsew signal input
flabel metal2 s 17912 0 17992 80 0 FreeSans 320 0 0 0 NN4END[8]
port 167 nsew signal input
flabel metal2 s 18104 0 18184 80 0 FreeSans 320 0 0 0 NN4END[9]
port 168 nsew signal input
flabel metal2 s 19640 0 19720 80 0 FreeSans 320 0 0 0 S1BEG[0]
port 169 nsew signal output
flabel metal2 s 19832 0 19912 80 0 FreeSans 320 0 0 0 S1BEG[1]
port 170 nsew signal output
flabel metal2 s 20024 0 20104 80 0 FreeSans 320 0 0 0 S1BEG[2]
port 171 nsew signal output
flabel metal2 s 20216 0 20296 80 0 FreeSans 320 0 0 0 S1BEG[3]
port 172 nsew signal output
flabel metal2 s 20408 0 20488 80 0 FreeSans 320 0 0 0 S2BEG[0]
port 173 nsew signal output
flabel metal2 s 20600 0 20680 80 0 FreeSans 320 0 0 0 S2BEG[1]
port 174 nsew signal output
flabel metal2 s 20792 0 20872 80 0 FreeSans 320 0 0 0 S2BEG[2]
port 175 nsew signal output
flabel metal2 s 20984 0 21064 80 0 FreeSans 320 0 0 0 S2BEG[3]
port 176 nsew signal output
flabel metal2 s 21176 0 21256 80 0 FreeSans 320 0 0 0 S2BEG[4]
port 177 nsew signal output
flabel metal2 s 21368 0 21448 80 0 FreeSans 320 0 0 0 S2BEG[5]
port 178 nsew signal output
flabel metal2 s 21560 0 21640 80 0 FreeSans 320 0 0 0 S2BEG[6]
port 179 nsew signal output
flabel metal2 s 21752 0 21832 80 0 FreeSans 320 0 0 0 S2BEG[7]
port 180 nsew signal output
flabel metal2 s 21944 0 22024 80 0 FreeSans 320 0 0 0 S2BEGb[0]
port 181 nsew signal output
flabel metal2 s 22136 0 22216 80 0 FreeSans 320 0 0 0 S2BEGb[1]
port 182 nsew signal output
flabel metal2 s 22328 0 22408 80 0 FreeSans 320 0 0 0 S2BEGb[2]
port 183 nsew signal output
flabel metal2 s 22520 0 22600 80 0 FreeSans 320 0 0 0 S2BEGb[3]
port 184 nsew signal output
flabel metal2 s 22712 0 22792 80 0 FreeSans 320 0 0 0 S2BEGb[4]
port 185 nsew signal output
flabel metal2 s 22904 0 22984 80 0 FreeSans 320 0 0 0 S2BEGb[5]
port 186 nsew signal output
flabel metal2 s 23096 0 23176 80 0 FreeSans 320 0 0 0 S2BEGb[6]
port 187 nsew signal output
flabel metal2 s 23288 0 23368 80 0 FreeSans 320 0 0 0 S2BEGb[7]
port 188 nsew signal output
flabel metal2 s 23480 0 23560 80 0 FreeSans 320 0 0 0 S4BEG[0]
port 189 nsew signal output
flabel metal2 s 25400 0 25480 80 0 FreeSans 320 0 0 0 S4BEG[10]
port 190 nsew signal output
flabel metal2 s 25592 0 25672 80 0 FreeSans 320 0 0 0 S4BEG[11]
port 191 nsew signal output
flabel metal2 s 25784 0 25864 80 0 FreeSans 320 0 0 0 S4BEG[12]
port 192 nsew signal output
flabel metal2 s 25976 0 26056 80 0 FreeSans 320 0 0 0 S4BEG[13]
port 193 nsew signal output
flabel metal2 s 26168 0 26248 80 0 FreeSans 320 0 0 0 S4BEG[14]
port 194 nsew signal output
flabel metal2 s 26360 0 26440 80 0 FreeSans 320 0 0 0 S4BEG[15]
port 195 nsew signal output
flabel metal2 s 23672 0 23752 80 0 FreeSans 320 0 0 0 S4BEG[1]
port 196 nsew signal output
flabel metal2 s 23864 0 23944 80 0 FreeSans 320 0 0 0 S4BEG[2]
port 197 nsew signal output
flabel metal2 s 24056 0 24136 80 0 FreeSans 320 0 0 0 S4BEG[3]
port 198 nsew signal output
flabel metal2 s 24248 0 24328 80 0 FreeSans 320 0 0 0 S4BEG[4]
port 199 nsew signal output
flabel metal2 s 24440 0 24520 80 0 FreeSans 320 0 0 0 S4BEG[5]
port 200 nsew signal output
flabel metal2 s 24632 0 24712 80 0 FreeSans 320 0 0 0 S4BEG[6]
port 201 nsew signal output
flabel metal2 s 24824 0 24904 80 0 FreeSans 320 0 0 0 S4BEG[7]
port 202 nsew signal output
flabel metal2 s 25016 0 25096 80 0 FreeSans 320 0 0 0 S4BEG[8]
port 203 nsew signal output
flabel metal2 s 25208 0 25288 80 0 FreeSans 320 0 0 0 S4BEG[9]
port 204 nsew signal output
flabel metal2 s 26552 0 26632 80 0 FreeSans 320 0 0 0 SS4BEG[0]
port 205 nsew signal output
flabel metal2 s 28472 0 28552 80 0 FreeSans 320 0 0 0 SS4BEG[10]
port 206 nsew signal output
flabel metal2 s 28664 0 28744 80 0 FreeSans 320 0 0 0 SS4BEG[11]
port 207 nsew signal output
flabel metal2 s 28856 0 28936 80 0 FreeSans 320 0 0 0 SS4BEG[12]
port 208 nsew signal output
flabel metal2 s 29048 0 29128 80 0 FreeSans 320 0 0 0 SS4BEG[13]
port 209 nsew signal output
flabel metal2 s 29240 0 29320 80 0 FreeSans 320 0 0 0 SS4BEG[14]
port 210 nsew signal output
flabel metal2 s 29432 0 29512 80 0 FreeSans 320 0 0 0 SS4BEG[15]
port 211 nsew signal output
flabel metal2 s 26744 0 26824 80 0 FreeSans 320 0 0 0 SS4BEG[1]
port 212 nsew signal output
flabel metal2 s 26936 0 27016 80 0 FreeSans 320 0 0 0 SS4BEG[2]
port 213 nsew signal output
flabel metal2 s 27128 0 27208 80 0 FreeSans 320 0 0 0 SS4BEG[3]
port 214 nsew signal output
flabel metal2 s 27320 0 27400 80 0 FreeSans 320 0 0 0 SS4BEG[4]
port 215 nsew signal output
flabel metal2 s 27512 0 27592 80 0 FreeSans 320 0 0 0 SS4BEG[5]
port 216 nsew signal output
flabel metal2 s 27704 0 27784 80 0 FreeSans 320 0 0 0 SS4BEG[6]
port 217 nsew signal output
flabel metal2 s 27896 0 27976 80 0 FreeSans 320 0 0 0 SS4BEG[7]
port 218 nsew signal output
flabel metal2 s 28088 0 28168 80 0 FreeSans 320 0 0 0 SS4BEG[8]
port 219 nsew signal output
flabel metal2 s 28280 0 28360 80 0 FreeSans 320 0 0 0 SS4BEG[9]
port 220 nsew signal output
flabel metal2 s 29624 0 29704 80 0 FreeSans 320 0 0 0 UserCLK
port 221 nsew signal input
flabel metal2 s 16760 10672 16840 10752 0 FreeSans 320 0 0 0 UserCLKo
port 222 nsew signal output
flabel metal6 s 4892 0 5332 10752 0 FreeSans 2624 90 0 0 VGND
port 223 nsew ground bidirectional
flabel metal6 s 4892 0 5332 328 0 FreeSans 2624 0 0 0 VGND
port 223 nsew ground bidirectional
flabel metal6 s 4892 10424 5332 10752 0 FreeSans 2624 0 0 0 VGND
port 223 nsew ground bidirectional
flabel metal6 s 20012 0 20452 10752 0 FreeSans 2624 90 0 0 VGND
port 223 nsew ground bidirectional
flabel metal6 s 20012 0 20452 328 0 FreeSans 2624 0 0 0 VGND
port 223 nsew ground bidirectional
flabel metal6 s 20012 10424 20452 10752 0 FreeSans 2624 0 0 0 VGND
port 223 nsew ground bidirectional
flabel metal6 s 35132 0 35572 10752 0 FreeSans 2624 90 0 0 VGND
port 223 nsew ground bidirectional
flabel metal6 s 35132 0 35572 328 0 FreeSans 2624 0 0 0 VGND
port 223 nsew ground bidirectional
flabel metal6 s 35132 10424 35572 10752 0 FreeSans 2624 0 0 0 VGND
port 223 nsew ground bidirectional
flabel metal6 s 3652 0 4092 10752 0 FreeSans 2624 90 0 0 VPWR
port 224 nsew power bidirectional
flabel metal6 s 3652 0 4092 328 0 FreeSans 2624 0 0 0 VPWR
port 224 nsew power bidirectional
flabel metal6 s 3652 10424 4092 10752 0 FreeSans 2624 0 0 0 VPWR
port 224 nsew power bidirectional
flabel metal6 s 18772 0 19212 10752 0 FreeSans 2624 90 0 0 VPWR
port 224 nsew power bidirectional
flabel metal6 s 18772 0 19212 328 0 FreeSans 2624 0 0 0 VPWR
port 224 nsew power bidirectional
flabel metal6 s 18772 10424 19212 10752 0 FreeSans 2624 0 0 0 VPWR
port 224 nsew power bidirectional
flabel metal6 s 33892 0 34332 10752 0 FreeSans 2624 90 0 0 VPWR
port 224 nsew power bidirectional
flabel metal6 s 33892 0 34332 328 0 FreeSans 2624 0 0 0 VPWR
port 224 nsew power bidirectional
flabel metal6 s 33892 10424 34332 10752 0 FreeSans 2624 0 0 0 VPWR
port 224 nsew power bidirectional
rlabel metal1 21504 9828 21504 9828 0 VGND
rlabel metal1 21504 9072 21504 9072 0 VPWR
rlabel metal2 10080 2100 10080 2100 0 A_I_top
rlabel metal3 18480 2604 18480 2604 0 A_O_top
rlabel metal2 3552 3780 3552 3780 0 A_T_top
rlabel metal3 8976 5460 8976 5460 0 B_I_top
rlabel metal2 37920 2646 37920 2646 0 B_O_top
rlabel metal2 1440 9912 1440 9912 0 B_T_top
rlabel metal2 11040 10386 11040 10386 0 C_I_top
rlabel metal3 19776 2436 19776 2436 0 C_O_top
rlabel metal2 11712 7518 11712 7518 0 C_T_top
rlabel metal2 14496 10008 14496 10008 0 D_I_top
rlabel metal2 38592 5754 38592 5754 0 D_O_top
rlabel metal2 15744 9114 15744 9114 0 D_T_top
rlabel metal2 41280 1008 41280 1008 0 FrameData[0]
rlabel metal2 1440 3906 1440 3906 0 FrameData[10]
rlabel metal2 36576 2646 36576 2646 0 FrameData[11]
rlabel metal2 41280 4410 41280 4410 0 FrameData[12]
rlabel metal3 222 4452 222 4452 0 FrameData[13]
rlabel metal2 38400 4872 38400 4872 0 FrameData[14]
rlabel metal2 37824 4494 37824 4494 0 FrameData[15]
rlabel metal3 990 5460 990 5460 0 FrameData[16]
rlabel metal3 1230 5796 1230 5796 0 FrameData[17]
rlabel metal3 798 6132 798 6132 0 FrameData[18]
rlabel metal3 894 6468 894 6468 0 FrameData[19]
rlabel metal4 20736 1134 20736 1134 0 FrameData[1]
rlabel metal2 1776 5628 1776 5628 0 FrameData[20]
rlabel metal3 1278 7140 1278 7140 0 FrameData[21]
rlabel metal2 41184 8442 41184 8442 0 FrameData[22]
rlabel metal3 654 7812 654 7812 0 FrameData[23]
rlabel metal2 18144 9408 18144 9408 0 FrameData[24]
rlabel metal3 558 8484 558 8484 0 FrameData[25]
rlabel metal3 39552 5712 39552 5712 0 FrameData[26]
rlabel metal2 41232 4872 41232 4872 0 FrameData[27]
rlabel metal3 750 9492 750 9492 0 FrameData[28]
rlabel metal2 40896 9576 40896 9576 0 FrameData[29]
rlabel metal2 38592 2016 38592 2016 0 FrameData[2]
rlabel metal3 270 10164 270 10164 0 FrameData[30]
rlabel metal3 39648 5880 39648 5880 0 FrameData[31]
rlabel metal2 39408 3360 39408 3360 0 FrameData[3]
rlabel metal2 39936 4032 39936 4032 0 FrameData[4]
rlabel metal2 1824 840 1824 840 0 FrameData[5]
rlabel metal2 39648 3066 39648 3066 0 FrameData[6]
rlabel metal2 1824 2730 1824 2730 0 FrameData[7]
rlabel metal4 1344 4872 1344 4872 0 FrameData[8]
rlabel metal2 1632 3570 1632 3570 0 FrameData[9]
rlabel metal2 41472 504 41472 504 0 FrameData_O[0]
rlabel metal2 40704 3360 40704 3360 0 FrameData_O[10]
rlabel metal2 41088 3696 41088 3696 0 FrameData_O[11]
rlabel metal2 41472 4032 41472 4032 0 FrameData_O[12]
rlabel metal2 41088 4410 41088 4410 0 FrameData_O[13]
rlabel metal3 41826 4788 41826 4788 0 FrameData_O[14]
rlabel metal2 41088 4956 41088 4956 0 FrameData_O[15]
rlabel metal3 41826 5460 41826 5460 0 FrameData_O[16]
rlabel metal3 42018 5796 42018 5796 0 FrameData_O[17]
rlabel metal3 41526 6216 41526 6216 0 FrameData_O[18]
rlabel metal2 41088 6384 41088 6384 0 FrameData_O[19]
rlabel metal2 40416 1806 40416 1806 0 FrameData_O[1]
rlabel metal2 41088 6888 41088 6888 0 FrameData_O[20]
rlabel metal2 41472 7056 41472 7056 0 FrameData_O[21]
rlabel metal2 41280 7602 41280 7602 0 FrameData_O[22]
rlabel metal3 42306 7812 42306 7812 0 FrameData_O[23]
rlabel metal2 41088 8316 41088 8316 0 FrameData_O[24]
rlabel metal3 42210 8484 42210 8484 0 FrameData_O[25]
rlabel metal3 41136 5880 41136 5880 0 FrameData_O[26]
rlabel metal2 41424 4788 41424 4788 0 FrameData_O[27]
rlabel metal2 41472 9408 41472 9408 0 FrameData_O[28]
rlabel metal2 41088 9744 41088 9744 0 FrameData_O[29]
rlabel metal2 40800 1974 40800 1974 0 FrameData_O[2]
rlabel metal2 40704 9912 40704 9912 0 FrameData_O[30]
rlabel metal2 40944 8148 40944 8148 0 FrameData_O[31]
rlabel metal2 40608 1848 40608 1848 0 FrameData_O[3]
rlabel metal4 40896 2478 40896 2478 0 FrameData_O[4]
rlabel metal2 41088 1470 41088 1470 0 FrameData_O[5]
rlabel metal3 42306 2100 42306 2100 0 FrameData_O[6]
rlabel metal2 41280 2268 41280 2268 0 FrameData_O[7]
rlabel metal3 42306 2772 42306 2772 0 FrameData_O[8]
rlabel metal3 41526 3192 41526 3192 0 FrameData_O[9]
rlabel metal2 15744 6300 15744 6300 0 FrameStrobe[0]
rlabel metal2 31776 366 31776 366 0 FrameStrobe[10]
rlabel metal2 31968 114 31968 114 0 FrameStrobe[11]
rlabel metal2 38640 8736 38640 8736 0 FrameStrobe[12]
rlabel metal2 32352 408 32352 408 0 FrameStrobe[13]
rlabel metal2 39552 7686 39552 7686 0 FrameStrobe[14]
rlabel metal2 32736 492 32736 492 0 FrameStrobe[15]
rlabel metal2 38352 7896 38352 7896 0 FrameStrobe[16]
rlabel metal2 38016 6804 38016 6804 0 FrameStrobe[17]
rlabel metal2 39936 2016 39936 2016 0 FrameStrobe[18]
rlabel metal2 39840 4536 39840 4536 0 FrameStrobe[19]
rlabel metal3 39456 1092 39456 1092 0 FrameStrobe[1]
rlabel metal3 21888 1092 21888 1092 0 FrameStrobe[2]
rlabel metal3 13776 1092 13776 1092 0 FrameStrobe[3]
rlabel metal2 30624 1290 30624 1290 0 FrameStrobe[4]
rlabel metal2 30816 618 30816 618 0 FrameStrobe[5]
rlabel metal2 31056 3192 31056 3192 0 FrameStrobe[6]
rlabel metal2 31200 954 31200 954 0 FrameStrobe[7]
rlabel metal2 31392 660 31392 660 0 FrameStrobe[8]
rlabel metal2 31584 954 31584 954 0 FrameStrobe[9]
rlabel metal2 15936 6678 15936 6678 0 FrameStrobe_O[0]
rlabel metal3 33408 9660 33408 9660 0 FrameStrobe_O[10]
rlabel metal2 32304 3612 32304 3612 0 FrameStrobe_O[11]
rlabel metal2 38592 8148 38592 8148 0 FrameStrobe_O[12]
rlabel metal3 33840 5880 33840 5880 0 FrameStrobe_O[13]
rlabel metal2 39360 9786 39360 9786 0 FrameStrobe_O[14]
rlabel metal2 35232 4956 35232 4956 0 FrameStrobe_O[15]
rlabel metal2 38208 8778 38208 8778 0 FrameStrobe_O[16]
rlabel metal2 37824 7434 37824 7434 0 FrameStrobe_O[17]
rlabel metal3 39216 9660 39216 9660 0 FrameStrobe_O[18]
rlabel metal2 40128 9828 40128 9828 0 FrameStrobe_O[19]
rlabel metal2 20016 6636 20016 6636 0 FrameStrobe_O[1]
rlabel metal2 20256 8862 20256 8862 0 FrameStrobe_O[2]
rlabel metal2 21120 9240 21120 9240 0 FrameStrobe_O[3]
rlabel metal2 22464 8694 22464 8694 0 FrameStrobe_O[4]
rlabel metal2 32352 8904 32352 8904 0 FrameStrobe_O[5]
rlabel metal2 31680 6468 31680 6468 0 FrameStrobe_O[6]
rlabel metal2 36576 10122 36576 10122 0 FrameStrobe_O[7]
rlabel metal2 36960 10080 36960 10080 0 FrameStrobe_O[8]
rlabel metal2 34560 9744 34560 9744 0 FrameStrobe_O[9]
rlabel metal2 18624 6342 18624 6342 0 Inst_A_IO_1_bidirectional_frame_config_pass.Q
rlabel metal2 11472 1932 11472 1932 0 Inst_B_IO_1_bidirectional_frame_config_pass.Q
rlabel metal2 39648 7812 39648 7812 0 Inst_C_IO_1_bidirectional_frame_config_pass.Q
rlabel metal2 11808 1932 11808 1932 0 Inst_D_IO_1_bidirectional_frame_config_pass.Q
rlabel metal2 28992 1596 28992 1596 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit0.Q
rlabel metal2 30528 1631 30528 1631 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit1.Q
rlabel metal2 3264 3066 3264 3066 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit10.Q
rlabel metal3 6720 3192 6720 3192 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit11.Q
rlabel via1 7680 5632 7680 5632 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit12.Q
rlabel metal2 7968 3486 7968 3486 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit13.Q
rlabel metal3 8928 5628 8928 5628 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit14.Q
rlabel metal3 1824 2268 1824 2268 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit15.Q
rlabel metal2 1680 1932 1680 1932 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit16.Q
rlabel metal2 1728 9534 1728 9534 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit17.Q
rlabel metal2 4224 7224 4224 7224 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit18.Q
rlabel metal2 1488 5964 1488 5964 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit19.Q
rlabel metal2 9408 2181 9408 2181 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit2.Q
rlabel metal2 1344 7014 1344 7014 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit20.Q
rlabel metal2 2880 8316 2880 8316 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit21.Q
rlabel metal2 10176 7896 10176 7896 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 10416 8148 10416 8148 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit23.Q
rlabel metal2 11328 9030 11328 9030 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit24.Q
rlabel metal2 6528 5964 6528 5964 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit25.Q
rlabel metal2 13536 7224 13536 7224 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit26.Q
rlabel metal3 8112 7980 8112 7980 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit27.Q
rlabel metal2 9120 9198 9120 9198 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit28.Q
rlabel metal3 13296 8652 13296 8652 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit29.Q
rlabel metal2 7872 1974 7872 1974 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit3.Q
rlabel metal2 15072 8612 15072 8612 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit30.Q
rlabel metal2 14544 9240 14544 9240 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit31.Q
rlabel metal2 1344 1050 1344 1050 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit4.Q
rlabel metal2 1632 966 1632 966 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit5.Q
rlabel metal2 14208 2856 14208 2856 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit6.Q
rlabel metal2 12864 2110 12864 2110 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit7.Q
rlabel metal2 1344 4032 1344 4032 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit8.Q
rlabel metal2 1632 2772 1632 2772 0 Inst_N_IO4_ConfigMem.Inst_frame0_bit9.Q
rlabel metal2 26208 2352 26208 2352 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit0.Q
rlabel metal3 27408 1260 27408 1260 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit1.Q
rlabel metal2 28176 2856 28176 2856 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit10.Q
rlabel metal2 29760 3143 29760 3143 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit11.Q
rlabel metal2 24576 3696 24576 3696 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit12.Q
rlabel metal2 25872 4204 25872 4204 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit13.Q
rlabel metal2 12672 5586 12672 5586 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit14.Q
rlabel metal2 14112 5124 14112 5124 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit15.Q
rlabel metal2 31632 7203 31632 7203 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit16.Q
rlabel metal2 30048 7434 30048 7434 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit17.Q
rlabel metal2 13584 6468 13584 6468 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit18.Q
rlabel via1 15216 6463 15216 6463 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit19.Q
rlabel metal3 34080 1260 34080 1260 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit2.Q
rlabel metal2 38688 6636 38688 6636 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit20.Q
rlabel metal3 40368 6636 40368 6636 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit21.Q
rlabel metal2 27072 6720 27072 6720 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit22.Q
rlabel metal2 28704 6720 28704 6720 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit23.Q
rlabel metal2 32352 6468 32352 6468 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit24.Q
rlabel metal2 33984 6927 33984 6927 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit25.Q
rlabel metal2 38784 8190 38784 8190 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit26.Q
rlabel via1 40368 7975 40368 7975 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit27.Q
rlabel metal2 28416 8607 28416 8607 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit28.Q
rlabel metal2 26880 8022 26880 8022 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit29.Q
rlabel metal2 35424 1428 35424 1428 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit3.Q
rlabel metal2 28128 4410 28128 4410 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit30.Q
rlabel metal2 29616 4130 29616 4130 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit31.Q
rlabel metal2 32208 1344 32208 1344 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit4.Q
rlabel metal2 33792 2181 33792 2181 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit5.Q
rlabel metal2 38736 1344 38736 1344 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit6.Q
rlabel metal2 40320 2181 40320 2181 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit7.Q
rlabel metal2 13152 3696 13152 3696 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit8.Q
rlabel metal2 14688 3693 14688 3693 0 Inst_N_IO4_ConfigMem.Inst_frame1_bit9.Q
rlabel metal2 21408 2184 21408 2184 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit0.Q
rlabel metal3 22176 1302 22176 1302 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit1.Q
rlabel metal2 38976 4071 38976 4071 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit10.Q
rlabel metal2 37440 3150 37440 3150 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit11.Q
rlabel metal3 25632 2772 25632 2772 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit12.Q
rlabel metal2 27072 3479 27072 3479 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit13.Q
rlabel metal3 37248 5040 37248 5040 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit14.Q
rlabel metal2 39216 4368 39216 4368 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit15.Q
rlabel metal2 23136 7098 23136 7098 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit16.Q
rlabel metal2 24720 7203 24720 7203 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit17.Q
rlabel metal2 33888 5761 33888 5761 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit18.Q
rlabel metal2 32352 5922 32352 5922 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit19.Q
rlabel metal2 24000 1638 24000 1638 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit2.Q
rlabel via1 19728 6463 19728 6463 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit20.Q
rlabel metal3 17856 6468 17856 6468 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit21.Q
rlabel metal2 25968 5691 25968 5691 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit22.Q
rlabel metal2 24384 5922 24384 5922 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit23.Q
rlabel metal2 23040 8736 23040 8736 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit24.Q
rlabel metal2 24624 8715 24624 8715 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit25.Q
rlabel metal2 35904 8190 35904 8190 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit26.Q
rlabel metal2 37440 7609 37440 7609 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit27.Q
rlabel metal2 25152 8946 25152 8946 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit28.Q
rlabel metal2 26688 8953 26688 8953 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit29.Q
rlabel metal2 25728 1344 25728 1344 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit3.Q
rlabel metal2 29376 5922 29376 5922 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit30.Q
rlabel metal2 31056 5124 31056 5124 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit31.Q
rlabel metal2 19632 1344 19632 1344 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit4.Q
rlabel metal2 18144 1974 18144 1974 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit5.Q
rlabel metal2 38304 2181 38304 2181 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit6.Q
rlabel metal2 36912 1344 36912 1344 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit7.Q
rlabel metal2 23760 1008 23760 1008 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit8.Q
rlabel metal2 21984 2898 21984 2898 0 Inst_N_IO4_ConfigMem.Inst_frame2_bit9.Q
rlabel metal3 9168 1092 9168 1092 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit0.Q
rlabel metal2 11232 1771 11232 1771 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit1.Q
rlabel metal3 30240 3444 30240 3444 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit10.Q
rlabel metal3 31680 2856 31680 2856 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit11.Q
rlabel metal2 16608 4998 16608 4998 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit12.Q
rlabel via2 18144 4953 18144 4953 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit13.Q
rlabel metal2 32352 4419 32352 4419 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit14.Q
rlabel metal3 34176 3612 34176 3612 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit15.Q
rlabel metal2 16608 8610 16608 8610 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit16.Q
rlabel metal2 18144 8229 18144 8229 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit17.Q
rlabel metal2 34656 5460 34656 5460 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit18.Q
rlabel metal2 36192 6169 36192 6169 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit19.Q
rlabel metal3 10128 1008 10128 1008 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit2.Q
rlabel metal2 15792 4179 15792 4179 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit20.Q
rlabel metal2 14208 4032 14208 4032 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit21.Q
rlabel metal2 19488 6307 19488 6307 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit22.Q
rlabel metal2 17952 5964 17952 5964 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit23.Q
rlabel metal2 19536 8715 19536 8715 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit24.Q
rlabel metal2 17904 8652 17904 8652 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit25.Q
rlabel metal2 22752 7137 22752 7137 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit26.Q
rlabel metal2 21216 7854 21216 7854 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit27.Q
rlabel metal2 22176 6685 22176 6685 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit28.Q
rlabel metal2 20640 6300 20640 6300 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit29.Q
rlabel metal2 13152 1008 13152 1008 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit3.Q
rlabel metal2 21792 4074 21792 4074 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit30.Q
rlabel metal2 23376 4179 23376 4179 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit31.Q
rlabel metal2 13920 2184 13920 2184 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit4.Q
rlabel metal3 15168 1260 15168 1260 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit5.Q
rlabel metal3 34848 3612 34848 3612 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit6.Q
rlabel metal2 36432 2772 36432 2772 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit7.Q
rlabel metal2 17520 3612 17520 3612 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit8.Q
rlabel metal2 19104 3866 19104 3866 0 Inst_N_IO4_ConfigMem.Inst_frame3_bit9.Q
rlabel metal2 12096 3157 12096 3157 0 Inst_N_IO4_ConfigMem.Inst_frame4_bit28.Q
rlabel metal2 10560 2730 10560 2730 0 Inst_N_IO4_ConfigMem.Inst_frame4_bit29.Q
rlabel metal2 10752 3486 10752 3486 0 Inst_N_IO4_ConfigMem.Inst_frame4_bit30.Q
rlabel metal2 12288 3567 12288 3567 0 Inst_N_IO4_ConfigMem.Inst_frame4_bit31.Q
rlabel metal2 12288 2604 12288 2604 0 Inst_N_IO4_switch_matrix.S1BEG0
rlabel metal3 12576 3360 12576 3360 0 Inst_N_IO4_switch_matrix.S1BEG1
rlabel metal2 15552 1092 15552 1092 0 Inst_N_IO4_switch_matrix.S1BEG2
rlabel metal3 14256 1848 14256 1848 0 Inst_N_IO4_switch_matrix.S1BEG3
rlabel metal2 15648 2142 15648 2142 0 Inst_N_IO4_switch_matrix.S2BEG0
rlabel metal2 37056 4116 37056 4116 0 Inst_N_IO4_switch_matrix.S2BEG1
rlabel metal2 19968 3654 19968 3654 0 Inst_N_IO4_switch_matrix.S2BEG2
rlabel metal2 32160 3906 32160 3906 0 Inst_N_IO4_switch_matrix.S2BEG3
rlabel metal2 18336 4956 18336 4956 0 Inst_N_IO4_switch_matrix.S2BEG4
rlabel metal2 34464 4116 34464 4116 0 Inst_N_IO4_switch_matrix.S2BEG5
rlabel metal2 20544 8442 20544 8442 0 Inst_N_IO4_switch_matrix.S2BEG6
rlabel metal2 36528 5712 36528 5712 0 Inst_N_IO4_switch_matrix.S2BEG7
rlabel metal2 20832 3738 20832 3738 0 Inst_N_IO4_switch_matrix.S2BEGb0
rlabel metal2 19680 5208 19680 5208 0 Inst_N_IO4_switch_matrix.S2BEGb1
rlabel metal2 19680 8190 19680 8190 0 Inst_N_IO4_switch_matrix.S2BEGb2
rlabel metal2 22848 6132 22848 6132 0 Inst_N_IO4_switch_matrix.S2BEGb3
rlabel metal3 22800 5712 22800 5712 0 Inst_N_IO4_switch_matrix.S2BEGb4
rlabel metal2 22752 3570 22752 3570 0 Inst_N_IO4_switch_matrix.S2BEGb5
rlabel metal3 23520 1848 23520 1848 0 Inst_N_IO4_switch_matrix.S2BEGb6
rlabel metal3 25632 2100 25632 2100 0 Inst_N_IO4_switch_matrix.S2BEGb7
rlabel metal2 23328 1932 23328 1932 0 Inst_N_IO4_switch_matrix.S4BEG0
rlabel metal3 37824 2100 37824 2100 0 Inst_N_IO4_switch_matrix.S4BEG1
rlabel metal2 25632 7854 25632 7854 0 Inst_N_IO4_switch_matrix.S4BEG10
rlabel metal2 37248 6342 37248 6342 0 Inst_N_IO4_switch_matrix.S4BEG11
rlabel metal2 27264 8694 27264 8694 0 Inst_N_IO4_switch_matrix.S4BEG12
rlabel metal2 31344 5712 31344 5712 0 Inst_N_IO4_switch_matrix.S4BEG13
rlabel metal2 31104 2142 31104 2142 0 Inst_N_IO4_switch_matrix.S4BEG14
rlabel metal2 36096 2184 36096 2184 0 Inst_N_IO4_switch_matrix.S4BEG15
rlabel metal2 23712 2604 23712 2604 0 Inst_N_IO4_switch_matrix.S4BEG2
rlabel metal2 40896 2184 40896 2184 0 Inst_N_IO4_switch_matrix.S4BEG3
rlabel metal3 27888 1848 27888 1848 0 Inst_N_IO4_switch_matrix.S4BEG4
rlabel metal2 39648 4368 39648 4368 0 Inst_N_IO4_switch_matrix.S4BEG5
rlabel metal3 25056 7224 25056 7224 0 Inst_N_IO4_switch_matrix.S4BEG6
rlabel metal2 35040 4452 35040 4452 0 Inst_N_IO4_switch_matrix.S4BEG7
rlabel metal2 23904 6132 23904 6132 0 Inst_N_IO4_switch_matrix.S4BEG8
rlabel metal3 26304 5712 26304 5712 0 Inst_N_IO4_switch_matrix.S4BEG9
rlabel metal2 33984 2142 33984 2142 0 Inst_N_IO4_switch_matrix.SS4BEG0
rlabel metal2 40512 1596 40512 1596 0 Inst_N_IO4_switch_matrix.SS4BEG1
rlabel metal2 35040 4956 35040 4956 0 Inst_N_IO4_switch_matrix.SS4BEG10
rlabel metal2 40656 7224 40656 7224 0 Inst_N_IO4_switch_matrix.SS4BEG11
rlabel metal2 29376 7644 29376 7644 0 Inst_N_IO4_switch_matrix.SS4BEG12
rlabel metal3 30816 1932 30816 1932 0 Inst_N_IO4_switch_matrix.SS4BEG13
rlabel metal3 31344 1848 31344 1848 0 Inst_N_IO4_switch_matrix.SS4BEG14
rlabel metal2 31488 1932 31488 1932 0 Inst_N_IO4_switch_matrix.SS4BEG15
rlabel metal2 27648 3444 27648 3444 0 Inst_N_IO4_switch_matrix.SS4BEG2
rlabel metal3 29712 3612 29712 3612 0 Inst_N_IO4_switch_matrix.SS4BEG3
rlabel metal2 28032 2100 28032 2100 0 Inst_N_IO4_switch_matrix.SS4BEG4
rlabel metal2 14400 4830 14400 4830 0 Inst_N_IO4_switch_matrix.SS4BEG5
rlabel metal3 31968 7224 31968 7224 0 Inst_N_IO4_switch_matrix.SS4BEG6
rlabel metal4 17760 6384 17760 6384 0 Inst_N_IO4_switch_matrix.SS4BEG7
rlabel metal2 40128 6006 40128 6006 0 Inst_N_IO4_switch_matrix.SS4BEG8
rlabel metal2 28752 4872 28752 4872 0 Inst_N_IO4_switch_matrix.SS4BEG9
rlabel metal2 9792 1260 9792 1260 0 N1END[0]
rlabel metal2 10176 966 10176 966 0 N1END[1]
rlabel metal2 9888 828 9888 828 0 N1END[2]
rlabel metal2 11328 1806 11328 1806 0 N1END[3]
rlabel metal2 24384 2184 24384 2184 0 N2END[0]
rlabel metal2 21504 1638 21504 1638 0 N2END[1]
rlabel metal2 12192 660 12192 660 0 N2END[2]
rlabel metal2 12384 583 12384 583 0 N2END[3]
rlabel metal2 1824 3612 1824 3612 0 N2END[4]
rlabel metal2 1776 4872 1776 4872 0 N2END[5]
rlabel metal2 1536 2058 1536 2058 0 N2END[6]
rlabel metal2 13488 1176 13488 1176 0 N2END[7]
rlabel metal4 28320 1470 28320 1470 0 N2MID[0]
rlabel metal2 11520 7140 11520 7140 0 N2MID[1]
rlabel metal3 29184 1848 29184 1848 0 N2MID[2]
rlabel metal2 13728 6174 13728 6174 0 N2MID[3]
rlabel metal3 23940 1470 23940 1470 0 N2MID[4]
rlabel metal2 14016 6384 14016 6384 0 N2MID[5]
rlabel via2 11424 72 11424 72 0 N2MID[6]
rlabel metal2 14016 1848 14016 1848 0 N2MID[7]
rlabel metal3 24768 1974 24768 1974 0 N4END[0]
rlabel metal2 39360 2352 39360 2352 0 N4END[10]
rlabel metal2 15456 576 15456 576 0 N4END[11]
rlabel metal2 15648 408 15648 408 0 N4END[12]
rlabel metal2 15840 240 15840 240 0 N4END[13]
rlabel metal3 21456 504 21456 504 0 N4END[14]
rlabel metal2 16224 408 16224 408 0 N4END[15]
rlabel metal2 21888 2142 21888 2142 0 N4END[1]
rlabel via2 13728 72 13728 72 0 N4END[2]
rlabel metal2 13920 366 13920 366 0 N4END[3]
rlabel metal2 14112 240 14112 240 0 N4END[4]
rlabel metal2 14304 1122 14304 1122 0 N4END[5]
rlabel metal2 38880 3528 38880 3528 0 N4END[6]
rlabel metal2 14400 1386 14400 1386 0 N4END[7]
rlabel metal2 39264 1806 39264 1806 0 N4END[8]
rlabel metal3 22032 1176 22032 1176 0 N4END[9]
rlabel metal2 24864 1722 24864 1722 0 NN4END[0]
rlabel metal2 38016 3780 38016 3780 0 NN4END[10]
rlabel metal2 17664 4830 17664 4830 0 NN4END[11]
rlabel metal2 18720 870 18720 870 0 NN4END[12]
rlabel metal2 18912 702 18912 702 0 NN4END[13]
rlabel metal3 19488 1512 19488 1512 0 NN4END[14]
rlabel metal2 18720 1806 18720 1806 0 NN4END[15]
rlabel metal2 21984 2100 21984 2100 0 NN4END[1]
rlabel metal2 16800 450 16800 450 0 NN4END[2]
rlabel metal2 17184 5208 17184 5208 0 NN4END[3]
rlabel metal2 17184 1290 17184 1290 0 NN4END[4]
rlabel metal2 17376 1164 17376 1164 0 NN4END[5]
rlabel metal2 17568 1290 17568 1290 0 NN4END[6]
rlabel metal2 17760 1080 17760 1080 0 NN4END[7]
rlabel metal2 25344 1890 25344 1890 0 NN4END[8]
rlabel metal2 22464 2016 22464 2016 0 NN4END[9]
rlabel metal2 15744 2352 15744 2352 0 S1BEG[0]
rlabel metal2 19872 156 19872 156 0 S1BEG[1]
rlabel metal2 20064 282 20064 282 0 S1BEG[2]
rlabel metal2 20256 324 20256 324 0 S1BEG[3]
rlabel metal2 20448 324 20448 324 0 S2BEG[0]
rlabel metal2 20640 618 20640 618 0 S2BEG[1]
rlabel metal2 20496 3192 20496 3192 0 S2BEG[2]
rlabel metal2 21024 282 21024 282 0 S2BEG[3]
rlabel metal2 21216 408 21216 408 0 S2BEG[4]
rlabel metal2 21408 324 21408 324 0 S2BEG[5]
rlabel metal2 21504 3864 21504 3864 0 S2BEG[6]
rlabel metal2 21792 492 21792 492 0 S2BEG[7]
rlabel metal2 21984 450 21984 450 0 S2BEGb[0]
rlabel metal2 22176 576 22176 576 0 S2BEGb[1]
rlabel metal2 22368 492 22368 492 0 S2BEGb[2]
rlabel metal2 22560 1248 22560 1248 0 S2BEGb[3]
rlabel metal2 22800 3192 22800 3192 0 S2BEGb[4]
rlabel metal2 22944 828 22944 828 0 S2BEGb[5]
rlabel metal2 23136 870 23136 870 0 S2BEGb[6]
rlabel metal2 23328 702 23328 702 0 S2BEGb[7]
rlabel metal2 23520 870 23520 870 0 S4BEG[0]
rlabel metal2 25440 492 25440 492 0 S4BEG[10]
rlabel metal2 25632 576 25632 576 0 S4BEG[11]
rlabel metal2 27072 8022 27072 8022 0 S4BEG[12]
rlabel metal2 26016 618 26016 618 0 S4BEG[13]
rlabel metal2 26208 744 26208 744 0 S4BEG[14]
rlabel metal2 26400 912 26400 912 0 S4BEG[15]
rlabel metal2 23712 282 23712 282 0 S4BEG[1]
rlabel metal2 23904 660 23904 660 0 S4BEG[2]
rlabel metal2 24096 450 24096 450 0 S4BEG[3]
rlabel metal2 24288 492 24288 492 0 S4BEG[4]
rlabel metal4 37824 1050 37824 1050 0 S4BEG[5]
rlabel metal2 24864 4788 24864 4788 0 S4BEG[6]
rlabel metal2 24864 114 24864 114 0 S4BEG[7]
rlabel metal3 24576 3024 24576 3024 0 S4BEG[8]
rlabel metal2 25248 996 25248 996 0 S4BEG[9]
rlabel metal2 37248 4662 37248 4662 0 SS4BEG[0]
rlabel metal2 28512 366 28512 366 0 SS4BEG[10]
rlabel metal3 40464 6972 40464 6972 0 SS4BEG[11]
rlabel metal2 28896 576 28896 576 0 SS4BEG[12]
rlabel metal2 29088 492 29088 492 0 SS4BEG[13]
rlabel metal2 29280 870 29280 870 0 SS4BEG[14]
rlabel metal2 29472 702 29472 702 0 SS4BEG[15]
rlabel metal2 40320 504 40320 504 0 SS4BEG[1]
rlabel metal2 26976 996 26976 996 0 SS4BEG[2]
rlabel metal2 27168 114 27168 114 0 SS4BEG[3]
rlabel metal2 27360 870 27360 870 0 SS4BEG[4]
rlabel metal2 27552 198 27552 198 0 SS4BEG[5]
rlabel metal2 27744 1290 27744 1290 0 SS4BEG[6]
rlabel metal2 27936 618 27936 618 0 SS4BEG[7]
rlabel metal4 37920 2856 37920 2856 0 SS4BEG[8]
rlabel metal2 28320 1206 28320 1206 0 SS4BEG[9]
rlabel metal2 31872 9114 31872 9114 0 UserCLK
rlabel metal2 35520 7434 35520 7434 0 UserCLK_regs
rlabel via2 16800 10680 16800 10680 0 UserCLKo
rlabel metal3 1872 1764 1872 1764 0 _000_
rlabel metal2 1200 5628 1200 5628 0 _001_
rlabel metal2 5088 9156 5088 9156 0 _002_
rlabel metal2 10272 5544 10272 5544 0 _003_
rlabel metal2 3360 3696 3360 3696 0 _004_
rlabel metal3 3312 2604 3312 2604 0 _005_
rlabel metal2 3360 5712 3360 5712 0 _006_
rlabel metal2 5424 2604 5424 2604 0 _007_
rlabel metal2 3456 3402 3456 3402 0 _008_
rlabel metal2 2976 9030 2976 9030 0 _009_
rlabel metal2 1344 1596 1344 1596 0 _010_
rlabel metal2 4512 7182 4512 7182 0 _011_
rlabel metal3 4320 1176 4320 1176 0 _012_
rlabel metal2 2016 7224 2016 7224 0 _013_
rlabel metal2 12768 8652 12768 8652 0 _014_
rlabel metal3 11904 6468 11904 6468 0 _015_
rlabel metal2 9792 8442 9792 8442 0 _016_
rlabel metal2 9936 8148 9936 8148 0 _017_
rlabel metal2 11616 7014 11616 7014 0 _018_
rlabel metal2 14112 7476 14112 7476 0 _019_
rlabel metal2 15408 8484 15408 8484 0 _020_
rlabel metal2 15744 7980 15744 7980 0 _021_
rlabel metal2 14304 7560 14304 7560 0 _022_
rlabel metal2 15696 8148 15696 8148 0 _023_
rlabel metal3 11664 7140 11664 7140 0 _024_
rlabel metal2 13728 8358 13728 8358 0 _025_
rlabel metal2 13632 7518 13632 7518 0 _026_
rlabel metal3 8448 7392 8448 7392 0 _027_
rlabel metal3 4896 4998 4896 4998 0 _028_
rlabel metal3 8208 9492 8208 9492 0 _029_
rlabel metal2 8221 7804 8221 7804 0 _030_
rlabel metal2 7968 8610 7968 8610 0 _031_
rlabel metal2 6768 6636 6768 6636 0 _032_
rlabel metal2 9408 8022 9408 8022 0 _033_
rlabel metal2 9504 8064 9504 8064 0 _034_
rlabel metal2 8832 7518 8832 7518 0 _035_
rlabel metal2 8880 6636 8880 6636 0 _036_
rlabel metal2 9264 9492 9264 9492 0 _037_
rlabel metal2 9408 9072 9408 9072 0 _038_
rlabel metal2 3504 4956 3504 4956 0 _039_
rlabel metal2 1392 6048 1392 6048 0 _040_
rlabel metal2 1296 6216 1296 6216 0 _041_
rlabel metal2 3168 5082 3168 5082 0 _042_
rlabel metal2 2016 8442 2016 8442 0 _043_
rlabel metal2 4512 9576 4512 9576 0 _044_
rlabel metal2 3744 5712 3744 5712 0 _045_
rlabel metal2 1344 5418 1344 5418 0 _046_
rlabel metal2 5376 8946 5376 8946 0 _047_
rlabel metal2 5520 6300 5520 6300 0 _048_
rlabel metal2 5232 7140 5232 7140 0 _049_
rlabel metal2 6048 7434 6048 7434 0 _050_
rlabel metal2 5472 7266 5472 7266 0 _051_
rlabel via2 5184 8482 5184 8482 0 _052_
rlabel metal3 8784 5040 8784 5040 0 _053_
rlabel metal2 10368 5712 10368 5712 0 _054_
rlabel metal3 5424 4116 5424 4116 0 _055_
rlabel metal3 6480 3276 6480 3276 0 _056_
rlabel metal3 7920 4116 7920 4116 0 _057_
rlabel metal2 9888 5712 9888 5712 0 _058_
rlabel metal2 9792 5838 9792 5838 0 _059_
rlabel metal2 8256 3612 8256 3612 0 _060_
rlabel metal2 8352 3738 8352 3738 0 _061_
rlabel metal2 9216 5040 9216 5040 0 _062_
rlabel metal2 9408 5544 9408 5544 0 _063_
rlabel metal2 4128 1260 4128 1260 0 _064_
rlabel metal2 12960 3066 12960 3066 0 _065_
rlabel metal2 1632 1386 1632 1386 0 _066_
rlabel metal3 7056 2352 7056 2352 0 _067_
rlabel metal2 14400 2688 14400 2688 0 _068_
rlabel metal2 14304 3192 14304 3192 0 _069_
rlabel metal2 1344 2982 1344 2982 0 _070_
rlabel metal2 15360 1764 15360 1764 0 _071_
rlabel metal3 14016 2268 14016 2268 0 _072_
rlabel metal3 13536 1932 13536 1932 0 _073_
rlabel metal3 12768 1974 12768 1974 0 _074_
rlabel metal3 7152 1092 7152 1092 0 _075_
rlabel metal2 7152 924 7152 924 0 _076_
rlabel metal2 10464 1596 10464 1596 0 _077_
rlabel metal3 10128 2100 10128 2100 0 _078_
rlabel metal2 37824 7728 37824 7728 0 _079_
rlabel metal2 36768 7224 36768 7224 0 _080_
rlabel metal2 29616 7308 29616 7308 0 _081_
rlabel metal2 36384 6468 36384 6468 0 _082_
rlabel metal2 31104 9030 31104 9030 0 clknet_0_UserCLK
rlabel metal2 34560 8022 34560 8022 0 clknet_0_UserCLK_regs
rlabel metal3 31680 8820 31680 8820 0 clknet_1_0__leaf_UserCLK
rlabel metal2 30240 8946 30240 8946 0 clknet_1_0__leaf_UserCLK_regs
rlabel metal3 35712 7980 35712 7980 0 clknet_1_1__leaf_UserCLK_regs
<< properties >>
string FIXED_BBOX 0 0 43008 10752
<< end >>
