* NGSPICE file created from heichips25_example_large.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_2 abstract view
.subckt sg13g2_a21oi_2 VSS VDD B1 Y A2 A1
.ends

.subckt heichips25_example_large VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2]
+ ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3]
+ uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3]
+ uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3]
+ uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3]
+ uo_out[4] uo_out[5] uo_out[6] uo_out[7]
XFILLER_95_851 VPWR VGND sg13g2_decap_8
XFILLER_67_553 VPWR VGND sg13g2_decap_8
XFILLER_94_350 VPWR VGND sg13g2_decap_8
XFILLER_27_417 VPWR VGND sg13g2_decap_8
XFILLER_39_277 VPWR VGND sg13g2_decap_8
XFILLER_54_214 VPWR VGND sg13g2_decap_8
XFILLER_82_567 VPWR VGND sg13g2_decap_8
XFILLER_70_707 VPWR VGND sg13g2_decap_8
XFILLER_36_973 VPWR VGND sg13g2_decap_8
XFILLER_63_770 VPWR VGND sg13g2_decap_8
XFILLER_51_921 VPWR VGND sg13g2_decap_8
XFILLER_23_623 VPWR VGND sg13g2_decap_8
XFILLER_35_483 VPWR VGND sg13g2_decap_8
XFILLER_62_280 VPWR VGND sg13g2_decap_8
XFILLER_50_420 VPWR VGND sg13g2_decap_8
XFILLER_51_998 VPWR VGND sg13g2_decap_8
XFILLER_22_144 VPWR VGND sg13g2_decap_8
XFILLER_50_497 VPWR VGND sg13g2_decap_8
XFILLER_105_945 VPWR VGND sg13g2_decap_8
XFILLER_104_455 VPWR VGND sg13g2_decap_8
XFILLER_89_133 VPWR VGND sg13g2_decap_8
XFILLER_78_818 VPWR VGND sg13g2_decap_8
XFILLER_86_851 VPWR VGND sg13g2_decap_8
XFILLER_100_672 VPWR VGND sg13g2_decap_8
XFILLER_85_350 VPWR VGND sg13g2_decap_8
XFILLER_73_501 VPWR VGND sg13g2_decap_8
XFILLER_58_553 VPWR VGND sg13g2_decap_8
XFILLER_46_704 VPWR VGND sg13g2_decap_8
XFILLER_18_406 VPWR VGND sg13g2_decap_8
XFILLER_93_47 VPWR VGND sg13g2_decap_8
XFILLER_45_203 VPWR VGND sg13g2_decap_8
XFILLER_73_578 VPWR VGND sg13g2_decap_8
XFILLER_61_718 VPWR VGND sg13g2_decap_8
XFILLER_60_228 VPWR VGND sg13g2_decap_8
XFILLER_54_781 VPWR VGND sg13g2_decap_8
XFILLER_42_921 VPWR VGND sg13g2_decap_8
XFILLER_14_623 VPWR VGND sg13g2_decap_8
XFILLER_26_63 VPWR VGND sg13g2_decap_8
XFILLER_26_483 VPWR VGND sg13g2_decap_8
XFILLER_27_984 VPWR VGND sg13g2_decap_8
XFILLER_53_280 VPWR VGND sg13g2_decap_8
XFILLER_13_133 VPWR VGND sg13g2_decap_8
XFILLER_41_420 VPWR VGND sg13g2_decap_8
XFILLER_42_998 VPWR VGND sg13g2_decap_8
XFILLER_9_126 VPWR VGND sg13g2_decap_8
XFILLER_41_497 VPWR VGND sg13g2_decap_8
XFILLER_42_95 VPWR VGND sg13g2_decap_8
XFILLER_10_851 VPWR VGND sg13g2_decap_8
XFILLER_6_833 VPWR VGND sg13g2_decap_8
XFILLER_5_354 VPWR VGND sg13g2_decap_8
XFILLER_96_637 VPWR VGND sg13g2_decap_8
XFILLER_68_306 VPWR VGND sg13g2_decap_8
XFILLER_3_56 VPWR VGND sg13g2_decap_8
XFILLER_1_560 VPWR VGND sg13g2_decap_8
XFILLER_77_840 VPWR VGND sg13g2_decap_8
XFILLER_95_158 VPWR VGND sg13g2_decap_8
XFILLER_76_361 VPWR VGND sg13g2_decap_8
XFILLER_67_70 VPWR VGND sg13g2_decap_8
XFILLER_64_501 VPWR VGND sg13g2_decap_8
XFILLER_49_564 VPWR VGND sg13g2_decap_8
XFILLER_37_704 VPWR VGND sg13g2_decap_8
XFILLER_36_203 VPWR VGND sg13g2_decap_8
XFILLER_92_854 VPWR VGND sg13g2_decap_8
XFILLER_64_578 VPWR VGND sg13g2_decap_8
XFILLER_52_707 VPWR VGND sg13g2_decap_8
XFILLER_18_973 VPWR VGND sg13g2_decap_8
XFILLER_91_364 VPWR VGND sg13g2_decap_8
XFILLER_51_228 VPWR VGND sg13g2_decap_8
XFILLER_45_770 VPWR VGND sg13g2_decap_8
XFILLER_33_910 VPWR VGND sg13g2_decap_8
XFILLER_44_291 VPWR VGND sg13g2_decap_8
XFILLER_17_494 VPWR VGND sg13g2_decap_8
XFILLER_32_431 VPWR VGND sg13g2_decap_8
XFILLER_33_987 VPWR VGND sg13g2_decap_8
XFILLER_60_795 VPWR VGND sg13g2_decap_8
XFILLER_20_648 VPWR VGND sg13g2_decap_8
XFILLER_9_693 VPWR VGND sg13g2_decap_8
XFILLER_99_420 VPWR VGND sg13g2_decap_8
XFILLER_99_497 VPWR VGND sg13g2_decap_8
XFILLER_87_637 VPWR VGND sg13g2_decap_8
XFILLER_59_306 VPWR VGND sg13g2_decap_8
XFILLER_102_959 VPWR VGND sg13g2_decap_8
XFILLER_101_469 VPWR VGND sg13g2_decap_8
XFILLER_86_158 VPWR VGND sg13g2_decap_8
XFILLER_74_309 VPWR VGND sg13g2_decap_8
XFILLER_68_873 VPWR VGND sg13g2_decap_8
XFILLER_67_350 VPWR VGND sg13g2_decap_8
XFILLER_27_214 VPWR VGND sg13g2_decap_8
XFILLER_103_35 VPWR VGND sg13g2_decap_8
XFILLER_83_865 VPWR VGND sg13g2_decap_8
XFILLER_55_567 VPWR VGND sg13g2_decap_8
XFILLER_43_707 VPWR VGND sg13g2_decap_8
XFILLER_82_364 VPWR VGND sg13g2_decap_8
XFILLER_70_504 VPWR VGND sg13g2_decap_8
XFILLER_63_28 VPWR VGND sg13g2_decap_8
XFILLER_42_228 VPWR VGND sg13g2_decap_8
XFILLER_24_921 VPWR VGND sg13g2_decap_8
XFILLER_36_770 VPWR VGND sg13g2_decap_8
XFILLER_23_420 VPWR VGND sg13g2_decap_8
XFILLER_35_280 VPWR VGND sg13g2_decap_8
XFILLER_24_998 VPWR VGND sg13g2_decap_8
XFILLER_51_795 VPWR VGND sg13g2_decap_8
XFILLER_50_294 VPWR VGND sg13g2_decap_8
XFILLER_11_637 VPWR VGND sg13g2_decap_8
XFILLER_23_497 VPWR VGND sg13g2_decap_8
XFILLER_10_158 VPWR VGND sg13g2_decap_8
XFILLER_12_32 VPWR VGND sg13g2_decap_8
XFILLER_88_25 VPWR VGND sg13g2_decap_8
XFILLER_3_847 VPWR VGND sg13g2_decap_8
XFILLER_105_742 VPWR VGND sg13g2_decap_8
XFILLER_5_4 VPWR VGND sg13g2_decap_8
XFILLER_104_252 VPWR VGND sg13g2_decap_8
XFILLER_78_615 VPWR VGND sg13g2_decap_8
XFILLER_2_368 VPWR VGND sg13g2_decap_8
XFILLER_77_147 VPWR VGND sg13g2_decap_8
XFILLER_93_607 VPWR VGND sg13g2_decap_8
XFILLER_59_873 VPWR VGND sg13g2_decap_8
XFILLER_58_350 VPWR VGND sg13g2_decap_8
XFILLER_46_501 VPWR VGND sg13g2_decap_8
XFILLER_18_203 VPWR VGND sg13g2_decap_8
XFILLER_74_876 VPWR VGND sg13g2_decap_8
XFILLER_73_375 VPWR VGND sg13g2_decap_8
XFILLER_61_515 VPWR VGND sg13g2_decap_8
XFILLER_46_578 VPWR VGND sg13g2_decap_8
XFILLER_15_921 VPWR VGND sg13g2_decap_8
XFILLER_27_781 VPWR VGND sg13g2_decap_8
XFILLER_33_217 VPWR VGND sg13g2_decap_8
XFILLER_34_718 VPWR VGND sg13g2_decap_8
XFILLER_37_95 VPWR VGND sg13g2_decap_8
XFILLER_14_420 VPWR VGND sg13g2_decap_8
XFILLER_26_280 VPWR VGND sg13g2_decap_8
XFILLER_15_998 VPWR VGND sg13g2_decap_8
XFILLER_18_1015 VPWR VGND sg13g2_decap_8
XFILLER_30_924 VPWR VGND sg13g2_decap_8
XFILLER_42_795 VPWR VGND sg13g2_decap_8
XFILLER_14_497 VPWR VGND sg13g2_decap_8
XFILLER_41_294 VPWR VGND sg13g2_decap_8
XFILLER_6_630 VPWR VGND sg13g2_decap_8
XFILLER_5_151 VPWR VGND sg13g2_decap_8
XFILLER_97_924 VPWR VGND sg13g2_decap_8
XFILLER_68_103 VPWR VGND sg13g2_decap_8
XFILLER_96_434 VPWR VGND sg13g2_decap_8
XFILLER_69_659 VPWR VGND sg13g2_decap_8
XFILLER_25_1008 VPWR VGND sg13g2_decap_8
XFILLER_49_361 VPWR VGND sg13g2_decap_8
XFILLER_37_501 VPWR VGND sg13g2_decap_8
XFILLER_92_651 VPWR VGND sg13g2_decap_8
XFILLER_65_854 VPWR VGND sg13g2_decap_8
XFILLER_25_707 VPWR VGND sg13g2_decap_8
XFILLER_91_161 VPWR VGND sg13g2_decap_8
XFILLER_64_375 VPWR VGND sg13g2_decap_8
XFILLER_52_504 VPWR VGND sg13g2_decap_8
XFILLER_18_770 VPWR VGND sg13g2_decap_8
XFILLER_37_578 VPWR VGND sg13g2_decap_8
XFILLER_80_868 VPWR VGND sg13g2_decap_8
XFILLER_17_291 VPWR VGND sg13g2_decap_8
XFILLER_24_228 VPWR VGND sg13g2_decap_8
XFILLER_71_1028 VPWR VGND sg13g2_fill_1
XFILLER_60_592 VPWR VGND sg13g2_decap_8
XFILLER_21_924 VPWR VGND sg13g2_decap_8
XFILLER_33_784 VPWR VGND sg13g2_decap_8
XFILLER_20_445 VPWR VGND sg13g2_decap_8
XFILLER_9_490 VPWR VGND sg13g2_decap_8
XFILLER_106_539 VPWR VGND sg13g2_decap_8
XFILLER_88_935 VPWR VGND sg13g2_decap_8
XFILLER_58_28 VPWR VGND sg13g2_decap_8
XFILLER_102_756 VPWR VGND sg13g2_decap_8
XFILLER_99_294 VPWR VGND sg13g2_decap_8
XFILLER_87_434 VPWR VGND sg13g2_decap_8
XFILLER_101_266 VPWR VGND sg13g2_decap_8
XFILLER_74_106 VPWR VGND sg13g2_decap_8
XFILLER_68_670 VPWR VGND sg13g2_decap_8
XFILLER_74_49 VPWR VGND sg13g2_decap_4
XFILLER_71_802 VPWR VGND sg13g2_decap_8
XFILLER_56_865 VPWR VGND sg13g2_decap_8
XFILLER_16_707 VPWR VGND sg13g2_decap_8
XFILLER_28_567 VPWR VGND sg13g2_decap_8
XFILLER_83_662 VPWR VGND sg13g2_decap_8
XFILLER_82_161 VPWR VGND sg13g2_decap_8
XFILLER_70_301 VPWR VGND sg13g2_decap_8
XFILLER_55_364 VPWR VGND sg13g2_decap_8
XFILLER_43_504 VPWR VGND sg13g2_decap_8
XFILLER_15_228 VPWR VGND sg13g2_decap_8
XFILLER_71_879 VPWR VGND sg13g2_decap_8
XFILLER_70_378 VPWR VGND sg13g2_decap_8
XFILLER_51_592 VPWR VGND sg13g2_decap_8
XFILLER_12_935 VPWR VGND sg13g2_decap_8
XFILLER_24_795 VPWR VGND sg13g2_decap_8
XFILLER_8_917 VPWR VGND sg13g2_decap_8
XFILLER_11_434 VPWR VGND sg13g2_decap_8
XFILLER_23_42 VPWR VGND sg13g2_decap_8
XFILLER_23_294 VPWR VGND sg13g2_decap_8
XFILLER_7_438 VPWR VGND sg13g2_decap_8
XFILLER_99_35 VPWR VGND sg13g2_decap_8
XFILLER_48_1008 VPWR VGND sg13g2_decap_8
XFILLER_3_644 VPWR VGND sg13g2_decap_8
XFILLER_79_935 VPWR VGND sg13g2_decap_8
XFILLER_78_412 VPWR VGND sg13g2_decap_8
XFILLER_2_165 VPWR VGND sg13g2_decap_8
XFILLER_93_404 VPWR VGND sg13g2_decap_8
XFILLER_94_938 VPWR VGND sg13g2_decap_8
XFILLER_78_489 VPWR VGND sg13g2_decap_8
XFILLER_66_629 VPWR VGND sg13g2_decap_8
XFILLER_59_670 VPWR VGND sg13g2_decap_8
XFILLER_47_854 VPWR VGND sg13g2_decap_8
XFILLER_0_35 VPWR VGND sg13g2_decap_8
XFILLER_74_673 VPWR VGND sg13g2_decap_8
XFILLER_46_375 VPWR VGND sg13g2_decap_8
XFILLER_19_567 VPWR VGND sg13g2_decap_8
XFILLER_34_515 VPWR VGND sg13g2_decap_8
XFILLER_73_172 VPWR VGND sg13g2_decap_8
XFILLER_64_60 VPWR VGND sg13g2_decap_8
XFILLER_62_868 VPWR VGND sg13g2_decap_8
XFILLER_61_312 VPWR VGND sg13g2_decap_8
XFILLER_61_389 VPWR VGND sg13g2_decap_8
XFILLER_42_592 VPWR VGND sg13g2_decap_8
XFILLER_15_795 VPWR VGND sg13g2_decap_8
XFILLER_30_721 VPWR VGND sg13g2_decap_8
XFILLER_9_77 VPWR VGND sg13g2_decap_8
XFILLER_14_294 VPWR VGND sg13g2_decap_8
XFILLER_80_70 VPWR VGND sg13g2_decap_8
XFILLER_30_798 VPWR VGND sg13g2_decap_8
XFILLER_31_1001 VPWR VGND sg13g2_decap_8
XFILLER_97_721 VPWR VGND sg13g2_decap_8
XFILLER_96_231 VPWR VGND sg13g2_decap_8
XFILLER_69_456 VPWR VGND sg13g2_decap_8
XFILLER_97_798 VPWR VGND sg13g2_decap_8
XFILLER_85_938 VPWR VGND sg13g2_decap_8
XFILLER_84_448 VPWR VGND sg13g2_decap_8
XFILLER_65_651 VPWR VGND sg13g2_decap_8
XFILLER_38_854 VPWR VGND sg13g2_decap_8
XFILLER_93_971 VPWR VGND sg13g2_decap_8
XFILLER_71_109 VPWR VGND sg13g2_decap_8
X_49_ _17_ _13_ _15_ VPWR VGND sg13g2_nand2_1
XFILLER_52_301 VPWR VGND sg13g2_decap_8
XFILLER_25_504 VPWR VGND sg13g2_decap_8
XFILLER_37_375 VPWR VGND sg13g2_decap_8
XFILLER_64_172 VPWR VGND sg13g2_decap_8
XFILLER_53_868 VPWR VGND sg13g2_decap_8
XFILLER_80_665 VPWR VGND sg13g2_decap_8
XFILLER_52_378 VPWR VGND sg13g2_decap_8
XFILLER_40_518 VPWR VGND sg13g2_decap_8
XFILLER_100_14 VPWR VGND sg13g2_decap_8
XFILLER_21_721 VPWR VGND sg13g2_decap_8
XFILLER_33_581 VPWR VGND sg13g2_decap_8
XFILLER_60_18 VPWR VGND sg13g2_fill_2
XFILLER_20_242 VPWR VGND sg13g2_decap_8
XFILLER_21_798 VPWR VGND sg13g2_decap_8
XFILLER_106_336 VPWR VGND sg13g2_decap_8
XFILLER_69_49 VPWR VGND sg13g2_decap_8
XFILLER_88_732 VPWR VGND sg13g2_decap_8
XFILLER_102_553 VPWR VGND sg13g2_decap_8
XFILLER_87_231 VPWR VGND sg13g2_decap_8
XFILLER_0_658 VPWR VGND sg13g2_decap_8
XFILLER_76_949 VPWR VGND sg13g2_decap_8
XFILLER_75_448 VPWR VGND sg13g2_decap_8
XFILLER_18_42 VPWR VGND sg13g2_decap_8
XFILLER_29_865 VPWR VGND sg13g2_decap_8
XFILLER_56_662 VPWR VGND sg13g2_decap_8
XFILLER_55_161 VPWR VGND sg13g2_decap_8
XFILLER_44_802 VPWR VGND sg13g2_decap_8
XFILLER_43_301 VPWR VGND sg13g2_decap_8
XFILLER_16_504 VPWR VGND sg13g2_decap_8
XFILLER_28_364 VPWR VGND sg13g2_decap_8
XFILLER_71_676 VPWR VGND sg13g2_decap_8
XFILLER_44_879 VPWR VGND sg13g2_decap_8
XFILLER_31_518 VPWR VGND sg13g2_decap_8
XFILLER_70_175 VPWR VGND sg13g2_decap_8
XFILLER_54_1012 VPWR VGND sg13g2_decap_8
XFILLER_43_378 VPWR VGND sg13g2_decap_8
XFILLER_11_231 VPWR VGND sg13g2_decap_8
XFILLER_12_732 VPWR VGND sg13g2_decap_8
XFILLER_24_592 VPWR VGND sg13g2_decap_8
XFILLER_34_74 VPWR VGND sg13g2_decap_8
XFILLER_8_714 VPWR VGND sg13g2_decap_8
XFILLER_7_235 VPWR VGND sg13g2_decap_8
XFILLER_50_84 VPWR VGND sg13g2_decap_8
XFILLER_4_931 VPWR VGND sg13g2_decap_8
XFILLER_98_529 VPWR VGND sg13g2_decap_8
XFILLER_3_441 VPWR VGND sg13g2_decap_8
XFILLER_79_732 VPWR VGND sg13g2_decap_8
XFILLER_59_71 VPWR VGND sg13g2_fill_1
XFILLER_59_60 VPWR VGND sg13g2_decap_8
XFILLER_61_1005 VPWR VGND sg13g2_decap_8
XFILLER_94_735 VPWR VGND sg13g2_decap_8
XFILLER_93_201 VPWR VGND sg13g2_decap_8
XFILLER_78_286 VPWR VGND sg13g2_decap_8
XFILLER_67_938 VPWR VGND sg13g2_decap_8
XFILLER_66_426 VPWR VGND sg13g2_decap_8
XFILLER_93_278 VPWR VGND sg13g2_decap_8
XFILLER_75_70 VPWR VGND sg13g2_decap_8
XFILLER_47_651 VPWR VGND sg13g2_decap_8
XFILLER_19_364 VPWR VGND sg13g2_decap_8
XFILLER_74_470 VPWR VGND sg13g2_decap_8
XFILLER_46_172 VPWR VGND sg13g2_decap_8
XFILLER_34_312 VPWR VGND sg13g2_decap_8
XFILLER_90_963 VPWR VGND sg13g2_decap_8
XFILLER_62_665 VPWR VGND sg13g2_decap_8
XFILLER_50_805 VPWR VGND sg13g2_decap_8
XFILLER_35_868 VPWR VGND sg13g2_decap_8
XFILLER_61_186 VPWR VGND sg13g2_decap_8
XFILLER_22_529 VPWR VGND sg13g2_decap_8
XFILLER_34_389 VPWR VGND sg13g2_decap_8
XFILLER_91_91 VPWR VGND sg13g2_decap_8
XFILLER_15_592 VPWR VGND sg13g2_decap_8
XFILLER_30_595 VPWR VGND sg13g2_decap_8
XFILLER_89_518 VPWR VGND sg13g2_decap_8
XFILLER_69_253 VPWR VGND sg13g2_decap_8
XFILLER_97_595 VPWR VGND sg13g2_decap_8
XFILLER_85_735 VPWR VGND sg13g2_decap_8
XFILLER_58_938 VPWR VGND sg13g2_decap_8
XFILLER_84_245 VPWR VGND sg13g2_decap_8
XFILLER_57_448 VPWR VGND sg13g2_decap_8
XFILLER_77_1001 VPWR VGND sg13g2_decap_8
XFILLER_44_109 VPWR VGND sg13g2_decap_8
XFILLER_38_651 VPWR VGND sg13g2_decap_8
XFILLER_66_993 VPWR VGND sg13g2_decap_8
XFILLER_25_301 VPWR VGND sg13g2_decap_8
XFILLER_37_172 VPWR VGND sg13g2_decap_8
XFILLER_81_963 VPWR VGND sg13g2_decap_8
XFILLER_80_462 VPWR VGND sg13g2_decap_8
XFILLER_53_665 VPWR VGND sg13g2_decap_8
XFILLER_41_805 VPWR VGND sg13g2_decap_8
XFILLER_26_868 VPWR VGND sg13g2_decap_8
XFILLER_52_175 VPWR VGND sg13g2_decap_8
XFILLER_13_518 VPWR VGND sg13g2_decap_8
XFILLER_25_378 VPWR VGND sg13g2_decap_8
XFILLER_40_315 VPWR VGND sg13g2_decap_8
XFILLER_71_39 VPWR VGND sg13g2_decap_8
XFILLER_21_595 VPWR VGND sg13g2_decap_8
XFILLER_5_739 VPWR VGND sg13g2_decap_8
XFILLER_106_133 VPWR VGND sg13g2_decap_8
XFILLER_4_238 VPWR VGND sg13g2_decap_8
XFILLER_20_32 VPWR VGND sg13g2_decap_8
XFILLER_96_14 VPWR VGND sg13g2_decap_8
XFILLER_1_945 VPWR VGND sg13g2_decap_8
XFILLER_103_840 VPWR VGND sg13g2_decap_8
XFILLER_0_455 VPWR VGND sg13g2_decap_8
XFILLER_102_350 VPWR VGND sg13g2_decap_8
XFILLER_49_949 VPWR VGND sg13g2_decap_8
XFILLER_76_746 VPWR VGND sg13g2_decap_8
XFILLER_75_245 VPWR VGND sg13g2_decap_8
XFILLER_48_448 VPWR VGND sg13g2_decap_8
XFILLER_29_74 VPWR VGND sg13g2_decap_8
XFILLER_17_802 VPWR VGND sg13g2_decap_8
XFILLER_21_1022 VPWR VGND sg13g2_decap_8
XFILLER_29_662 VPWR VGND sg13g2_decap_8
XFILLER_91_749 VPWR VGND sg13g2_decap_8
XFILLER_16_301 VPWR VGND sg13g2_decap_8
XFILLER_28_161 VPWR VGND sg13g2_decap_8
XFILLER_72_952 VPWR VGND sg13g2_decap_8
XFILLER_44_676 VPWR VGND sg13g2_decap_8
XFILLER_17_879 VPWR VGND sg13g2_decap_8
XFILLER_32_816 VPWR VGND sg13g2_decap_8
XFILLER_71_473 VPWR VGND sg13g2_decap_8
XFILLER_45_84 VPWR VGND sg13g2_decap_8
XFILLER_43_175 VPWR VGND sg13g2_decap_8
XFILLER_16_378 VPWR VGND sg13g2_decap_8
XFILLER_31_315 VPWR VGND sg13g2_decap_8
XFILLER_8_511 VPWR VGND sg13g2_decap_8
XFILLER_40_882 VPWR VGND sg13g2_decap_8
XFILLER_8_588 VPWR VGND sg13g2_decap_8
XFILLER_6_56 VPWR VGND sg13g2_decap_8
XFILLER_99_805 VPWR VGND sg13g2_decap_8
XFILLER_98_326 VPWR VGND sg13g2_decap_8
XFILLER_67_735 VPWR VGND sg13g2_decap_8
XFILLER_20_4 VPWR VGND sg13g2_decap_8
XFILLER_94_532 VPWR VGND sg13g2_decap_8
XFILLER_66_223 VPWR VGND sg13g2_decap_8
XFILLER_39_459 VPWR VGND sg13g2_decap_8
XFILLER_82_749 VPWR VGND sg13g2_decap_8
XFILLER_19_161 VPWR VGND sg13g2_decap_8
XFILLER_90_760 VPWR VGND sg13g2_decap_8
XFILLER_63_952 VPWR VGND sg13g2_decap_8
XFILLER_23_805 VPWR VGND sg13g2_decap_8
XFILLER_35_665 VPWR VGND sg13g2_decap_8
XFILLER_62_462 VPWR VGND sg13g2_decap_8
XFILLER_50_602 VPWR VGND sg13g2_decap_8
XFILLER_96_0 VPWR VGND sg13g2_decap_8
XFILLER_22_326 VPWR VGND sg13g2_decap_8
XFILLER_34_186 VPWR VGND sg13g2_decap_8
XFILLER_50_679 VPWR VGND sg13g2_decap_8
XFILLER_31_882 VPWR VGND sg13g2_decap_8
XFILLER_30_392 VPWR VGND sg13g2_decap_8
XFILLER_104_637 VPWR VGND sg13g2_decap_8
XFILLER_89_315 VPWR VGND sg13g2_decap_8
XFILLER_106_35 VPWR VGND sg13g2_decap_8
XFILLER_103_147 VPWR VGND sg13g2_decap_8
XFILLER_98_893 VPWR VGND sg13g2_decap_8
XFILLER_58_735 VPWR VGND sg13g2_decap_8
XFILLER_100_854 VPWR VGND sg13g2_decap_8
XFILLER_97_392 VPWR VGND sg13g2_decap_8
XFILLER_85_532 VPWR VGND sg13g2_decap_8
XFILLER_57_245 VPWR VGND sg13g2_decap_8
XFILLER_17_109 VPWR VGND sg13g2_decap_8
XFILLER_66_790 VPWR VGND sg13g2_decap_8
XFILLER_81_760 VPWR VGND sg13g2_decap_8
XFILLER_72_259 VPWR VGND sg13g2_decap_8
XFILLER_54_963 VPWR VGND sg13g2_decap_8
XFILLER_14_805 VPWR VGND sg13g2_decap_8
XFILLER_26_665 VPWR VGND sg13g2_decap_8
XFILLER_82_49 VPWR VGND sg13g2_decap_8
XFILLER_53_462 VPWR VGND sg13g2_decap_8
XFILLER_41_602 VPWR VGND sg13g2_decap_8
XFILLER_13_315 VPWR VGND sg13g2_decap_8
XFILLER_15_32 VPWR VGND sg13g2_decap_8
XFILLER_25_175 VPWR VGND sg13g2_decap_8
XFILLER_40_112 VPWR VGND sg13g2_decap_8
XFILLER_41_679 VPWR VGND sg13g2_decap_8
XFILLER_9_308 VPWR VGND sg13g2_decap_8
XFILLER_51_1026 VPWR VGND sg13g2_fill_2
XFILLER_22_893 VPWR VGND sg13g2_decap_8
XFILLER_40_189 VPWR VGND sg13g2_decap_8
XFILLER_21_392 VPWR VGND sg13g2_decap_8
XFILLER_31_42 VPWR VGND sg13g2_decap_8
XFILLER_5_536 VPWR VGND sg13g2_decap_8
Xoutput20 net20 uo_out[3] VPWR VGND sg13g2_buf_1
XFILLER_96_819 VPWR VGND sg13g2_decap_8
XFILLER_1_742 VPWR VGND sg13g2_decap_8
XFILLER_89_882 VPWR VGND sg13g2_decap_8
XFILLER_0_252 VPWR VGND sg13g2_decap_8
XFILLER_76_543 VPWR VGND sg13g2_decap_8
XFILLER_49_746 VPWR VGND sg13g2_decap_8
XFILLER_48_245 VPWR VGND sg13g2_decap_8
XFILLER_91_546 VPWR VGND sg13g2_decap_8
XFILLER_63_259 VPWR VGND sg13g2_decap_8
XFILLER_60_900 VPWR VGND sg13g2_decap_8
XFILLER_45_952 VPWR VGND sg13g2_decap_8
XFILLER_44_473 VPWR VGND sg13g2_decap_8
XFILLER_16_175 VPWR VGND sg13g2_decap_8
XFILLER_17_676 VPWR VGND sg13g2_decap_8
XFILLER_32_613 VPWR VGND sg13g2_decap_8
XFILLER_71_270 VPWR VGND sg13g2_decap_8
XFILLER_31_112 VPWR VGND sg13g2_decap_8
XFILLER_60_977 VPWR VGND sg13g2_decap_8
XFILLER_13_882 VPWR VGND sg13g2_decap_8
XFILLER_31_189 VPWR VGND sg13g2_decap_8
XFILLER_9_875 VPWR VGND sg13g2_decap_8
XFILLER_68_4 VPWR VGND sg13g2_decap_8
XFILLER_8_385 VPWR VGND sg13g2_decap_8
XFILLER_99_602 VPWR VGND sg13g2_decap_8
XFILLER_67_1022 VPWR VGND sg13g2_decap_8
XFILLER_99_679 VPWR VGND sg13g2_decap_8
XFILLER_98_123 VPWR VGND sg13g2_decap_8
XFILLER_87_819 VPWR VGND sg13g2_decap_8
XFILLER_95_830 VPWR VGND sg13g2_decap_8
XFILLER_67_532 VPWR VGND sg13g2_decap_8
XFILLER_11_0 VPWR VGND sg13g2_decap_8
XFILLER_39_256 VPWR VGND sg13g2_decap_8
XFILLER_55_749 VPWR VGND sg13g2_decap_8
XFILLER_82_546 VPWR VGND sg13g2_decap_8
XFILLER_36_952 VPWR VGND sg13g2_decap_8
XFILLER_51_900 VPWR VGND sg13g2_decap_8
XFILLER_23_602 VPWR VGND sg13g2_decap_8
XFILLER_35_462 VPWR VGND sg13g2_decap_8
XFILLER_22_123 VPWR VGND sg13g2_decap_8
XFILLER_51_977 VPWR VGND sg13g2_decap_8
XFILLER_50_476 VPWR VGND sg13g2_decap_8
XFILLER_11_819 VPWR VGND sg13g2_decap_8
XFILLER_23_679 VPWR VGND sg13g2_decap_8
XFILLER_105_924 VPWR VGND sg13g2_decap_8
XFILLER_89_112 VPWR VGND sg13g2_decap_8
XFILLER_104_434 VPWR VGND sg13g2_decap_8
XFILLER_81_1019 VPWR VGND sg13g2_decap_8
XFILLER_89_189 VPWR VGND sg13g2_decap_8
XFILLER_77_329 VPWR VGND sg13g2_decap_8
XFILLER_77_49 VPWR VGND sg13g2_decap_8
XFILLER_98_690 VPWR VGND sg13g2_decap_8
XFILLER_86_830 VPWR VGND sg13g2_decap_8
XFILLER_58_532 VPWR VGND sg13g2_decap_8
XFILLER_100_651 VPWR VGND sg13g2_decap_8
XFILLER_93_26 VPWR VGND sg13g2_decap_8
XFILLER_73_557 VPWR VGND sg13g2_decap_8
XFILLER_45_259 VPWR VGND sg13g2_decap_8
XFILLER_26_42 VPWR VGND sg13g2_decap_8
XFILLER_27_963 VPWR VGND sg13g2_decap_8
XFILLER_60_207 VPWR VGND sg13g2_decap_8
XFILLER_54_760 VPWR VGND sg13g2_decap_8
XFILLER_42_900 VPWR VGND sg13g2_decap_8
XFILLER_14_602 VPWR VGND sg13g2_decap_8
XFILLER_26_462 VPWR VGND sg13g2_decap_8
XFILLER_13_112 VPWR VGND sg13g2_decap_8
XFILLER_42_977 VPWR VGND sg13g2_decap_8
XFILLER_9_105 VPWR VGND sg13g2_decap_8
XFILLER_14_679 VPWR VGND sg13g2_decap_8
XFILLER_41_476 VPWR VGND sg13g2_decap_8
XFILLER_10_830 VPWR VGND sg13g2_decap_8
XFILLER_13_189 VPWR VGND sg13g2_decap_8
XFILLER_42_74 VPWR VGND sg13g2_decap_8
XFILLER_6_812 VPWR VGND sg13g2_decap_8
XFILLER_22_690 VPWR VGND sg13g2_decap_8
XFILLER_5_333 VPWR VGND sg13g2_decap_8
XFILLER_6_889 VPWR VGND sg13g2_decap_8
XFILLER_96_616 VPWR VGND sg13g2_decap_8
XFILLER_3_35 VPWR VGND sg13g2_decap_8
XFILLER_95_137 VPWR VGND sg13g2_decap_8
XFILLER_76_340 VPWR VGND sg13g2_decap_8
XFILLER_49_543 VPWR VGND sg13g2_decap_8
XFILLER_3_1008 VPWR VGND sg13g2_decap_8
XFILLER_97_1015 VPWR VGND sg13g2_decap_8
XFILLER_92_833 VPWR VGND sg13g2_decap_8
XFILLER_77_896 VPWR VGND sg13g2_decap_8
XFILLER_91_343 VPWR VGND sg13g2_decap_8
XFILLER_64_557 VPWR VGND sg13g2_decap_8
XFILLER_18_952 VPWR VGND sg13g2_decap_8
XFILLER_36_259 VPWR VGND sg13g2_decap_8
XFILLER_51_207 VPWR VGND sg13g2_decap_8
XFILLER_17_473 VPWR VGND sg13g2_decap_8
XFILLER_83_81 VPWR VGND sg13g2_decap_8
XFILLER_44_270 VPWR VGND sg13g2_decap_8
XFILLER_32_410 VPWR VGND sg13g2_decap_8
XFILLER_60_774 VPWR VGND sg13g2_decap_8
XFILLER_33_966 VPWR VGND sg13g2_decap_8
XFILLER_20_627 VPWR VGND sg13g2_decap_8
XFILLER_32_487 VPWR VGND sg13g2_decap_8
XFILLER_9_672 VPWR VGND sg13g2_decap_8
XFILLER_8_182 VPWR VGND sg13g2_decap_8
XFILLER_102_938 VPWR VGND sg13g2_decap_8
XFILLER_99_476 VPWR VGND sg13g2_decap_8
XFILLER_87_616 VPWR VGND sg13g2_decap_8
XFILLER_101_448 VPWR VGND sg13g2_decap_8
XFILLER_86_137 VPWR VGND sg13g2_decap_8
XFILLER_68_852 VPWR VGND sg13g2_decap_8
XFILLER_103_14 VPWR VGND sg13g2_decap_8
XFILLER_83_844 VPWR VGND sg13g2_decap_8
XFILLER_28_749 VPWR VGND sg13g2_decap_8
XFILLER_82_343 VPWR VGND sg13g2_decap_8
XFILLER_55_546 VPWR VGND sg13g2_decap_8
XFILLER_42_207 VPWR VGND sg13g2_decap_8
XFILLER_24_900 VPWR VGND sg13g2_decap_8
XFILLER_51_774 VPWR VGND sg13g2_decap_8
XFILLER_24_977 VPWR VGND sg13g2_decap_8
XFILLER_50_273 VPWR VGND sg13g2_decap_8
XFILLER_11_616 VPWR VGND sg13g2_decap_8
XFILLER_23_476 VPWR VGND sg13g2_decap_8
XFILLER_10_137 VPWR VGND sg13g2_decap_8
XFILLER_12_11 VPWR VGND sg13g2_decap_8
XFILLER_6_119 VPWR VGND sg13g2_decap_8
XFILLER_12_88 VPWR VGND sg13g2_decap_8
XFILLER_105_721 VPWR VGND sg13g2_decap_8
XFILLER_3_826 VPWR VGND sg13g2_decap_8
XFILLER_104_231 VPWR VGND sg13g2_decap_8
XFILLER_2_347 VPWR VGND sg13g2_decap_8
XFILLER_105_798 VPWR VGND sg13g2_decap_8
XFILLER_77_126 VPWR VGND sg13g2_decap_8
XFILLER_59_852 VPWR VGND sg13g2_decap_8
XFILLER_19_749 VPWR VGND sg13g2_decap_8
XFILLER_74_855 VPWR VGND sg13g2_decap_8
XFILLER_46_557 VPWR VGND sg13g2_decap_8
XFILLER_18_259 VPWR VGND sg13g2_decap_8
XFILLER_37_74 VPWR VGND sg13g2_decap_8
XFILLER_73_354 VPWR VGND sg13g2_decap_8
XFILLER_15_900 VPWR VGND sg13g2_decap_8
XFILLER_27_760 VPWR VGND sg13g2_decap_8
XFILLER_42_774 VPWR VGND sg13g2_decap_8
XFILLER_15_977 VPWR VGND sg13g2_decap_8
XFILLER_30_903 VPWR VGND sg13g2_decap_8
XFILLER_105_1008 VPWR VGND sg13g2_decap_8
XFILLER_53_84 VPWR VGND sg13g2_decap_8
XFILLER_14_476 VPWR VGND sg13g2_decap_8
XFILLER_41_273 VPWR VGND sg13g2_decap_8
XFILLER_5_130 VPWR VGND sg13g2_decap_8
XFILLER_52_7 VPWR VGND sg13g2_decap_8
XFILLER_6_686 VPWR VGND sg13g2_decap_8
XFILLER_97_903 VPWR VGND sg13g2_decap_8
XFILLER_96_413 VPWR VGND sg13g2_decap_8
XFILLER_69_638 VPWR VGND sg13g2_decap_8
XFILLER_68_159 VPWR VGND sg13g2_decap_8
XFILLER_49_340 VPWR VGND sg13g2_decap_8
XFILLER_77_693 VPWR VGND sg13g2_decap_8
XFILLER_65_833 VPWR VGND sg13g2_decap_8
XFILLER_92_630 VPWR VGND sg13g2_decap_8
X_65_ net9 net1 net17 VPWR VGND sg13g2_xor2_1
XFILLER_37_557 VPWR VGND sg13g2_decap_8
XFILLER_94_91 VPWR VGND sg13g2_decap_8
XFILLER_91_140 VPWR VGND sg13g2_decap_8
XFILLER_64_354 VPWR VGND sg13g2_decap_8
XFILLER_24_207 VPWR VGND sg13g2_decap_8
XFILLER_80_847 VPWR VGND sg13g2_decap_8
XFILLER_17_270 VPWR VGND sg13g2_decap_8
XFILLER_21_903 VPWR VGND sg13g2_decap_8
XFILLER_33_763 VPWR VGND sg13g2_decap_8
XFILLER_60_571 VPWR VGND sg13g2_decap_8
XFILLER_20_424 VPWR VGND sg13g2_decap_8
XFILLER_32_284 VPWR VGND sg13g2_decap_8
XFILLER_106_518 VPWR VGND sg13g2_decap_8
XFILLER_88_914 VPWR VGND sg13g2_decap_8
XFILLER_102_735 VPWR VGND sg13g2_decap_8
XFILLER_99_273 VPWR VGND sg13g2_decap_8
XFILLER_87_413 VPWR VGND sg13g2_decap_8
XFILLER_101_245 VPWR VGND sg13g2_decap_8
XFILLER_59_159 VPWR VGND sg13g2_decap_8
XFILLER_96_980 VPWR VGND sg13g2_decap_8
XFILLER_83_641 VPWR VGND sg13g2_decap_8
XFILLER_74_28 VPWR VGND sg13g2_decap_8
XFILLER_56_844 VPWR VGND sg13g2_decap_8
XFILLER_55_343 VPWR VGND sg13g2_decap_8
XFILLER_28_546 VPWR VGND sg13g2_decap_8
XFILLER_82_140 VPWR VGND sg13g2_decap_8
XFILLER_15_207 VPWR VGND sg13g2_decap_8
XFILLER_71_858 VPWR VGND sg13g2_decap_8
XFILLER_70_357 VPWR VGND sg13g2_decap_8
XFILLER_12_914 VPWR VGND sg13g2_decap_8
XFILLER_51_571 VPWR VGND sg13g2_decap_8
XFILLER_11_413 VPWR VGND sg13g2_decap_8
XFILLER_23_21 VPWR VGND sg13g2_decap_8
XFILLER_23_273 VPWR VGND sg13g2_decap_8
XFILLER_24_774 VPWR VGND sg13g2_decap_8
XFILLER_7_417 VPWR VGND sg13g2_decap_8
XFILLER_99_14 VPWR VGND sg13g2_decap_8
XFILLER_20_991 VPWR VGND sg13g2_decap_8
XFILLER_23_98 VPWR VGND sg13g2_decap_8
XFILLER_3_623 VPWR VGND sg13g2_decap_8
XFILLER_79_914 VPWR VGND sg13g2_decap_8
XFILLER_2_144 VPWR VGND sg13g2_decap_8
XFILLER_105_595 VPWR VGND sg13g2_decap_8
XFILLER_94_917 VPWR VGND sg13g2_decap_8
XFILLER_78_468 VPWR VGND sg13g2_decap_8
XFILLER_66_608 VPWR VGND sg13g2_decap_8
XFILLER_87_980 VPWR VGND sg13g2_decap_8
XFILLER_47_833 VPWR VGND sg13g2_decap_8
XFILLER_48_84 VPWR VGND sg13g2_decap_8
XFILLER_74_652 VPWR VGND sg13g2_decap_8
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_19_546 VPWR VGND sg13g2_decap_8
XFILLER_73_151 VPWR VGND sg13g2_decap_8
XFILLER_46_354 VPWR VGND sg13g2_decap_8
XFILLER_62_847 VPWR VGND sg13g2_decap_8
XFILLER_61_368 VPWR VGND sg13g2_decap_8
XFILLER_42_571 VPWR VGND sg13g2_decap_8
XFILLER_14_273 VPWR VGND sg13g2_decap_8
XFILLER_15_774 VPWR VGND sg13g2_decap_8
XFILLER_30_700 VPWR VGND sg13g2_decap_8
XFILLER_9_56 VPWR VGND sg13g2_decap_8
XFILLER_30_777 VPWR VGND sg13g2_decap_8
XFILLER_11_980 VPWR VGND sg13g2_decap_8
XFILLER_7_984 VPWR VGND sg13g2_decap_8
XFILLER_6_483 VPWR VGND sg13g2_decap_8
XFILLER_97_700 VPWR VGND sg13g2_decap_8
XFILLER_89_91 VPWR VGND sg13g2_decap_8
XFILLER_96_210 VPWR VGND sg13g2_decap_8
XFILLER_69_435 VPWR VGND sg13g2_decap_8
XFILLER_97_777 VPWR VGND sg13g2_decap_8
XFILLER_85_917 VPWR VGND sg13g2_decap_8
XFILLER_96_287 VPWR VGND sg13g2_decap_8
XFILLER_84_427 VPWR VGND sg13g2_decap_8
XFILLER_93_950 VPWR VGND sg13g2_decap_8
XFILLER_77_490 VPWR VGND sg13g2_decap_8
XFILLER_65_630 VPWR VGND sg13g2_decap_8
XFILLER_38_833 VPWR VGND sg13g2_decap_8
X_48_ VPWR _16_ _15_ VGND sg13g2_inv_1
XFILLER_64_151 VPWR VGND sg13g2_decap_8
XFILLER_37_354 VPWR VGND sg13g2_decap_8
XFILLER_80_644 VPWR VGND sg13g2_decap_8
XFILLER_53_847 VPWR VGND sg13g2_decap_8
XFILLER_52_357 VPWR VGND sg13g2_decap_8
XFILLER_21_700 VPWR VGND sg13g2_decap_8
XFILLER_33_560 VPWR VGND sg13g2_decap_8
XFILLER_20_221 VPWR VGND sg13g2_decap_8
XFILLER_21_777 VPWR VGND sg13g2_decap_8
XFILLER_20_298 VPWR VGND sg13g2_decap_8
XFILLER_106_315 VPWR VGND sg13g2_decap_8
XFILLER_69_28 VPWR VGND sg13g2_decap_8
XFILLER_88_711 VPWR VGND sg13g2_decap_8
XFILLER_87_210 VPWR VGND sg13g2_decap_8
XFILLER_0_637 VPWR VGND sg13g2_decap_8
XFILLER_102_532 VPWR VGND sg13g2_decap_8
XFILLER_88_788 VPWR VGND sg13g2_decap_8
XFILLER_87_287 VPWR VGND sg13g2_decap_8
XFILLER_85_49 VPWR VGND sg13g2_decap_8
XFILLER_76_928 VPWR VGND sg13g2_decap_8
XFILLER_75_427 VPWR VGND sg13g2_decap_8
XFILLER_56_641 VPWR VGND sg13g2_decap_8
XFILLER_18_21 VPWR VGND sg13g2_decap_8
XFILLER_29_844 VPWR VGND sg13g2_decap_8
XFILLER_55_140 VPWR VGND sg13g2_decap_8
XFILLER_28_343 VPWR VGND sg13g2_decap_8
XFILLER_84_994 VPWR VGND sg13g2_decap_8
XFILLER_44_858 VPWR VGND sg13g2_decap_8
XFILLER_18_98 VPWR VGND sg13g2_decap_8
XFILLER_71_655 VPWR VGND sg13g2_decap_8
XFILLER_70_154 VPWR VGND sg13g2_decap_8
XFILLER_43_357 VPWR VGND sg13g2_decap_8
XFILLER_12_711 VPWR VGND sg13g2_decap_8
XFILLER_24_571 VPWR VGND sg13g2_decap_8
XFILLER_34_53 VPWR VGND sg13g2_decap_8
XFILLER_11_210 VPWR VGND sg13g2_decap_8
XFILLER_15_1019 VPWR VGND sg13g2_decap_8
XFILLER_7_214 VPWR VGND sg13g2_decap_8
XFILLER_12_788 VPWR VGND sg13g2_decap_8
XFILLER_11_287 VPWR VGND sg13g2_decap_8
XFILLER_50_63 VPWR VGND sg13g2_decap_8
XFILLER_4_910 VPWR VGND sg13g2_decap_8
XFILLER_3_420 VPWR VGND sg13g2_decap_8
XFILLER_98_508 VPWR VGND sg13g2_decap_8
XFILLER_4_987 VPWR VGND sg13g2_decap_8
XFILLER_106_882 VPWR VGND sg13g2_decap_8
XFILLER_79_711 VPWR VGND sg13g2_decap_8
XFILLER_3_497 VPWR VGND sg13g2_decap_8
XFILLER_105_392 VPWR VGND sg13g2_decap_8
XFILLER_67_917 VPWR VGND sg13g2_decap_8
XFILLER_61_1028 VPWR VGND sg13g2_fill_1
XFILLER_94_714 VPWR VGND sg13g2_decap_8
XFILLER_79_788 VPWR VGND sg13g2_decap_8
XFILLER_78_265 VPWR VGND sg13g2_decap_8
XFILLER_66_405 VPWR VGND sg13g2_decap_8
XFILLER_47_630 VPWR VGND sg13g2_decap_8
XFILLER_93_257 VPWR VGND sg13g2_decap_8
XFILLER_46_151 VPWR VGND sg13g2_decap_8
XFILLER_19_343 VPWR VGND sg13g2_decap_8
XFILLER_90_942 VPWR VGND sg13g2_decap_8
XFILLER_75_994 VPWR VGND sg13g2_decap_8
XFILLER_35_847 VPWR VGND sg13g2_decap_8
XFILLER_62_644 VPWR VGND sg13g2_decap_8
XFILLER_22_508 VPWR VGND sg13g2_decap_8
XFILLER_34_368 VPWR VGND sg13g2_decap_8
XFILLER_61_165 VPWR VGND sg13g2_decap_8
XFILLER_15_571 VPWR VGND sg13g2_decap_8
XFILLER_98_4 VPWR VGND sg13g2_decap_8
XFILLER_91_70 VPWR VGND sg13g2_decap_8
XFILLER_30_574 VPWR VGND sg13g2_decap_8
XFILLER_7_781 VPWR VGND sg13g2_decap_8
XFILLER_6_280 VPWR VGND sg13g2_decap_8
XFILLER_104_819 VPWR VGND sg13g2_decap_8
XFILLER_103_329 VPWR VGND sg13g2_decap_8
XFILLER_41_0 VPWR VGND sg13g2_decap_8
XFILLER_69_232 VPWR VGND sg13g2_decap_8
XFILLER_58_917 VPWR VGND sg13g2_decap_8
XFILLER_97_574 VPWR VGND sg13g2_decap_8
XFILLER_85_714 VPWR VGND sg13g2_decap_8
XFILLER_57_427 VPWR VGND sg13g2_decap_8
XFILLER_84_224 VPWR VGND sg13g2_decap_8
XFILLER_38_630 VPWR VGND sg13g2_decap_8
XFILLER_66_972 VPWR VGND sg13g2_decap_8
XFILLER_37_151 VPWR VGND sg13g2_decap_8
XFILLER_81_942 VPWR VGND sg13g2_decap_8
XFILLER_26_847 VPWR VGND sg13g2_decap_8
XFILLER_80_441 VPWR VGND sg13g2_decap_8
XFILLER_53_644 VPWR VGND sg13g2_decap_8
XFILLER_25_357 VPWR VGND sg13g2_decap_8
XFILLER_38_1008 VPWR VGND sg13g2_decap_8
XFILLER_71_18 VPWR VGND sg13g2_decap_8
XFILLER_52_154 VPWR VGND sg13g2_decap_8
XFILLER_21_574 VPWR VGND sg13g2_decap_8
XFILLER_101_1022 VPWR VGND sg13g2_decap_8
XFILLER_5_718 VPWR VGND sg13g2_decap_8
XFILLER_106_112 VPWR VGND sg13g2_decap_8
XFILLER_4_217 VPWR VGND sg13g2_decap_8
XFILLER_20_11 VPWR VGND sg13g2_decap_8
XFILLER_106_189 VPWR VGND sg13g2_decap_8
XFILLER_1_924 VPWR VGND sg13g2_decap_8
XFILLER_20_88 VPWR VGND sg13g2_decap_8
XFILLER_0_434 VPWR VGND sg13g2_decap_8
XFILLER_103_896 VPWR VGND sg13g2_decap_8
XFILLER_88_585 VPWR VGND sg13g2_decap_8
XFILLER_76_725 VPWR VGND sg13g2_decap_8
XFILLER_49_928 VPWR VGND sg13g2_decap_8
XFILLER_48_427 VPWR VGND sg13g2_decap_8
XFILLER_29_53 VPWR VGND sg13g2_decap_8
XFILLER_75_224 VPWR VGND sg13g2_decap_8
XFILLER_21_1001 VPWR VGND sg13g2_decap_8
XFILLER_91_728 VPWR VGND sg13g2_decap_8
XFILLER_28_140 VPWR VGND sg13g2_decap_8
XFILLER_29_641 VPWR VGND sg13g2_decap_8
XFILLER_84_791 VPWR VGND sg13g2_decap_8
XFILLER_72_931 VPWR VGND sg13g2_decap_8
XFILLER_57_994 VPWR VGND sg13g2_decap_8
XFILLER_90_249 VPWR VGND sg13g2_decap_8
XFILLER_71_452 VPWR VGND sg13g2_decap_8
XFILLER_45_63 VPWR VGND sg13g2_decap_8
XFILLER_44_655 VPWR VGND sg13g2_decap_8
XFILLER_16_357 VPWR VGND sg13g2_decap_8
XFILLER_17_858 VPWR VGND sg13g2_decap_8
XFILLER_43_154 VPWR VGND sg13g2_decap_8
XFILLER_101_91 VPWR VGND sg13g2_decap_8
XFILLER_40_861 VPWR VGND sg13g2_decap_8
XFILLER_61_95 VPWR VGND sg13g2_decap_8
XFILLER_12_585 VPWR VGND sg13g2_decap_8
XFILLER_8_567 VPWR VGND sg13g2_decap_8
XFILLER_6_35 VPWR VGND sg13g2_decap_8
XFILLER_98_305 VPWR VGND sg13g2_decap_8
XFILLER_4_784 VPWR VGND sg13g2_decap_8
XFILLER_3_294 VPWR VGND sg13g2_decap_8
XFILLER_94_511 VPWR VGND sg13g2_decap_8
XFILLER_79_585 VPWR VGND sg13g2_decap_8
XFILLER_67_714 VPWR VGND sg13g2_decap_8
XFILLER_66_202 VPWR VGND sg13g2_decap_8
XFILLER_86_81 VPWR VGND sg13g2_decap_8
XFILLER_39_438 VPWR VGND sg13g2_decap_8
XFILLER_94_588 VPWR VGND sg13g2_decap_8
XFILLER_82_728 VPWR VGND sg13g2_decap_8
XFILLER_66_279 VPWR VGND sg13g2_decap_8
XFILLER_19_140 VPWR VGND sg13g2_decap_8
XFILLER_75_791 VPWR VGND sg13g2_decap_8
XFILLER_63_931 VPWR VGND sg13g2_decap_8
XFILLER_48_994 VPWR VGND sg13g2_decap_8
XFILLER_81_249 VPWR VGND sg13g2_decap_8
XFILLER_62_441 VPWR VGND sg13g2_decap_8
XFILLER_35_644 VPWR VGND sg13g2_decap_8
XFILLER_22_305 VPWR VGND sg13g2_decap_8
XFILLER_34_165 VPWR VGND sg13g2_decap_8
XFILLER_50_658 VPWR VGND sg13g2_decap_8
XFILLER_89_0 VPWR VGND sg13g2_decap_8
XFILLER_31_861 VPWR VGND sg13g2_decap_8
XFILLER_30_371 VPWR VGND sg13g2_decap_8
XFILLER_104_616 VPWR VGND sg13g2_decap_8
XFILLER_106_14 VPWR VGND sg13g2_decap_8
XFILLER_103_126 VPWR VGND sg13g2_decap_8
XFILLER_44_1012 VPWR VGND sg13g2_decap_8
XFILLER_98_872 VPWR VGND sg13g2_decap_8
XFILLER_97_371 VPWR VGND sg13g2_decap_8
XFILLER_85_511 VPWR VGND sg13g2_decap_8
XFILLER_66_18 VPWR VGND sg13g2_fill_1
XFILLER_58_714 VPWR VGND sg13g2_decap_8
XFILLER_100_833 VPWR VGND sg13g2_decap_8
XFILLER_57_224 VPWR VGND sg13g2_decap_8
XFILLER_85_588 VPWR VGND sg13g2_decap_8
XFILLER_73_739 VPWR VGND sg13g2_decap_8
XFILLER_82_28 VPWR VGND sg13g2_decap_8
XFILLER_72_238 VPWR VGND sg13g2_decap_8
XFILLER_54_942 VPWR VGND sg13g2_decap_8
XFILLER_53_441 VPWR VGND sg13g2_decap_8
XFILLER_26_644 VPWR VGND sg13g2_decap_8
XFILLER_15_11 VPWR VGND sg13g2_decap_8
XFILLER_25_154 VPWR VGND sg13g2_decap_8
XFILLER_41_658 VPWR VGND sg13g2_decap_8
XFILLER_51_1005 VPWR VGND sg13g2_decap_8
XFILLER_15_88 VPWR VGND sg13g2_decap_8
XFILLER_22_872 VPWR VGND sg13g2_decap_8
XFILLER_40_168 VPWR VGND sg13g2_decap_8
XFILLER_21_371 VPWR VGND sg13g2_decap_8
XFILLER_31_21 VPWR VGND sg13g2_decap_8
XFILLER_5_515 VPWR VGND sg13g2_decap_8
XFILLER_31_98 VPWR VGND sg13g2_decap_8
Xoutput21 net21 uo_out[4] VPWR VGND sg13g2_buf_1
XFILLER_1_721 VPWR VGND sg13g2_decap_8
XFILLER_95_319 VPWR VGND sg13g2_decap_8
XFILLER_89_861 VPWR VGND sg13g2_decap_8
XFILLER_49_725 VPWR VGND sg13g2_decap_8
XFILLER_0_231 VPWR VGND sg13g2_decap_8
XFILLER_103_693 VPWR VGND sg13g2_decap_8
XFILLER_88_382 VPWR VGND sg13g2_decap_8
XFILLER_76_522 VPWR VGND sg13g2_decap_8
XFILLER_48_224 VPWR VGND sg13g2_decap_8
XFILLER_1_798 VPWR VGND sg13g2_decap_8
XFILLER_91_525 VPWR VGND sg13g2_decap_8
XFILLER_76_599 VPWR VGND sg13g2_decap_8
XFILLER_64_739 VPWR VGND sg13g2_decap_8
XFILLER_57_791 VPWR VGND sg13g2_decap_8
XFILLER_45_931 VPWR VGND sg13g2_decap_8
XFILLER_63_238 VPWR VGND sg13g2_decap_8
XFILLER_56_95 VPWR VGND sg13g2_decap_8
XFILLER_17_655 VPWR VGND sg13g2_decap_8
XFILLER_44_452 VPWR VGND sg13g2_decap_8
XFILLER_16_154 VPWR VGND sg13g2_decap_8
XFILLER_60_956 VPWR VGND sg13g2_decap_8
XFILLER_13_861 VPWR VGND sg13g2_decap_8
XFILLER_20_809 VPWR VGND sg13g2_decap_8
XFILLER_31_168 VPWR VGND sg13g2_decap_8
XFILLER_32_669 VPWR VGND sg13g2_decap_8
XFILLER_82_7 VPWR VGND sg13g2_decap_8
XFILLER_9_854 VPWR VGND sg13g2_decap_8
XFILLER_12_382 VPWR VGND sg13g2_decap_8
XFILLER_8_364 VPWR VGND sg13g2_decap_8
XFILLER_67_1001 VPWR VGND sg13g2_decap_8
XFILLER_98_102 VPWR VGND sg13g2_decap_8
XFILLER_99_658 VPWR VGND sg13g2_decap_8
XFILLER_4_581 VPWR VGND sg13g2_decap_8
XFILLER_98_179 VPWR VGND sg13g2_decap_8
XFILLER_97_91 VPWR VGND sg13g2_decap_8
XFILLER_86_319 VPWR VGND sg13g2_decap_8
XFILLER_79_382 VPWR VGND sg13g2_decap_8
XFILLER_67_511 VPWR VGND sg13g2_decap_8
XFILLER_95_886 VPWR VGND sg13g2_decap_8
XFILLER_39_235 VPWR VGND sg13g2_decap_8
XFILLER_94_385 VPWR VGND sg13g2_decap_8
XFILLER_82_525 VPWR VGND sg13g2_decap_8
XFILLER_67_588 VPWR VGND sg13g2_decap_8
XFILLER_55_728 VPWR VGND sg13g2_decap_8
XFILLER_48_791 VPWR VGND sg13g2_decap_8
XFILLER_36_931 VPWR VGND sg13g2_decap_8
XFILLER_54_249 VPWR VGND sg13g2_decap_8
XFILLER_35_441 VPWR VGND sg13g2_decap_8
XFILLER_74_1016 VPWR VGND sg13g2_decap_8
XFILLER_74_1027 VPWR VGND sg13g2_fill_2
XFILLER_51_956 VPWR VGND sg13g2_decap_8
XFILLER_22_102 VPWR VGND sg13g2_decap_8
XFILLER_50_455 VPWR VGND sg13g2_decap_8
XFILLER_23_658 VPWR VGND sg13g2_decap_8
XFILLER_10_319 VPWR VGND sg13g2_decap_8
XFILLER_22_179 VPWR VGND sg13g2_decap_8
XFILLER_11_1022 VPWR VGND sg13g2_decap_8
XFILLER_105_903 VPWR VGND sg13g2_decap_8
XFILLER_104_413 VPWR VGND sg13g2_decap_8
XFILLER_2_529 VPWR VGND sg13g2_decap_8
XFILLER_77_28 VPWR VGND sg13g2_decap_8
XFILLER_89_168 VPWR VGND sg13g2_decap_8
XFILLER_77_308 VPWR VGND sg13g2_decap_8
XFILLER_58_511 VPWR VGND sg13g2_decap_8
XFILLER_100_630 VPWR VGND sg13g2_decap_8
XFILLER_86_886 VPWR VGND sg13g2_decap_8
XFILLER_85_385 VPWR VGND sg13g2_decap_8
XFILLER_73_536 VPWR VGND sg13g2_decap_8
XFILLER_58_588 VPWR VGND sg13g2_decap_8
XFILLER_46_739 VPWR VGND sg13g2_decap_8
XFILLER_45_238 VPWR VGND sg13g2_decap_8
XFILLER_26_21 VPWR VGND sg13g2_decap_8
XFILLER_27_942 VPWR VGND sg13g2_decap_8
XFILLER_26_441 VPWR VGND sg13g2_decap_8
XFILLER_42_956 VPWR VGND sg13g2_decap_8
XFILLER_26_98 VPWR VGND sg13g2_decap_8
XFILLER_14_658 VPWR VGND sg13g2_decap_8
XFILLER_41_455 VPWR VGND sg13g2_decap_8
XFILLER_42_53 VPWR VGND sg13g2_decap_8
XFILLER_13_168 VPWR VGND sg13g2_decap_8
XFILLER_5_312 VPWR VGND sg13g2_decap_8
XFILLER_10_886 VPWR VGND sg13g2_decap_8
XFILLER_6_868 VPWR VGND sg13g2_decap_8
XFILLER_5_389 VPWR VGND sg13g2_decap_8
XFILLER_3_14 VPWR VGND sg13g2_decap_8
XFILLER_104_980 VPWR VGND sg13g2_decap_8
XFILLER_95_116 VPWR VGND sg13g2_decap_8
XFILLER_49_522 VPWR VGND sg13g2_decap_8
XFILLER_1_595 VPWR VGND sg13g2_decap_8
XFILLER_103_490 VPWR VGND sg13g2_decap_8
XFILLER_77_875 VPWR VGND sg13g2_decap_8
XFILLER_92_812 VPWR VGND sg13g2_decap_8
XFILLER_49_599 VPWR VGND sg13g2_decap_8
XFILLER_37_739 VPWR VGND sg13g2_decap_8
XFILLER_91_322 VPWR VGND sg13g2_decap_8
XFILLER_76_396 VPWR VGND sg13g2_decap_8
XFILLER_64_536 VPWR VGND sg13g2_decap_8
XFILLER_18_931 VPWR VGND sg13g2_decap_8
XFILLER_36_238 VPWR VGND sg13g2_decap_8
XFILLER_92_889 VPWR VGND sg13g2_decap_8
XFILLER_83_60 VPWR VGND sg13g2_decap_8
XFILLER_17_452 VPWR VGND sg13g2_decap_8
XFILLER_91_399 VPWR VGND sg13g2_decap_8
XFILLER_33_945 VPWR VGND sg13g2_decap_8
XFILLER_60_753 VPWR VGND sg13g2_decap_8
XFILLER_20_606 VPWR VGND sg13g2_decap_8
XFILLER_32_466 VPWR VGND sg13g2_decap_8
XFILLER_9_651 VPWR VGND sg13g2_decap_8
XFILLER_8_161 VPWR VGND sg13g2_decap_8
XFILLER_102_917 VPWR VGND sg13g2_decap_8
XFILLER_99_455 VPWR VGND sg13g2_decap_8
XFILLER_101_427 VPWR VGND sg13g2_decap_8
XFILLER_86_116 VPWR VGND sg13g2_decap_8
XFILLER_68_831 VPWR VGND sg13g2_decap_8
XFILLER_41_1015 VPWR VGND sg13g2_decap_8
XFILLER_95_683 VPWR VGND sg13g2_decap_8
XFILLER_83_823 VPWR VGND sg13g2_decap_8
XFILLER_67_385 VPWR VGND sg13g2_decap_8
XFILLER_55_525 VPWR VGND sg13g2_decap_8
XFILLER_28_728 VPWR VGND sg13g2_decap_8
XFILLER_94_182 VPWR VGND sg13g2_decap_8
XFILLER_82_322 VPWR VGND sg13g2_decap_8
XFILLER_27_249 VPWR VGND sg13g2_decap_8
XFILLER_82_399 VPWR VGND sg13g2_decap_8
XFILLER_70_539 VPWR VGND sg13g2_decap_8
XFILLER_24_956 VPWR VGND sg13g2_decap_8
XFILLER_51_753 VPWR VGND sg13g2_decap_8
XFILLER_23_455 VPWR VGND sg13g2_decap_8
XFILLER_50_252 VPWR VGND sg13g2_decap_8
XFILLER_10_116 VPWR VGND sg13g2_decap_8
XFILLER_12_67 VPWR VGND sg13g2_decap_8
XFILLER_105_700 VPWR VGND sg13g2_decap_8
XFILLER_3_805 VPWR VGND sg13g2_decap_8
XFILLER_104_210 VPWR VGND sg13g2_decap_8
XFILLER_2_326 VPWR VGND sg13g2_decap_8
XFILLER_105_777 VPWR VGND sg13g2_decap_8
XFILLER_104_287 VPWR VGND sg13g2_decap_8
XFILLER_77_105 VPWR VGND sg13g2_decap_8
XFILLER_59_831 VPWR VGND sg13g2_decap_8
XFILLER_101_994 VPWR VGND sg13g2_decap_8
XFILLER_92_119 VPWR VGND sg13g2_decap_8
XFILLER_86_683 VPWR VGND sg13g2_decap_8
XFILLER_74_834 VPWR VGND sg13g2_decap_8
XFILLER_58_385 VPWR VGND sg13g2_decap_8
XFILLER_19_728 VPWR VGND sg13g2_decap_8
XFILLER_85_182 VPWR VGND sg13g2_decap_8
XFILLER_73_333 VPWR VGND sg13g2_decap_8
XFILLER_46_536 VPWR VGND sg13g2_decap_8
XFILLER_18_238 VPWR VGND sg13g2_decap_8
XFILLER_37_53 VPWR VGND sg13g2_decap_8
XFILLER_57_1022 VPWR VGND sg13g2_decap_8
XFILLER_53_63 VPWR VGND sg13g2_decap_8
XFILLER_42_753 VPWR VGND sg13g2_decap_8
XFILLER_14_455 VPWR VGND sg13g2_decap_8
XFILLER_15_956 VPWR VGND sg13g2_decap_8
XFILLER_41_252 VPWR VGND sg13g2_decap_8
XFILLER_30_959 VPWR VGND sg13g2_decap_8
XFILLER_10_683 VPWR VGND sg13g2_decap_8
XFILLER_6_665 VPWR VGND sg13g2_decap_8
XFILLER_45_7 VPWR VGND sg13g2_decap_8
XFILLER_5_186 VPWR VGND sg13g2_decap_8
XFILLER_78_60 VPWR VGND sg13g2_fill_1
XFILLER_69_617 VPWR VGND sg13g2_decap_8
XFILLER_64_1026 VPWR VGND sg13g2_fill_2
XFILLER_97_959 VPWR VGND sg13g2_decap_8
XFILLER_2_893 VPWR VGND sg13g2_decap_8
XFILLER_96_469 VPWR VGND sg13g2_decap_8
XFILLER_84_609 VPWR VGND sg13g2_decap_8
XFILLER_68_138 VPWR VGND sg13g2_decap_8
XFILLER_1_392 VPWR VGND sg13g2_decap_8
X_64_ net24 _27_ _28_ VPWR VGND sg13g2_xnor2_1
XFILLER_77_672 VPWR VGND sg13g2_decap_8
XFILLER_65_812 VPWR VGND sg13g2_decap_8
XFILLER_94_70 VPWR VGND sg13g2_decap_8
XFILLER_76_193 VPWR VGND sg13g2_decap_8
XFILLER_64_333 VPWR VGND sg13g2_decap_8
XFILLER_49_396 VPWR VGND sg13g2_decap_8
XFILLER_37_536 VPWR VGND sg13g2_decap_8
XFILLER_92_686 VPWR VGND sg13g2_decap_8
XFILLER_80_826 VPWR VGND sg13g2_decap_8
XFILLER_65_889 VPWR VGND sg13g2_decap_8
XFILLER_91_196 VPWR VGND sg13g2_decap_8
XFILLER_52_539 VPWR VGND sg13g2_decap_8
XFILLER_60_550 VPWR VGND sg13g2_decap_8
XFILLER_33_742 VPWR VGND sg13g2_decap_8
XFILLER_71_1019 VPWR VGND sg13g2_decap_8
XFILLER_20_403 VPWR VGND sg13g2_decap_8
XFILLER_32_263 VPWR VGND sg13g2_decap_8
XFILLER_21_959 VPWR VGND sg13g2_decap_8
XFILLER_99_252 VPWR VGND sg13g2_decap_8
XFILLER_0_819 VPWR VGND sg13g2_decap_8
XFILLER_102_714 VPWR VGND sg13g2_decap_8
XFILLER_59_127 VPWR VGND sg13g2_decap_8
XFILLER_101_224 VPWR VGND sg13g2_decap_8
XFILLER_87_469 VPWR VGND sg13g2_decap_8
XFILLER_75_609 VPWR VGND sg13g2_decap_8
XFILLER_59_138 VPWR VGND sg13g2_fill_2
XFILLER_56_823 VPWR VGND sg13g2_decap_8
XFILLER_95_480 VPWR VGND sg13g2_decap_8
XFILLER_83_620 VPWR VGND sg13g2_decap_8
XFILLER_67_182 VPWR VGND sg13g2_decap_8
XFILLER_55_322 VPWR VGND sg13g2_decap_8
XFILLER_28_525 VPWR VGND sg13g2_decap_8
XFILLER_83_697 VPWR VGND sg13g2_decap_8
XFILLER_82_196 VPWR VGND sg13g2_decap_8
XFILLER_71_837 VPWR VGND sg13g2_decap_8
XFILLER_70_336 VPWR VGND sg13g2_decap_8
XFILLER_55_399 VPWR VGND sg13g2_decap_8
XFILLER_43_539 VPWR VGND sg13g2_decap_8
XFILLER_51_550 VPWR VGND sg13g2_decap_8
XFILLER_24_753 VPWR VGND sg13g2_decap_8
XFILLER_90_39 VPWR VGND sg13g2_decap_8
XFILLER_23_252 VPWR VGND sg13g2_decap_8
XFILLER_11_469 VPWR VGND sg13g2_decap_8
XFILLER_20_970 VPWR VGND sg13g2_decap_8
XFILLER_23_77 VPWR VGND sg13g2_decap_8
XFILLER_87_1015 VPWR VGND sg13g2_decap_8
XFILLER_3_602 VPWR VGND sg13g2_decap_8
XFILLER_3_679 VPWR VGND sg13g2_decap_8
XFILLER_2_123 VPWR VGND sg13g2_decap_8
XFILLER_105_574 VPWR VGND sg13g2_decap_8
XFILLER_78_447 VPWR VGND sg13g2_decap_8
XFILLER_65_119 VPWR VGND sg13g2_decap_8
XFILLER_47_812 VPWR VGND sg13g2_decap_8
XFILLER_48_63 VPWR VGND sg13g2_decap_8
XFILLER_101_791 VPWR VGND sg13g2_decap_8
XFILLER_93_439 VPWR VGND sg13g2_decap_8
XFILLER_86_480 VPWR VGND sg13g2_decap_8
XFILLER_74_631 VPWR VGND sg13g2_decap_8
XFILLER_58_182 VPWR VGND sg13g2_decap_8
XFILLER_46_333 VPWR VGND sg13g2_decap_8
XFILLER_19_525 VPWR VGND sg13g2_decap_8
XFILLER_94_1008 VPWR VGND sg13g2_decap_8
XFILLER_73_130 VPWR VGND sg13g2_decap_8
XFILLER_62_826 VPWR VGND sg13g2_decap_8
XFILLER_47_889 VPWR VGND sg13g2_decap_8
XFILLER_104_91 VPWR VGND sg13g2_decap_8
XFILLER_64_95 VPWR VGND sg13g2_decap_8
XFILLER_61_347 VPWR VGND sg13g2_decap_8
XFILLER_15_753 VPWR VGND sg13g2_decap_8
XFILLER_42_550 VPWR VGND sg13g2_decap_8
XFILLER_9_35 VPWR VGND sg13g2_decap_8
XFILLER_14_252 VPWR VGND sg13g2_decap_8
XFILLER_30_756 VPWR VGND sg13g2_decap_8
XFILLER_10_480 VPWR VGND sg13g2_decap_8
XFILLER_7_963 VPWR VGND sg13g2_decap_8
XFILLER_6_462 VPWR VGND sg13g2_decap_8
XFILLER_89_70 VPWR VGND sg13g2_decap_8
XFILLER_69_414 VPWR VGND sg13g2_decap_8
XFILLER_9_1015 VPWR VGND sg13g2_decap_8
XFILLER_97_756 VPWR VGND sg13g2_decap_8
XFILLER_57_609 VPWR VGND sg13g2_decap_8
XFILLER_2_690 VPWR VGND sg13g2_decap_8
XFILLER_96_266 VPWR VGND sg13g2_decap_8
XFILLER_84_406 VPWR VGND sg13g2_decap_8
XFILLER_38_812 VPWR VGND sg13g2_decap_8
XFILLER_49_193 VPWR VGND sg13g2_decap_8
XFILLER_37_333 VPWR VGND sg13g2_decap_8
X_47_ net13 net5 _15_ VPWR VGND sg13g2_xor2_1
XFILLER_64_130 VPWR VGND sg13g2_decap_8
XFILLER_38_889 VPWR VGND sg13g2_decap_8
XFILLER_92_483 VPWR VGND sg13g2_decap_8
XFILLER_80_623 VPWR VGND sg13g2_decap_8
XFILLER_65_686 VPWR VGND sg13g2_decap_8
XFILLER_53_826 VPWR VGND sg13g2_decap_8
XFILLER_25_539 VPWR VGND sg13g2_decap_8
XFILLER_52_336 VPWR VGND sg13g2_decap_8
XFILLER_100_49 VPWR VGND sg13g2_decap_8
XFILLER_20_200 VPWR VGND sg13g2_decap_8
XFILLER_21_756 VPWR VGND sg13g2_decap_8
XFILLER_20_277 VPWR VGND sg13g2_decap_8
XFILLER_102_511 VPWR VGND sg13g2_decap_8
XFILLER_0_616 VPWR VGND sg13g2_decap_8
XFILLER_88_767 VPWR VGND sg13g2_decap_8
XFILLER_76_907 VPWR VGND sg13g2_decap_8
XFILLER_48_609 VPWR VGND sg13g2_decap_8
XFILLER_102_588 VPWR VGND sg13g2_decap_8
XFILLER_87_266 VPWR VGND sg13g2_decap_8
XFILLER_85_28 VPWR VGND sg13g2_decap_8
XFILLER_75_406 VPWR VGND sg13g2_decap_8
XFILLER_69_981 VPWR VGND sg13g2_decap_8
XFILLER_47_119 VPWR VGND sg13g2_decap_8
XFILLER_29_823 VPWR VGND sg13g2_decap_8
XFILLER_56_620 VPWR VGND sg13g2_decap_8
XFILLER_28_322 VPWR VGND sg13g2_decap_8
XFILLER_84_973 VPWR VGND sg13g2_decap_8
XFILLER_18_77 VPWR VGND sg13g2_decap_8
XFILLER_83_494 VPWR VGND sg13g2_decap_8
XFILLER_71_634 VPWR VGND sg13g2_decap_8
XFILLER_56_697 VPWR VGND sg13g2_decap_8
XFILLER_44_837 VPWR VGND sg13g2_decap_8
XFILLER_16_539 VPWR VGND sg13g2_decap_8
XFILLER_28_399 VPWR VGND sg13g2_decap_8
XFILLER_70_133 VPWR VGND sg13g2_decap_8
XFILLER_55_196 VPWR VGND sg13g2_decap_8
XFILLER_43_336 VPWR VGND sg13g2_decap_8
XFILLER_24_550 VPWR VGND sg13g2_decap_8
XFILLER_34_32 VPWR VGND sg13g2_decap_8
XFILLER_11_266 VPWR VGND sg13g2_decap_8
XFILLER_12_767 VPWR VGND sg13g2_decap_8
XFILLER_50_42 VPWR VGND sg13g2_decap_8
XFILLER_8_749 VPWR VGND sg13g2_decap_8
XFILLER_106_861 VPWR VGND sg13g2_decap_8
XFILLER_4_966 VPWR VGND sg13g2_decap_8
XFILLER_105_371 VPWR VGND sg13g2_decap_8
XFILLER_3_476 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_decap_8
XFILLER_79_767 VPWR VGND sg13g2_decap_8
XFILLER_78_244 VPWR VGND sg13g2_decap_8
XFILLER_38_119 VPWR VGND sg13g2_decap_8
XFILLER_93_236 VPWR VGND sg13g2_decap_8
XFILLER_19_322 VPWR VGND sg13g2_decap_8
XFILLER_75_973 VPWR VGND sg13g2_decap_8
XFILLER_46_130 VPWR VGND sg13g2_decap_8
XFILLER_90_921 VPWR VGND sg13g2_decap_8
XFILLER_62_623 VPWR VGND sg13g2_decap_8
XFILLER_47_686 VPWR VGND sg13g2_decap_8
XFILLER_19_399 VPWR VGND sg13g2_decap_8
XFILLER_35_826 VPWR VGND sg13g2_decap_8
XFILLER_34_347 VPWR VGND sg13g2_decap_8
XFILLER_90_998 VPWR VGND sg13g2_decap_8
XFILLER_15_550 VPWR VGND sg13g2_decap_8
XFILLER_30_553 VPWR VGND sg13g2_decap_8
XFILLER_7_760 VPWR VGND sg13g2_decap_8
XFILLER_103_308 VPWR VGND sg13g2_decap_8
XFILLER_69_211 VPWR VGND sg13g2_decap_8
XFILLER_97_553 VPWR VGND sg13g2_decap_8
XFILLER_84_203 VPWR VGND sg13g2_decap_8
XFILLER_57_406 VPWR VGND sg13g2_decap_8
XFILLER_69_288 VPWR VGND sg13g2_decap_8
XFILLER_66_951 VPWR VGND sg13g2_decap_8
XFILLER_37_130 VPWR VGND sg13g2_decap_8
XFILLER_81_921 VPWR VGND sg13g2_decap_8
XFILLER_65_483 VPWR VGND sg13g2_decap_8
XFILLER_53_623 VPWR VGND sg13g2_decap_8
XFILLER_1_91 VPWR VGND sg13g2_decap_8
XFILLER_26_826 VPWR VGND sg13g2_decap_8
XFILLER_38_686 VPWR VGND sg13g2_decap_8
XFILLER_92_280 VPWR VGND sg13g2_decap_8
XFILLER_80_420 VPWR VGND sg13g2_decap_8
XFILLER_52_133 VPWR VGND sg13g2_decap_8
XFILLER_25_336 VPWR VGND sg13g2_decap_8
XFILLER_81_998 VPWR VGND sg13g2_decap_8
XFILLER_80_497 VPWR VGND sg13g2_decap_8
XFILLER_21_553 VPWR VGND sg13g2_decap_8
XFILLER_101_1001 VPWR VGND sg13g2_decap_8
XFILLER_1_903 VPWR VGND sg13g2_decap_8
XFILLER_20_67 VPWR VGND sg13g2_decap_8
XFILLER_106_168 VPWR VGND sg13g2_decap_8
XFILLER_0_413 VPWR VGND sg13g2_decap_8
XFILLER_96_49 VPWR VGND sg13g2_decap_8
XFILLER_49_907 VPWR VGND sg13g2_decap_8
XFILLER_103_875 VPWR VGND sg13g2_decap_8
XFILLER_88_564 VPWR VGND sg13g2_decap_8
XFILLER_76_704 VPWR VGND sg13g2_decap_8
XFILLER_75_203 VPWR VGND sg13g2_decap_8
XFILLER_48_406 VPWR VGND sg13g2_decap_8
XFILLER_29_32 VPWR VGND sg13g2_decap_8
XFILLER_102_385 VPWR VGND sg13g2_decap_8
XFILLER_29_620 VPWR VGND sg13g2_decap_8
XFILLER_91_707 VPWR VGND sg13g2_decap_8
XFILLER_57_973 VPWR VGND sg13g2_decap_8
XFILLER_90_228 VPWR VGND sg13g2_decap_8
XFILLER_84_770 VPWR VGND sg13g2_decap_8
XFILLER_72_910 VPWR VGND sg13g2_decap_8
XFILLER_17_837 VPWR VGND sg13g2_decap_8
XFILLER_29_697 VPWR VGND sg13g2_decap_8
XFILLER_83_291 VPWR VGND sg13g2_decap_8
XFILLER_71_431 VPWR VGND sg13g2_decap_8
XFILLER_56_494 VPWR VGND sg13g2_decap_8
XFILLER_45_42 VPWR VGND sg13g2_decap_8
XFILLER_44_634 VPWR VGND sg13g2_decap_8
XFILLER_43_133 VPWR VGND sg13g2_decap_8
XFILLER_16_336 VPWR VGND sg13g2_decap_8
XFILLER_28_196 VPWR VGND sg13g2_decap_8
XFILLER_72_987 VPWR VGND sg13g2_decap_8
XFILLER_101_70 VPWR VGND sg13g2_decap_8
XFILLER_12_564 VPWR VGND sg13g2_decap_8
XFILLER_40_840 VPWR VGND sg13g2_decap_8
XFILLER_61_74 VPWR VGND sg13g2_decap_8
XFILLER_8_546 VPWR VGND sg13g2_decap_8
XFILLER_6_14 VPWR VGND sg13g2_decap_8
XFILLER_4_763 VPWR VGND sg13g2_decap_8
XFILLER_3_273 VPWR VGND sg13g2_decap_8
XFILLER_79_564 VPWR VGND sg13g2_decap_8
XFILLER_39_417 VPWR VGND sg13g2_decap_8
XFILLER_86_60 VPWR VGND sg13g2_decap_8
XFILLER_0_980 VPWR VGND sg13g2_decap_8
XFILLER_94_567 VPWR VGND sg13g2_decap_8
XFILLER_82_707 VPWR VGND sg13g2_decap_8
XFILLER_66_258 VPWR VGND sg13g2_decap_8
XFILLER_48_973 VPWR VGND sg13g2_decap_8
XFILLER_81_228 VPWR VGND sg13g2_decap_8
XFILLER_75_770 VPWR VGND sg13g2_decap_8
XFILLER_63_910 VPWR VGND sg13g2_decap_8
XFILLER_47_483 VPWR VGND sg13g2_decap_8
XFILLER_35_623 VPWR VGND sg13g2_decap_8
XFILLER_62_420 VPWR VGND sg13g2_decap_8
XFILLER_19_196 VPWR VGND sg13g2_decap_8
XFILLER_63_987 VPWR VGND sg13g2_decap_8
XFILLER_34_144 VPWR VGND sg13g2_decap_8
XFILLER_90_795 VPWR VGND sg13g2_decap_8
XFILLER_62_497 VPWR VGND sg13g2_decap_8
XFILLER_50_637 VPWR VGND sg13g2_decap_8
XFILLER_31_840 VPWR VGND sg13g2_decap_8
XFILLER_30_350 VPWR VGND sg13g2_decap_8
XFILLER_103_105 VPWR VGND sg13g2_decap_8
XFILLER_98_851 VPWR VGND sg13g2_decap_8
XFILLER_100_812 VPWR VGND sg13g2_decap_8
XFILLER_97_350 VPWR VGND sg13g2_decap_8
XFILLER_57_203 VPWR VGND sg13g2_decap_8
XFILLER_85_567 VPWR VGND sg13g2_decap_8
XFILLER_73_718 VPWR VGND sg13g2_decap_8
XFILLER_100_889 VPWR VGND sg13g2_decap_8
XFILLER_72_217 VPWR VGND sg13g2_decap_8
XFILLER_54_921 VPWR VGND sg13g2_decap_8
XFILLER_26_623 VPWR VGND sg13g2_decap_8
XFILLER_38_483 VPWR VGND sg13g2_decap_8
XFILLER_39_984 VPWR VGND sg13g2_decap_8
XFILLER_65_280 VPWR VGND sg13g2_decap_8
XFILLER_53_420 VPWR VGND sg13g2_decap_8
XFILLER_25_133 VPWR VGND sg13g2_decap_8
XFILLER_54_998 VPWR VGND sg13g2_decap_8
XFILLER_81_795 VPWR VGND sg13g2_decap_8
XFILLER_80_294 VPWR VGND sg13g2_decap_8
XFILLER_53_497 VPWR VGND sg13g2_decap_8
XFILLER_41_637 VPWR VGND sg13g2_decap_8
XFILLER_15_67 VPWR VGND sg13g2_decap_8
XFILLER_22_851 VPWR VGND sg13g2_decap_8
XFILLER_40_147 VPWR VGND sg13g2_decap_8
XFILLER_51_1028 VPWR VGND sg13g2_fill_1
XFILLER_21_350 VPWR VGND sg13g2_decap_8
XFILLER_31_77 VPWR VGND sg13g2_decap_8
XFILLER_1_700 VPWR VGND sg13g2_decap_8
Xoutput22 net22 uo_out[5] VPWR VGND sg13g2_buf_1
XFILLER_89_840 VPWR VGND sg13g2_decap_8
XFILLER_0_210 VPWR VGND sg13g2_decap_8
XFILLER_88_361 VPWR VGND sg13g2_decap_8
XFILLER_76_501 VPWR VGND sg13g2_decap_8
XFILLER_49_704 VPWR VGND sg13g2_decap_8
XFILLER_1_777 VPWR VGND sg13g2_decap_8
XFILLER_103_672 VPWR VGND sg13g2_decap_8
XFILLER_48_203 VPWR VGND sg13g2_decap_8
XFILLER_0_287 VPWR VGND sg13g2_decap_8
XFILLER_102_182 VPWR VGND sg13g2_decap_8
XFILLER_76_578 VPWR VGND sg13g2_decap_8
XFILLER_64_718 VPWR VGND sg13g2_decap_8
XFILLER_91_504 VPWR VGND sg13g2_decap_8
XFILLER_63_217 VPWR VGND sg13g2_decap_8
XFILLER_57_770 VPWR VGND sg13g2_decap_8
XFILLER_56_74 VPWR VGND sg13g2_decap_8
XFILLER_45_910 VPWR VGND sg13g2_decap_8
XFILLER_56_291 VPWR VGND sg13g2_decap_8
XFILLER_44_431 VPWR VGND sg13g2_decap_8
XFILLER_17_634 VPWR VGND sg13g2_decap_8
XFILLER_29_494 VPWR VGND sg13g2_decap_8
XFILLER_72_784 VPWR VGND sg13g2_decap_8
XFILLER_45_987 VPWR VGND sg13g2_decap_8
XFILLER_16_133 VPWR VGND sg13g2_decap_8
XFILLER_60_935 VPWR VGND sg13g2_decap_8
XFILLER_32_648 VPWR VGND sg13g2_decap_8
XFILLER_72_84 VPWR VGND sg13g2_decap_8
XFILLER_13_840 VPWR VGND sg13g2_decap_8
XFILLER_31_147 VPWR VGND sg13g2_decap_8
XFILLER_9_833 VPWR VGND sg13g2_decap_8
XFILLER_12_361 VPWR VGND sg13g2_decap_8
XFILLER_75_7 VPWR VGND sg13g2_decap_8
XFILLER_8_343 VPWR VGND sg13g2_decap_8
XFILLER_99_637 VPWR VGND sg13g2_decap_8
XFILLER_4_560 VPWR VGND sg13g2_decap_8
XFILLER_28_1008 VPWR VGND sg13g2_decap_8
XFILLER_101_609 VPWR VGND sg13g2_decap_8
XFILLER_98_158 VPWR VGND sg13g2_decap_8
XFILLER_97_70 VPWR VGND sg13g2_decap_8
XFILLER_79_361 VPWR VGND sg13g2_decap_8
XFILLER_100_119 VPWR VGND sg13g2_decap_8
XFILLER_39_214 VPWR VGND sg13g2_decap_8
XFILLER_95_865 VPWR VGND sg13g2_decap_8
XFILLER_67_567 VPWR VGND sg13g2_decap_8
XFILLER_55_707 VPWR VGND sg13g2_decap_8
XFILLER_94_364 VPWR VGND sg13g2_decap_8
XFILLER_82_504 VPWR VGND sg13g2_decap_8
XFILLER_48_770 VPWR VGND sg13g2_decap_8
XFILLER_36_910 VPWR VGND sg13g2_decap_8
XFILLER_54_228 VPWR VGND sg13g2_decap_8
XFILLER_47_280 VPWR VGND sg13g2_decap_8
XFILLER_35_420 VPWR VGND sg13g2_decap_8
XFILLER_63_784 VPWR VGND sg13g2_decap_8
XFILLER_36_987 VPWR VGND sg13g2_decap_8
XFILLER_90_592 VPWR VGND sg13g2_decap_8
XFILLER_51_935 VPWR VGND sg13g2_decap_8
XFILLER_50_434 VPWR VGND sg13g2_decap_8
XFILLER_23_637 VPWR VGND sg13g2_decap_8
XFILLER_35_497 VPWR VGND sg13g2_decap_8
XFILLER_62_294 VPWR VGND sg13g2_decap_8
XFILLER_22_158 VPWR VGND sg13g2_decap_8
XFILLER_11_1001 VPWR VGND sg13g2_decap_8
XFILLER_2_508 VPWR VGND sg13g2_decap_8
XFILLER_105_959 VPWR VGND sg13g2_decap_8
XFILLER_104_469 VPWR VGND sg13g2_decap_8
XFILLER_89_147 VPWR VGND sg13g2_decap_8
XFILLER_86_865 VPWR VGND sg13g2_decap_8
XFILLER_58_567 VPWR VGND sg13g2_decap_8
XFILLER_100_686 VPWR VGND sg13g2_decap_8
XFILLER_85_364 VPWR VGND sg13g2_decap_8
XFILLER_73_515 VPWR VGND sg13g2_decap_8
XFILLER_46_718 VPWR VGND sg13g2_decap_8
XFILLER_45_217 VPWR VGND sg13g2_decap_8
XFILLER_27_921 VPWR VGND sg13g2_decap_8
XFILLER_39_781 VPWR VGND sg13g2_decap_8
XFILLER_26_420 VPWR VGND sg13g2_decap_8
XFILLER_38_280 VPWR VGND sg13g2_decap_8
XFILLER_27_998 VPWR VGND sg13g2_decap_8
XFILLER_81_592 VPWR VGND sg13g2_decap_8
XFILLER_54_795 VPWR VGND sg13g2_decap_8
XFILLER_42_935 VPWR VGND sg13g2_decap_8
XFILLER_14_637 VPWR VGND sg13g2_decap_8
XFILLER_26_77 VPWR VGND sg13g2_decap_8
XFILLER_26_497 VPWR VGND sg13g2_decap_8
XFILLER_53_294 VPWR VGND sg13g2_decap_8
XFILLER_13_147 VPWR VGND sg13g2_decap_8
XFILLER_41_434 VPWR VGND sg13g2_decap_8
XFILLER_42_32 VPWR VGND sg13g2_decap_8
XFILLER_10_865 VPWR VGND sg13g2_decap_8
XFILLER_6_847 VPWR VGND sg13g2_decap_8
XFILLER_101_0 VPWR VGND sg13g2_decap_8
XFILLER_5_368 VPWR VGND sg13g2_decap_8
XFILLER_49_501 VPWR VGND sg13g2_decap_8
XFILLER_1_574 VPWR VGND sg13g2_decap_8
XFILLER_77_854 VPWR VGND sg13g2_decap_8
XFILLER_67_84 VPWR VGND sg13g2_decap_8
XFILLER_91_301 VPWR VGND sg13g2_decap_8
XFILLER_76_375 VPWR VGND sg13g2_decap_8
XFILLER_64_515 VPWR VGND sg13g2_decap_8
XFILLER_49_578 VPWR VGND sg13g2_decap_8
XFILLER_18_910 VPWR VGND sg13g2_decap_8
XFILLER_36_217 VPWR VGND sg13g2_decap_8
XFILLER_37_718 VPWR VGND sg13g2_decap_8
XFILLER_92_868 VPWR VGND sg13g2_decap_8
XFILLER_17_431 VPWR VGND sg13g2_decap_8
XFILLER_29_291 VPWR VGND sg13g2_decap_8
XFILLER_91_378 VPWR VGND sg13g2_decap_8
XFILLER_18_987 VPWR VGND sg13g2_decap_8
XFILLER_72_581 VPWR VGND sg13g2_decap_8
XFILLER_60_732 VPWR VGND sg13g2_decap_8
XFILLER_45_784 VPWR VGND sg13g2_decap_8
XFILLER_33_924 VPWR VGND sg13g2_decap_8
XFILLER_32_445 VPWR VGND sg13g2_decap_8
XFILLER_34_1012 VPWR VGND sg13g2_decap_8
XFILLER_9_630 VPWR VGND sg13g2_decap_8
XFILLER_73_4 VPWR VGND sg13g2_decap_8
XFILLER_8_140 VPWR VGND sg13g2_decap_8
XFILLER_99_434 VPWR VGND sg13g2_decap_8
XFILLER_101_406 VPWR VGND sg13g2_decap_8
XFILLER_68_810 VPWR VGND sg13g2_decap_8
XFILLER_28_707 VPWR VGND sg13g2_decap_8
XFILLER_95_662 VPWR VGND sg13g2_decap_8
XFILLER_94_161 VPWR VGND sg13g2_decap_8
XFILLER_83_802 VPWR VGND sg13g2_decap_8
XFILLER_82_301 VPWR VGND sg13g2_decap_8
XFILLER_68_887 VPWR VGND sg13g2_decap_8
XFILLER_67_364 VPWR VGND sg13g2_decap_8
XFILLER_55_504 VPWR VGND sg13g2_decap_8
XFILLER_103_49 VPWR VGND sg13g2_decap_8
XFILLER_27_228 VPWR VGND sg13g2_decap_8
XFILLER_83_879 VPWR VGND sg13g2_decap_8
XFILLER_82_378 VPWR VGND sg13g2_decap_8
XFILLER_70_518 VPWR VGND sg13g2_decap_8
XFILLER_63_581 VPWR VGND sg13g2_decap_8
XFILLER_51_732 VPWR VGND sg13g2_decap_8
XFILLER_24_935 VPWR VGND sg13g2_decap_8
XFILLER_36_784 VPWR VGND sg13g2_decap_8
XFILLER_50_231 VPWR VGND sg13g2_decap_8
XFILLER_23_434 VPWR VGND sg13g2_decap_8
XFILLER_35_294 VPWR VGND sg13g2_decap_8
XFILLER_12_46 VPWR VGND sg13g2_decap_8
XFILLER_2_305 VPWR VGND sg13g2_decap_8
XFILLER_88_39 VPWR VGND sg13g2_decap_8
XFILLER_105_756 VPWR VGND sg13g2_decap_8
XFILLER_104_266 VPWR VGND sg13g2_decap_8
XFILLER_78_629 VPWR VGND sg13g2_decap_8
XFILLER_59_810 VPWR VGND sg13g2_decap_8
XFILLER_101_973 VPWR VGND sg13g2_decap_8
XFILLER_86_662 VPWR VGND sg13g2_decap_8
XFILLER_85_161 VPWR VGND sg13g2_decap_8
XFILLER_74_813 VPWR VGND sg13g2_decap_8
XFILLER_59_887 VPWR VGND sg13g2_decap_8
XFILLER_58_364 VPWR VGND sg13g2_decap_8
XFILLER_46_515 VPWR VGND sg13g2_decap_8
XFILLER_19_707 VPWR VGND sg13g2_decap_8
XFILLER_37_32 VPWR VGND sg13g2_decap_8
XFILLER_100_483 VPWR VGND sg13g2_decap_8
XFILLER_73_312 VPWR VGND sg13g2_decap_8
XFILLER_18_217 VPWR VGND sg13g2_decap_8
XFILLER_57_1001 VPWR VGND sg13g2_decap_8
XFILLER_73_389 VPWR VGND sg13g2_decap_8
XFILLER_61_529 VPWR VGND sg13g2_decap_8
XFILLER_42_732 VPWR VGND sg13g2_decap_8
XFILLER_15_935 VPWR VGND sg13g2_decap_8
XFILLER_27_795 VPWR VGND sg13g2_decap_8
XFILLER_54_592 VPWR VGND sg13g2_decap_8
XFILLER_53_42 VPWR VGND sg13g2_decap_8
XFILLER_14_434 VPWR VGND sg13g2_decap_8
XFILLER_26_294 VPWR VGND sg13g2_decap_8
XFILLER_41_231 VPWR VGND sg13g2_decap_8
XFILLER_30_938 VPWR VGND sg13g2_decap_8
XFILLER_10_662 VPWR VGND sg13g2_decap_8
XFILLER_6_644 VPWR VGND sg13g2_decap_8
XFILLER_64_1005 VPWR VGND sg13g2_decap_8
XFILLER_5_165 VPWR VGND sg13g2_decap_8
XFILLER_97_938 VPWR VGND sg13g2_decap_8
XFILLER_78_83 VPWR VGND sg13g2_decap_8
XFILLER_68_117 VPWR VGND sg13g2_decap_8
XFILLER_2_872 VPWR VGND sg13g2_decap_8
XFILLER_1_371 VPWR VGND sg13g2_decap_8
XFILLER_38_7 VPWR VGND sg13g2_decap_8
XFILLER_96_448 VPWR VGND sg13g2_decap_8
XFILLER_77_651 VPWR VGND sg13g2_decap_8
XFILLER_83_109 VPWR VGND sg13g2_decap_8
X_63_ _28_ net8 net16 VPWR VGND sg13g2_xnor2_1
XFILLER_49_375 VPWR VGND sg13g2_decap_8
XFILLER_37_515 VPWR VGND sg13g2_decap_8
XFILLER_76_172 VPWR VGND sg13g2_decap_8
XFILLER_64_312 VPWR VGND sg13g2_decap_8
XFILLER_92_665 VPWR VGND sg13g2_decap_8
XFILLER_80_805 VPWR VGND sg13g2_decap_8
XFILLER_65_868 VPWR VGND sg13g2_decap_8
XFILLER_52_518 VPWR VGND sg13g2_decap_8
XFILLER_91_175 VPWR VGND sg13g2_decap_8
XFILLER_64_389 VPWR VGND sg13g2_decap_8
XFILLER_45_581 VPWR VGND sg13g2_decap_8
XFILLER_18_784 VPWR VGND sg13g2_decap_8
XFILLER_33_721 VPWR VGND sg13g2_decap_8
XFILLER_21_938 VPWR VGND sg13g2_decap_8
XFILLER_32_242 VPWR VGND sg13g2_decap_8
XFILLER_33_798 VPWR VGND sg13g2_decap_8
XFILLER_20_459 VPWR VGND sg13g2_decap_8
XFILLER_99_231 VPWR VGND sg13g2_decap_8
XFILLER_101_203 VPWR VGND sg13g2_decap_8
XFILLER_88_949 VPWR VGND sg13g2_decap_8
XFILLER_59_106 VPWR VGND sg13g2_decap_8
XFILLER_87_448 VPWR VGND sg13g2_decap_8
XFILLER_4_91 VPWR VGND sg13g2_decap_8
XFILLER_68_684 VPWR VGND sg13g2_decap_8
XFILLER_56_802 VPWR VGND sg13g2_decap_8
XFILLER_55_301 VPWR VGND sg13g2_decap_8
XFILLER_28_504 VPWR VGND sg13g2_decap_8
XFILLER_67_161 VPWR VGND sg13g2_decap_8
XFILLER_83_676 VPWR VGND sg13g2_decap_8
XFILLER_71_816 VPWR VGND sg13g2_decap_8
XFILLER_56_879 VPWR VGND sg13g2_decap_8
XFILLER_82_175 VPWR VGND sg13g2_decap_8
XFILLER_70_315 VPWR VGND sg13g2_decap_8
XFILLER_55_378 VPWR VGND sg13g2_decap_8
XFILLER_43_518 VPWR VGND sg13g2_decap_8
XFILLER_36_581 VPWR VGND sg13g2_decap_8
XFILLER_90_18 VPWR VGND sg13g2_decap_8
XFILLER_23_231 VPWR VGND sg13g2_decap_8
XFILLER_24_732 VPWR VGND sg13g2_decap_8
XFILLER_11_448 VPWR VGND sg13g2_decap_8
XFILLER_12_949 VPWR VGND sg13g2_decap_8
XFILLER_23_56 VPWR VGND sg13g2_decap_8
XFILLER_99_49 VPWR VGND sg13g2_decap_8
XFILLER_2_102 VPWR VGND sg13g2_decap_8
XFILLER_105_553 VPWR VGND sg13g2_decap_8
XFILLER_3_658 VPWR VGND sg13g2_decap_8
XFILLER_79_949 VPWR VGND sg13g2_decap_8
XFILLER_78_426 VPWR VGND sg13g2_decap_8
XFILLER_2_179 VPWR VGND sg13g2_decap_8
XFILLER_48_42 VPWR VGND sg13g2_decap_8
XFILLER_101_770 VPWR VGND sg13g2_decap_8
XFILLER_93_418 VPWR VGND sg13g2_decap_8
XFILLER_19_504 VPWR VGND sg13g2_decap_8
XFILLER_100_280 VPWR VGND sg13g2_decap_8
XFILLER_74_610 VPWR VGND sg13g2_decap_8
XFILLER_59_684 VPWR VGND sg13g2_decap_8
XFILLER_58_161 VPWR VGND sg13g2_decap_8
XFILLER_46_312 VPWR VGND sg13g2_decap_8
XFILLER_104_70 VPWR VGND sg13g2_decap_8
XFILLER_62_805 VPWR VGND sg13g2_decap_8
XFILLER_47_868 VPWR VGND sg13g2_decap_8
XFILLER_0_49 VPWR VGND sg13g2_decap_8
XFILLER_74_687 VPWR VGND sg13g2_decap_8
XFILLER_73_186 VPWR VGND sg13g2_decap_8
XFILLER_61_326 VPWR VGND sg13g2_decap_8
XFILLER_46_389 VPWR VGND sg13g2_decap_8
XFILLER_34_529 VPWR VGND sg13g2_decap_8
XFILLER_64_74 VPWR VGND sg13g2_decap_8
XFILLER_14_231 VPWR VGND sg13g2_decap_8
XFILLER_15_732 VPWR VGND sg13g2_decap_8
XFILLER_27_592 VPWR VGND sg13g2_decap_8
XFILLER_70_882 VPWR VGND sg13g2_decap_8
XFILLER_9_14 VPWR VGND sg13g2_decap_8
XFILLER_30_735 VPWR VGND sg13g2_decap_8
XFILLER_80_84 VPWR VGND sg13g2_decap_8
XFILLER_31_1015 VPWR VGND sg13g2_decap_8
XFILLER_7_942 VPWR VGND sg13g2_decap_8
XFILLER_6_441 VPWR VGND sg13g2_decap_8
XFILLER_97_735 VPWR VGND sg13g2_decap_8
XFILLER_96_245 VPWR VGND sg13g2_decap_8
XFILLER_56_109 VPWR VGND sg13g2_decap_8
XFILLER_78_993 VPWR VGND sg13g2_decap_8
XFILLER_49_172 VPWR VGND sg13g2_decap_8
XFILLER_37_312 VPWR VGND sg13g2_decap_8
XFILLER_93_985 VPWR VGND sg13g2_decap_8
X_46_ _14_ net5 net13 VPWR VGND sg13g2_nand2_1
XFILLER_65_665 VPWR VGND sg13g2_decap_8
XFILLER_53_805 VPWR VGND sg13g2_decap_8
XFILLER_38_868 VPWR VGND sg13g2_decap_8
XFILLER_92_462 VPWR VGND sg13g2_decap_8
XFILLER_80_602 VPWR VGND sg13g2_decap_8
XFILLER_64_186 VPWR VGND sg13g2_decap_8
XFILLER_52_315 VPWR VGND sg13g2_decap_8
XFILLER_25_518 VPWR VGND sg13g2_decap_8
XFILLER_37_389 VPWR VGND sg13g2_decap_8
XFILLER_18_581 VPWR VGND sg13g2_decap_8
XFILLER_100_28 VPWR VGND sg13g2_decap_8
XFILLER_80_679 VPWR VGND sg13g2_decap_8
XFILLER_61_893 VPWR VGND sg13g2_decap_8
XFILLER_21_735 VPWR VGND sg13g2_decap_8
XFILLER_33_595 VPWR VGND sg13g2_decap_8
XFILLER_20_256 VPWR VGND sg13g2_decap_8
XFILLER_47_1022 VPWR VGND sg13g2_decap_8
XFILLER_88_746 VPWR VGND sg13g2_decap_8
XFILLER_87_245 VPWR VGND sg13g2_decap_8
XFILLER_102_567 VPWR VGND sg13g2_decap_8
XFILLER_69_960 VPWR VGND sg13g2_decap_8
XFILLER_29_802 VPWR VGND sg13g2_decap_8
XFILLER_68_481 VPWR VGND sg13g2_decap_8
XFILLER_28_301 VPWR VGND sg13g2_decap_8
XFILLER_84_952 VPWR VGND sg13g2_decap_8
XFILLER_44_816 VPWR VGND sg13g2_decap_8
XFILLER_18_56 VPWR VGND sg13g2_decap_8
XFILLER_29_879 VPWR VGND sg13g2_decap_8
XFILLER_83_473 VPWR VGND sg13g2_decap_8
XFILLER_71_613 VPWR VGND sg13g2_decap_8
XFILLER_56_676 VPWR VGND sg13g2_decap_8
XFILLER_55_175 VPWR VGND sg13g2_decap_8
XFILLER_43_315 VPWR VGND sg13g2_decap_8
XFILLER_16_518 VPWR VGND sg13g2_decap_8
XFILLER_28_378 VPWR VGND sg13g2_decap_8
XFILLER_93_1020 VPWR VGND sg13g2_decap_8
XFILLER_70_112 VPWR VGND sg13g2_decap_8
XFILLER_34_11 VPWR VGND sg13g2_decap_8
XFILLER_52_882 VPWR VGND sg13g2_decap_8
XFILLER_70_189 VPWR VGND sg13g2_decap_8
XFILLER_54_1026 VPWR VGND sg13g2_fill_2
XFILLER_12_746 VPWR VGND sg13g2_decap_8
XFILLER_34_88 VPWR VGND sg13g2_decap_8
XFILLER_8_728 VPWR VGND sg13g2_decap_8
XFILLER_11_245 VPWR VGND sg13g2_decap_8
XFILLER_50_21 VPWR VGND sg13g2_decap_8
XFILLER_7_249 VPWR VGND sg13g2_decap_8
XFILLER_50_98 VPWR VGND sg13g2_decap_8
XFILLER_106_840 VPWR VGND sg13g2_decap_8
XFILLER_4_945 VPWR VGND sg13g2_decap_8
XFILLER_105_350 VPWR VGND sg13g2_decap_8
XFILLER_3_455 VPWR VGND sg13g2_decap_8
XFILLER_79_746 VPWR VGND sg13g2_decap_8
XFILLER_78_223 VPWR VGND sg13g2_decap_8
XFILLER_61_1019 VPWR VGND sg13g2_decap_8
XFILLER_59_85 VPWR VGND sg13g2_decap_8
XFILLER_94_749 VPWR VGND sg13g2_decap_8
XFILLER_93_215 VPWR VGND sg13g2_decap_8
XFILLER_59_481 VPWR VGND sg13g2_decap_8
XFILLER_19_301 VPWR VGND sg13g2_decap_8
XFILLER_90_900 VPWR VGND sg13g2_decap_8
XFILLER_75_952 VPWR VGND sg13g2_decap_8
XFILLER_47_665 VPWR VGND sg13g2_decap_8
XFILLER_35_805 VPWR VGND sg13g2_decap_8
XFILLER_75_84 VPWR VGND sg13g2_decap_8
XFILLER_74_484 VPWR VGND sg13g2_decap_8
XFILLER_62_602 VPWR VGND sg13g2_decap_8
XFILLER_19_378 VPWR VGND sg13g2_decap_8
XFILLER_90_977 VPWR VGND sg13g2_decap_8
XFILLER_61_123 VPWR VGND sg13g2_decap_8
XFILLER_46_186 VPWR VGND sg13g2_decap_8
XFILLER_34_326 VPWR VGND sg13g2_decap_8
XFILLER_62_679 VPWR VGND sg13g2_decap_8
XFILLER_50_819 VPWR VGND sg13g2_decap_8
XFILLER_43_882 VPWR VGND sg13g2_decap_8
XFILLER_30_532 VPWR VGND sg13g2_decap_8
XFILLER_97_532 VPWR VGND sg13g2_decap_8
XFILLER_69_267 VPWR VGND sg13g2_decap_8
XFILLER_29_109 VPWR VGND sg13g2_decap_8
XFILLER_85_749 VPWR VGND sg13g2_decap_8
XFILLER_78_790 VPWR VGND sg13g2_decap_8
XFILLER_66_930 VPWR VGND sg13g2_decap_8
XFILLER_84_259 VPWR VGND sg13g2_decap_8
XFILLER_81_900 VPWR VGND sg13g2_decap_8
XFILLER_26_805 VPWR VGND sg13g2_decap_8
XFILLER_38_665 VPWR VGND sg13g2_decap_8
XFILLER_93_782 VPWR VGND sg13g2_decap_8
XFILLER_77_1015 VPWR VGND sg13g2_decap_8
XFILLER_65_462 VPWR VGND sg13g2_decap_8
X_29_ net1 net9 _00_ VPWR VGND sg13g2_and2_1
XFILLER_53_602 VPWR VGND sg13g2_decap_8
XFILLER_1_70 VPWR VGND sg13g2_decap_8
XFILLER_25_315 VPWR VGND sg13g2_decap_8
XFILLER_52_112 VPWR VGND sg13g2_decap_8
XFILLER_37_186 VPWR VGND sg13g2_decap_8
XFILLER_81_977 VPWR VGND sg13g2_decap_8
XFILLER_80_476 VPWR VGND sg13g2_decap_8
XFILLER_53_679 VPWR VGND sg13g2_decap_8
XFILLER_41_819 VPWR VGND sg13g2_decap_8
XFILLER_61_690 VPWR VGND sg13g2_decap_8
XFILLER_52_189 VPWR VGND sg13g2_decap_8
XFILLER_34_893 VPWR VGND sg13g2_decap_8
XFILLER_40_329 VPWR VGND sg13g2_decap_8
XFILLER_21_532 VPWR VGND sg13g2_decap_8
XFILLER_33_392 VPWR VGND sg13g2_decap_8
XFILLER_106_147 VPWR VGND sg13g2_decap_8
XFILLER_105_7 VPWR VGND sg13g2_decap_8
XFILLER_84_1008 VPWR VGND sg13g2_decap_8
XFILLER_20_46 VPWR VGND sg13g2_decap_8
XFILLER_103_854 VPWR VGND sg13g2_decap_8
XFILLER_96_28 VPWR VGND sg13g2_decap_8
XFILLER_88_543 VPWR VGND sg13g2_decap_8
XFILLER_1_959 VPWR VGND sg13g2_decap_8
XFILLER_29_11 VPWR VGND sg13g2_decap_8
XFILLER_102_364 VPWR VGND sg13g2_decap_8
XFILLER_0_469 VPWR VGND sg13g2_decap_8
XFILLER_75_259 VPWR VGND sg13g2_decap_8
XFILLER_57_952 VPWR VGND sg13g2_decap_8
XFILLER_29_88 VPWR VGND sg13g2_decap_8
XFILLER_90_207 VPWR VGND sg13g2_decap_8
XFILLER_56_473 VPWR VGND sg13g2_decap_8
XFILLER_45_21 VPWR VGND sg13g2_decap_8
XFILLER_44_613 VPWR VGND sg13g2_decap_8
XFILLER_16_315 VPWR VGND sg13g2_decap_8
XFILLER_17_816 VPWR VGND sg13g2_decap_8
XFILLER_28_175 VPWR VGND sg13g2_decap_8
XFILLER_29_676 VPWR VGND sg13g2_decap_8
XFILLER_83_270 VPWR VGND sg13g2_decap_8
XFILLER_72_966 VPWR VGND sg13g2_decap_8
XFILLER_71_410 VPWR VGND sg13g2_decap_8
XFILLER_43_112 VPWR VGND sg13g2_decap_8
XFILLER_45_98 VPWR VGND sg13g2_decap_8
XFILLER_71_487 VPWR VGND sg13g2_decap_8
XFILLER_43_189 VPWR VGND sg13g2_decap_8
XFILLER_25_882 VPWR VGND sg13g2_decap_8
XFILLER_31_329 VPWR VGND sg13g2_decap_8
XFILLER_61_31 VPWR VGND sg13g2_fill_1
XFILLER_12_543 VPWR VGND sg13g2_decap_8
XFILLER_8_525 VPWR VGND sg13g2_decap_8
XFILLER_40_896 VPWR VGND sg13g2_decap_8
XFILLER_99_819 VPWR VGND sg13g2_decap_8
XFILLER_4_742 VPWR VGND sg13g2_decap_8
XFILLER_3_252 VPWR VGND sg13g2_decap_8
XFILLER_79_543 VPWR VGND sg13g2_decap_8
XFILLER_6_1008 VPWR VGND sg13g2_decap_8
XFILLER_67_749 VPWR VGND sg13g2_decap_8
XFILLER_94_546 VPWR VGND sg13g2_decap_8
XFILLER_66_237 VPWR VGND sg13g2_decap_8
XFILLER_48_952 VPWR VGND sg13g2_decap_8
XFILLER_81_207 VPWR VGND sg13g2_decap_8
XFILLER_47_462 VPWR VGND sg13g2_decap_8
XFILLER_35_602 VPWR VGND sg13g2_decap_8
XFILLER_74_281 VPWR VGND sg13g2_decap_8
XFILLER_63_966 VPWR VGND sg13g2_decap_8
XFILLER_19_175 VPWR VGND sg13g2_decap_8
XFILLER_34_123 VPWR VGND sg13g2_decap_8
XFILLER_90_774 VPWR VGND sg13g2_decap_8
XFILLER_62_476 VPWR VGND sg13g2_decap_8
XFILLER_50_616 VPWR VGND sg13g2_decap_8
XFILLER_23_819 VPWR VGND sg13g2_decap_8
XFILLER_35_679 VPWR VGND sg13g2_decap_8
XFILLER_16_882 VPWR VGND sg13g2_decap_8
XFILLER_31_896 VPWR VGND sg13g2_decap_8
XFILLER_89_329 VPWR VGND sg13g2_decap_8
XFILLER_98_830 VPWR VGND sg13g2_decap_8
XFILLER_106_49 VPWR VGND sg13g2_decap_8
XFILLER_58_749 VPWR VGND sg13g2_decap_8
XFILLER_100_868 VPWR VGND sg13g2_decap_8
XFILLER_85_546 VPWR VGND sg13g2_decap_8
XFILLER_57_259 VPWR VGND sg13g2_decap_8
XFILLER_39_963 VPWR VGND sg13g2_decap_8
XFILLER_54_900 VPWR VGND sg13g2_decap_8
XFILLER_26_602 VPWR VGND sg13g2_decap_8
XFILLER_38_462 VPWR VGND sg13g2_decap_8
XFILLER_25_112 VPWR VGND sg13g2_decap_8
XFILLER_81_774 VPWR VGND sg13g2_decap_8
XFILLER_54_977 VPWR VGND sg13g2_decap_8
XFILLER_53_476 VPWR VGND sg13g2_decap_8
XFILLER_41_616 VPWR VGND sg13g2_decap_8
XFILLER_14_819 VPWR VGND sg13g2_decap_8
XFILLER_26_679 VPWR VGND sg13g2_decap_8
XFILLER_90_1012 VPWR VGND sg13g2_decap_8
XFILLER_80_273 VPWR VGND sg13g2_decap_8
XFILLER_13_329 VPWR VGND sg13g2_decap_8
XFILLER_15_46 VPWR VGND sg13g2_decap_8
XFILLER_25_189 VPWR VGND sg13g2_decap_8
XFILLER_40_126 VPWR VGND sg13g2_decap_8
XFILLER_22_830 VPWR VGND sg13g2_decap_8
XFILLER_34_690 VPWR VGND sg13g2_decap_8
XFILLER_31_56 VPWR VGND sg13g2_decap_8
Xoutput23 net23 uo_out[6] VPWR VGND sg13g2_buf_1
XFILLER_103_651 VPWR VGND sg13g2_decap_8
XFILLER_88_340 VPWR VGND sg13g2_decap_8
XFILLER_1_756 VPWR VGND sg13g2_decap_8
XFILLER_102_161 VPWR VGND sg13g2_decap_8
XFILLER_89_896 VPWR VGND sg13g2_decap_8
XFILLER_0_266 VPWR VGND sg13g2_decap_8
XFILLER_76_557 VPWR VGND sg13g2_decap_8
XFILLER_48_259 VPWR VGND sg13g2_decap_8
XFILLER_56_53 VPWR VGND sg13g2_decap_8
XFILLER_17_613 VPWR VGND sg13g2_decap_8
XFILLER_29_473 VPWR VGND sg13g2_decap_8
XFILLER_56_270 VPWR VGND sg13g2_decap_8
XFILLER_44_410 VPWR VGND sg13g2_decap_8
XFILLER_16_112 VPWR VGND sg13g2_decap_8
XFILLER_72_763 VPWR VGND sg13g2_decap_8
XFILLER_60_914 VPWR VGND sg13g2_decap_8
XFILLER_45_966 VPWR VGND sg13g2_decap_8
XFILLER_71_284 VPWR VGND sg13g2_decap_8
XFILLER_44_487 VPWR VGND sg13g2_decap_8
XFILLER_16_189 VPWR VGND sg13g2_decap_8
XFILLER_32_627 VPWR VGND sg13g2_decap_8
XFILLER_72_63 VPWR VGND sg13g2_decap_8
XFILLER_31_126 VPWR VGND sg13g2_decap_8
XFILLER_9_812 VPWR VGND sg13g2_decap_8
XFILLER_12_340 VPWR VGND sg13g2_decap_8
XFILLER_13_896 VPWR VGND sg13g2_decap_8
XFILLER_8_322 VPWR VGND sg13g2_decap_8
XFILLER_40_693 VPWR VGND sg13g2_decap_8
XFILLER_9_889 VPWR VGND sg13g2_decap_8
XFILLER_8_399 VPWR VGND sg13g2_decap_8
XFILLER_99_616 VPWR VGND sg13g2_decap_8
XFILLER_98_137 VPWR VGND sg13g2_decap_8
XFILLER_79_340 VPWR VGND sg13g2_decap_8
XFILLER_95_844 VPWR VGND sg13g2_decap_8
XFILLER_94_343 VPWR VGND sg13g2_decap_8
XFILLER_67_546 VPWR VGND sg13g2_decap_8
XFILLER_54_207 VPWR VGND sg13g2_decap_8
XFILLER_63_763 VPWR VGND sg13g2_decap_8
XFILLER_51_914 VPWR VGND sg13g2_decap_8
XFILLER_36_966 VPWR VGND sg13g2_decap_8
XFILLER_90_571 VPWR VGND sg13g2_decap_8
XFILLER_62_273 VPWR VGND sg13g2_decap_8
XFILLER_50_413 VPWR VGND sg13g2_decap_8
XFILLER_23_616 VPWR VGND sg13g2_decap_8
XFILLER_35_476 VPWR VGND sg13g2_decap_8
XFILLER_94_0 VPWR VGND sg13g2_decap_8
XFILLER_22_137 VPWR VGND sg13g2_decap_8
XFILLER_31_693 VPWR VGND sg13g2_decap_8
XFILLER_105_938 VPWR VGND sg13g2_decap_8
XFILLER_89_126 VPWR VGND sg13g2_decap_8
XFILLER_104_448 VPWR VGND sg13g2_decap_8
XFILLER_86_844 VPWR VGND sg13g2_decap_8
XFILLER_85_343 VPWR VGND sg13g2_decap_8
XFILLER_58_546 VPWR VGND sg13g2_decap_8
XFILLER_100_665 VPWR VGND sg13g2_decap_8
XFILLER_27_900 VPWR VGND sg13g2_decap_8
XFILLER_39_760 VPWR VGND sg13g2_decap_8
XFILLER_54_774 VPWR VGND sg13g2_decap_8
XFILLER_42_914 VPWR VGND sg13g2_decap_8
XFILLER_26_56 VPWR VGND sg13g2_decap_8
XFILLER_27_977 VPWR VGND sg13g2_decap_8
XFILLER_81_571 VPWR VGND sg13g2_decap_8
XFILLER_53_273 VPWR VGND sg13g2_decap_8
XFILLER_14_616 VPWR VGND sg13g2_decap_8
XFILLER_26_476 VPWR VGND sg13g2_decap_8
XFILLER_41_413 VPWR VGND sg13g2_decap_8
XFILLER_42_11 VPWR VGND sg13g2_decap_8
XFILLER_13_126 VPWR VGND sg13g2_decap_8
XFILLER_50_980 VPWR VGND sg13g2_decap_8
XFILLER_9_119 VPWR VGND sg13g2_decap_8
XFILLER_10_844 VPWR VGND sg13g2_decap_8
XFILLER_42_88 VPWR VGND sg13g2_decap_8
XFILLER_6_826 VPWR VGND sg13g2_decap_8
XFILLER_5_347 VPWR VGND sg13g2_decap_8
XFILLER_1_553 VPWR VGND sg13g2_decap_8
XFILLER_89_693 VPWR VGND sg13g2_decap_8
XFILLER_77_833 VPWR VGND sg13g2_decap_8
XFILLER_3_49 VPWR VGND sg13g2_decap_8
XFILLER_49_557 VPWR VGND sg13g2_decap_8
XFILLER_76_354 VPWR VGND sg13g2_decap_8
XFILLER_92_847 VPWR VGND sg13g2_decap_8
XFILLER_17_410 VPWR VGND sg13g2_decap_8
XFILLER_29_270 VPWR VGND sg13g2_decap_8
XFILLER_91_357 VPWR VGND sg13g2_decap_8
XFILLER_45_763 VPWR VGND sg13g2_decap_8
XFILLER_18_966 VPWR VGND sg13g2_decap_8
XFILLER_33_903 VPWR VGND sg13g2_decap_8
XFILLER_83_95 VPWR VGND sg13g2_decap_8
XFILLER_72_560 VPWR VGND sg13g2_decap_8
XFILLER_60_711 VPWR VGND sg13g2_decap_8
XFILLER_17_487 VPWR VGND sg13g2_decap_8
XFILLER_32_424 VPWR VGND sg13g2_decap_8
XFILLER_44_284 VPWR VGND sg13g2_decap_8
XFILLER_60_788 VPWR VGND sg13g2_decap_8
XFILLER_41_980 VPWR VGND sg13g2_decap_8
XFILLER_13_693 VPWR VGND sg13g2_decap_8
XFILLER_40_490 VPWR VGND sg13g2_decap_8
XFILLER_9_686 VPWR VGND sg13g2_decap_8
XFILLER_66_4 VPWR VGND sg13g2_decap_8
XFILLER_8_196 VPWR VGND sg13g2_decap_8
XFILLER_99_413 VPWR VGND sg13g2_decap_8
XFILLER_80_1022 VPWR VGND sg13g2_decap_8
XFILLER_95_641 VPWR VGND sg13g2_decap_8
XFILLER_68_866 VPWR VGND sg13g2_decap_8
XFILLER_67_343 VPWR VGND sg13g2_decap_8
XFILLER_94_140 VPWR VGND sg13g2_decap_8
XFILLER_27_207 VPWR VGND sg13g2_decap_8
XFILLER_103_28 VPWR VGND sg13g2_decap_8
XFILLER_83_858 VPWR VGND sg13g2_decap_8
XFILLER_82_357 VPWR VGND sg13g2_decap_8
XFILLER_36_763 VPWR VGND sg13g2_decap_8
XFILLER_63_560 VPWR VGND sg13g2_decap_8
XFILLER_51_711 VPWR VGND sg13g2_decap_8
XFILLER_23_413 VPWR VGND sg13g2_decap_8
XFILLER_24_914 VPWR VGND sg13g2_decap_8
XFILLER_35_273 VPWR VGND sg13g2_decap_8
XFILLER_50_210 VPWR VGND sg13g2_decap_8
XFILLER_51_788 VPWR VGND sg13g2_decap_8
XFILLER_50_287 VPWR VGND sg13g2_decap_8
XFILLER_32_991 VPWR VGND sg13g2_decap_8
XFILLER_12_25 VPWR VGND sg13g2_decap_8
XFILLER_31_490 VPWR VGND sg13g2_decap_8
XFILLER_88_18 VPWR VGND sg13g2_decap_8
XFILLER_105_735 VPWR VGND sg13g2_decap_8
XFILLER_104_245 VPWR VGND sg13g2_decap_8
XFILLER_78_608 VPWR VGND sg13g2_decap_8
XFILLER_99_980 VPWR VGND sg13g2_decap_8
XFILLER_101_952 VPWR VGND sg13g2_decap_8
XFILLER_86_641 VPWR VGND sg13g2_decap_8
XFILLER_59_866 VPWR VGND sg13g2_decap_8
XFILLER_100_462 VPWR VGND sg13g2_decap_8
XFILLER_85_140 VPWR VGND sg13g2_decap_8
XFILLER_58_343 VPWR VGND sg13g2_decap_8
XFILLER_37_11 VPWR VGND sg13g2_decap_8
XFILLER_74_869 VPWR VGND sg13g2_decap_8
XFILLER_73_368 VPWR VGND sg13g2_decap_8
XFILLER_61_508 VPWR VGND sg13g2_decap_8
XFILLER_37_88 VPWR VGND sg13g2_decap_8
XFILLER_54_571 VPWR VGND sg13g2_decap_8
XFILLER_42_711 VPWR VGND sg13g2_decap_8
XFILLER_14_413 VPWR VGND sg13g2_decap_8
XFILLER_15_914 VPWR VGND sg13g2_decap_8
XFILLER_26_273 VPWR VGND sg13g2_decap_8
XFILLER_27_774 VPWR VGND sg13g2_decap_8
XFILLER_53_21 VPWR VGND sg13g2_decap_8
XFILLER_18_1008 VPWR VGND sg13g2_decap_8
XFILLER_41_210 VPWR VGND sg13g2_decap_8
XFILLER_42_788 VPWR VGND sg13g2_decap_8
XFILLER_30_917 VPWR VGND sg13g2_decap_8
XFILLER_53_98 VPWR VGND sg13g2_decap_8
XFILLER_23_980 VPWR VGND sg13g2_decap_8
XFILLER_41_287 VPWR VGND sg13g2_decap_8
XFILLER_10_641 VPWR VGND sg13g2_decap_8
XFILLER_6_623 VPWR VGND sg13g2_decap_8
XFILLER_5_144 VPWR VGND sg13g2_decap_8
XFILLER_97_917 VPWR VGND sg13g2_decap_8
XFILLER_64_1028 VPWR VGND sg13g2_fill_1
XFILLER_2_851 VPWR VGND sg13g2_decap_8
XFILLER_96_427 VPWR VGND sg13g2_decap_8
XFILLER_1_350 VPWR VGND sg13g2_decap_8
XFILLER_89_490 VPWR VGND sg13g2_decap_8
XFILLER_77_630 VPWR VGND sg13g2_decap_8
XFILLER_76_151 VPWR VGND sg13g2_decap_8
X_62_ _24_ VPWR _27_ VGND _23_ _25_ sg13g2_o21ai_1
XFILLER_49_354 VPWR VGND sg13g2_decap_8
XFILLER_92_644 VPWR VGND sg13g2_decap_8
XFILLER_65_847 VPWR VGND sg13g2_decap_8
XFILLER_91_154 VPWR VGND sg13g2_decap_8
XFILLER_64_368 VPWR VGND sg13g2_decap_8
XFILLER_18_763 VPWR VGND sg13g2_decap_8
XFILLER_45_560 VPWR VGND sg13g2_decap_8
XFILLER_33_700 VPWR VGND sg13g2_decap_8
XFILLER_17_284 VPWR VGND sg13g2_decap_8
XFILLER_32_221 VPWR VGND sg13g2_decap_8
XFILLER_21_917 VPWR VGND sg13g2_decap_8
XFILLER_33_777 VPWR VGND sg13g2_decap_8
XFILLER_60_585 VPWR VGND sg13g2_decap_8
XFILLER_14_980 VPWR VGND sg13g2_decap_8
XFILLER_20_438 VPWR VGND sg13g2_decap_8
XFILLER_32_298 VPWR VGND sg13g2_decap_8
XFILLER_13_490 VPWR VGND sg13g2_decap_8
XFILLER_9_483 VPWR VGND sg13g2_decap_8
XFILLER_99_210 VPWR VGND sg13g2_decap_8
XFILLER_57_0 VPWR VGND sg13g2_decap_8
XFILLER_99_287 VPWR VGND sg13g2_decap_8
XFILLER_88_928 VPWR VGND sg13g2_decap_8
XFILLER_87_427 VPWR VGND sg13g2_decap_8
XFILLER_4_70 VPWR VGND sg13g2_decap_8
XFILLER_102_749 VPWR VGND sg13g2_decap_8
XFILLER_101_259 VPWR VGND sg13g2_decap_8
XFILLER_68_663 VPWR VGND sg13g2_decap_8
XFILLER_67_140 VPWR VGND sg13g2_decap_8
XFILLER_96_994 VPWR VGND sg13g2_decap_8
XFILLER_56_858 VPWR VGND sg13g2_decap_8
XFILLER_83_655 VPWR VGND sg13g2_decap_8
XFILLER_55_357 VPWR VGND sg13g2_decap_8
XFILLER_82_154 VPWR VGND sg13g2_decap_8
XFILLER_24_711 VPWR VGND sg13g2_decap_8
XFILLER_36_560 VPWR VGND sg13g2_decap_8
XFILLER_23_210 VPWR VGND sg13g2_decap_8
XFILLER_12_928 VPWR VGND sg13g2_decap_8
XFILLER_24_788 VPWR VGND sg13g2_decap_8
XFILLER_51_585 VPWR VGND sg13g2_decap_8
XFILLER_11_427 VPWR VGND sg13g2_decap_8
XFILLER_23_35 VPWR VGND sg13g2_decap_8
XFILLER_23_287 VPWR VGND sg13g2_decap_8
XFILLER_104_1022 VPWR VGND sg13g2_decap_8
XFILLER_99_28 VPWR VGND sg13g2_decap_8
XFILLER_3_637 VPWR VGND sg13g2_decap_8
XFILLER_105_532 VPWR VGND sg13g2_decap_8
XFILLER_79_928 VPWR VGND sg13g2_decap_8
XFILLER_78_405 VPWR VGND sg13g2_decap_8
XFILLER_2_158 VPWR VGND sg13g2_decap_8
XFILLER_48_21 VPWR VGND sg13g2_decap_8
XFILLER_24_1012 VPWR VGND sg13g2_decap_8
XFILLER_59_663 VPWR VGND sg13g2_decap_8
XFILLER_87_994 VPWR VGND sg13g2_decap_8
XFILLER_47_847 VPWR VGND sg13g2_decap_8
XFILLER_48_98 VPWR VGND sg13g2_decap_8
XFILLER_74_666 VPWR VGND sg13g2_decap_8
XFILLER_0_28 VPWR VGND sg13g2_decap_8
XFILLER_34_508 VPWR VGND sg13g2_decap_8
XFILLER_73_165 VPWR VGND sg13g2_decap_8
XFILLER_64_53 VPWR VGND sg13g2_decap_8
XFILLER_61_305 VPWR VGND sg13g2_decap_8
XFILLER_46_368 VPWR VGND sg13g2_decap_8
XFILLER_15_711 VPWR VGND sg13g2_decap_8
XFILLER_27_571 VPWR VGND sg13g2_decap_8
XFILLER_14_210 VPWR VGND sg13g2_decap_8
XFILLER_70_861 VPWR VGND sg13g2_decap_8
XFILLER_15_788 VPWR VGND sg13g2_decap_8
XFILLER_30_714 VPWR VGND sg13g2_decap_8
XFILLER_42_585 VPWR VGND sg13g2_decap_8
XFILLER_14_287 VPWR VGND sg13g2_decap_8
XFILLER_80_63 VPWR VGND sg13g2_decap_8
XFILLER_7_921 VPWR VGND sg13g2_decap_8
XFILLER_6_420 VPWR VGND sg13g2_decap_8
XFILLER_11_994 VPWR VGND sg13g2_decap_8
XFILLER_50_7 VPWR VGND sg13g2_decap_8
XFILLER_7_998 VPWR VGND sg13g2_decap_8
XFILLER_6_497 VPWR VGND sg13g2_decap_8
XFILLER_97_714 VPWR VGND sg13g2_decap_8
XFILLER_96_224 VPWR VGND sg13g2_decap_8
XFILLER_69_449 VPWR VGND sg13g2_decap_8
XFILLER_78_972 VPWR VGND sg13g2_decap_8
XFILLER_29_4 VPWR VGND sg13g2_decap_8
XFILLER_49_151 VPWR VGND sg13g2_decap_8
XFILLER_38_847 VPWR VGND sg13g2_decap_8
XFILLER_93_964 VPWR VGND sg13g2_decap_8
XFILLER_92_441 VPWR VGND sg13g2_decap_8
XFILLER_65_644 VPWR VGND sg13g2_decap_8
X_45_ _12_ VPWR _13_ VGND _03_ _11_ sg13g2_o21ai_1
XFILLER_64_165 VPWR VGND sg13g2_decap_8
XFILLER_18_560 VPWR VGND sg13g2_decap_8
XFILLER_37_368 VPWR VGND sg13g2_decap_8
XFILLER_80_658 VPWR VGND sg13g2_decap_8
XFILLER_61_872 VPWR VGND sg13g2_decap_8
XFILLER_21_714 VPWR VGND sg13g2_decap_8
XFILLER_60_382 VPWR VGND sg13g2_decap_8
XFILLER_33_574 VPWR VGND sg13g2_decap_8
XFILLER_20_235 VPWR VGND sg13g2_decap_8
XFILLER_9_280 VPWR VGND sg13g2_decap_8
XFILLER_106_329 VPWR VGND sg13g2_decap_8
XFILLER_47_1001 VPWR VGND sg13g2_decap_8
XFILLER_88_725 VPWR VGND sg13g2_decap_8
XFILLER_102_546 VPWR VGND sg13g2_decap_8
XFILLER_87_224 VPWR VGND sg13g2_decap_8
XFILLER_96_791 VPWR VGND sg13g2_decap_8
XFILLER_84_931 VPWR VGND sg13g2_decap_8
XFILLER_68_460 VPWR VGND sg13g2_decap_8
XFILLER_18_35 VPWR VGND sg13g2_decap_8
XFILLER_83_452 VPWR VGND sg13g2_decap_8
XFILLER_56_655 VPWR VGND sg13g2_decap_8
XFILLER_28_357 VPWR VGND sg13g2_decap_8
XFILLER_29_858 VPWR VGND sg13g2_decap_8
XFILLER_55_154 VPWR VGND sg13g2_decap_8
XFILLER_71_669 VPWR VGND sg13g2_decap_8
XFILLER_70_168 VPWR VGND sg13g2_decap_8
XFILLER_54_1005 VPWR VGND sg13g2_decap_8
XFILLER_52_861 VPWR VGND sg13g2_decap_8
XFILLER_51_382 VPWR VGND sg13g2_decap_8
XFILLER_12_725 VPWR VGND sg13g2_decap_8
XFILLER_24_585 VPWR VGND sg13g2_decap_8
XFILLER_34_67 VPWR VGND sg13g2_decap_8
XFILLER_8_707 VPWR VGND sg13g2_decap_8
XFILLER_11_224 VPWR VGND sg13g2_decap_8
XFILLER_7_228 VPWR VGND sg13g2_decap_8
XFILLER_50_77 VPWR VGND sg13g2_decap_8
XFILLER_4_924 VPWR VGND sg13g2_decap_8
XFILLER_3_434 VPWR VGND sg13g2_decap_8
XFILLER_79_725 VPWR VGND sg13g2_decap_8
XFILLER_78_202 VPWR VGND sg13g2_decap_8
XFILLER_106_896 VPWR VGND sg13g2_decap_8
XFILLER_59_53 VPWR VGND sg13g2_decap_8
XFILLER_94_728 VPWR VGND sg13g2_decap_8
XFILLER_66_419 VPWR VGND sg13g2_decap_8
XFILLER_87_791 VPWR VGND sg13g2_decap_8
XFILLER_78_279 VPWR VGND sg13g2_decap_8
XFILLER_75_931 VPWR VGND sg13g2_decap_8
XFILLER_59_460 VPWR VGND sg13g2_decap_8
XFILLER_75_63 VPWR VGND sg13g2_decap_8
XFILLER_47_644 VPWR VGND sg13g2_decap_8
XFILLER_19_357 VPWR VGND sg13g2_decap_8
XFILLER_74_463 VPWR VGND sg13g2_decap_8
XFILLER_46_165 VPWR VGND sg13g2_decap_8
XFILLER_34_305 VPWR VGND sg13g2_decap_8
XFILLER_90_956 VPWR VGND sg13g2_decap_8
XFILLER_62_658 VPWR VGND sg13g2_decap_8
XFILLER_61_102 VPWR VGND sg13g2_decap_8
XFILLER_43_861 VPWR VGND sg13g2_decap_8
XFILLER_91_84 VPWR VGND sg13g2_decap_8
XFILLER_61_179 VPWR VGND sg13g2_decap_8
XFILLER_42_382 VPWR VGND sg13g2_decap_8
XFILLER_15_585 VPWR VGND sg13g2_decap_8
XFILLER_30_511 VPWR VGND sg13g2_decap_8
XFILLER_30_588 VPWR VGND sg13g2_decap_8
XFILLER_11_791 VPWR VGND sg13g2_decap_8
XFILLER_7_795 VPWR VGND sg13g2_decap_8
XFILLER_6_294 VPWR VGND sg13g2_decap_8
XFILLER_97_511 VPWR VGND sg13g2_decap_8
XFILLER_69_246 VPWR VGND sg13g2_decap_8
XFILLER_97_588 VPWR VGND sg13g2_decap_8
XFILLER_85_728 VPWR VGND sg13g2_decap_8
XFILLER_84_238 VPWR VGND sg13g2_decap_8
XFILLER_65_441 VPWR VGND sg13g2_decap_8
XFILLER_38_644 VPWR VGND sg13g2_decap_8
XFILLER_93_761 VPWR VGND sg13g2_decap_8
XFILLER_66_986 VPWR VGND sg13g2_decap_8
XFILLER_37_165 VPWR VGND sg13g2_decap_8
XFILLER_81_956 VPWR VGND sg13g2_decap_8
XFILLER_53_658 VPWR VGND sg13g2_decap_8
XFILLER_80_455 VPWR VGND sg13g2_decap_8
XFILLER_52_168 VPWR VGND sg13g2_decap_8
XFILLER_34_872 VPWR VGND sg13g2_decap_8
XFILLER_40_308 VPWR VGND sg13g2_decap_8
XFILLER_21_511 VPWR VGND sg13g2_decap_8
XFILLER_33_371 VPWR VGND sg13g2_decap_8
XFILLER_14_1022 VPWR VGND sg13g2_decap_8
XFILLER_21_588 VPWR VGND sg13g2_decap_8
XFILLER_20_25 VPWR VGND sg13g2_decap_8
XFILLER_106_126 VPWR VGND sg13g2_decap_8
XFILLER_103_833 VPWR VGND sg13g2_decap_8
XFILLER_88_522 VPWR VGND sg13g2_decap_8
XFILLER_1_938 VPWR VGND sg13g2_decap_8
XFILLER_102_343 VPWR VGND sg13g2_decap_8
XFILLER_0_448 VPWR VGND sg13g2_decap_8
XFILLER_88_599 VPWR VGND sg13g2_decap_8
XFILLER_76_739 VPWR VGND sg13g2_decap_8
XFILLER_57_931 VPWR VGND sg13g2_decap_8
XFILLER_29_67 VPWR VGND sg13g2_decap_8
XFILLER_75_238 VPWR VGND sg13g2_decap_8
XFILLER_21_1015 VPWR VGND sg13g2_decap_8
XFILLER_29_655 VPWR VGND sg13g2_decap_8
XFILLER_56_452 VPWR VGND sg13g2_decap_8
XFILLER_28_154 VPWR VGND sg13g2_decap_8
XFILLER_72_945 VPWR VGND sg13g2_decap_8
XFILLER_71_466 VPWR VGND sg13g2_decap_8
XFILLER_45_77 VPWR VGND sg13g2_decap_8
XFILLER_44_669 VPWR VGND sg13g2_decap_8
XFILLER_43_168 VPWR VGND sg13g2_decap_8
XFILLER_25_861 VPWR VGND sg13g2_decap_8
XFILLER_31_308 VPWR VGND sg13g2_decap_8
XFILLER_32_809 VPWR VGND sg13g2_decap_8
XFILLER_8_504 VPWR VGND sg13g2_decap_8
XFILLER_12_522 VPWR VGND sg13g2_decap_8
XFILLER_24_382 VPWR VGND sg13g2_decap_8
XFILLER_40_875 VPWR VGND sg13g2_decap_8
XFILLER_12_599 VPWR VGND sg13g2_decap_8
XFILLER_6_49 VPWR VGND sg13g2_decap_8
XFILLER_4_721 VPWR VGND sg13g2_decap_8
XFILLER_98_319 VPWR VGND sg13g2_decap_8
XFILLER_3_231 VPWR VGND sg13g2_decap_8
XFILLER_106_693 VPWR VGND sg13g2_decap_8
XFILLER_79_522 VPWR VGND sg13g2_decap_8
XFILLER_4_798 VPWR VGND sg13g2_decap_8
XFILLER_94_525 VPWR VGND sg13g2_decap_8
XFILLER_79_599 VPWR VGND sg13g2_decap_8
XFILLER_67_728 VPWR VGND sg13g2_decap_8
XFILLER_66_216 VPWR VGND sg13g2_decap_8
XFILLER_48_931 VPWR VGND sg13g2_decap_8
XFILLER_86_95 VPWR VGND sg13g2_decap_8
XFILLER_47_441 VPWR VGND sg13g2_decap_8
XFILLER_13_7 VPWR VGND sg13g2_decap_8
XFILLER_74_260 VPWR VGND sg13g2_decap_8
XFILLER_19_154 VPWR VGND sg13g2_decap_8
XFILLER_63_945 VPWR VGND sg13g2_decap_8
XFILLER_34_102 VPWR VGND sg13g2_decap_8
XFILLER_90_753 VPWR VGND sg13g2_decap_8
XFILLER_62_455 VPWR VGND sg13g2_decap_8
XFILLER_16_861 VPWR VGND sg13g2_decap_8
XFILLER_35_658 VPWR VGND sg13g2_decap_8
XFILLER_22_319 VPWR VGND sg13g2_decap_8
XFILLER_34_179 VPWR VGND sg13g2_decap_8
XFILLER_15_382 VPWR VGND sg13g2_decap_8
XFILLER_31_875 VPWR VGND sg13g2_decap_8
XFILLER_30_385 VPWR VGND sg13g2_decap_8
XFILLER_7_592 VPWR VGND sg13g2_decap_8
XFILLER_89_308 VPWR VGND sg13g2_decap_8
XFILLER_106_28 VPWR VGND sg13g2_decap_8
XFILLER_44_1026 VPWR VGND sg13g2_fill_2
XFILLER_98_886 VPWR VGND sg13g2_decap_8
XFILLER_97_385 VPWR VGND sg13g2_decap_8
XFILLER_85_525 VPWR VGND sg13g2_decap_8
XFILLER_58_728 VPWR VGND sg13g2_decap_8
XFILLER_100_847 VPWR VGND sg13g2_decap_8
XFILLER_57_238 VPWR VGND sg13g2_decap_8
XFILLER_39_942 VPWR VGND sg13g2_decap_8
XFILLER_66_783 VPWR VGND sg13g2_decap_8
XFILLER_38_441 VPWR VGND sg13g2_decap_8
XFILLER_54_956 VPWR VGND sg13g2_decap_8
XFILLER_81_753 VPWR VGND sg13g2_decap_8
XFILLER_80_252 VPWR VGND sg13g2_decap_8
XFILLER_53_455 VPWR VGND sg13g2_decap_8
XFILLER_26_658 VPWR VGND sg13g2_decap_8
XFILLER_13_308 VPWR VGND sg13g2_decap_8
XFILLER_15_25 VPWR VGND sg13g2_decap_8
XFILLER_25_168 VPWR VGND sg13g2_decap_8
XFILLER_40_105 VPWR VGND sg13g2_decap_8
XFILLER_51_1019 VPWR VGND sg13g2_decap_8
XFILLER_22_886 VPWR VGND sg13g2_decap_8
XFILLER_21_385 VPWR VGND sg13g2_decap_8
XFILLER_31_35 VPWR VGND sg13g2_decap_8
XFILLER_5_529 VPWR VGND sg13g2_decap_8
Xoutput24 net24 uo_out[7] VPWR VGND sg13g2_buf_1
XFILLER_1_735 VPWR VGND sg13g2_decap_8
XFILLER_103_630 VPWR VGND sg13g2_decap_8
XFILLER_89_875 VPWR VGND sg13g2_decap_8
XFILLER_0_245 VPWR VGND sg13g2_decap_8
XFILLER_102_140 VPWR VGND sg13g2_decap_8
XFILLER_49_739 VPWR VGND sg13g2_decap_8
XFILLER_88_396 VPWR VGND sg13g2_decap_8
XFILLER_76_536 VPWR VGND sg13g2_decap_8
XFILLER_56_32 VPWR VGND sg13g2_decap_8
XFILLER_48_238 VPWR VGND sg13g2_decap_8
XFILLER_29_452 VPWR VGND sg13g2_decap_8
XFILLER_91_539 VPWR VGND sg13g2_decap_8
XFILLER_45_945 VPWR VGND sg13g2_decap_8
XFILLER_72_742 VPWR VGND sg13g2_decap_8
XFILLER_44_466 VPWR VGND sg13g2_decap_8
XFILLER_17_669 VPWR VGND sg13g2_decap_8
XFILLER_32_606 VPWR VGND sg13g2_decap_8
XFILLER_72_42 VPWR VGND sg13g2_decap_8
XFILLER_71_263 VPWR VGND sg13g2_decap_8
XFILLER_16_168 VPWR VGND sg13g2_decap_8
XFILLER_31_105 VPWR VGND sg13g2_decap_8
XFILLER_8_301 VPWR VGND sg13g2_decap_8
XFILLER_13_875 VPWR VGND sg13g2_decap_8
XFILLER_40_672 VPWR VGND sg13g2_decap_8
XFILLER_9_868 VPWR VGND sg13g2_decap_8
XFILLER_12_396 VPWR VGND sg13g2_decap_8
XFILLER_8_378 VPWR VGND sg13g2_decap_8
XFILLER_67_1015 VPWR VGND sg13g2_decap_8
XFILLER_98_116 VPWR VGND sg13g2_decap_8
XFILLER_4_595 VPWR VGND sg13g2_decap_8
XFILLER_106_490 VPWR VGND sg13g2_decap_8
XFILLER_95_823 VPWR VGND sg13g2_decap_8
XFILLER_67_525 VPWR VGND sg13g2_decap_8
XFILLER_94_322 VPWR VGND sg13g2_decap_8
XFILLER_79_396 VPWR VGND sg13g2_decap_8
XFILLER_39_249 VPWR VGND sg13g2_decap_8
XFILLER_94_399 VPWR VGND sg13g2_decap_8
XFILLER_82_539 VPWR VGND sg13g2_decap_8
XFILLER_36_945 VPWR VGND sg13g2_decap_8
XFILLER_90_550 VPWR VGND sg13g2_decap_8
XFILLER_63_742 VPWR VGND sg13g2_decap_8
XFILLER_35_455 VPWR VGND sg13g2_decap_8
XFILLER_62_252 VPWR VGND sg13g2_decap_8
XFILLER_22_116 VPWR VGND sg13g2_decap_8
XFILLER_87_0 VPWR VGND sg13g2_decap_8
XFILLER_50_469 VPWR VGND sg13g2_decap_8
XFILLER_31_672 VPWR VGND sg13g2_decap_8
XFILLER_30_182 VPWR VGND sg13g2_decap_8
XFILLER_7_81 VPWR VGND sg13g2_decap_8
XFILLER_105_917 VPWR VGND sg13g2_decap_8
XFILLER_104_427 VPWR VGND sg13g2_decap_8
XFILLER_89_105 VPWR VGND sg13g2_decap_8
XFILLER_98_683 VPWR VGND sg13g2_decap_8
XFILLER_86_823 VPWR VGND sg13g2_decap_8
XFILLER_58_525 VPWR VGND sg13g2_decap_8
XFILLER_100_644 VPWR VGND sg13g2_decap_8
XFILLER_97_182 VPWR VGND sg13g2_decap_8
XFILLER_85_322 VPWR VGND sg13g2_decap_8
XFILLER_93_19 VPWR VGND sg13g2_decap_8
XFILLER_85_399 VPWR VGND sg13g2_decap_8
XFILLER_66_580 VPWR VGND sg13g2_decap_8
XFILLER_81_550 VPWR VGND sg13g2_decap_8
XFILLER_54_753 VPWR VGND sg13g2_decap_8
XFILLER_26_35 VPWR VGND sg13g2_decap_8
XFILLER_26_455 VPWR VGND sg13g2_decap_8
XFILLER_27_956 VPWR VGND sg13g2_decap_8
XFILLER_53_252 VPWR VGND sg13g2_decap_8
XFILLER_13_105 VPWR VGND sg13g2_decap_8
XFILLER_41_469 VPWR VGND sg13g2_decap_8
XFILLER_42_67 VPWR VGND sg13g2_decap_8
XFILLER_10_823 VPWR VGND sg13g2_decap_8
XFILLER_22_683 VPWR VGND sg13g2_decap_8
XFILLER_6_805 VPWR VGND sg13g2_decap_8
XFILLER_21_182 VPWR VGND sg13g2_decap_8
XFILLER_5_326 VPWR VGND sg13g2_decap_8
XFILLER_96_609 VPWR VGND sg13g2_decap_8
XFILLER_3_28 VPWR VGND sg13g2_decap_8
XFILLER_1_532 VPWR VGND sg13g2_decap_8
XFILLER_104_994 VPWR VGND sg13g2_decap_8
XFILLER_89_672 VPWR VGND sg13g2_decap_8
XFILLER_77_812 VPWR VGND sg13g2_decap_8
XFILLER_67_31 VPWR VGND sg13g2_fill_2
XFILLER_88_193 VPWR VGND sg13g2_decap_8
XFILLER_76_333 VPWR VGND sg13g2_decap_8
XFILLER_49_536 VPWR VGND sg13g2_decap_8
XFILLER_97_1008 VPWR VGND sg13g2_decap_8
XFILLER_92_826 VPWR VGND sg13g2_decap_8
XFILLER_77_889 VPWR VGND sg13g2_decap_8
XFILLER_91_336 VPWR VGND sg13g2_decap_8
XFILLER_18_945 VPWR VGND sg13g2_decap_8
XFILLER_45_742 VPWR VGND sg13g2_decap_8
XFILLER_83_74 VPWR VGND sg13g2_decap_8
XFILLER_44_263 VPWR VGND sg13g2_decap_8
XFILLER_17_466 VPWR VGND sg13g2_decap_8
XFILLER_32_403 VPWR VGND sg13g2_decap_8
XFILLER_33_959 VPWR VGND sg13g2_decap_8
XFILLER_60_767 VPWR VGND sg13g2_decap_8
XFILLER_80_7 VPWR VGND sg13g2_decap_8
XFILLER_13_672 VPWR VGND sg13g2_decap_8
XFILLER_9_665 VPWR VGND sg13g2_decap_8
XFILLER_12_193 VPWR VGND sg13g2_decap_8
XFILLER_8_175 VPWR VGND sg13g2_decap_8
XFILLER_59_4 VPWR VGND sg13g2_decap_8
XFILLER_5_893 VPWR VGND sg13g2_decap_8
XFILLER_99_469 VPWR VGND sg13g2_decap_8
XFILLER_87_609 VPWR VGND sg13g2_decap_8
XFILLER_4_392 VPWR VGND sg13g2_decap_8
XFILLER_80_1001 VPWR VGND sg13g2_decap_8
XFILLER_95_620 VPWR VGND sg13g2_decap_8
XFILLER_79_193 VPWR VGND sg13g2_decap_8
XFILLER_68_845 VPWR VGND sg13g2_decap_8
XFILLER_67_322 VPWR VGND sg13g2_decap_8
XFILLER_95_697 VPWR VGND sg13g2_decap_8
XFILLER_83_837 VPWR VGND sg13g2_decap_8
XFILLER_82_336 VPWR VGND sg13g2_decap_8
XFILLER_67_399 VPWR VGND sg13g2_decap_8
XFILLER_55_539 VPWR VGND sg13g2_decap_8
XFILLER_94_196 VPWR VGND sg13g2_decap_8
XFILLER_36_742 VPWR VGND sg13g2_decap_8
XFILLER_35_252 VPWR VGND sg13g2_decap_8
XFILLER_51_767 VPWR VGND sg13g2_decap_8
XFILLER_50_266 VPWR VGND sg13g2_decap_8
XFILLER_11_609 VPWR VGND sg13g2_decap_8
XFILLER_23_469 VPWR VGND sg13g2_decap_8
XFILLER_32_970 VPWR VGND sg13g2_decap_8
XFILLER_3_819 VPWR VGND sg13g2_decap_8
XFILLER_105_714 VPWR VGND sg13g2_decap_8
XFILLER_104_224 VPWR VGND sg13g2_decap_8
XFILLER_77_119 VPWR VGND sg13g2_decap_8
XFILLER_101_931 VPWR VGND sg13g2_decap_8
XFILLER_98_480 VPWR VGND sg13g2_decap_8
XFILLER_86_620 VPWR VGND sg13g2_decap_8
XFILLER_59_845 VPWR VGND sg13g2_decap_8
XFILLER_58_322 VPWR VGND sg13g2_decap_8
XFILLER_100_441 VPWR VGND sg13g2_decap_8
XFILLER_86_697 VPWR VGND sg13g2_decap_8
XFILLER_74_848 VPWR VGND sg13g2_decap_8
XFILLER_58_399 VPWR VGND sg13g2_decap_8
XFILLER_2_1012 VPWR VGND sg13g2_decap_8
XFILLER_37_67 VPWR VGND sg13g2_decap_8
XFILLER_85_196 VPWR VGND sg13g2_decap_8
XFILLER_73_347 VPWR VGND sg13g2_decap_8
XFILLER_27_753 VPWR VGND sg13g2_decap_8
XFILLER_54_550 VPWR VGND sg13g2_decap_8
XFILLER_26_252 VPWR VGND sg13g2_decap_8
XFILLER_53_77 VPWR VGND sg13g2_decap_8
XFILLER_42_767 VPWR VGND sg13g2_decap_8
XFILLER_14_469 VPWR VGND sg13g2_decap_8
XFILLER_41_266 VPWR VGND sg13g2_decap_8
XFILLER_10_620 VPWR VGND sg13g2_decap_8
XFILLER_22_480 VPWR VGND sg13g2_decap_8
XFILLER_6_602 VPWR VGND sg13g2_decap_8
XFILLER_10_697 VPWR VGND sg13g2_decap_8
XFILLER_6_679 VPWR VGND sg13g2_decap_8
XFILLER_5_123 VPWR VGND sg13g2_decap_8
XFILLER_2_830 VPWR VGND sg13g2_decap_8
XFILLER_96_406 VPWR VGND sg13g2_decap_8
XFILLER_104_791 VPWR VGND sg13g2_decap_8
XFILLER_49_333 VPWR VGND sg13g2_decap_8
XFILLER_76_130 VPWR VGND sg13g2_decap_8
X_61_ net23 _23_ _26_ VPWR VGND sg13g2_xnor2_1
XFILLER_92_623 VPWR VGND sg13g2_decap_8
XFILLER_77_686 VPWR VGND sg13g2_decap_8
XFILLER_65_826 VPWR VGND sg13g2_decap_8
XFILLER_94_84 VPWR VGND sg13g2_decap_8
XFILLER_91_133 VPWR VGND sg13g2_decap_8
XFILLER_64_347 VPWR VGND sg13g2_decap_8
XFILLER_18_742 VPWR VGND sg13g2_decap_8
XFILLER_17_263 VPWR VGND sg13g2_decap_8
XFILLER_32_200 VPWR VGND sg13g2_decap_8
XFILLER_33_756 VPWR VGND sg13g2_decap_8
XFILLER_60_564 VPWR VGND sg13g2_decap_8
XFILLER_20_417 VPWR VGND sg13g2_decap_8
XFILLER_32_277 VPWR VGND sg13g2_decap_8
XFILLER_9_462 VPWR VGND sg13g2_decap_8
XFILLER_88_907 VPWR VGND sg13g2_decap_8
XFILLER_5_690 VPWR VGND sg13g2_decap_8
XFILLER_102_728 VPWR VGND sg13g2_decap_8
XFILLER_99_266 VPWR VGND sg13g2_decap_8
XFILLER_87_406 VPWR VGND sg13g2_decap_8
XFILLER_101_238 VPWR VGND sg13g2_decap_8
XFILLER_96_973 VPWR VGND sg13g2_decap_8
XFILLER_68_642 VPWR VGND sg13g2_decap_8
XFILLER_95_494 VPWR VGND sg13g2_decap_8
XFILLER_83_634 VPWR VGND sg13g2_decap_8
XFILLER_56_837 VPWR VGND sg13g2_decap_8
XFILLER_28_539 VPWR VGND sg13g2_decap_8
XFILLER_82_133 VPWR VGND sg13g2_decap_8
XFILLER_67_196 VPWR VGND sg13g2_decap_8
XFILLER_55_336 VPWR VGND sg13g2_decap_8
XFILLER_51_564 VPWR VGND sg13g2_decap_8
XFILLER_11_406 VPWR VGND sg13g2_decap_8
XFILLER_12_907 VPWR VGND sg13g2_decap_8
XFILLER_24_767 VPWR VGND sg13g2_decap_8
XFILLER_23_14 VPWR VGND sg13g2_decap_8
XFILLER_23_266 VPWR VGND sg13g2_decap_8
XFILLER_104_1001 VPWR VGND sg13g2_decap_8
XFILLER_20_984 VPWR VGND sg13g2_decap_8
XFILLER_105_511 VPWR VGND sg13g2_decap_8
XFILLER_3_616 VPWR VGND sg13g2_decap_8
XFILLER_79_907 VPWR VGND sg13g2_decap_8
XFILLER_2_137 VPWR VGND sg13g2_decap_8
XFILLER_105_588 VPWR VGND sg13g2_decap_8
XFILLER_87_973 VPWR VGND sg13g2_decap_8
XFILLER_59_642 VPWR VGND sg13g2_decap_8
XFILLER_47_826 VPWR VGND sg13g2_decap_8
XFILLER_48_77 VPWR VGND sg13g2_decap_8
XFILLER_19_539 VPWR VGND sg13g2_decap_8
XFILLER_86_494 VPWR VGND sg13g2_decap_8
XFILLER_74_645 VPWR VGND sg13g2_decap_8
XFILLER_73_144 VPWR VGND sg13g2_decap_8
XFILLER_58_196 VPWR VGND sg13g2_decap_8
XFILLER_46_347 VPWR VGND sg13g2_decap_8
XFILLER_64_32 VPWR VGND sg13g2_decap_8
XFILLER_27_550 VPWR VGND sg13g2_decap_8
XFILLER_70_840 VPWR VGND sg13g2_decap_8
XFILLER_42_564 VPWR VGND sg13g2_decap_8
XFILLER_15_767 VPWR VGND sg13g2_decap_8
XFILLER_80_42 VPWR VGND sg13g2_decap_8
XFILLER_9_49 VPWR VGND sg13g2_decap_8
XFILLER_14_266 VPWR VGND sg13g2_decap_8
XFILLER_70_1022 VPWR VGND sg13g2_decap_8
XFILLER_7_900 VPWR VGND sg13g2_decap_8
XFILLER_11_973 VPWR VGND sg13g2_decap_8
XFILLER_10_494 VPWR VGND sg13g2_decap_8
XFILLER_7_977 VPWR VGND sg13g2_decap_8
XFILLER_13_91 VPWR VGND sg13g2_decap_8
XFILLER_6_476 VPWR VGND sg13g2_decap_8
XFILLER_89_84 VPWR VGND sg13g2_decap_8
XFILLER_96_203 VPWR VGND sg13g2_decap_8
XFILLER_43_7 VPWR VGND sg13g2_decap_8
XFILLER_69_428 VPWR VGND sg13g2_decap_8
XFILLER_78_951 VPWR VGND sg13g2_decap_8
XFILLER_49_130 VPWR VGND sg13g2_decap_8
XFILLER_77_483 VPWR VGND sg13g2_decap_8
XFILLER_65_623 VPWR VGND sg13g2_decap_8
XFILLER_38_826 VPWR VGND sg13g2_decap_8
XFILLER_93_943 VPWR VGND sg13g2_decap_8
XFILLER_92_420 VPWR VGND sg13g2_decap_8
X_44_ VGND VPWR _04_ _07_ _12_ _08_ sg13g2_a21oi_1
XFILLER_37_347 VPWR VGND sg13g2_decap_8
XFILLER_64_144 VPWR VGND sg13g2_decap_8
XFILLER_92_497 VPWR VGND sg13g2_decap_8
XFILLER_80_637 VPWR VGND sg13g2_decap_8
XFILLER_61_851 VPWR VGND sg13g2_decap_8
XFILLER_33_553 VPWR VGND sg13g2_decap_8
XFILLER_60_361 VPWR VGND sg13g2_decap_8
XFILLER_20_214 VPWR VGND sg13g2_decap_8
XFILLER_106_308 VPWR VGND sg13g2_decap_8
XFILLER_88_704 VPWR VGND sg13g2_decap_8
XFILLER_87_203 VPWR VGND sg13g2_decap_8
XFILLER_102_525 VPWR VGND sg13g2_decap_8
XFILLER_96_770 VPWR VGND sg13g2_decap_8
XFILLER_84_910 VPWR VGND sg13g2_decap_8
XFILLER_69_995 VPWR VGND sg13g2_decap_8
XFILLER_18_14 VPWR VGND sg13g2_decap_8
XFILLER_29_837 VPWR VGND sg13g2_decap_8
XFILLER_95_291 VPWR VGND sg13g2_decap_8
XFILLER_83_431 VPWR VGND sg13g2_decap_8
XFILLER_56_634 VPWR VGND sg13g2_decap_8
XFILLER_55_133 VPWR VGND sg13g2_decap_8
XFILLER_28_336 VPWR VGND sg13g2_decap_8
XFILLER_84_987 VPWR VGND sg13g2_decap_8
XFILLER_71_648 VPWR VGND sg13g2_decap_8
XFILLER_70_147 VPWR VGND sg13g2_decap_8
XFILLER_52_840 VPWR VGND sg13g2_decap_8
XFILLER_12_704 VPWR VGND sg13g2_decap_8
XFILLER_24_564 VPWR VGND sg13g2_decap_8
XFILLER_34_46 VPWR VGND sg13g2_decap_8
XFILLER_54_1028 VPWR VGND sg13g2_fill_1
XFILLER_51_361 VPWR VGND sg13g2_decap_8
XFILLER_11_203 VPWR VGND sg13g2_decap_8
XFILLER_7_207 VPWR VGND sg13g2_decap_8
XFILLER_50_56 VPWR VGND sg13g2_decap_8
XFILLER_20_781 VPWR VGND sg13g2_decap_8
XFILLER_4_903 VPWR VGND sg13g2_decap_8
XFILLER_3_413 VPWR VGND sg13g2_decap_8
XFILLER_106_875 VPWR VGND sg13g2_decap_8
XFILLER_79_704 VPWR VGND sg13g2_decap_8
XFILLER_59_32 VPWR VGND sg13g2_decap_8
XFILLER_105_385 VPWR VGND sg13g2_decap_8
XFILLER_94_707 VPWR VGND sg13g2_decap_8
XFILLER_78_258 VPWR VGND sg13g2_decap_8
XFILLER_87_770 VPWR VGND sg13g2_decap_8
XFILLER_75_910 VPWR VGND sg13g2_decap_8
XFILLER_47_623 VPWR VGND sg13g2_decap_8
XFILLER_86_291 VPWR VGND sg13g2_decap_8
XFILLER_75_42 VPWR VGND sg13g2_decap_8
XFILLER_74_442 VPWR VGND sg13g2_decap_8
XFILLER_19_336 VPWR VGND sg13g2_decap_8
XFILLER_75_987 VPWR VGND sg13g2_decap_8
XFILLER_46_144 VPWR VGND sg13g2_decap_8
XFILLER_90_935 VPWR VGND sg13g2_decap_8
XFILLER_62_637 VPWR VGND sg13g2_decap_8
XFILLER_61_158 VPWR VGND sg13g2_decap_8
XFILLER_43_840 VPWR VGND sg13g2_decap_8
XFILLER_91_63 VPWR VGND sg13g2_decap_8
XFILLER_42_361 VPWR VGND sg13g2_decap_8
XFILLER_15_564 VPWR VGND sg13g2_decap_8
XFILLER_11_770 VPWR VGND sg13g2_decap_8
XFILLER_30_567 VPWR VGND sg13g2_decap_8
XFILLER_10_291 VPWR VGND sg13g2_decap_8
XFILLER_7_774 VPWR VGND sg13g2_decap_8
XFILLER_6_273 VPWR VGND sg13g2_decap_8
XFILLER_69_225 VPWR VGND sg13g2_decap_8
XFILLER_3_980 VPWR VGND sg13g2_decap_8
XFILLER_97_567 VPWR VGND sg13g2_decap_8
XFILLER_85_707 VPWR VGND sg13g2_decap_8
XFILLER_84_217 VPWR VGND sg13g2_decap_8
XFILLER_38_623 VPWR VGND sg13g2_decap_8
XFILLER_93_740 VPWR VGND sg13g2_decap_8
XFILLER_77_280 VPWR VGND sg13g2_decap_8
XFILLER_66_965 VPWR VGND sg13g2_decap_8
XFILLER_65_420 VPWR VGND sg13g2_decap_8
XFILLER_37_144 VPWR VGND sg13g2_decap_8
XFILLER_92_294 VPWR VGND sg13g2_decap_8
XFILLER_81_935 VPWR VGND sg13g2_decap_8
XFILLER_80_434 VPWR VGND sg13g2_decap_8
XFILLER_65_497 VPWR VGND sg13g2_decap_8
XFILLER_53_637 VPWR VGND sg13g2_decap_8
XFILLER_52_147 VPWR VGND sg13g2_decap_8
XFILLER_34_851 VPWR VGND sg13g2_decap_8
XFILLER_33_350 VPWR VGND sg13g2_decap_8
XFILLER_14_1001 VPWR VGND sg13g2_decap_8
XFILLER_21_567 VPWR VGND sg13g2_decap_8
XFILLER_106_105 VPWR VGND sg13g2_decap_8
XFILLER_101_1015 VPWR VGND sg13g2_decap_8
XFILLER_88_501 VPWR VGND sg13g2_decap_8
XFILLER_1_917 VPWR VGND sg13g2_decap_8
XFILLER_103_812 VPWR VGND sg13g2_decap_8
XFILLER_0_427 VPWR VGND sg13g2_decap_8
XFILLER_102_322 VPWR VGND sg13g2_decap_8
XFILLER_76_718 VPWR VGND sg13g2_decap_8
XFILLER_103_889 VPWR VGND sg13g2_decap_8
XFILLER_88_578 VPWR VGND sg13g2_decap_8
XFILLER_75_217 VPWR VGND sg13g2_decap_8
XFILLER_57_910 VPWR VGND sg13g2_decap_8
XFILLER_29_46 VPWR VGND sg13g2_decap_8
XFILLER_102_399 VPWR VGND sg13g2_decap_8
XFILLER_69_792 VPWR VGND sg13g2_decap_8
XFILLER_56_431 VPWR VGND sg13g2_decap_8
XFILLER_29_634 VPWR VGND sg13g2_decap_8
XFILLER_84_784 VPWR VGND sg13g2_decap_8
XFILLER_72_924 VPWR VGND sg13g2_decap_8
XFILLER_57_987 VPWR VGND sg13g2_decap_8
XFILLER_28_133 VPWR VGND sg13g2_decap_8
XFILLER_45_56 VPWR VGND sg13g2_decap_8
XFILLER_44_648 VPWR VGND sg13g2_decap_8
XFILLER_71_445 VPWR VGND sg13g2_decap_8
XFILLER_43_147 VPWR VGND sg13g2_decap_8
XFILLER_25_840 VPWR VGND sg13g2_decap_8
XFILLER_12_501 VPWR VGND sg13g2_decap_8
XFILLER_24_361 VPWR VGND sg13g2_decap_8
XFILLER_101_84 VPWR VGND sg13g2_decap_8
XFILLER_61_11 VPWR VGND sg13g2_fill_2
XFILLER_40_854 VPWR VGND sg13g2_decap_8
XFILLER_61_44 VPWR VGND sg13g2_decap_8
XFILLER_12_578 VPWR VGND sg13g2_decap_8
XFILLER_61_88 VPWR VGND sg13g2_decap_8
XFILLER_6_28 VPWR VGND sg13g2_decap_8
XFILLER_4_700 VPWR VGND sg13g2_decap_8
XFILLER_3_210 VPWR VGND sg13g2_decap_8
XFILLER_79_501 VPWR VGND sg13g2_decap_8
XFILLER_4_777 VPWR VGND sg13g2_decap_8
XFILLER_106_672 VPWR VGND sg13g2_decap_8
XFILLER_10_81 VPWR VGND sg13g2_decap_8
XFILLER_3_287 VPWR VGND sg13g2_decap_8
XFILLER_105_182 VPWR VGND sg13g2_decap_8
XFILLER_67_707 VPWR VGND sg13g2_decap_8
XFILLER_94_504 VPWR VGND sg13g2_decap_8
XFILLER_86_74 VPWR VGND sg13g2_decap_8
XFILLER_79_578 VPWR VGND sg13g2_decap_8
XFILLER_48_910 VPWR VGND sg13g2_decap_8
XFILLER_47_420 VPWR VGND sg13g2_decap_8
XFILLER_0_994 VPWR VGND sg13g2_decap_8
XFILLER_48_987 VPWR VGND sg13g2_decap_8
XFILLER_19_133 VPWR VGND sg13g2_decap_8
XFILLER_90_732 VPWR VGND sg13g2_decap_8
XFILLER_75_784 VPWR VGND sg13g2_decap_8
XFILLER_63_924 VPWR VGND sg13g2_decap_8
XFILLER_47_497 VPWR VGND sg13g2_decap_8
XFILLER_35_637 VPWR VGND sg13g2_decap_8
XFILLER_62_434 VPWR VGND sg13g2_decap_8
XFILLER_16_840 VPWR VGND sg13g2_decap_8
XFILLER_34_158 VPWR VGND sg13g2_decap_8
XFILLER_15_361 VPWR VGND sg13g2_decap_8
XFILLER_37_1012 VPWR VGND sg13g2_decap_8
XFILLER_31_854 VPWR VGND sg13g2_decap_8
XFILLER_30_364 VPWR VGND sg13g2_decap_8
XFILLER_7_571 VPWR VGND sg13g2_decap_8
XFILLER_104_609 VPWR VGND sg13g2_decap_8
XFILLER_103_119 VPWR VGND sg13g2_decap_8
XFILLER_98_865 VPWR VGND sg13g2_decap_8
XFILLER_58_707 VPWR VGND sg13g2_decap_8
XFILLER_44_1005 VPWR VGND sg13g2_decap_8
XFILLER_100_826 VPWR VGND sg13g2_decap_8
XFILLER_97_364 VPWR VGND sg13g2_decap_8
XFILLER_85_504 VPWR VGND sg13g2_decap_8
XFILLER_57_217 VPWR VGND sg13g2_decap_8
XFILLER_39_921 VPWR VGND sg13g2_decap_8
XFILLER_38_420 VPWR VGND sg13g2_decap_8
XFILLER_66_762 VPWR VGND sg13g2_decap_8
XFILLER_81_732 VPWR VGND sg13g2_decap_8
XFILLER_54_935 VPWR VGND sg13g2_decap_8
XFILLER_26_637 VPWR VGND sg13g2_decap_8
XFILLER_38_497 VPWR VGND sg13g2_decap_8
XFILLER_39_998 VPWR VGND sg13g2_decap_8
XFILLER_80_231 VPWR VGND sg13g2_decap_8
XFILLER_65_294 VPWR VGND sg13g2_decap_8
XFILLER_53_434 VPWR VGND sg13g2_decap_8
XFILLER_25_147 VPWR VGND sg13g2_decap_8
XFILLER_21_364 VPWR VGND sg13g2_decap_8
XFILLER_22_865 VPWR VGND sg13g2_decap_8
XFILLER_31_14 VPWR VGND sg13g2_decap_8
XFILLER_5_508 VPWR VGND sg13g2_decap_8
XFILLER_1_714 VPWR VGND sg13g2_decap_8
XFILLER_89_854 VPWR VGND sg13g2_decap_8
XFILLER_0_224 VPWR VGND sg13g2_decap_8
XFILLER_103_686 VPWR VGND sg13g2_decap_8
XFILLER_88_375 VPWR VGND sg13g2_decap_8
XFILLER_76_515 VPWR VGND sg13g2_decap_8
XFILLER_49_718 VPWR VGND sg13g2_decap_8
XFILLER_48_217 VPWR VGND sg13g2_decap_8
XFILLER_102_196 VPWR VGND sg13g2_decap_8
XFILLER_56_11 VPWR VGND sg13g2_decap_8
XFILLER_29_431 VPWR VGND sg13g2_decap_8
XFILLER_91_518 VPWR VGND sg13g2_decap_8
XFILLER_84_581 VPWR VGND sg13g2_decap_8
XFILLER_72_721 VPWR VGND sg13g2_decap_8
XFILLER_57_784 VPWR VGND sg13g2_decap_8
XFILLER_56_88 VPWR VGND sg13g2_decap_8
XFILLER_45_924 VPWR VGND sg13g2_decap_8
XFILLER_71_242 VPWR VGND sg13g2_decap_8
XFILLER_44_445 VPWR VGND sg13g2_decap_8
XFILLER_16_147 VPWR VGND sg13g2_decap_8
XFILLER_17_648 VPWR VGND sg13g2_decap_8
XFILLER_72_798 VPWR VGND sg13g2_decap_8
XFILLER_72_21 VPWR VGND sg13g2_decap_8
XFILLER_60_949 VPWR VGND sg13g2_decap_8
XFILLER_13_854 VPWR VGND sg13g2_decap_8
XFILLER_72_98 VPWR VGND sg13g2_decap_8
XFILLER_40_651 VPWR VGND sg13g2_decap_8
XFILLER_9_847 VPWR VGND sg13g2_decap_8
XFILLER_12_375 VPWR VGND sg13g2_decap_8
XFILLER_8_357 VPWR VGND sg13g2_decap_8
XFILLER_21_91 VPWR VGND sg13g2_decap_8
XFILLER_4_574 VPWR VGND sg13g2_decap_8
XFILLER_97_84 VPWR VGND sg13g2_decap_8
XFILLER_95_802 VPWR VGND sg13g2_decap_8
XFILLER_94_301 VPWR VGND sg13g2_decap_8
XFILLER_79_375 VPWR VGND sg13g2_decap_8
XFILLER_67_504 VPWR VGND sg13g2_decap_8
XFILLER_0_791 VPWR VGND sg13g2_decap_8
XFILLER_39_228 VPWR VGND sg13g2_decap_8
XFILLER_95_879 VPWR VGND sg13g2_decap_8
XFILLER_94_378 VPWR VGND sg13g2_decap_8
XFILLER_82_518 VPWR VGND sg13g2_decap_8
XFILLER_75_581 VPWR VGND sg13g2_decap_8
XFILLER_63_721 VPWR VGND sg13g2_decap_8
XFILLER_48_784 VPWR VGND sg13g2_decap_8
XFILLER_36_924 VPWR VGND sg13g2_decap_8
XFILLER_62_231 VPWR VGND sg13g2_decap_8
XFILLER_47_294 VPWR VGND sg13g2_decap_8
XFILLER_35_434 VPWR VGND sg13g2_decap_8
XFILLER_74_1009 VPWR VGND sg13g2_decap_8
XFILLER_63_798 VPWR VGND sg13g2_decap_8
XFILLER_51_949 VPWR VGND sg13g2_decap_8
XFILLER_50_448 VPWR VGND sg13g2_decap_8
XFILLER_31_651 VPWR VGND sg13g2_decap_8
XFILLER_30_161 VPWR VGND sg13g2_decap_8
XFILLER_7_60 VPWR VGND sg13g2_decap_8
XFILLER_11_1015 VPWR VGND sg13g2_decap_8
XFILLER_104_406 VPWR VGND sg13g2_decap_8
XFILLER_98_662 VPWR VGND sg13g2_decap_8
XFILLER_97_161 VPWR VGND sg13g2_decap_8
XFILLER_86_802 VPWR VGND sg13g2_decap_8
XFILLER_85_301 VPWR VGND sg13g2_decap_8
XFILLER_58_504 VPWR VGND sg13g2_decap_8
XFILLER_100_623 VPWR VGND sg13g2_decap_8
XFILLER_86_879 VPWR VGND sg13g2_decap_8
XFILLER_85_378 VPWR VGND sg13g2_decap_8
XFILLER_73_529 VPWR VGND sg13g2_decap_8
XFILLER_26_14 VPWR VGND sg13g2_decap_8
XFILLER_27_935 VPWR VGND sg13g2_decap_8
XFILLER_39_795 VPWR VGND sg13g2_decap_8
XFILLER_54_732 VPWR VGND sg13g2_decap_8
XFILLER_53_231 VPWR VGND sg13g2_decap_8
XFILLER_26_434 VPWR VGND sg13g2_decap_8
XFILLER_38_294 VPWR VGND sg13g2_decap_8
XFILLER_42_949 VPWR VGND sg13g2_decap_8
XFILLER_41_448 VPWR VGND sg13g2_decap_8
XFILLER_10_802 VPWR VGND sg13g2_decap_8
XFILLER_22_662 VPWR VGND sg13g2_decap_8
XFILLER_42_46 VPWR VGND sg13g2_decap_8
XFILLER_21_161 VPWR VGND sg13g2_decap_8
XFILLER_10_879 VPWR VGND sg13g2_decap_8
XFILLER_5_305 VPWR VGND sg13g2_decap_8
XFILLER_1_511 VPWR VGND sg13g2_decap_8
XFILLER_104_973 VPWR VGND sg13g2_decap_8
XFILLER_95_109 VPWR VGND sg13g2_decap_8
XFILLER_89_651 VPWR VGND sg13g2_decap_8
XFILLER_49_515 VPWR VGND sg13g2_decap_8
XFILLER_103_483 VPWR VGND sg13g2_decap_8
XFILLER_88_172 VPWR VGND sg13g2_decap_8
XFILLER_76_312 VPWR VGND sg13g2_decap_8
XFILLER_1_588 VPWR VGND sg13g2_decap_8
XFILLER_92_805 VPWR VGND sg13g2_decap_8
XFILLER_77_868 VPWR VGND sg13g2_decap_8
XFILLER_67_98 VPWR VGND sg13g2_decap_8
XFILLER_91_315 VPWR VGND sg13g2_decap_8
XFILLER_76_389 VPWR VGND sg13g2_decap_8
XFILLER_64_529 VPWR VGND sg13g2_decap_8
XFILLER_57_581 VPWR VGND sg13g2_decap_8
XFILLER_45_721 VPWR VGND sg13g2_decap_8
XFILLER_18_924 VPWR VGND sg13g2_decap_8
XFILLER_83_53 VPWR VGND sg13g2_decap_8
XFILLER_17_445 VPWR VGND sg13g2_decap_8
XFILLER_45_798 VPWR VGND sg13g2_decap_8
XFILLER_44_242 VPWR VGND sg13g2_decap_8
XFILLER_33_938 VPWR VGND sg13g2_decap_8
XFILLER_72_595 VPWR VGND sg13g2_decap_8
XFILLER_60_746 VPWR VGND sg13g2_decap_8
XFILLER_13_651 VPWR VGND sg13g2_decap_8
XFILLER_16_91 VPWR VGND sg13g2_decap_8
XFILLER_32_459 VPWR VGND sg13g2_decap_8
XFILLER_9_644 VPWR VGND sg13g2_decap_8
XFILLER_12_172 VPWR VGND sg13g2_decap_8
XFILLER_34_1026 VPWR VGND sg13g2_fill_2
XFILLER_8_154 VPWR VGND sg13g2_decap_8
XFILLER_5_872 VPWR VGND sg13g2_decap_8
XFILLER_99_448 VPWR VGND sg13g2_decap_8
XFILLER_4_371 VPWR VGND sg13g2_decap_8
XFILLER_86_109 VPWR VGND sg13g2_decap_8
XFILLER_68_824 VPWR VGND sg13g2_decap_8
XFILLER_79_172 VPWR VGND sg13g2_decap_8
XFILLER_67_301 VPWR VGND sg13g2_decap_8
XFILLER_41_1008 VPWR VGND sg13g2_decap_8
XFILLER_95_676 VPWR VGND sg13g2_decap_8
XFILLER_83_816 VPWR VGND sg13g2_decap_8
XFILLER_94_175 VPWR VGND sg13g2_decap_8
XFILLER_82_315 VPWR VGND sg13g2_decap_8
XFILLER_67_378 VPWR VGND sg13g2_decap_8
XFILLER_55_518 VPWR VGND sg13g2_decap_8
XFILLER_48_581 VPWR VGND sg13g2_decap_8
XFILLER_36_721 VPWR VGND sg13g2_decap_8
XFILLER_35_231 VPWR VGND sg13g2_decap_8
XFILLER_91_882 VPWR VGND sg13g2_decap_8
XFILLER_36_798 VPWR VGND sg13g2_decap_8
XFILLER_63_595 VPWR VGND sg13g2_decap_8
XFILLER_51_746 VPWR VGND sg13g2_decap_8
XFILLER_23_448 VPWR VGND sg13g2_decap_8
XFILLER_24_949 VPWR VGND sg13g2_decap_8
XFILLER_50_245 VPWR VGND sg13g2_decap_8
XFILLER_10_109 VPWR VGND sg13g2_decap_8
XFILLER_104_203 VPWR VGND sg13g2_decap_8
XFILLER_2_319 VPWR VGND sg13g2_decap_8
XFILLER_101_910 VPWR VGND sg13g2_decap_8
XFILLER_100_420 VPWR VGND sg13g2_decap_8
XFILLER_59_824 VPWR VGND sg13g2_decap_8
XFILLER_58_301 VPWR VGND sg13g2_decap_8
XFILLER_86_676 VPWR VGND sg13g2_decap_8
XFILLER_101_987 VPWR VGND sg13g2_decap_8
XFILLER_85_175 VPWR VGND sg13g2_decap_8
XFILLER_74_827 VPWR VGND sg13g2_decap_8
XFILLER_73_326 VPWR VGND sg13g2_decap_8
XFILLER_58_378 VPWR VGND sg13g2_decap_8
XFILLER_46_529 VPWR VGND sg13g2_decap_8
XFILLER_37_46 VPWR VGND sg13g2_decap_8
XFILLER_100_497 VPWR VGND sg13g2_decap_8
XFILLER_26_231 VPWR VGND sg13g2_decap_8
XFILLER_27_732 VPWR VGND sg13g2_decap_8
XFILLER_39_592 VPWR VGND sg13g2_decap_8
XFILLER_82_882 VPWR VGND sg13g2_decap_8
XFILLER_57_1015 VPWR VGND sg13g2_decap_8
XFILLER_42_746 VPWR VGND sg13g2_decap_8
XFILLER_15_949 VPWR VGND sg13g2_decap_8
XFILLER_53_56 VPWR VGND sg13g2_decap_8
XFILLER_14_448 VPWR VGND sg13g2_decap_8
XFILLER_41_245 VPWR VGND sg13g2_decap_8
XFILLER_10_676 VPWR VGND sg13g2_decap_8
XFILLER_5_102 VPWR VGND sg13g2_decap_8
XFILLER_6_658 VPWR VGND sg13g2_decap_8
XFILLER_5_179 VPWR VGND sg13g2_decap_8
XFILLER_64_1019 VPWR VGND sg13g2_decap_8
XFILLER_78_53 VPWR VGND sg13g2_decap_8
XFILLER_104_770 VPWR VGND sg13g2_decap_8
XFILLER_78_97 VPWR VGND sg13g2_decap_8
XFILLER_49_312 VPWR VGND sg13g2_decap_8
XFILLER_2_886 VPWR VGND sg13g2_decap_8
XFILLER_1_385 VPWR VGND sg13g2_decap_8
XFILLER_103_280 VPWR VGND sg13g2_decap_8
XFILLER_77_665 VPWR VGND sg13g2_decap_8
X_60_ net15 net7 _26_ VPWR VGND sg13g2_xor2_1
XFILLER_65_805 VPWR VGND sg13g2_decap_8
XFILLER_94_63 VPWR VGND sg13g2_decap_8
XFILLER_92_602 VPWR VGND sg13g2_decap_8
XFILLER_64_326 VPWR VGND sg13g2_decap_8
XFILLER_49_389 VPWR VGND sg13g2_decap_8
XFILLER_37_529 VPWR VGND sg13g2_decap_8
XFILLER_91_112 VPWR VGND sg13g2_decap_8
XFILLER_76_186 VPWR VGND sg13g2_decap_8
XFILLER_18_721 VPWR VGND sg13g2_decap_8
XFILLER_92_679 VPWR VGND sg13g2_decap_8
XFILLER_80_819 VPWR VGND sg13g2_decap_8
XFILLER_17_242 VPWR VGND sg13g2_decap_8
XFILLER_91_189 VPWR VGND sg13g2_decap_8
XFILLER_73_893 VPWR VGND sg13g2_decap_8
XFILLER_72_392 VPWR VGND sg13g2_decap_8
XFILLER_45_595 VPWR VGND sg13g2_decap_8
XFILLER_18_798 VPWR VGND sg13g2_decap_8
XFILLER_33_735 VPWR VGND sg13g2_decap_8
XFILLER_60_543 VPWR VGND sg13g2_decap_8
XFILLER_32_256 VPWR VGND sg13g2_decap_8
XFILLER_9_441 VPWR VGND sg13g2_decap_8
XFILLER_71_4 VPWR VGND sg13g2_decap_8
XFILLER_99_245 VPWR VGND sg13g2_decap_8
XFILLER_102_707 VPWR VGND sg13g2_decap_8
XFILLER_101_217 VPWR VGND sg13g2_decap_8
XFILLER_68_621 VPWR VGND sg13g2_decap_8
XFILLER_96_952 VPWR VGND sg13g2_decap_8
XFILLER_95_473 VPWR VGND sg13g2_decap_8
XFILLER_83_613 VPWR VGND sg13g2_decap_8
XFILLER_68_698 VPWR VGND sg13g2_decap_8
XFILLER_67_175 VPWR VGND sg13g2_decap_8
XFILLER_56_816 VPWR VGND sg13g2_decap_8
XFILLER_55_315 VPWR VGND sg13g2_decap_8
XFILLER_28_518 VPWR VGND sg13g2_decap_8
XFILLER_82_112 VPWR VGND sg13g2_decap_8
XFILLER_82_189 VPWR VGND sg13g2_decap_8
XFILLER_70_329 VPWR VGND sg13g2_decap_8
XFILLER_64_893 VPWR VGND sg13g2_decap_8
XFILLER_24_746 VPWR VGND sg13g2_decap_8
XFILLER_36_595 VPWR VGND sg13g2_decap_8
XFILLER_63_392 VPWR VGND sg13g2_decap_8
XFILLER_51_543 VPWR VGND sg13g2_decap_8
XFILLER_23_245 VPWR VGND sg13g2_decap_8
XFILLER_20_963 VPWR VGND sg13g2_decap_8
XFILLER_87_1008 VPWR VGND sg13g2_decap_8
XFILLER_3_7 VPWR VGND sg13g2_decap_8
XFILLER_2_116 VPWR VGND sg13g2_decap_8
XFILLER_105_567 VPWR VGND sg13g2_decap_8
XFILLER_59_621 VPWR VGND sg13g2_decap_8
XFILLER_87_952 VPWR VGND sg13g2_decap_8
XFILLER_47_805 VPWR VGND sg13g2_decap_8
XFILLER_48_56 VPWR VGND sg13g2_decap_8
XFILLER_101_784 VPWR VGND sg13g2_decap_8
XFILLER_86_473 VPWR VGND sg13g2_decap_8
XFILLER_74_624 VPWR VGND sg13g2_decap_8
XFILLER_59_698 VPWR VGND sg13g2_decap_8
XFILLER_58_175 VPWR VGND sg13g2_decap_8
XFILLER_19_518 VPWR VGND sg13g2_decap_8
XFILLER_100_294 VPWR VGND sg13g2_decap_8
XFILLER_73_123 VPWR VGND sg13g2_decap_8
XFILLER_64_11 VPWR VGND sg13g2_decap_8
XFILLER_46_326 VPWR VGND sg13g2_decap_8
XFILLER_104_84 VPWR VGND sg13g2_decap_8
XFILLER_62_819 VPWR VGND sg13g2_decap_8
XFILLER_64_88 VPWR VGND sg13g2_decap_8
XFILLER_55_882 VPWR VGND sg13g2_decap_8
XFILLER_15_746 VPWR VGND sg13g2_decap_8
XFILLER_42_543 VPWR VGND sg13g2_decap_8
XFILLER_14_245 VPWR VGND sg13g2_decap_8
XFILLER_80_21 VPWR VGND sg13g2_decap_8
XFILLER_70_1001 VPWR VGND sg13g2_decap_8
XFILLER_70_896 VPWR VGND sg13g2_decap_8
XFILLER_9_28 VPWR VGND sg13g2_decap_8
XFILLER_11_952 VPWR VGND sg13g2_decap_8
XFILLER_30_749 VPWR VGND sg13g2_decap_8
XFILLER_80_98 VPWR VGND sg13g2_decap_8
XFILLER_10_473 VPWR VGND sg13g2_decap_8
XFILLER_7_956 VPWR VGND sg13g2_decap_8
XFILLER_13_70 VPWR VGND sg13g2_decap_8
XFILLER_6_455 VPWR VGND sg13g2_decap_8
XFILLER_89_63 VPWR VGND sg13g2_decap_8
XFILLER_69_407 VPWR VGND sg13g2_decap_8
XFILLER_9_1008 VPWR VGND sg13g2_decap_8
XFILLER_97_749 VPWR VGND sg13g2_decap_8
XFILLER_78_930 VPWR VGND sg13g2_decap_8
XFILLER_2_683 VPWR VGND sg13g2_decap_8
XFILLER_36_7 VPWR VGND sg13g2_decap_8
XFILLER_96_259 VPWR VGND sg13g2_decap_8
XFILLER_1_182 VPWR VGND sg13g2_decap_8
XFILLER_38_805 VPWR VGND sg13g2_decap_8
XFILLER_93_922 VPWR VGND sg13g2_decap_8
XFILLER_77_462 VPWR VGND sg13g2_decap_8
XFILLER_65_602 VPWR VGND sg13g2_decap_8
X_43_ _11_ _09_ _05_ VPWR VGND sg13g2_nand2b_1
XFILLER_64_123 VPWR VGND sg13g2_decap_8
XFILLER_49_186 VPWR VGND sg13g2_decap_8
XFILLER_37_326 VPWR VGND sg13g2_decap_8
XFILLER_93_999 VPWR VGND sg13g2_decap_8
XFILLER_92_476 VPWR VGND sg13g2_decap_8
XFILLER_80_616 VPWR VGND sg13g2_decap_8
XFILLER_65_679 VPWR VGND sg13g2_decap_8
XFILLER_53_819 VPWR VGND sg13g2_decap_8
XFILLER_73_690 VPWR VGND sg13g2_decap_8
XFILLER_61_830 VPWR VGND sg13g2_decap_8
XFILLER_52_329 VPWR VGND sg13g2_decap_8
XFILLER_46_893 VPWR VGND sg13g2_decap_8
XFILLER_18_595 VPWR VGND sg13g2_decap_8
XFILLER_60_340 VPWR VGND sg13g2_decap_8
XFILLER_45_392 VPWR VGND sg13g2_decap_8
XFILLER_33_532 VPWR VGND sg13g2_decap_8
XFILLER_21_749 VPWR VGND sg13g2_decap_8
XFILLER_62_0 VPWR VGND sg13g2_decap_8
XFILLER_102_504 VPWR VGND sg13g2_decap_8
XFILLER_0_609 VPWR VGND sg13g2_decap_8
XFILLER_87_259 VPWR VGND sg13g2_decap_8
XFILLER_69_974 VPWR VGND sg13g2_decap_8
XFILLER_56_613 VPWR VGND sg13g2_decap_8
XFILLER_28_315 VPWR VGND sg13g2_decap_8
XFILLER_29_816 VPWR VGND sg13g2_decap_8
XFILLER_95_270 VPWR VGND sg13g2_decap_8
XFILLER_84_966 VPWR VGND sg13g2_decap_8
XFILLER_83_410 VPWR VGND sg13g2_decap_8
XFILLER_68_495 VPWR VGND sg13g2_decap_8
XFILLER_55_112 VPWR VGND sg13g2_decap_8
XFILLER_83_487 VPWR VGND sg13g2_decap_8
XFILLER_71_627 VPWR VGND sg13g2_decap_8
XFILLER_70_126 VPWR VGND sg13g2_decap_8
XFILLER_64_690 VPWR VGND sg13g2_decap_8
XFILLER_55_189 VPWR VGND sg13g2_decap_8
XFILLER_43_329 VPWR VGND sg13g2_decap_8
XFILLER_37_893 VPWR VGND sg13g2_decap_8
XFILLER_51_340 VPWR VGND sg13g2_decap_8
XFILLER_24_543 VPWR VGND sg13g2_decap_8
XFILLER_34_25 VPWR VGND sg13g2_decap_8
XFILLER_36_392 VPWR VGND sg13g2_decap_8
XFILLER_52_896 VPWR VGND sg13g2_decap_8
XFILLER_11_259 VPWR VGND sg13g2_decap_8
XFILLER_20_760 VPWR VGND sg13g2_decap_8
XFILLER_50_35 VPWR VGND sg13g2_decap_8
XFILLER_4_959 VPWR VGND sg13g2_decap_8
XFILLER_106_854 VPWR VGND sg13g2_decap_8
XFILLER_59_11 VPWR VGND sg13g2_decap_8
XFILLER_3_469 VPWR VGND sg13g2_decap_8
XFILLER_105_364 VPWR VGND sg13g2_decap_8
XFILLER_78_237 VPWR VGND sg13g2_decap_8
XFILLER_59_99 VPWR VGND sg13g2_decap_8
XFILLER_93_229 VPWR VGND sg13g2_decap_8
XFILLER_75_21 VPWR VGND sg13g2_decap_8
XFILLER_47_602 VPWR VGND sg13g2_decap_8
XFILLER_101_581 VPWR VGND sg13g2_decap_8
XFILLER_86_270 VPWR VGND sg13g2_decap_8
XFILLER_75_966 VPWR VGND sg13g2_decap_8
XFILLER_74_421 VPWR VGND sg13g2_decap_8
XFILLER_59_495 VPWR VGND sg13g2_decap_8
XFILLER_46_123 VPWR VGND sg13g2_decap_8
XFILLER_19_315 VPWR VGND sg13g2_decap_8
XFILLER_90_914 VPWR VGND sg13g2_decap_8
XFILLER_75_98 VPWR VGND sg13g2_decap_8
XFILLER_62_616 VPWR VGND sg13g2_decap_8
XFILLER_47_679 VPWR VGND sg13g2_decap_8
XFILLER_35_819 VPWR VGND sg13g2_decap_8
XFILLER_74_498 VPWR VGND sg13g2_decap_8
XFILLER_28_882 VPWR VGND sg13g2_decap_8
XFILLER_91_42 VPWR VGND sg13g2_decap_8
XFILLER_42_340 VPWR VGND sg13g2_decap_8
XFILLER_15_543 VPWR VGND sg13g2_decap_8
XFILLER_43_896 VPWR VGND sg13g2_decap_8
XFILLER_70_693 VPWR VGND sg13g2_decap_8
XFILLER_30_546 VPWR VGND sg13g2_decap_8
XFILLER_10_270 VPWR VGND sg13g2_decap_8
XFILLER_7_753 VPWR VGND sg13g2_decap_8
XFILLER_6_252 VPWR VGND sg13g2_decap_8
XFILLER_69_204 VPWR VGND sg13g2_decap_8
XFILLER_34_4 VPWR VGND sg13g2_decap_8
XFILLER_97_546 VPWR VGND sg13g2_decap_8
XFILLER_2_480 VPWR VGND sg13g2_decap_8
XFILLER_38_602 VPWR VGND sg13g2_decap_8
XFILLER_66_944 VPWR VGND sg13g2_decap_8
XFILLER_37_123 VPWR VGND sg13g2_decap_8
XFILLER_81_914 VPWR VGND sg13g2_decap_8
XFILLER_26_819 VPWR VGND sg13g2_decap_8
XFILLER_38_679 VPWR VGND sg13g2_decap_8
XFILLER_93_796 VPWR VGND sg13g2_decap_8
XFILLER_92_273 VPWR VGND sg13g2_decap_8
XFILLER_80_413 VPWR VGND sg13g2_decap_8
XFILLER_65_476 VPWR VGND sg13g2_decap_8
XFILLER_53_616 VPWR VGND sg13g2_decap_8
XFILLER_1_84 VPWR VGND sg13g2_decap_8
XFILLER_19_882 VPWR VGND sg13g2_decap_8
XFILLER_25_329 VPWR VGND sg13g2_decap_8
XFILLER_52_126 VPWR VGND sg13g2_decap_8
XFILLER_46_690 VPWR VGND sg13g2_decap_8
XFILLER_18_392 VPWR VGND sg13g2_decap_8
XFILLER_34_830 VPWR VGND sg13g2_decap_8
XFILLER_21_546 VPWR VGND sg13g2_decap_8
XFILLER_102_301 VPWR VGND sg13g2_decap_8
XFILLER_0_406 VPWR VGND sg13g2_decap_8
XFILLER_103_868 VPWR VGND sg13g2_decap_8
XFILLER_88_557 VPWR VGND sg13g2_decap_8
XFILLER_29_25 VPWR VGND sg13g2_decap_8
XFILLER_102_378 VPWR VGND sg13g2_decap_8
XFILLER_69_771 VPWR VGND sg13g2_decap_8
XFILLER_29_613 VPWR VGND sg13g2_decap_8
XFILLER_68_292 VPWR VGND sg13g2_decap_8
XFILLER_56_410 VPWR VGND sg13g2_decap_8
XFILLER_28_112 VPWR VGND sg13g2_decap_8
XFILLER_84_763 VPWR VGND sg13g2_decap_8
XFILLER_72_903 VPWR VGND sg13g2_decap_8
XFILLER_57_966 VPWR VGND sg13g2_decap_8
XFILLER_83_284 VPWR VGND sg13g2_decap_8
XFILLER_71_424 VPWR VGND sg13g2_decap_8
XFILLER_56_487 VPWR VGND sg13g2_decap_8
XFILLER_45_35 VPWR VGND sg13g2_decap_8
XFILLER_44_627 VPWR VGND sg13g2_decap_8
XFILLER_16_329 VPWR VGND sg13g2_decap_8
XFILLER_28_189 VPWR VGND sg13g2_decap_8
XFILLER_43_126 VPWR VGND sg13g2_decap_8
XFILLER_37_690 VPWR VGND sg13g2_decap_8
XFILLER_80_980 VPWR VGND sg13g2_decap_8
XFILLER_24_340 VPWR VGND sg13g2_decap_8
XFILLER_25_896 VPWR VGND sg13g2_decap_8
XFILLER_101_63 VPWR VGND sg13g2_decap_8
XFILLER_52_693 VPWR VGND sg13g2_decap_8
XFILLER_40_833 VPWR VGND sg13g2_decap_8
XFILLER_12_557 VPWR VGND sg13g2_decap_8
XFILLER_8_539 VPWR VGND sg13g2_decap_8
XFILLER_106_651 VPWR VGND sg13g2_decap_8
XFILLER_4_756 VPWR VGND sg13g2_decap_8
XFILLER_105_161 VPWR VGND sg13g2_decap_8
XFILLER_10_60 VPWR VGND sg13g2_decap_8
XFILLER_3_266 VPWR VGND sg13g2_decap_8
XFILLER_79_557 VPWR VGND sg13g2_decap_8
XFILLER_86_53 VPWR VGND sg13g2_decap_8
XFILLER_0_973 VPWR VGND sg13g2_decap_8
XFILLER_19_112 VPWR VGND sg13g2_decap_8
XFILLER_75_763 VPWR VGND sg13g2_decap_8
XFILLER_63_903 VPWR VGND sg13g2_decap_8
XFILLER_59_292 VPWR VGND sg13g2_decap_8
XFILLER_48_966 VPWR VGND sg13g2_decap_8
XFILLER_19_91 VPWR VGND sg13g2_decap_8
XFILLER_90_711 VPWR VGND sg13g2_decap_8
XFILLER_62_413 VPWR VGND sg13g2_decap_8
XFILLER_47_476 VPWR VGND sg13g2_decap_8
XFILLER_19_189 VPWR VGND sg13g2_decap_8
XFILLER_35_616 VPWR VGND sg13g2_decap_8
XFILLER_74_295 VPWR VGND sg13g2_decap_8
XFILLER_34_137 VPWR VGND sg13g2_decap_8
XFILLER_90_788 VPWR VGND sg13g2_decap_8
XFILLER_15_340 VPWR VGND sg13g2_decap_8
XFILLER_71_991 VPWR VGND sg13g2_decap_8
XFILLER_70_490 VPWR VGND sg13g2_decap_8
XFILLER_43_693 VPWR VGND sg13g2_decap_8
XFILLER_16_896 VPWR VGND sg13g2_decap_8
XFILLER_31_833 VPWR VGND sg13g2_decap_8
XFILLER_30_343 VPWR VGND sg13g2_decap_8
XFILLER_7_550 VPWR VGND sg13g2_decap_8
XFILLER_98_844 VPWR VGND sg13g2_decap_8
XFILLER_97_343 VPWR VGND sg13g2_decap_8
XFILLER_44_1028 VPWR VGND sg13g2_fill_1
XFILLER_100_805 VPWR VGND sg13g2_decap_8
XFILLER_25_0 VPWR VGND sg13g2_decap_8
XFILLER_39_900 VPWR VGND sg13g2_decap_8
XFILLER_66_741 VPWR VGND sg13g2_decap_8
XFILLER_54_914 VPWR VGND sg13g2_decap_8
XFILLER_39_977 VPWR VGND sg13g2_decap_8
XFILLER_93_593 VPWR VGND sg13g2_decap_8
XFILLER_81_711 VPWR VGND sg13g2_decap_8
XFILLER_65_273 VPWR VGND sg13g2_decap_8
XFILLER_53_413 VPWR VGND sg13g2_decap_8
XFILLER_26_616 VPWR VGND sg13g2_decap_8
XFILLER_38_476 VPWR VGND sg13g2_decap_8
XFILLER_80_210 VPWR VGND sg13g2_decap_8
XFILLER_25_126 VPWR VGND sg13g2_decap_8
XFILLER_81_788 VPWR VGND sg13g2_decap_8
XFILLER_62_980 VPWR VGND sg13g2_decap_8
XFILLER_90_1026 VPWR VGND sg13g2_fill_2
XFILLER_80_287 VPWR VGND sg13g2_decap_8
XFILLER_22_844 VPWR VGND sg13g2_decap_8
XFILLER_21_343 VPWR VGND sg13g2_decap_8
XFILLER_103_7 VPWR VGND sg13g2_decap_8
XFILLER_89_833 VPWR VGND sg13g2_decap_8
XFILLER_0_203 VPWR VGND sg13g2_decap_8
XFILLER_103_665 VPWR VGND sg13g2_decap_8
XFILLER_88_354 VPWR VGND sg13g2_decap_8
XFILLER_102_175 VPWR VGND sg13g2_decap_8
XFILLER_29_410 VPWR VGND sg13g2_decap_8
XFILLER_57_763 VPWR VGND sg13g2_decap_8
XFILLER_45_903 VPWR VGND sg13g2_decap_8
XFILLER_84_560 VPWR VGND sg13g2_decap_8
XFILLER_72_700 VPWR VGND sg13g2_decap_8
XFILLER_56_67 VPWR VGND sg13g2_decap_8
XFILLER_17_627 VPWR VGND sg13g2_decap_8
XFILLER_29_487 VPWR VGND sg13g2_decap_8
XFILLER_71_221 VPWR VGND sg13g2_decap_8
XFILLER_56_284 VPWR VGND sg13g2_decap_8
XFILLER_44_424 VPWR VGND sg13g2_decap_8
XFILLER_16_126 VPWR VGND sg13g2_decap_8
XFILLER_72_777 VPWR VGND sg13g2_decap_8
XFILLER_60_928 VPWR VGND sg13g2_decap_8
XFILLER_53_980 VPWR VGND sg13g2_decap_8
XFILLER_72_77 VPWR VGND sg13g2_decap_8
XFILLER_71_298 VPWR VGND sg13g2_decap_8
XFILLER_52_490 VPWR VGND sg13g2_decap_8
XFILLER_13_833 VPWR VGND sg13g2_decap_8
XFILLER_25_693 VPWR VGND sg13g2_decap_8
XFILLER_40_630 VPWR VGND sg13g2_decap_8
XFILLER_9_826 VPWR VGND sg13g2_decap_8
XFILLER_12_354 VPWR VGND sg13g2_decap_8
XFILLER_8_336 VPWR VGND sg13g2_decap_8
XFILLER_21_70 VPWR VGND sg13g2_decap_8
XFILLER_4_553 VPWR VGND sg13g2_decap_8
XFILLER_97_63 VPWR VGND sg13g2_decap_8
XFILLER_79_354 VPWR VGND sg13g2_decap_8
XFILLER_39_207 VPWR VGND sg13g2_decap_8
XFILLER_95_858 VPWR VGND sg13g2_decap_8
XFILLER_0_770 VPWR VGND sg13g2_decap_8
XFILLER_94_357 VPWR VGND sg13g2_decap_8
XFILLER_48_763 VPWR VGND sg13g2_decap_8
XFILLER_36_903 VPWR VGND sg13g2_decap_8
XFILLER_75_560 VPWR VGND sg13g2_decap_8
XFILLER_63_700 VPWR VGND sg13g2_decap_8
XFILLER_47_273 VPWR VGND sg13g2_decap_8
XFILLER_35_413 VPWR VGND sg13g2_decap_8
XFILLER_62_210 VPWR VGND sg13g2_decap_8
XFILLER_63_777 VPWR VGND sg13g2_decap_8
XFILLER_51_928 VPWR VGND sg13g2_decap_8
XFILLER_90_585 VPWR VGND sg13g2_decap_8
XFILLER_62_287 VPWR VGND sg13g2_decap_8
XFILLER_50_427 VPWR VGND sg13g2_decap_8
XFILLER_44_991 VPWR VGND sg13g2_decap_8
XFILLER_16_693 VPWR VGND sg13g2_decap_8
XFILLER_43_490 VPWR VGND sg13g2_decap_8
XFILLER_31_630 VPWR VGND sg13g2_decap_8
XFILLER_30_140 VPWR VGND sg13g2_decap_8
XFILLER_98_641 VPWR VGND sg13g2_decap_8
XFILLER_100_602 VPWR VGND sg13g2_decap_8
XFILLER_97_140 VPWR VGND sg13g2_decap_8
XFILLER_86_858 VPWR VGND sg13g2_decap_8
XFILLER_85_357 VPWR VGND sg13g2_decap_8
XFILLER_73_508 VPWR VGND sg13g2_decap_8
XFILLER_100_679 VPWR VGND sg13g2_decap_8
XFILLER_54_711 VPWR VGND sg13g2_decap_8
XFILLER_26_413 VPWR VGND sg13g2_decap_8
XFILLER_27_914 VPWR VGND sg13g2_decap_8
XFILLER_38_273 VPWR VGND sg13g2_decap_8
XFILLER_39_774 VPWR VGND sg13g2_decap_8
XFILLER_93_390 VPWR VGND sg13g2_decap_8
XFILLER_53_210 VPWR VGND sg13g2_decap_8
XFILLER_54_788 VPWR VGND sg13g2_decap_8
XFILLER_42_928 VPWR VGND sg13g2_decap_8
XFILLER_81_585 VPWR VGND sg13g2_decap_8
XFILLER_53_287 VPWR VGND sg13g2_decap_8
XFILLER_35_980 VPWR VGND sg13g2_decap_8
XFILLER_41_427 VPWR VGND sg13g2_decap_8
XFILLER_42_25 VPWR VGND sg13g2_decap_8
XFILLER_22_641 VPWR VGND sg13g2_decap_8
XFILLER_50_994 VPWR VGND sg13g2_decap_8
XFILLER_21_140 VPWR VGND sg13g2_decap_8
XFILLER_10_858 VPWR VGND sg13g2_decap_8
XFILLER_89_630 VPWR VGND sg13g2_decap_8
XFILLER_27_1012 VPWR VGND sg13g2_decap_8
XFILLER_104_952 VPWR VGND sg13g2_decap_8
XFILLER_88_151 VPWR VGND sg13g2_decap_8
XFILLER_1_567 VPWR VGND sg13g2_decap_8
XFILLER_103_462 VPWR VGND sg13g2_decap_8
XFILLER_77_847 VPWR VGND sg13g2_decap_8
XFILLER_67_55 VPWR VGND sg13g2_fill_2
XFILLER_67_33 VPWR VGND sg13g2_fill_1
XFILLER_76_368 VPWR VGND sg13g2_decap_8
XFILLER_67_77 VPWR VGND sg13g2_decap_8
XFILLER_64_508 VPWR VGND sg13g2_decap_8
XFILLER_18_903 VPWR VGND sg13g2_decap_8
XFILLER_57_560 VPWR VGND sg13g2_decap_8
XFILLER_45_700 VPWR VGND sg13g2_decap_8
XFILLER_83_32 VPWR VGND sg13g2_decap_8
XFILLER_44_221 VPWR VGND sg13g2_decap_8
XFILLER_17_424 VPWR VGND sg13g2_decap_8
XFILLER_29_284 VPWR VGND sg13g2_decap_8
XFILLER_72_574 VPWR VGND sg13g2_decap_8
XFILLER_45_777 VPWR VGND sg13g2_decap_8
XFILLER_33_917 VPWR VGND sg13g2_decap_8
XFILLER_60_725 VPWR VGND sg13g2_decap_8
XFILLER_44_298 VPWR VGND sg13g2_decap_8
XFILLER_16_70 VPWR VGND sg13g2_decap_8
XFILLER_26_980 VPWR VGND sg13g2_decap_8
XFILLER_32_438 VPWR VGND sg13g2_decap_8
XFILLER_13_630 VPWR VGND sg13g2_decap_8
XFILLER_25_490 VPWR VGND sg13g2_decap_8
XFILLER_34_1005 VPWR VGND sg13g2_decap_8
XFILLER_41_994 VPWR VGND sg13g2_decap_8
XFILLER_9_623 VPWR VGND sg13g2_decap_8
XFILLER_12_151 VPWR VGND sg13g2_decap_8
XFILLER_8_133 VPWR VGND sg13g2_decap_8
XFILLER_5_851 VPWR VGND sg13g2_decap_8
XFILLER_99_427 VPWR VGND sg13g2_decap_8
XFILLER_4_350 VPWR VGND sg13g2_decap_8
XFILLER_79_151 VPWR VGND sg13g2_decap_8
XFILLER_68_803 VPWR VGND sg13g2_decap_8
XFILLER_95_655 VPWR VGND sg13g2_decap_8
XFILLER_67_357 VPWR VGND sg13g2_decap_8
XFILLER_94_154 VPWR VGND sg13g2_decap_8
XFILLER_48_560 VPWR VGND sg13g2_decap_8
XFILLER_36_700 VPWR VGND sg13g2_decap_8
XFILLER_35_210 VPWR VGND sg13g2_decap_8
XFILLER_91_861 VPWR VGND sg13g2_decap_8
XFILLER_63_574 VPWR VGND sg13g2_decap_8
XFILLER_24_928 VPWR VGND sg13g2_decap_8
XFILLER_36_777 VPWR VGND sg13g2_decap_8
XFILLER_90_382 VPWR VGND sg13g2_decap_8
XFILLER_51_725 VPWR VGND sg13g2_decap_8
XFILLER_50_224 VPWR VGND sg13g2_decap_8
XFILLER_17_991 VPWR VGND sg13g2_decap_8
XFILLER_23_427 VPWR VGND sg13g2_decap_8
XFILLER_35_287 VPWR VGND sg13g2_decap_8
XFILLER_92_0 VPWR VGND sg13g2_decap_8
XFILLER_16_490 VPWR VGND sg13g2_decap_8
XFILLER_12_39 VPWR VGND sg13g2_decap_8
XFILLER_105_749 VPWR VGND sg13g2_decap_8
XFILLER_104_259 VPWR VGND sg13g2_decap_8
XFILLER_59_803 VPWR VGND sg13g2_decap_8
XFILLER_99_994 VPWR VGND sg13g2_decap_8
XFILLER_101_966 VPWR VGND sg13g2_decap_8
XFILLER_86_655 VPWR VGND sg13g2_decap_8
XFILLER_74_806 VPWR VGND sg13g2_decap_8
XFILLER_58_357 VPWR VGND sg13g2_decap_8
XFILLER_100_476 VPWR VGND sg13g2_decap_8
XFILLER_85_154 VPWR VGND sg13g2_decap_8
XFILLER_73_305 VPWR VGND sg13g2_decap_8
XFILLER_46_508 VPWR VGND sg13g2_decap_8
XFILLER_27_711 VPWR VGND sg13g2_decap_8
XFILLER_37_25 VPWR VGND sg13g2_decap_8
XFILLER_39_571 VPWR VGND sg13g2_decap_8
XFILLER_26_210 VPWR VGND sg13g2_decap_8
XFILLER_82_861 VPWR VGND sg13g2_decap_8
XFILLER_15_928 VPWR VGND sg13g2_decap_8
XFILLER_27_788 VPWR VGND sg13g2_decap_8
XFILLER_81_382 VPWR VGND sg13g2_decap_8
XFILLER_54_585 VPWR VGND sg13g2_decap_8
XFILLER_53_35 VPWR VGND sg13g2_decap_8
XFILLER_42_725 VPWR VGND sg13g2_decap_8
XFILLER_14_427 VPWR VGND sg13g2_decap_8
XFILLER_26_287 VPWR VGND sg13g2_decap_8
XFILLER_41_224 VPWR VGND sg13g2_decap_8
XFILLER_23_994 VPWR VGND sg13g2_decap_8
XFILLER_50_791 VPWR VGND sg13g2_decap_8
XFILLER_10_655 VPWR VGND sg13g2_decap_8
XFILLER_6_637 VPWR VGND sg13g2_decap_8
XFILLER_5_158 VPWR VGND sg13g2_decap_8
XFILLER_78_32 VPWR VGND sg13g2_decap_8
XFILLER_78_76 VPWR VGND sg13g2_decap_8
XFILLER_2_865 VPWR VGND sg13g2_decap_8
XFILLER_1_364 VPWR VGND sg13g2_decap_8
XFILLER_77_644 VPWR VGND sg13g2_decap_8
XFILLER_94_42 VPWR VGND sg13g2_decap_8
XFILLER_76_165 VPWR VGND sg13g2_decap_8
XFILLER_64_305 VPWR VGND sg13g2_decap_8
XFILLER_49_368 VPWR VGND sg13g2_decap_8
XFILLER_18_700 VPWR VGND sg13g2_decap_8
XFILLER_37_508 VPWR VGND sg13g2_decap_8
XFILLER_92_658 VPWR VGND sg13g2_decap_8
XFILLER_17_221 VPWR VGND sg13g2_decap_8
XFILLER_91_168 VPWR VGND sg13g2_decap_8
XFILLER_73_872 VPWR VGND sg13g2_decap_8
XFILLER_18_777 VPWR VGND sg13g2_decap_8
XFILLER_72_371 VPWR VGND sg13g2_decap_8
XFILLER_60_522 VPWR VGND sg13g2_decap_8
XFILLER_45_574 VPWR VGND sg13g2_decap_8
XFILLER_33_714 VPWR VGND sg13g2_decap_8
XFILLER_17_298 VPWR VGND sg13g2_decap_8
XFILLER_32_235 VPWR VGND sg13g2_decap_8
XFILLER_60_599 VPWR VGND sg13g2_decap_8
XFILLER_14_994 VPWR VGND sg13g2_decap_8
XFILLER_41_791 VPWR VGND sg13g2_decap_8
XFILLER_9_420 VPWR VGND sg13g2_decap_8
XFILLER_64_4 VPWR VGND sg13g2_decap_8
XFILLER_9_497 VPWR VGND sg13g2_decap_8
XFILLER_99_224 VPWR VGND sg13g2_decap_8
XFILLER_96_931 VPWR VGND sg13g2_decap_8
XFILLER_68_600 VPWR VGND sg13g2_decap_8
XFILLER_4_84 VPWR VGND sg13g2_decap_8
XFILLER_95_452 VPWR VGND sg13g2_decap_8
XFILLER_68_677 VPWR VGND sg13g2_decap_8
XFILLER_67_154 VPWR VGND sg13g2_decap_8
XFILLER_83_669 VPWR VGND sg13g2_decap_8
XFILLER_82_168 VPWR VGND sg13g2_decap_8
XFILLER_71_809 VPWR VGND sg13g2_decap_8
XFILLER_70_308 VPWR VGND sg13g2_decap_8
XFILLER_64_872 VPWR VGND sg13g2_decap_8
XFILLER_63_371 VPWR VGND sg13g2_decap_8
XFILLER_51_522 VPWR VGND sg13g2_decap_8
XFILLER_24_725 VPWR VGND sg13g2_decap_8
XFILLER_36_574 VPWR VGND sg13g2_decap_8
XFILLER_23_224 VPWR VGND sg13g2_decap_8
XFILLER_51_599 VPWR VGND sg13g2_decap_8
XFILLER_20_942 VPWR VGND sg13g2_decap_8
XFILLER_23_49 VPWR VGND sg13g2_decap_8
XFILLER_105_546 VPWR VGND sg13g2_decap_8
XFILLER_99_791 VPWR VGND sg13g2_decap_8
XFILLER_87_931 VPWR VGND sg13g2_decap_8
XFILLER_78_419 VPWR VGND sg13g2_decap_8
XFILLER_59_600 VPWR VGND sg13g2_decap_8
XFILLER_48_35 VPWR VGND sg13g2_decap_8
XFILLER_24_1026 VPWR VGND sg13g2_fill_2
XFILLER_101_763 VPWR VGND sg13g2_decap_8
XFILLER_86_452 VPWR VGND sg13g2_decap_8
XFILLER_74_603 VPWR VGND sg13g2_decap_8
XFILLER_59_677 VPWR VGND sg13g2_decap_8
XFILLER_58_154 VPWR VGND sg13g2_decap_8
XFILLER_46_305 VPWR VGND sg13g2_decap_8
XFILLER_104_63 VPWR VGND sg13g2_decap_8
XFILLER_100_273 VPWR VGND sg13g2_decap_8
XFILLER_73_102 VPWR VGND sg13g2_decap_8
XFILLER_55_861 VPWR VGND sg13g2_decap_8
XFILLER_73_179 VPWR VGND sg13g2_decap_8
XFILLER_64_67 VPWR VGND sg13g2_decap_8
XFILLER_61_319 VPWR VGND sg13g2_decap_8
XFILLER_54_382 VPWR VGND sg13g2_decap_8
XFILLER_42_522 VPWR VGND sg13g2_decap_8
XFILLER_15_725 VPWR VGND sg13g2_decap_8
XFILLER_27_585 VPWR VGND sg13g2_decap_8
XFILLER_14_224 VPWR VGND sg13g2_decap_8
XFILLER_70_875 VPWR VGND sg13g2_decap_8
XFILLER_30_728 VPWR VGND sg13g2_decap_8
XFILLER_42_599 VPWR VGND sg13g2_decap_8
XFILLER_11_931 VPWR VGND sg13g2_decap_8
XFILLER_23_791 VPWR VGND sg13g2_decap_8
XFILLER_80_77 VPWR VGND sg13g2_decap_8
XFILLER_10_452 VPWR VGND sg13g2_decap_8
XFILLER_7_935 VPWR VGND sg13g2_decap_8
XFILLER_31_1008 VPWR VGND sg13g2_decap_8
XFILLER_6_434 VPWR VGND sg13g2_decap_8
XFILLER_89_42 VPWR VGND sg13g2_decap_8
XFILLER_97_728 VPWR VGND sg13g2_decap_8
XFILLER_2_662 VPWR VGND sg13g2_decap_8
XFILLER_1_161 VPWR VGND sg13g2_decap_8
XFILLER_96_238 VPWR VGND sg13g2_decap_8
XFILLER_77_441 VPWR VGND sg13g2_decap_8
XFILLER_93_901 VPWR VGND sg13g2_decap_8
XFILLER_78_986 VPWR VGND sg13g2_decap_8
X_42_ net20 _09_ _10_ VPWR VGND sg13g2_xnor2_1
XFILLER_49_165 VPWR VGND sg13g2_decap_8
XFILLER_37_305 VPWR VGND sg13g2_decap_8
XFILLER_65_658 VPWR VGND sg13g2_decap_8
XFILLER_64_102 VPWR VGND sg13g2_decap_8
XFILLER_93_978 VPWR VGND sg13g2_decap_8
XFILLER_92_455 VPWR VGND sg13g2_decap_8
XFILLER_52_308 VPWR VGND sg13g2_decap_8
XFILLER_64_179 VPWR VGND sg13g2_decap_8
XFILLER_46_872 VPWR VGND sg13g2_decap_8
XFILLER_45_371 VPWR VGND sg13g2_decap_8
XFILLER_18_574 VPWR VGND sg13g2_decap_8
XFILLER_33_511 VPWR VGND sg13g2_decap_8
XFILLER_61_886 VPWR VGND sg13g2_decap_8
XFILLER_21_728 VPWR VGND sg13g2_decap_8
XFILLER_33_588 VPWR VGND sg13g2_decap_8
XFILLER_60_396 VPWR VGND sg13g2_decap_8
XFILLER_14_791 VPWR VGND sg13g2_decap_8
XFILLER_20_249 VPWR VGND sg13g2_decap_8
XFILLER_9_294 VPWR VGND sg13g2_decap_8
XFILLER_55_0 VPWR VGND sg13g2_decap_8
XFILLER_47_1015 VPWR VGND sg13g2_decap_8
XFILLER_88_739 VPWR VGND sg13g2_decap_8
XFILLER_87_238 VPWR VGND sg13g2_decap_8
XFILLER_69_953 VPWR VGND sg13g2_decap_8
XFILLER_68_474 VPWR VGND sg13g2_decap_8
XFILLER_84_945 VPWR VGND sg13g2_decap_8
XFILLER_18_49 VPWR VGND sg13g2_decap_8
XFILLER_83_466 VPWR VGND sg13g2_decap_8
XFILLER_71_606 VPWR VGND sg13g2_decap_8
XFILLER_56_669 VPWR VGND sg13g2_decap_8
XFILLER_44_809 VPWR VGND sg13g2_decap_8
XFILLER_43_308 VPWR VGND sg13g2_decap_8
XFILLER_93_1013 VPWR VGND sg13g2_decap_8
XFILLER_70_105 VPWR VGND sg13g2_decap_8
XFILLER_55_168 VPWR VGND sg13g2_decap_8
XFILLER_36_371 VPWR VGND sg13g2_decap_8
XFILLER_37_872 VPWR VGND sg13g2_decap_8
XFILLER_24_522 VPWR VGND sg13g2_decap_8
XFILLER_54_1019 VPWR VGND sg13g2_decap_8
XFILLER_52_875 VPWR VGND sg13g2_decap_8
XFILLER_51_396 VPWR VGND sg13g2_decap_8
XFILLER_11_238 VPWR VGND sg13g2_decap_8
XFILLER_12_739 VPWR VGND sg13g2_decap_8
XFILLER_24_599 VPWR VGND sg13g2_decap_8
XFILLER_50_14 VPWR VGND sg13g2_decap_8
XFILLER_106_833 VPWR VGND sg13g2_decap_8
XFILLER_4_938 VPWR VGND sg13g2_decap_8
XFILLER_105_343 VPWR VGND sg13g2_decap_8
XFILLER_3_448 VPWR VGND sg13g2_decap_8
XFILLER_79_739 VPWR VGND sg13g2_decap_8
XFILLER_78_216 VPWR VGND sg13g2_decap_8
XFILLER_59_67 VPWR VGND sg13g2_decap_4
XFILLER_101_560 VPWR VGND sg13g2_decap_8
XFILLER_93_208 VPWR VGND sg13g2_decap_8
XFILLER_59_474 VPWR VGND sg13g2_decap_8
XFILLER_75_945 VPWR VGND sg13g2_decap_8
XFILLER_74_400 VPWR VGND sg13g2_decap_8
XFILLER_46_102 VPWR VGND sg13g2_decap_8
XFILLER_75_77 VPWR VGND sg13g2_decap_8
XFILLER_47_658 VPWR VGND sg13g2_decap_8
XFILLER_28_861 VPWR VGND sg13g2_decap_8
XFILLER_74_477 VPWR VGND sg13g2_decap_8
XFILLER_61_116 VPWR VGND sg13g2_decap_8
XFILLER_46_179 VPWR VGND sg13g2_decap_8
XFILLER_34_319 VPWR VGND sg13g2_decap_8
XFILLER_91_21 VPWR VGND sg13g2_decap_8
XFILLER_15_522 VPWR VGND sg13g2_decap_8
XFILLER_27_382 VPWR VGND sg13g2_decap_8
XFILLER_70_672 VPWR VGND sg13g2_decap_8
XFILLER_43_875 VPWR VGND sg13g2_decap_8
XFILLER_91_98 VPWR VGND sg13g2_decap_8
XFILLER_42_396 VPWR VGND sg13g2_decap_8
XFILLER_15_599 VPWR VGND sg13g2_decap_8
XFILLER_30_525 VPWR VGND sg13g2_decap_8
XFILLER_24_81 VPWR VGND sg13g2_decap_8
XFILLER_7_732 VPWR VGND sg13g2_decap_8
XFILLER_6_231 VPWR VGND sg13g2_decap_8
XFILLER_40_91 VPWR VGND sg13g2_decap_8
XFILLER_97_525 VPWR VGND sg13g2_decap_8
XFILLER_66_923 VPWR VGND sg13g2_decap_8
XFILLER_27_4 VPWR VGND sg13g2_decap_8
XFILLER_78_783 VPWR VGND sg13g2_decap_8
XFILLER_37_102 VPWR VGND sg13g2_decap_8
XFILLER_93_775 VPWR VGND sg13g2_decap_8
XFILLER_92_252 VPWR VGND sg13g2_decap_8
XFILLER_77_1008 VPWR VGND sg13g2_decap_8
XFILLER_65_455 VPWR VGND sg13g2_decap_8
XFILLER_1_63 VPWR VGND sg13g2_decap_8
XFILLER_19_861 VPWR VGND sg13g2_decap_8
XFILLER_38_658 VPWR VGND sg13g2_decap_8
XFILLER_52_105 VPWR VGND sg13g2_decap_8
XFILLER_18_371 VPWR VGND sg13g2_decap_8
XFILLER_25_308 VPWR VGND sg13g2_decap_8
XFILLER_37_179 VPWR VGND sg13g2_decap_8
XFILLER_80_469 VPWR VGND sg13g2_decap_8
XFILLER_34_886 VPWR VGND sg13g2_decap_8
XFILLER_61_683 VPWR VGND sg13g2_decap_8
XFILLER_21_525 VPWR VGND sg13g2_decap_8
XFILLER_33_385 VPWR VGND sg13g2_decap_8
XFILLER_60_193 VPWR VGND sg13g2_decap_8
XFILLER_20_39 VPWR VGND sg13g2_decap_8
XFILLER_103_847 VPWR VGND sg13g2_decap_8
XFILLER_88_536 VPWR VGND sg13g2_decap_8
XFILLER_102_357 VPWR VGND sg13g2_decap_8
XFILLER_69_750 VPWR VGND sg13g2_decap_8
XFILLER_60_1012 VPWR VGND sg13g2_decap_8
XFILLER_68_271 VPWR VGND sg13g2_decap_8
XFILLER_57_945 VPWR VGND sg13g2_decap_8
XFILLER_84_742 VPWR VGND sg13g2_decap_8
XFILLER_56_466 VPWR VGND sg13g2_decap_8
XFILLER_44_606 VPWR VGND sg13g2_decap_8
XFILLER_17_809 VPWR VGND sg13g2_decap_8
XFILLER_29_669 VPWR VGND sg13g2_decap_8
XFILLER_83_263 VPWR VGND sg13g2_decap_8
XFILLER_71_403 VPWR VGND sg13g2_decap_8
XFILLER_45_14 VPWR VGND sg13g2_decap_8
XFILLER_43_105 VPWR VGND sg13g2_decap_8
XFILLER_16_308 VPWR VGND sg13g2_decap_8
XFILLER_28_168 VPWR VGND sg13g2_decap_8
XFILLER_72_959 VPWR VGND sg13g2_decap_8
XFILLER_101_42 VPWR VGND sg13g2_decap_8
XFILLER_52_672 VPWR VGND sg13g2_decap_8
XFILLER_25_875 VPWR VGND sg13g2_decap_8
XFILLER_40_812 VPWR VGND sg13g2_decap_8
XFILLER_61_13 VPWR VGND sg13g2_fill_1
XFILLER_12_536 VPWR VGND sg13g2_decap_8
XFILLER_24_396 VPWR VGND sg13g2_decap_8
XFILLER_61_68 VPWR VGND sg13g2_fill_2
XFILLER_51_193 VPWR VGND sg13g2_decap_8
XFILLER_8_518 VPWR VGND sg13g2_decap_8
XFILLER_40_889 VPWR VGND sg13g2_decap_8
XFILLER_4_735 VPWR VGND sg13g2_decap_8
XFILLER_106_630 VPWR VGND sg13g2_decap_8
XFILLER_3_245 VPWR VGND sg13g2_decap_8
XFILLER_105_140 VPWR VGND sg13g2_decap_8
XFILLER_79_536 VPWR VGND sg13g2_decap_8
XFILLER_86_32 VPWR VGND sg13g2_decap_8
XFILLER_0_952 VPWR VGND sg13g2_decap_8
XFILLER_94_539 VPWR VGND sg13g2_decap_8
XFILLER_59_271 VPWR VGND sg13g2_decap_8
XFILLER_48_945 VPWR VGND sg13g2_decap_8
XFILLER_75_742 VPWR VGND sg13g2_decap_8
XFILLER_47_455 VPWR VGND sg13g2_decap_8
XFILLER_19_70 VPWR VGND sg13g2_decap_8
XFILLER_74_274 VPWR VGND sg13g2_decap_8
XFILLER_19_168 VPWR VGND sg13g2_decap_8
XFILLER_90_767 VPWR VGND sg13g2_decap_8
XFILLER_63_959 VPWR VGND sg13g2_decap_8
XFILLER_34_116 VPWR VGND sg13g2_decap_8
XFILLER_71_970 VPWR VGND sg13g2_decap_8
XFILLER_62_469 VPWR VGND sg13g2_decap_8
XFILLER_50_609 VPWR VGND sg13g2_decap_8
XFILLER_43_672 VPWR VGND sg13g2_decap_8
XFILLER_16_875 VPWR VGND sg13g2_decap_8
XFILLER_31_812 VPWR VGND sg13g2_decap_8
XFILLER_96_7 VPWR VGND sg13g2_decap_8
XFILLER_15_396 VPWR VGND sg13g2_decap_8
XFILLER_30_322 VPWR VGND sg13g2_decap_8
XFILLER_35_91 VPWR VGND sg13g2_decap_8
XFILLER_42_193 VPWR VGND sg13g2_decap_8
XFILLER_31_889 VPWR VGND sg13g2_decap_8
XFILLER_30_399 VPWR VGND sg13g2_decap_8
XFILLER_98_823 VPWR VGND sg13g2_decap_8
XFILLER_83_1012 VPWR VGND sg13g2_decap_8
XFILLER_97_322 VPWR VGND sg13g2_decap_8
XFILLER_97_399 VPWR VGND sg13g2_decap_8
XFILLER_85_539 VPWR VGND sg13g2_decap_8
XFILLER_78_580 VPWR VGND sg13g2_decap_8
XFILLER_66_720 VPWR VGND sg13g2_decap_8
XFILLER_18_0 VPWR VGND sg13g2_decap_8
XFILLER_38_455 VPWR VGND sg13g2_decap_8
XFILLER_39_956 VPWR VGND sg13g2_decap_8
XFILLER_93_572 VPWR VGND sg13g2_decap_8
XFILLER_66_797 VPWR VGND sg13g2_decap_8
XFILLER_65_252 VPWR VGND sg13g2_decap_8
XFILLER_25_105 VPWR VGND sg13g2_decap_8
XFILLER_81_767 VPWR VGND sg13g2_decap_8
XFILLER_80_266 VPWR VGND sg13g2_decap_8
XFILLER_53_469 VPWR VGND sg13g2_decap_8
XFILLER_41_609 VPWR VGND sg13g2_decap_8
XFILLER_15_39 VPWR VGND sg13g2_decap_8
XFILLER_90_1005 VPWR VGND sg13g2_decap_8
XFILLER_61_480 VPWR VGND sg13g2_decap_8
XFILLER_22_823 VPWR VGND sg13g2_decap_8
XFILLER_34_683 VPWR VGND sg13g2_decap_8
XFILLER_40_119 VPWR VGND sg13g2_decap_8
XFILLER_21_322 VPWR VGND sg13g2_decap_8
XFILLER_33_182 VPWR VGND sg13g2_decap_8
XFILLER_21_399 VPWR VGND sg13g2_decap_8
XFILLER_31_49 VPWR VGND sg13g2_decap_8
XFILLER_89_812 VPWR VGND sg13g2_decap_8
XFILLER_103_644 VPWR VGND sg13g2_decap_8
XFILLER_88_333 VPWR VGND sg13g2_decap_8
XFILLER_1_749 VPWR VGND sg13g2_decap_8
XFILLER_102_154 VPWR VGND sg13g2_decap_8
XFILLER_89_889 VPWR VGND sg13g2_decap_8
XFILLER_0_259 VPWR VGND sg13g2_decap_8
XFILLER_5_1012 VPWR VGND sg13g2_decap_8
XFILLER_57_742 VPWR VGND sg13g2_decap_8
XFILLER_56_46 VPWR VGND sg13g2_decap_8
XFILLER_71_200 VPWR VGND sg13g2_decap_8
XFILLER_56_263 VPWR VGND sg13g2_decap_8
XFILLER_44_403 VPWR VGND sg13g2_decap_8
XFILLER_16_105 VPWR VGND sg13g2_decap_8
XFILLER_17_606 VPWR VGND sg13g2_decap_8
XFILLER_29_466 VPWR VGND sg13g2_decap_8
XFILLER_72_756 VPWR VGND sg13g2_decap_8
XFILLER_45_959 VPWR VGND sg13g2_decap_8
XFILLER_60_907 VPWR VGND sg13g2_decap_8
XFILLER_72_56 VPWR VGND sg13g2_decap_8
XFILLER_71_277 VPWR VGND sg13g2_decap_8
XFILLER_13_812 VPWR VGND sg13g2_decap_8
XFILLER_25_672 VPWR VGND sg13g2_decap_8
XFILLER_31_119 VPWR VGND sg13g2_decap_8
XFILLER_9_805 VPWR VGND sg13g2_decap_8
XFILLER_12_333 VPWR VGND sg13g2_decap_8
XFILLER_24_193 VPWR VGND sg13g2_decap_8
XFILLER_8_315 VPWR VGND sg13g2_decap_8
XFILLER_13_889 VPWR VGND sg13g2_decap_8
XFILLER_40_686 VPWR VGND sg13g2_decap_8
XFILLER_99_609 VPWR VGND sg13g2_decap_8
XFILLER_4_532 VPWR VGND sg13g2_decap_8
XFILLER_97_42 VPWR VGND sg13g2_decap_8
XFILLER_79_333 VPWR VGND sg13g2_decap_8
XFILLER_95_837 VPWR VGND sg13g2_decap_8
XFILLER_67_539 VPWR VGND sg13g2_decap_8
XFILLER_94_336 VPWR VGND sg13g2_decap_8
XFILLER_48_742 VPWR VGND sg13g2_decap_8
XFILLER_11_7 VPWR VGND sg13g2_decap_8
XFILLER_47_252 VPWR VGND sg13g2_decap_8
XFILLER_63_756 VPWR VGND sg13g2_decap_8
XFILLER_36_959 VPWR VGND sg13g2_decap_8
XFILLER_90_564 VPWR VGND sg13g2_decap_8
XFILLER_62_266 VPWR VGND sg13g2_decap_8
XFILLER_51_907 VPWR VGND sg13g2_decap_8
XFILLER_50_406 VPWR VGND sg13g2_decap_8
XFILLER_44_970 VPWR VGND sg13g2_decap_8
XFILLER_23_609 VPWR VGND sg13g2_decap_8
XFILLER_35_469 VPWR VGND sg13g2_decap_8
XFILLER_16_672 VPWR VGND sg13g2_decap_8
XFILLER_15_193 VPWR VGND sg13g2_decap_8
XFILLER_31_686 VPWR VGND sg13g2_decap_8
XFILLER_50_1022 VPWR VGND sg13g2_decap_8
XFILLER_30_196 VPWR VGND sg13g2_decap_8
XFILLER_8_882 VPWR VGND sg13g2_decap_8
XFILLER_7_95 VPWR VGND sg13g2_decap_8
XFILLER_89_119 VPWR VGND sg13g2_decap_8
XFILLER_98_620 VPWR VGND sg13g2_decap_8
XFILLER_98_697 VPWR VGND sg13g2_decap_8
XFILLER_86_837 VPWR VGND sg13g2_decap_8
XFILLER_58_539 VPWR VGND sg13g2_decap_8
XFILLER_100_658 VPWR VGND sg13g2_decap_8
XFILLER_97_196 VPWR VGND sg13g2_decap_8
XFILLER_85_336 VPWR VGND sg13g2_decap_8
XFILLER_39_753 VPWR VGND sg13g2_decap_8
XFILLER_38_252 VPWR VGND sg13g2_decap_8
XFILLER_66_594 VPWR VGND sg13g2_decap_8
XFILLER_81_564 VPWR VGND sg13g2_decap_8
XFILLER_54_767 VPWR VGND sg13g2_decap_8
XFILLER_53_266 VPWR VGND sg13g2_decap_8
XFILLER_42_907 VPWR VGND sg13g2_decap_8
XFILLER_14_609 VPWR VGND sg13g2_decap_8
XFILLER_26_49 VPWR VGND sg13g2_decap_8
XFILLER_26_469 VPWR VGND sg13g2_decap_8
XFILLER_41_406 VPWR VGND sg13g2_decap_8
XFILLER_13_119 VPWR VGND sg13g2_decap_8
XFILLER_22_620 VPWR VGND sg13g2_decap_8
XFILLER_34_480 VPWR VGND sg13g2_decap_8
XFILLER_50_973 VPWR VGND sg13g2_decap_8
XFILLER_6_819 VPWR VGND sg13g2_decap_8
XFILLER_10_837 VPWR VGND sg13g2_decap_8
XFILLER_21_196 VPWR VGND sg13g2_decap_8
XFILLER_22_697 VPWR VGND sg13g2_decap_8
XFILLER_104_931 VPWR VGND sg13g2_decap_8
XFILLER_103_441 VPWR VGND sg13g2_decap_8
XFILLER_88_130 VPWR VGND sg13g2_decap_8
XFILLER_1_546 VPWR VGND sg13g2_decap_8
XFILLER_89_686 VPWR VGND sg13g2_decap_8
XFILLER_77_826 VPWR VGND sg13g2_decap_8
XFILLER_67_45 VPWR VGND sg13g2_fill_2
XFILLER_76_347 VPWR VGND sg13g2_decap_8
XFILLER_17_403 VPWR VGND sg13g2_decap_8
XFILLER_29_263 VPWR VGND sg13g2_decap_8
XFILLER_83_11 VPWR VGND sg13g2_decap_8
XFILLER_44_200 VPWR VGND sg13g2_decap_8
XFILLER_18_959 VPWR VGND sg13g2_decap_8
XFILLER_72_553 VPWR VGND sg13g2_decap_8
XFILLER_60_704 VPWR VGND sg13g2_decap_8
XFILLER_45_756 VPWR VGND sg13g2_decap_8
XFILLER_83_88 VPWR VGND sg13g2_decap_8
XFILLER_44_277 VPWR VGND sg13g2_decap_8
XFILLER_32_417 VPWR VGND sg13g2_decap_8
XFILLER_9_602 VPWR VGND sg13g2_decap_8
XFILLER_41_973 VPWR VGND sg13g2_decap_8
XFILLER_8_112 VPWR VGND sg13g2_decap_8
XFILLER_12_130 VPWR VGND sg13g2_decap_8
XFILLER_13_686 VPWR VGND sg13g2_decap_8
XFILLER_34_1028 VPWR VGND sg13g2_fill_1
XFILLER_40_483 VPWR VGND sg13g2_decap_8
XFILLER_9_679 VPWR VGND sg13g2_decap_8
XFILLER_32_81 VPWR VGND sg13g2_decap_8
XFILLER_8_189 VPWR VGND sg13g2_decap_8
XFILLER_5_830 VPWR VGND sg13g2_decap_8
XFILLER_99_406 VPWR VGND sg13g2_decap_8
XFILLER_80_1015 VPWR VGND sg13g2_decap_8
XFILLER_79_130 VPWR VGND sg13g2_decap_8
XFILLER_95_634 VPWR VGND sg13g2_decap_8
XFILLER_94_133 VPWR VGND sg13g2_decap_8
XFILLER_68_859 VPWR VGND sg13g2_decap_8
XFILLER_67_336 VPWR VGND sg13g2_decap_8
XFILLER_91_840 VPWR VGND sg13g2_decap_8
XFILLER_63_553 VPWR VGND sg13g2_decap_8
XFILLER_51_704 VPWR VGND sg13g2_decap_8
XFILLER_24_907 VPWR VGND sg13g2_decap_8
XFILLER_36_756 VPWR VGND sg13g2_decap_8
XFILLER_90_361 VPWR VGND sg13g2_decap_8
XFILLER_50_203 VPWR VGND sg13g2_decap_8
XFILLER_17_970 VPWR VGND sg13g2_decap_8
XFILLER_23_406 VPWR VGND sg13g2_decap_8
XFILLER_35_266 VPWR VGND sg13g2_decap_8
XFILLER_85_0 VPWR VGND sg13g2_decap_8
XFILLER_32_984 VPWR VGND sg13g2_decap_8
XFILLER_12_18 VPWR VGND sg13g2_decap_8
XFILLER_31_483 VPWR VGND sg13g2_decap_8
XFILLER_105_728 VPWR VGND sg13g2_decap_8
XFILLER_104_238 VPWR VGND sg13g2_decap_8
XFILLER_99_973 VPWR VGND sg13g2_decap_8
XFILLER_101_945 VPWR VGND sg13g2_decap_8
XFILLER_98_494 VPWR VGND sg13g2_decap_8
XFILLER_86_634 VPWR VGND sg13g2_decap_8
XFILLER_85_133 VPWR VGND sg13g2_decap_8
XFILLER_59_859 VPWR VGND sg13g2_decap_8
XFILLER_58_336 VPWR VGND sg13g2_decap_8
XFILLER_100_455 VPWR VGND sg13g2_decap_8
XFILLER_39_550 VPWR VGND sg13g2_decap_8
XFILLER_96_1022 VPWR VGND sg13g2_decap_8
XFILLER_82_840 VPWR VGND sg13g2_decap_8
XFILLER_2_1026 VPWR VGND sg13g2_fill_2
XFILLER_66_391 VPWR VGND sg13g2_decap_8
XFILLER_54_564 VPWR VGND sg13g2_decap_8
XFILLER_42_704 VPWR VGND sg13g2_decap_8
XFILLER_15_907 VPWR VGND sg13g2_decap_8
XFILLER_27_767 VPWR VGND sg13g2_decap_8
XFILLER_81_361 VPWR VGND sg13g2_decap_8
XFILLER_53_14 VPWR VGND sg13g2_decap_8
XFILLER_14_406 VPWR VGND sg13g2_decap_8
XFILLER_26_266 VPWR VGND sg13g2_decap_8
XFILLER_41_203 VPWR VGND sg13g2_decap_8
XFILLER_50_770 VPWR VGND sg13g2_decap_8
XFILLER_23_973 VPWR VGND sg13g2_decap_8
XFILLER_10_634 VPWR VGND sg13g2_decap_8
XFILLER_22_494 VPWR VGND sg13g2_decap_8
XFILLER_6_616 VPWR VGND sg13g2_decap_8
XFILLER_5_137 VPWR VGND sg13g2_decap_8
XFILLER_78_11 VPWR VGND sg13g2_decap_8
XFILLER_2_844 VPWR VGND sg13g2_decap_8
XFILLER_1_343 VPWR VGND sg13g2_decap_8
XFILLER_89_483 VPWR VGND sg13g2_decap_8
XFILLER_77_623 VPWR VGND sg13g2_decap_8
XFILLER_49_347 VPWR VGND sg13g2_decap_8
XFILLER_94_21 VPWR VGND sg13g2_decap_8
XFILLER_76_144 VPWR VGND sg13g2_decap_8
XFILLER_92_637 VPWR VGND sg13g2_decap_8
XFILLER_17_200 VPWR VGND sg13g2_decap_8
XFILLER_94_98 VPWR VGND sg13g2_decap_8
XFILLER_91_147 VPWR VGND sg13g2_decap_8
XFILLER_73_851 VPWR VGND sg13g2_decap_8
XFILLER_45_553 VPWR VGND sg13g2_decap_8
XFILLER_18_756 VPWR VGND sg13g2_decap_8
XFILLER_27_81 VPWR VGND sg13g2_decap_8
XFILLER_72_350 VPWR VGND sg13g2_decap_8
XFILLER_60_501 VPWR VGND sg13g2_decap_8
XFILLER_17_277 VPWR VGND sg13g2_decap_8
XFILLER_32_214 VPWR VGND sg13g2_decap_8
XFILLER_60_578 VPWR VGND sg13g2_decap_8
XFILLER_41_770 VPWR VGND sg13g2_decap_8
XFILLER_14_973 VPWR VGND sg13g2_decap_8
XFILLER_43_91 VPWR VGND sg13g2_decap_8
XFILLER_13_483 VPWR VGND sg13g2_decap_8
XFILLER_40_280 VPWR VGND sg13g2_decap_8
XFILLER_9_476 VPWR VGND sg13g2_decap_8
XFILLER_99_203 VPWR VGND sg13g2_decap_8
XFILLER_96_910 VPWR VGND sg13g2_decap_8
XFILLER_4_63 VPWR VGND sg13g2_decap_8
XFILLER_95_431 VPWR VGND sg13g2_decap_8
XFILLER_68_656 VPWR VGND sg13g2_decap_8
XFILLER_67_133 VPWR VGND sg13g2_decap_8
XFILLER_96_987 VPWR VGND sg13g2_decap_8
XFILLER_83_648 VPWR VGND sg13g2_decap_8
XFILLER_82_147 VPWR VGND sg13g2_decap_8
XFILLER_64_851 VPWR VGND sg13g2_decap_8
XFILLER_24_704 VPWR VGND sg13g2_decap_8
XFILLER_36_553 VPWR VGND sg13g2_decap_8
XFILLER_63_350 VPWR VGND sg13g2_decap_8
XFILLER_51_501 VPWR VGND sg13g2_decap_8
XFILLER_23_203 VPWR VGND sg13g2_decap_8
XFILLER_51_578 VPWR VGND sg13g2_decap_8
XFILLER_17_1012 VPWR VGND sg13g2_decap_8
XFILLER_23_28 VPWR VGND sg13g2_decap_8
XFILLER_104_1015 VPWR VGND sg13g2_decap_8
XFILLER_20_921 VPWR VGND sg13g2_decap_8
XFILLER_31_280 VPWR VGND sg13g2_decap_8
XFILLER_32_781 VPWR VGND sg13g2_decap_8
XFILLER_20_998 VPWR VGND sg13g2_decap_8
XFILLER_105_525 VPWR VGND sg13g2_decap_8
XFILLER_99_770 VPWR VGND sg13g2_decap_8
XFILLER_87_910 VPWR VGND sg13g2_decap_8
XFILLER_48_14 VPWR VGND sg13g2_decap_8
XFILLER_101_742 VPWR VGND sg13g2_decap_8
XFILLER_98_291 VPWR VGND sg13g2_decap_8
XFILLER_86_431 VPWR VGND sg13g2_decap_8
XFILLER_59_656 VPWR VGND sg13g2_decap_8
XFILLER_58_133 VPWR VGND sg13g2_decap_4
XFILLER_24_1005 VPWR VGND sg13g2_decap_8
XFILLER_100_252 VPWR VGND sg13g2_decap_8
XFILLER_87_987 VPWR VGND sg13g2_decap_8
XFILLER_104_42 VPWR VGND sg13g2_decap_8
XFILLER_74_659 VPWR VGND sg13g2_decap_8
XFILLER_73_158 VPWR VGND sg13g2_decap_8
XFILLER_55_840 VPWR VGND sg13g2_decap_8
XFILLER_64_46 VPWR VGND sg13g2_decap_8
XFILLER_54_361 VPWR VGND sg13g2_decap_8
XFILLER_42_501 VPWR VGND sg13g2_decap_8
XFILLER_14_203 VPWR VGND sg13g2_decap_8
XFILLER_15_704 VPWR VGND sg13g2_decap_8
XFILLER_27_564 VPWR VGND sg13g2_decap_8
XFILLER_70_854 VPWR VGND sg13g2_decap_8
XFILLER_42_578 VPWR VGND sg13g2_decap_8
XFILLER_11_910 VPWR VGND sg13g2_decap_8
XFILLER_30_707 VPWR VGND sg13g2_decap_8
XFILLER_80_56 VPWR VGND sg13g2_decap_8
XFILLER_23_770 VPWR VGND sg13g2_decap_8
XFILLER_10_431 VPWR VGND sg13g2_decap_8
XFILLER_7_914 VPWR VGND sg13g2_decap_8
XFILLER_22_291 VPWR VGND sg13g2_decap_8
XFILLER_6_413 VPWR VGND sg13g2_decap_8
XFILLER_11_987 VPWR VGND sg13g2_decap_8
XFILLER_89_21 VPWR VGND sg13g2_decap_8
XFILLER_97_707 VPWR VGND sg13g2_decap_8
XFILLER_89_98 VPWR VGND sg13g2_decap_8
XFILLER_2_641 VPWR VGND sg13g2_decap_8
XFILLER_96_217 VPWR VGND sg13g2_decap_8
XFILLER_1_140 VPWR VGND sg13g2_decap_8
XFILLER_89_280 VPWR VGND sg13g2_decap_8
XFILLER_78_965 VPWR VGND sg13g2_decap_8
XFILLER_77_420 VPWR VGND sg13g2_decap_8
X_41_ _04_ _06_ _10_ VPWR VGND sg13g2_nor2_1
XFILLER_49_144 VPWR VGND sg13g2_decap_8
XFILLER_93_957 VPWR VGND sg13g2_decap_8
XFILLER_92_434 VPWR VGND sg13g2_decap_8
XFILLER_77_497 VPWR VGND sg13g2_decap_8
XFILLER_65_637 VPWR VGND sg13g2_decap_8
XFILLER_64_158 VPWR VGND sg13g2_decap_8
XFILLER_46_851 VPWR VGND sg13g2_decap_8
XFILLER_18_553 VPWR VGND sg13g2_decap_8
XFILLER_38_91 VPWR VGND sg13g2_decap_8
XFILLER_45_350 VPWR VGND sg13g2_decap_8
XFILLER_61_865 VPWR VGND sg13g2_decap_8
XFILLER_21_707 VPWR VGND sg13g2_decap_8
XFILLER_33_567 VPWR VGND sg13g2_decap_8
XFILLER_60_375 VPWR VGND sg13g2_decap_8
XFILLER_14_770 VPWR VGND sg13g2_decap_8
XFILLER_20_228 VPWR VGND sg13g2_decap_8
XFILLER_13_280 VPWR VGND sg13g2_decap_8
XFILLER_9_273 VPWR VGND sg13g2_decap_8
XFILLER_6_980 VPWR VGND sg13g2_decap_8
XFILLER_48_0 VPWR VGND sg13g2_decap_8
XFILLER_88_718 VPWR VGND sg13g2_decap_8
XFILLER_87_217 VPWR VGND sg13g2_decap_8
XFILLER_102_539 VPWR VGND sg13g2_decap_8
XFILLER_69_932 VPWR VGND sg13g2_decap_8
XFILLER_84_924 VPWR VGND sg13g2_decap_8
XFILLER_68_453 VPWR VGND sg13g2_decap_8
XFILLER_96_784 VPWR VGND sg13g2_decap_8
XFILLER_56_648 VPWR VGND sg13g2_decap_8
XFILLER_18_28 VPWR VGND sg13g2_decap_8
XFILLER_83_445 VPWR VGND sg13g2_decap_8
XFILLER_55_147 VPWR VGND sg13g2_decap_8
XFILLER_37_851 VPWR VGND sg13g2_decap_8
XFILLER_24_501 VPWR VGND sg13g2_decap_8
XFILLER_36_350 VPWR VGND sg13g2_decap_8
XFILLER_52_854 VPWR VGND sg13g2_decap_8
XFILLER_12_718 VPWR VGND sg13g2_decap_8
XFILLER_24_578 VPWR VGND sg13g2_decap_8
XFILLER_51_375 VPWR VGND sg13g2_decap_8
XFILLER_11_217 VPWR VGND sg13g2_decap_8
XFILLER_20_795 VPWR VGND sg13g2_decap_8
XFILLER_4_917 VPWR VGND sg13g2_decap_8
XFILLER_106_812 VPWR VGND sg13g2_decap_8
XFILLER_3_427 VPWR VGND sg13g2_decap_8
XFILLER_105_322 VPWR VGND sg13g2_decap_8
XFILLER_106_889 VPWR VGND sg13g2_decap_8
XFILLER_79_718 VPWR VGND sg13g2_decap_8
XFILLER_59_46 VPWR VGND sg13g2_decap_8
XFILLER_105_399 VPWR VGND sg13g2_decap_8
XFILLER_59_453 VPWR VGND sg13g2_decap_8
XFILLER_87_784 VPWR VGND sg13g2_decap_8
XFILLER_75_924 VPWR VGND sg13g2_decap_8
XFILLER_47_637 VPWR VGND sg13g2_decap_8
XFILLER_75_56 VPWR VGND sg13g2_fill_2
XFILLER_74_456 VPWR VGND sg13g2_decap_8
XFILLER_46_158 VPWR VGND sg13g2_decap_8
XFILLER_28_840 VPWR VGND sg13g2_decap_8
XFILLER_90_949 VPWR VGND sg13g2_decap_8
XFILLER_15_501 VPWR VGND sg13g2_decap_8
XFILLER_27_361 VPWR VGND sg13g2_decap_8
XFILLER_43_854 VPWR VGND sg13g2_decap_8
XFILLER_70_651 VPWR VGND sg13g2_decap_8
XFILLER_15_578 VPWR VGND sg13g2_decap_8
XFILLER_30_504 VPWR VGND sg13g2_decap_8
XFILLER_91_77 VPWR VGND sg13g2_decap_8
XFILLER_42_375 VPWR VGND sg13g2_decap_8
XFILLER_24_60 VPWR VGND sg13g2_decap_8
XFILLER_7_711 VPWR VGND sg13g2_decap_8
XFILLER_6_210 VPWR VGND sg13g2_decap_8
XFILLER_11_784 VPWR VGND sg13g2_decap_8
XFILLER_7_788 VPWR VGND sg13g2_decap_8
XFILLER_6_287 VPWR VGND sg13g2_decap_8
XFILLER_40_70 VPWR VGND sg13g2_decap_8
XFILLER_97_504 VPWR VGND sg13g2_decap_8
XFILLER_41_7 VPWR VGND sg13g2_decap_8
XFILLER_69_239 VPWR VGND sg13g2_decap_8
XFILLER_3_994 VPWR VGND sg13g2_decap_8
XFILLER_78_762 VPWR VGND sg13g2_decap_8
XFILLER_66_902 VPWR VGND sg13g2_decap_8
XFILLER_38_637 VPWR VGND sg13g2_decap_8
XFILLER_93_754 VPWR VGND sg13g2_decap_8
XFILLER_92_231 VPWR VGND sg13g2_decap_8
XFILLER_77_294 VPWR VGND sg13g2_decap_8
XFILLER_66_979 VPWR VGND sg13g2_decap_8
XFILLER_65_434 VPWR VGND sg13g2_decap_8
XFILLER_1_42 VPWR VGND sg13g2_decap_8
XFILLER_19_840 VPWR VGND sg13g2_decap_8
XFILLER_81_949 VPWR VGND sg13g2_decap_8
XFILLER_18_350 VPWR VGND sg13g2_decap_8
XFILLER_37_158 VPWR VGND sg13g2_decap_8
XFILLER_80_448 VPWR VGND sg13g2_decap_8
XFILLER_61_662 VPWR VGND sg13g2_decap_8
XFILLER_21_504 VPWR VGND sg13g2_decap_8
XFILLER_33_364 VPWR VGND sg13g2_decap_8
XFILLER_34_865 VPWR VGND sg13g2_decap_8
XFILLER_60_172 VPWR VGND sg13g2_decap_8
XFILLER_14_1015 VPWR VGND sg13g2_decap_8
XFILLER_106_119 VPWR VGND sg13g2_decap_8
XFILLER_20_18 VPWR VGND sg13g2_decap_8
XFILLER_103_826 VPWR VGND sg13g2_decap_8
XFILLER_88_515 VPWR VGND sg13g2_decap_8
XFILLER_102_336 VPWR VGND sg13g2_decap_8
XFILLER_96_581 VPWR VGND sg13g2_decap_8
XFILLER_84_721 VPWR VGND sg13g2_decap_8
XFILLER_68_250 VPWR VGND sg13g2_decap_8
XFILLER_57_924 VPWR VGND sg13g2_decap_8
XFILLER_21_1008 VPWR VGND sg13g2_decap_8
XFILLER_83_242 VPWR VGND sg13g2_decap_8
XFILLER_56_445 VPWR VGND sg13g2_decap_8
XFILLER_28_147 VPWR VGND sg13g2_decap_8
XFILLER_29_648 VPWR VGND sg13g2_decap_8
XFILLER_84_798 VPWR VGND sg13g2_decap_8
XFILLER_72_938 VPWR VGND sg13g2_decap_8
XFILLER_71_459 VPWR VGND sg13g2_decap_8
XFILLER_101_21 VPWR VGND sg13g2_decap_8
XFILLER_52_651 VPWR VGND sg13g2_decap_8
XFILLER_25_854 VPWR VGND sg13g2_decap_8
XFILLER_51_172 VPWR VGND sg13g2_decap_8
XFILLER_12_515 VPWR VGND sg13g2_decap_8
XFILLER_24_375 VPWR VGND sg13g2_decap_8
XFILLER_101_98 VPWR VGND sg13g2_decap_8
XFILLER_40_868 VPWR VGND sg13g2_decap_8
XFILLER_20_592 VPWR VGND sg13g2_decap_8
XFILLER_4_714 VPWR VGND sg13g2_decap_8
XFILLER_3_224 VPWR VGND sg13g2_decap_8
XFILLER_106_686 VPWR VGND sg13g2_decap_8
XFILLER_79_515 VPWR VGND sg13g2_decap_8
XFILLER_105_196 VPWR VGND sg13g2_decap_8
XFILLER_86_11 VPWR VGND sg13g2_decap_8
XFILLER_10_95 VPWR VGND sg13g2_decap_8
XFILLER_0_931 VPWR VGND sg13g2_decap_8
XFILLER_94_518 VPWR VGND sg13g2_decap_8
XFILLER_66_209 VPWR VGND sg13g2_decap_8
XFILLER_87_581 VPWR VGND sg13g2_decap_8
XFILLER_86_88 VPWR VGND sg13g2_decap_8
XFILLER_75_721 VPWR VGND sg13g2_decap_8
XFILLER_59_250 VPWR VGND sg13g2_decap_8
XFILLER_48_924 VPWR VGND sg13g2_decap_8
XFILLER_47_434 VPWR VGND sg13g2_decap_8
XFILLER_19_147 VPWR VGND sg13g2_decap_8
XFILLER_75_798 VPWR VGND sg13g2_decap_8
XFILLER_74_253 VPWR VGND sg13g2_decap_8
XFILLER_63_938 VPWR VGND sg13g2_decap_8
XFILLER_90_746 VPWR VGND sg13g2_decap_8
XFILLER_62_448 VPWR VGND sg13g2_decap_8
XFILLER_43_651 VPWR VGND sg13g2_decap_8
XFILLER_16_854 VPWR VGND sg13g2_decap_8
XFILLER_35_70 VPWR VGND sg13g2_decap_8
XFILLER_42_172 VPWR VGND sg13g2_decap_8
XFILLER_15_375 VPWR VGND sg13g2_decap_8
XFILLER_30_301 VPWR VGND sg13g2_decap_8
XFILLER_37_1026 VPWR VGND sg13g2_fill_2
XFILLER_89_7 VPWR VGND sg13g2_decap_8
XFILLER_31_868 VPWR VGND sg13g2_decap_8
XFILLER_30_378 VPWR VGND sg13g2_decap_8
XFILLER_11_581 VPWR VGND sg13g2_decap_8
XFILLER_7_585 VPWR VGND sg13g2_decap_8
XFILLER_98_802 VPWR VGND sg13g2_decap_8
XFILLER_97_301 VPWR VGND sg13g2_decap_8
XFILLER_44_1019 VPWR VGND sg13g2_decap_8
XFILLER_3_791 VPWR VGND sg13g2_decap_8
XFILLER_98_879 VPWR VGND sg13g2_decap_8
XFILLER_97_378 VPWR VGND sg13g2_decap_8
XFILLER_85_518 VPWR VGND sg13g2_decap_8
XFILLER_39_935 VPWR VGND sg13g2_decap_8
XFILLER_65_231 VPWR VGND sg13g2_decap_8
XFILLER_38_434 VPWR VGND sg13g2_decap_8
XFILLER_93_551 VPWR VGND sg13g2_decap_8
XFILLER_66_776 VPWR VGND sg13g2_decap_8
XFILLER_81_746 VPWR VGND sg13g2_decap_8
XFILLER_54_949 VPWR VGND sg13g2_decap_8
XFILLER_53_448 VPWR VGND sg13g2_decap_8
XFILLER_80_245 VPWR VGND sg13g2_decap_8
XFILLER_15_18 VPWR VGND sg13g2_decap_8
XFILLER_22_802 VPWR VGND sg13g2_decap_8
XFILLER_34_662 VPWR VGND sg13g2_decap_8
XFILLER_90_1028 VPWR VGND sg13g2_fill_1
XFILLER_21_301 VPWR VGND sg13g2_decap_8
XFILLER_33_161 VPWR VGND sg13g2_decap_8
XFILLER_22_879 VPWR VGND sg13g2_decap_8
XFILLER_21_378 VPWR VGND sg13g2_decap_8
XFILLER_31_28 VPWR VGND sg13g2_decap_8
Xoutput17 net17 uo_out[0] VPWR VGND sg13g2_buf_1
XFILLER_103_623 VPWR VGND sg13g2_decap_8
XFILLER_88_312 VPWR VGND sg13g2_decap_8
XFILLER_1_728 VPWR VGND sg13g2_decap_8
XFILLER_102_133 VPWR VGND sg13g2_decap_8
XFILLER_89_868 VPWR VGND sg13g2_decap_8
XFILLER_0_238 VPWR VGND sg13g2_decap_8
XFILLER_88_389 VPWR VGND sg13g2_decap_8
XFILLER_76_529 VPWR VGND sg13g2_decap_8
XFILLER_57_721 VPWR VGND sg13g2_decap_8
XFILLER_56_25 VPWR VGND sg13g2_decap_8
XFILLER_29_445 VPWR VGND sg13g2_decap_8
XFILLER_57_798 VPWR VGND sg13g2_decap_8
XFILLER_56_242 VPWR VGND sg13g2_decap_8
XFILLER_45_938 VPWR VGND sg13g2_decap_8
XFILLER_84_595 VPWR VGND sg13g2_decap_8
XFILLER_72_735 VPWR VGND sg13g2_decap_8
XFILLER_71_256 VPWR VGND sg13g2_decap_8
XFILLER_44_459 VPWR VGND sg13g2_decap_8
XFILLER_25_651 VPWR VGND sg13g2_decap_8
XFILLER_72_35 VPWR VGND sg13g2_decap_8
XFILLER_12_312 VPWR VGND sg13g2_decap_8
XFILLER_24_172 VPWR VGND sg13g2_decap_8
XFILLER_13_868 VPWR VGND sg13g2_decap_8
XFILLER_40_665 VPWR VGND sg13g2_decap_8
XFILLER_12_389 VPWR VGND sg13g2_decap_8
XFILLER_67_1008 VPWR VGND sg13g2_decap_8
XFILLER_4_511 VPWR VGND sg13g2_decap_8
XFILLER_98_109 VPWR VGND sg13g2_decap_8
XFILLER_97_21 VPWR VGND sg13g2_decap_8
XFILLER_106_483 VPWR VGND sg13g2_decap_8
XFILLER_79_312 VPWR VGND sg13g2_decap_8
XFILLER_4_588 VPWR VGND sg13g2_decap_8
XFILLER_97_98 VPWR VGND sg13g2_decap_8
XFILLER_95_816 VPWR VGND sg13g2_decap_8
XFILLER_94_315 VPWR VGND sg13g2_decap_8
XFILLER_79_389 VPWR VGND sg13g2_decap_8
XFILLER_67_518 VPWR VGND sg13g2_decap_8
XFILLER_48_721 VPWR VGND sg13g2_decap_8
XFILLER_47_231 VPWR VGND sg13g2_decap_8
XFILLER_36_938 VPWR VGND sg13g2_decap_8
XFILLER_75_595 VPWR VGND sg13g2_decap_8
XFILLER_63_735 VPWR VGND sg13g2_decap_8
XFILLER_48_798 VPWR VGND sg13g2_decap_8
XFILLER_90_543 VPWR VGND sg13g2_decap_8
XFILLER_62_245 VPWR VGND sg13g2_decap_8
XFILLER_16_651 VPWR VGND sg13g2_decap_8
XFILLER_35_448 VPWR VGND sg13g2_decap_8
XFILLER_22_109 VPWR VGND sg13g2_decap_8
XFILLER_15_172 VPWR VGND sg13g2_decap_8
XFILLER_50_1001 VPWR VGND sg13g2_decap_8
XFILLER_31_665 VPWR VGND sg13g2_decap_8
XFILLER_30_175 VPWR VGND sg13g2_decap_8
XFILLER_8_861 VPWR VGND sg13g2_decap_8
XFILLER_7_382 VPWR VGND sg13g2_decap_8
XFILLER_7_74 VPWR VGND sg13g2_decap_8
XFILLER_98_676 VPWR VGND sg13g2_decap_8
XFILLER_86_816 VPWR VGND sg13g2_decap_8
XFILLER_30_0 VPWR VGND sg13g2_decap_8
XFILLER_97_175 VPWR VGND sg13g2_decap_8
XFILLER_85_315 VPWR VGND sg13g2_decap_8
XFILLER_58_518 VPWR VGND sg13g2_decap_8
XFILLER_100_637 VPWR VGND sg13g2_decap_8
XFILLER_39_732 VPWR VGND sg13g2_decap_8
XFILLER_94_882 VPWR VGND sg13g2_decap_8
XFILLER_66_573 VPWR VGND sg13g2_decap_8
XFILLER_38_231 VPWR VGND sg13g2_decap_8
XFILLER_54_746 VPWR VGND sg13g2_decap_8
XFILLER_26_28 VPWR VGND sg13g2_decap_8
XFILLER_27_949 VPWR VGND sg13g2_decap_8
XFILLER_81_543 VPWR VGND sg13g2_decap_8
XFILLER_53_245 VPWR VGND sg13g2_decap_8
XFILLER_26_448 VPWR VGND sg13g2_decap_8
XFILLER_50_952 VPWR VGND sg13g2_decap_8
XFILLER_10_816 VPWR VGND sg13g2_decap_8
XFILLER_22_676 VPWR VGND sg13g2_decap_8
XFILLER_21_175 VPWR VGND sg13g2_decap_8
XFILLER_5_319 VPWR VGND sg13g2_decap_8
XFILLER_104_910 VPWR VGND sg13g2_decap_8
XFILLER_1_525 VPWR VGND sg13g2_decap_8
XFILLER_103_420 VPWR VGND sg13g2_decap_8
XFILLER_89_665 VPWR VGND sg13g2_decap_8
XFILLER_77_805 VPWR VGND sg13g2_decap_8
XFILLER_104_987 VPWR VGND sg13g2_decap_8
XFILLER_67_57 VPWR VGND sg13g2_fill_1
XFILLER_49_529 VPWR VGND sg13g2_decap_8
XFILLER_103_497 VPWR VGND sg13g2_decap_8
XFILLER_88_186 VPWR VGND sg13g2_decap_8
XFILLER_76_326 VPWR VGND sg13g2_decap_8
XFILLER_92_819 VPWR VGND sg13g2_decap_8
XFILLER_29_242 VPWR VGND sg13g2_decap_8
XFILLER_91_329 VPWR VGND sg13g2_decap_8
XFILLER_85_882 VPWR VGND sg13g2_decap_8
XFILLER_72_532 VPWR VGND sg13g2_decap_8
XFILLER_57_595 VPWR VGND sg13g2_decap_8
XFILLER_45_735 VPWR VGND sg13g2_decap_8
XFILLER_18_938 VPWR VGND sg13g2_decap_8
XFILLER_84_392 VPWR VGND sg13g2_decap_8
XFILLER_83_67 VPWR VGND sg13g2_decap_8
XFILLER_44_256 VPWR VGND sg13g2_decap_8
XFILLER_17_459 VPWR VGND sg13g2_decap_8
XFILLER_73_1012 VPWR VGND sg13g2_decap_8
XFILLER_41_952 VPWR VGND sg13g2_decap_8
XFILLER_13_665 VPWR VGND sg13g2_decap_8
XFILLER_40_462 VPWR VGND sg13g2_decap_8
XFILLER_9_658 VPWR VGND sg13g2_decap_8
XFILLER_12_186 VPWR VGND sg13g2_decap_8
XFILLER_8_168 VPWR VGND sg13g2_decap_8
XFILLER_32_60 VPWR VGND sg13g2_decap_8
XFILLER_5_886 VPWR VGND sg13g2_decap_8
XFILLER_4_385 VPWR VGND sg13g2_decap_8
XFILLER_106_280 VPWR VGND sg13g2_decap_8
XFILLER_95_613 VPWR VGND sg13g2_decap_8
XFILLER_68_838 VPWR VGND sg13g2_decap_8
XFILLER_67_315 VPWR VGND sg13g2_decap_8
XFILLER_94_112 VPWR VGND sg13g2_decap_8
XFILLER_79_186 VPWR VGND sg13g2_decap_8
XFILLER_94_189 VPWR VGND sg13g2_decap_8
XFILLER_82_329 VPWR VGND sg13g2_decap_8
XFILLER_76_893 VPWR VGND sg13g2_decap_8
XFILLER_48_595 VPWR VGND sg13g2_decap_8
XFILLER_36_735 VPWR VGND sg13g2_decap_8
XFILLER_90_340 VPWR VGND sg13g2_decap_8
XFILLER_75_392 VPWR VGND sg13g2_decap_8
XFILLER_63_532 VPWR VGND sg13g2_decap_8
XFILLER_35_245 VPWR VGND sg13g2_decap_8
XFILLER_91_896 VPWR VGND sg13g2_decap_8
XFILLER_50_259 VPWR VGND sg13g2_decap_8
XFILLER_31_462 VPWR VGND sg13g2_decap_8
XFILLER_32_963 VPWR VGND sg13g2_decap_8
XFILLER_105_707 VPWR VGND sg13g2_decap_8
XFILLER_104_217 VPWR VGND sg13g2_decap_8
XFILLER_99_952 VPWR VGND sg13g2_decap_8
XFILLER_101_924 VPWR VGND sg13g2_decap_8
XFILLER_98_473 VPWR VGND sg13g2_decap_8
XFILLER_86_613 VPWR VGND sg13g2_decap_8
XFILLER_59_838 VPWR VGND sg13g2_decap_8
XFILLER_58_315 VPWR VGND sg13g2_decap_8
XFILLER_100_434 VPWR VGND sg13g2_decap_8
XFILLER_85_112 VPWR VGND sg13g2_decap_8
XFILLER_2_1005 VPWR VGND sg13g2_decap_8
XFILLER_96_1001 VPWR VGND sg13g2_decap_8
XFILLER_85_189 VPWR VGND sg13g2_decap_8
XFILLER_67_882 VPWR VGND sg13g2_decap_8
XFILLER_66_370 VPWR VGND sg13g2_decap_8
XFILLER_81_340 VPWR VGND sg13g2_decap_8
XFILLER_54_543 VPWR VGND sg13g2_decap_8
XFILLER_26_245 VPWR VGND sg13g2_decap_8
XFILLER_27_746 VPWR VGND sg13g2_decap_8
XFILLER_82_896 VPWR VGND sg13g2_decap_8
XFILLER_23_952 VPWR VGND sg13g2_decap_8
XFILLER_41_259 VPWR VGND sg13g2_decap_8
XFILLER_10_613 VPWR VGND sg13g2_decap_8
XFILLER_22_473 VPWR VGND sg13g2_decap_8
XFILLER_5_116 VPWR VGND sg13g2_decap_8
XFILLER_2_823 VPWR VGND sg13g2_decap_8
XFILLER_1_322 VPWR VGND sg13g2_decap_8
XFILLER_104_784 VPWR VGND sg13g2_decap_8
XFILLER_89_462 VPWR VGND sg13g2_decap_8
XFILLER_77_602 VPWR VGND sg13g2_decap_8
XFILLER_103_294 VPWR VGND sg13g2_decap_8
XFILLER_76_123 VPWR VGND sg13g2_decap_8
XFILLER_49_326 VPWR VGND sg13g2_decap_8
XFILLER_1_399 VPWR VGND sg13g2_decap_8
XFILLER_92_616 VPWR VGND sg13g2_decap_8
XFILLER_77_679 VPWR VGND sg13g2_decap_8
XFILLER_65_819 VPWR VGND sg13g2_decap_8
XFILLER_40_1022 VPWR VGND sg13g2_decap_8
XFILLER_94_77 VPWR VGND sg13g2_decap_8
XFILLER_91_126 VPWR VGND sg13g2_decap_8
XFILLER_73_830 VPWR VGND sg13g2_decap_8
XFILLER_58_882 VPWR VGND sg13g2_decap_8
XFILLER_18_735 VPWR VGND sg13g2_decap_8
XFILLER_57_392 VPWR VGND sg13g2_decap_8
XFILLER_45_532 VPWR VGND sg13g2_decap_8
XFILLER_27_60 VPWR VGND sg13g2_decap_8
XFILLER_17_256 VPWR VGND sg13g2_decap_8
XFILLER_60_557 VPWR VGND sg13g2_decap_8
XFILLER_33_749 VPWR VGND sg13g2_decap_8
XFILLER_14_952 VPWR VGND sg13g2_decap_8
XFILLER_43_70 VPWR VGND sg13g2_decap_8
XFILLER_13_462 VPWR VGND sg13g2_decap_8
XFILLER_9_455 VPWR VGND sg13g2_decap_8
XFILLER_5_683 VPWR VGND sg13g2_decap_8
XFILLER_99_259 VPWR VGND sg13g2_decap_8
XFILLER_4_182 VPWR VGND sg13g2_decap_8
XFILLER_4_42 VPWR VGND sg13g2_decap_8
XFILLER_96_966 VPWR VGND sg13g2_decap_8
XFILLER_95_410 VPWR VGND sg13g2_decap_8
XFILLER_68_635 VPWR VGND sg13g2_decap_8
XFILLER_67_112 VPWR VGND sg13g2_decap_8
XFILLER_95_487 VPWR VGND sg13g2_decap_8
XFILLER_83_627 VPWR VGND sg13g2_decap_8
XFILLER_82_126 VPWR VGND sg13g2_decap_8
XFILLER_67_189 VPWR VGND sg13g2_decap_8
XFILLER_64_830 VPWR VGND sg13g2_decap_8
XFILLER_55_329 VPWR VGND sg13g2_decap_8
XFILLER_49_893 VPWR VGND sg13g2_decap_8
XFILLER_76_690 VPWR VGND sg13g2_decap_8
XFILLER_48_392 VPWR VGND sg13g2_decap_8
XFILLER_36_532 VPWR VGND sg13g2_decap_8
XFILLER_91_693 VPWR VGND sg13g2_decap_8
XFILLER_51_557 VPWR VGND sg13g2_decap_8
XFILLER_20_900 VPWR VGND sg13g2_decap_8
XFILLER_23_259 VPWR VGND sg13g2_decap_8
XFILLER_32_760 VPWR VGND sg13g2_decap_8
XFILLER_20_977 VPWR VGND sg13g2_decap_8
XFILLER_3_609 VPWR VGND sg13g2_decap_8
XFILLER_105_504 VPWR VGND sg13g2_decap_8
XFILLER_63_1022 VPWR VGND sg13g2_decap_8
XFILLER_101_721 VPWR VGND sg13g2_decap_8
XFILLER_98_270 VPWR VGND sg13g2_decap_8
XFILLER_86_410 VPWR VGND sg13g2_decap_8
XFILLER_59_635 VPWR VGND sg13g2_decap_8
XFILLER_58_112 VPWR VGND sg13g2_decap_8
XFILLER_104_21 VPWR VGND sg13g2_decap_8
XFILLER_100_231 VPWR VGND sg13g2_decap_8
XFILLER_87_966 VPWR VGND sg13g2_decap_8
XFILLER_47_819 VPWR VGND sg13g2_decap_8
XFILLER_24_1028 VPWR VGND sg13g2_fill_1
XFILLER_101_798 VPWR VGND sg13g2_decap_8
XFILLER_86_487 VPWR VGND sg13g2_decap_8
XFILLER_74_638 VPWR VGND sg13g2_decap_8
XFILLER_58_189 VPWR VGND sg13g2_decap_8
XFILLER_73_137 VPWR VGND sg13g2_decap_8
XFILLER_64_25 VPWR VGND sg13g2_decap_8
XFILLER_27_543 VPWR VGND sg13g2_decap_8
XFILLER_104_98 VPWR VGND sg13g2_decap_8
XFILLER_55_896 VPWR VGND sg13g2_decap_8
XFILLER_54_340 VPWR VGND sg13g2_decap_8
XFILLER_82_693 VPWR VGND sg13g2_decap_8
XFILLER_70_833 VPWR VGND sg13g2_decap_8
XFILLER_42_557 VPWR VGND sg13g2_decap_8
XFILLER_14_259 VPWR VGND sg13g2_decap_8
XFILLER_80_35 VPWR VGND sg13g2_decap_8
XFILLER_70_1015 VPWR VGND sg13g2_decap_8
XFILLER_10_410 VPWR VGND sg13g2_decap_8
XFILLER_22_270 VPWR VGND sg13g2_decap_8
XFILLER_11_966 VPWR VGND sg13g2_decap_8
XFILLER_10_487 VPWR VGND sg13g2_decap_8
XFILLER_13_84 VPWR VGND sg13g2_decap_8
XFILLER_6_469 VPWR VGND sg13g2_decap_8
XFILLER_89_77 VPWR VGND sg13g2_decap_8
XFILLER_8_0 VPWR VGND sg13g2_decap_8
XFILLER_2_620 VPWR VGND sg13g2_decap_8
XFILLER_104_581 VPWR VGND sg13g2_decap_8
XFILLER_78_944 VPWR VGND sg13g2_decap_8
XFILLER_49_123 VPWR VGND sg13g2_decap_8
XFILLER_2_697 VPWR VGND sg13g2_decap_8
X_40_ net12 net4 _09_ VPWR VGND sg13g2_xor2_1
XFILLER_1_196 VPWR VGND sg13g2_decap_8
XFILLER_38_819 VPWR VGND sg13g2_decap_8
XFILLER_93_936 VPWR VGND sg13g2_decap_8
XFILLER_92_413 VPWR VGND sg13g2_decap_8
XFILLER_77_476 VPWR VGND sg13g2_decap_8
XFILLER_65_616 VPWR VGND sg13g2_decap_8
XFILLER_38_70 VPWR VGND sg13g2_decap_8
XFILLER_64_137 VPWR VGND sg13g2_decap_8
XFILLER_46_830 VPWR VGND sg13g2_decap_8
XFILLER_18_532 VPWR VGND sg13g2_decap_8
XFILLER_61_844 VPWR VGND sg13g2_decap_8
XFILLER_33_546 VPWR VGND sg13g2_decap_8
XFILLER_60_354 VPWR VGND sg13g2_decap_8
XFILLER_20_207 VPWR VGND sg13g2_decap_8
XFILLER_9_252 VPWR VGND sg13g2_decap_8
XFILLER_5_480 VPWR VGND sg13g2_decap_8
XFILLER_102_518 VPWR VGND sg13g2_decap_8
XFILLER_69_911 VPWR VGND sg13g2_decap_8
XFILLER_68_432 VPWR VGND sg13g2_decap_8
XFILLER_96_763 VPWR VGND sg13g2_decap_8
XFILLER_84_903 VPWR VGND sg13g2_decap_8
XFILLER_69_988 VPWR VGND sg13g2_decap_8
XFILLER_95_284 VPWR VGND sg13g2_decap_8
XFILLER_83_424 VPWR VGND sg13g2_decap_8
XFILLER_56_627 VPWR VGND sg13g2_decap_8
XFILLER_28_329 VPWR VGND sg13g2_decap_8
XFILLER_55_126 VPWR VGND sg13g2_decap_8
XFILLER_49_690 VPWR VGND sg13g2_decap_8
XFILLER_37_830 VPWR VGND sg13g2_decap_8
XFILLER_92_980 VPWR VGND sg13g2_decap_8
XFILLER_91_490 VPWR VGND sg13g2_decap_8
XFILLER_52_833 VPWR VGND sg13g2_decap_8
XFILLER_51_354 VPWR VGND sg13g2_decap_8
XFILLER_24_557 VPWR VGND sg13g2_decap_8
XFILLER_34_39 VPWR VGND sg13g2_decap_8
XFILLER_50_49 VPWR VGND sg13g2_decap_8
XFILLER_20_774 VPWR VGND sg13g2_decap_8
XFILLER_105_301 VPWR VGND sg13g2_decap_8
XFILLER_3_406 VPWR VGND sg13g2_decap_8
XFILLER_106_868 VPWR VGND sg13g2_decap_8
XFILLER_59_25 VPWR VGND sg13g2_decap_8
XFILLER_105_378 VPWR VGND sg13g2_decap_8
XFILLER_1_7 VPWR VGND sg13g2_decap_8
XFILLER_8_1022 VPWR VGND sg13g2_decap_8
XFILLER_87_763 VPWR VGND sg13g2_decap_8
XFILLER_75_903 VPWR VGND sg13g2_decap_8
XFILLER_59_432 VPWR VGND sg13g2_decap_8
XFILLER_86_284 VPWR VGND sg13g2_decap_8
XFILLER_75_35 VPWR VGND sg13g2_decap_8
XFILLER_47_616 VPWR VGND sg13g2_decap_8
XFILLER_19_329 VPWR VGND sg13g2_decap_8
XFILLER_101_595 VPWR VGND sg13g2_decap_8
XFILLER_74_435 VPWR VGND sg13g2_decap_8
XFILLER_46_137 VPWR VGND sg13g2_decap_8
XFILLER_90_928 VPWR VGND sg13g2_decap_8
XFILLER_27_340 VPWR VGND sg13g2_decap_8
XFILLER_83_991 VPWR VGND sg13g2_decap_8
XFILLER_82_490 VPWR VGND sg13g2_decap_8
XFILLER_70_630 VPWR VGND sg13g2_decap_8
XFILLER_55_693 VPWR VGND sg13g2_decap_8
XFILLER_43_833 VPWR VGND sg13g2_decap_8
XFILLER_28_896 VPWR VGND sg13g2_decap_8
XFILLER_91_56 VPWR VGND sg13g2_decap_8
XFILLER_42_354 VPWR VGND sg13g2_decap_8
XFILLER_15_557 VPWR VGND sg13g2_decap_8
XFILLER_11_763 VPWR VGND sg13g2_decap_8
XFILLER_10_284 VPWR VGND sg13g2_decap_8
XFILLER_7_767 VPWR VGND sg13g2_decap_8
XFILLER_6_266 VPWR VGND sg13g2_decap_8
XFILLER_3_973 VPWR VGND sg13g2_decap_8
XFILLER_69_218 VPWR VGND sg13g2_decap_8
XFILLER_78_741 VPWR VGND sg13g2_decap_8
XFILLER_2_494 VPWR VGND sg13g2_decap_8
XFILLER_93_733 VPWR VGND sg13g2_decap_8
XFILLER_77_273 VPWR VGND sg13g2_decap_8
XFILLER_65_413 VPWR VGND sg13g2_decap_8
XFILLER_1_21 VPWR VGND sg13g2_decap_8
XFILLER_38_616 VPWR VGND sg13g2_decap_8
XFILLER_92_210 VPWR VGND sg13g2_decap_8
XFILLER_66_958 VPWR VGND sg13g2_decap_8
XFILLER_37_137 VPWR VGND sg13g2_decap_8
XFILLER_81_928 VPWR VGND sg13g2_decap_8
XFILLER_1_98 VPWR VGND sg13g2_decap_8
XFILLER_92_287 VPWR VGND sg13g2_decap_8
XFILLER_80_427 VPWR VGND sg13g2_decap_8
XFILLER_19_896 VPWR VGND sg13g2_decap_8
XFILLER_34_844 VPWR VGND sg13g2_decap_8
XFILLER_61_641 VPWR VGND sg13g2_decap_8
XFILLER_33_343 VPWR VGND sg13g2_decap_8
XFILLER_60_151 VPWR VGND sg13g2_decap_8
XFILLER_101_1008 VPWR VGND sg13g2_decap_8
XFILLER_60_0 VPWR VGND sg13g2_decap_8
XFILLER_103_805 VPWR VGND sg13g2_decap_8
XFILLER_102_315 VPWR VGND sg13g2_decap_8
XFILLER_57_903 VPWR VGND sg13g2_decap_8
XFILLER_29_39 VPWR VGND sg13g2_decap_8
XFILLER_96_560 VPWR VGND sg13g2_decap_8
XFILLER_84_700 VPWR VGND sg13g2_decap_8
XFILLER_69_785 VPWR VGND sg13g2_decap_8
XFILLER_29_627 VPWR VGND sg13g2_decap_8
XFILLER_83_221 VPWR VGND sg13g2_decap_8
XFILLER_56_424 VPWR VGND sg13g2_decap_8
XFILLER_28_126 VPWR VGND sg13g2_decap_8
XFILLER_84_777 VPWR VGND sg13g2_decap_8
XFILLER_72_917 VPWR VGND sg13g2_decap_8
XFILLER_83_298 VPWR VGND sg13g2_decap_8
XFILLER_71_438 VPWR VGND sg13g2_decap_8
XFILLER_65_980 VPWR VGND sg13g2_decap_8
XFILLER_45_49 VPWR VGND sg13g2_decap_8
XFILLER_25_833 VPWR VGND sg13g2_decap_8
XFILLER_52_630 VPWR VGND sg13g2_decap_8
XFILLER_24_354 VPWR VGND sg13g2_decap_8
XFILLER_80_994 VPWR VGND sg13g2_decap_8
XFILLER_51_151 VPWR VGND sg13g2_decap_8
XFILLER_101_77 VPWR VGND sg13g2_decap_8
XFILLER_61_37 VPWR VGND sg13g2_decap_8
XFILLER_40_847 VPWR VGND sg13g2_decap_8
XFILLER_20_571 VPWR VGND sg13g2_decap_8
XFILLER_3_203 VPWR VGND sg13g2_decap_8
XFILLER_106_665 VPWR VGND sg13g2_decap_8
XFILLER_105_175 VPWR VGND sg13g2_decap_8
XFILLER_10_74 VPWR VGND sg13g2_decap_8
XFILLER_0_910 VPWR VGND sg13g2_decap_8
XFILLER_48_903 VPWR VGND sg13g2_decap_8
XFILLER_102_882 VPWR VGND sg13g2_decap_8
XFILLER_87_560 VPWR VGND sg13g2_decap_8
XFILLER_86_67 VPWR VGND sg13g2_decap_8
XFILLER_75_700 VPWR VGND sg13g2_decap_8
XFILLER_47_413 VPWR VGND sg13g2_decap_8
XFILLER_0_987 VPWR VGND sg13g2_decap_8
XFILLER_101_392 VPWR VGND sg13g2_decap_8
XFILLER_74_232 VPWR VGND sg13g2_decap_8
XFILLER_19_126 VPWR VGND sg13g2_decap_8
XFILLER_75_777 VPWR VGND sg13g2_decap_8
XFILLER_63_917 VPWR VGND sg13g2_decap_8
XFILLER_90_725 VPWR VGND sg13g2_decap_8
XFILLER_62_427 VPWR VGND sg13g2_decap_8
XFILLER_56_991 VPWR VGND sg13g2_decap_8
XFILLER_16_833 VPWR VGND sg13g2_decap_8
XFILLER_28_693 VPWR VGND sg13g2_decap_8
XFILLER_55_490 VPWR VGND sg13g2_decap_8
XFILLER_43_630 VPWR VGND sg13g2_decap_8
XFILLER_15_354 VPWR VGND sg13g2_decap_8
XFILLER_37_1005 VPWR VGND sg13g2_decap_8
XFILLER_42_151 VPWR VGND sg13g2_decap_8
XFILLER_31_847 VPWR VGND sg13g2_decap_8
XFILLER_11_560 VPWR VGND sg13g2_decap_8
XFILLER_30_357 VPWR VGND sg13g2_decap_8
XFILLER_51_81 VPWR VGND sg13g2_decap_8
XFILLER_7_564 VPWR VGND sg13g2_decap_8
XFILLER_98_858 VPWR VGND sg13g2_decap_8
XFILLER_3_770 VPWR VGND sg13g2_decap_8
XFILLER_97_357 VPWR VGND sg13g2_decap_8
XFILLER_2_291 VPWR VGND sg13g2_decap_8
XFILLER_32_4 VPWR VGND sg13g2_decap_8
XFILLER_100_819 VPWR VGND sg13g2_decap_8
XFILLER_38_413 VPWR VGND sg13g2_decap_8
XFILLER_39_914 VPWR VGND sg13g2_decap_8
XFILLER_93_530 VPWR VGND sg13g2_decap_8
XFILLER_66_755 VPWR VGND sg13g2_decap_8
XFILLER_65_210 VPWR VGND sg13g2_decap_8
XFILLER_54_928 VPWR VGND sg13g2_decap_8
XFILLER_81_725 VPWR VGND sg13g2_decap_8
XFILLER_80_224 VPWR VGND sg13g2_decap_8
XFILLER_65_287 VPWR VGND sg13g2_decap_8
XFILLER_53_427 VPWR VGND sg13g2_decap_8
XFILLER_47_980 VPWR VGND sg13g2_decap_8
XFILLER_19_693 VPWR VGND sg13g2_decap_8
XFILLER_34_641 VPWR VGND sg13g2_decap_8
XFILLER_62_994 VPWR VGND sg13g2_decap_8
XFILLER_33_140 VPWR VGND sg13g2_decap_8
XFILLER_22_858 VPWR VGND sg13g2_decap_8
XFILLER_21_357 VPWR VGND sg13g2_decap_8
Xoutput18 net18 uo_out[1] VPWR VGND sg13g2_buf_1
XFILLER_1_707 VPWR VGND sg13g2_decap_8
XFILLER_103_602 VPWR VGND sg13g2_decap_8
XFILLER_89_847 VPWR VGND sg13g2_decap_8
XFILLER_0_217 VPWR VGND sg13g2_decap_8
XFILLER_102_112 VPWR VGND sg13g2_decap_8
XFILLER_88_368 VPWR VGND sg13g2_decap_8
XFILLER_76_508 VPWR VGND sg13g2_decap_8
XFILLER_103_679 VPWR VGND sg13g2_decap_8
XFILLER_57_700 VPWR VGND sg13g2_decap_8
XFILLER_102_189 VPWR VGND sg13g2_decap_8
XFILLER_69_582 VPWR VGND sg13g2_decap_8
XFILLER_56_221 VPWR VGND sg13g2_decap_8
XFILLER_29_424 VPWR VGND sg13g2_decap_8
XFILLER_84_574 VPWR VGND sg13g2_decap_8
XFILLER_72_714 VPWR VGND sg13g2_decap_8
XFILLER_57_777 VPWR VGND sg13g2_decap_8
XFILLER_45_917 VPWR VGND sg13g2_decap_8
XFILLER_56_298 VPWR VGND sg13g2_decap_8
XFILLER_44_438 VPWR VGND sg13g2_decap_8
XFILLER_38_980 VPWR VGND sg13g2_decap_8
XFILLER_72_14 VPWR VGND sg13g2_decap_8
XFILLER_71_235 VPWR VGND sg13g2_decap_8
XFILLER_25_630 VPWR VGND sg13g2_decap_8
XFILLER_53_994 VPWR VGND sg13g2_decap_8
XFILLER_24_151 VPWR VGND sg13g2_decap_8
XFILLER_80_791 VPWR VGND sg13g2_decap_8
XFILLER_13_847 VPWR VGND sg13g2_decap_8
XFILLER_40_644 VPWR VGND sg13g2_decap_8
XFILLER_12_368 VPWR VGND sg13g2_decap_8
XFILLER_4_567 VPWR VGND sg13g2_decap_8
XFILLER_21_84 VPWR VGND sg13g2_decap_8
XFILLER_106_462 VPWR VGND sg13g2_decap_8
XFILLER_97_77 VPWR VGND sg13g2_decap_8
XFILLER_79_368 VPWR VGND sg13g2_decap_8
XFILLER_48_700 VPWR VGND sg13g2_decap_8
XFILLER_47_210 VPWR VGND sg13g2_decap_8
XFILLER_0_784 VPWR VGND sg13g2_decap_8
XFILLER_75_574 VPWR VGND sg13g2_decap_8
XFILLER_63_714 VPWR VGND sg13g2_decap_8
XFILLER_48_777 VPWR VGND sg13g2_decap_8
XFILLER_36_917 VPWR VGND sg13g2_decap_8
XFILLER_90_522 VPWR VGND sg13g2_decap_8
XFILLER_62_224 VPWR VGND sg13g2_decap_8
XFILLER_47_287 VPWR VGND sg13g2_decap_8
XFILLER_29_991 VPWR VGND sg13g2_decap_8
XFILLER_35_427 VPWR VGND sg13g2_decap_8
XFILLER_46_81 VPWR VGND sg13g2_decap_8
XFILLER_16_630 VPWR VGND sg13g2_decap_8
XFILLER_28_490 VPWR VGND sg13g2_decap_8
XFILLER_90_599 VPWR VGND sg13g2_decap_8
XFILLER_15_151 VPWR VGND sg13g2_decap_8
XFILLER_31_644 VPWR VGND sg13g2_decap_8
XFILLER_30_154 VPWR VGND sg13g2_decap_8
XFILLER_8_840 VPWR VGND sg13g2_decap_8
XFILLER_7_53 VPWR VGND sg13g2_decap_8
XFILLER_11_1008 VPWR VGND sg13g2_decap_8
XFILLER_7_361 VPWR VGND sg13g2_decap_8
XFILLER_98_655 VPWR VGND sg13g2_decap_8
XFILLER_100_616 VPWR VGND sg13g2_decap_8
XFILLER_97_154 VPWR VGND sg13g2_decap_8
XFILLER_23_0 VPWR VGND sg13g2_decap_8
XFILLER_39_711 VPWR VGND sg13g2_decap_8
XFILLER_38_210 VPWR VGND sg13g2_decap_8
XFILLER_94_861 VPWR VGND sg13g2_decap_8
XFILLER_66_552 VPWR VGND sg13g2_decap_8
XFILLER_27_928 VPWR VGND sg13g2_decap_8
XFILLER_39_788 VPWR VGND sg13g2_decap_8
XFILLER_81_522 VPWR VGND sg13g2_decap_8
XFILLER_54_725 VPWR VGND sg13g2_decap_8
XFILLER_26_427 VPWR VGND sg13g2_decap_8
XFILLER_38_287 VPWR VGND sg13g2_decap_8
XFILLER_53_224 VPWR VGND sg13g2_decap_8
XFILLER_19_490 VPWR VGND sg13g2_decap_8
XFILLER_81_599 VPWR VGND sg13g2_decap_8
XFILLER_35_994 VPWR VGND sg13g2_decap_8
XFILLER_62_791 VPWR VGND sg13g2_decap_8
XFILLER_50_931 VPWR VGND sg13g2_decap_8
XFILLER_42_39 VPWR VGND sg13g2_decap_8
XFILLER_21_154 VPWR VGND sg13g2_decap_8
XFILLER_22_655 VPWR VGND sg13g2_decap_8
XFILLER_101_7 VPWR VGND sg13g2_decap_8
XFILLER_1_504 VPWR VGND sg13g2_decap_8
XFILLER_104_966 VPWR VGND sg13g2_decap_8
XFILLER_89_644 VPWR VGND sg13g2_decap_8
XFILLER_67_14 VPWR VGND sg13g2_fill_1
XFILLER_27_1026 VPWR VGND sg13g2_fill_2
XFILLER_103_476 VPWR VGND sg13g2_decap_8
XFILLER_88_165 VPWR VGND sg13g2_decap_8
XFILLER_76_305 VPWR VGND sg13g2_decap_8
XFILLER_67_47 VPWR VGND sg13g2_fill_1
XFILLER_49_508 VPWR VGND sg13g2_decap_8
XFILLER_29_221 VPWR VGND sg13g2_decap_8
XFILLER_91_308 VPWR VGND sg13g2_decap_8
XFILLER_85_861 VPWR VGND sg13g2_decap_8
XFILLER_18_917 VPWR VGND sg13g2_decap_8
XFILLER_84_371 VPWR VGND sg13g2_decap_8
XFILLER_72_511 VPWR VGND sg13g2_decap_8
XFILLER_57_574 VPWR VGND sg13g2_decap_8
XFILLER_45_714 VPWR VGND sg13g2_decap_8
XFILLER_83_46 VPWR VGND sg13g2_decap_8
XFILLER_44_235 VPWR VGND sg13g2_decap_8
XFILLER_17_438 VPWR VGND sg13g2_decap_8
XFILLER_29_298 VPWR VGND sg13g2_decap_8
XFILLER_72_588 VPWR VGND sg13g2_decap_8
XFILLER_60_739 VPWR VGND sg13g2_decap_8
XFILLER_26_994 VPWR VGND sg13g2_decap_8
XFILLER_53_791 VPWR VGND sg13g2_decap_8
XFILLER_41_931 VPWR VGND sg13g2_decap_8
XFILLER_13_644 VPWR VGND sg13g2_decap_8
XFILLER_16_84 VPWR VGND sg13g2_decap_8
XFILLER_34_1019 VPWR VGND sg13g2_decap_8
XFILLER_40_441 VPWR VGND sg13g2_decap_8
XFILLER_9_637 VPWR VGND sg13g2_decap_8
XFILLER_12_165 VPWR VGND sg13g2_decap_8
XFILLER_8_147 VPWR VGND sg13g2_decap_8
XFILLER_5_865 VPWR VGND sg13g2_decap_8
XFILLER_4_364 VPWR VGND sg13g2_decap_8
XFILLER_79_165 VPWR VGND sg13g2_decap_8
XFILLER_68_817 VPWR VGND sg13g2_decap_8
XFILLER_0_581 VPWR VGND sg13g2_decap_8
XFILLER_95_669 VPWR VGND sg13g2_decap_8
XFILLER_94_168 VPWR VGND sg13g2_decap_8
XFILLER_83_809 VPWR VGND sg13g2_decap_8
XFILLER_82_308 VPWR VGND sg13g2_decap_8
XFILLER_76_872 VPWR VGND sg13g2_decap_8
XFILLER_75_371 VPWR VGND sg13g2_decap_8
XFILLER_63_511 VPWR VGND sg13g2_decap_8
XFILLER_57_91 VPWR VGND sg13g2_decap_8
XFILLER_48_574 VPWR VGND sg13g2_decap_8
XFILLER_36_714 VPWR VGND sg13g2_decap_8
XFILLER_35_224 VPWR VGND sg13g2_decap_8
XFILLER_91_875 VPWR VGND sg13g2_decap_8
XFILLER_63_588 VPWR VGND sg13g2_decap_8
XFILLER_51_739 VPWR VGND sg13g2_decap_8
XFILLER_90_396 VPWR VGND sg13g2_decap_8
XFILLER_50_238 VPWR VGND sg13g2_decap_8
XFILLER_32_942 VPWR VGND sg13g2_decap_8
XFILLER_31_441 VPWR VGND sg13g2_decap_8
XFILLER_99_931 VPWR VGND sg13g2_decap_8
XFILLER_101_903 VPWR VGND sg13g2_decap_8
XFILLER_98_452 VPWR VGND sg13g2_decap_8
XFILLER_59_817 VPWR VGND sg13g2_decap_8
XFILLER_100_413 VPWR VGND sg13g2_decap_8
XFILLER_86_669 VPWR VGND sg13g2_decap_8
XFILLER_85_168 VPWR VGND sg13g2_decap_8
XFILLER_67_861 VPWR VGND sg13g2_decap_8
XFILLER_37_39 VPWR VGND sg13g2_decap_8
XFILLER_73_319 VPWR VGND sg13g2_decap_8
XFILLER_54_522 VPWR VGND sg13g2_decap_8
XFILLER_2_1028 VPWR VGND sg13g2_fill_1
XFILLER_27_725 VPWR VGND sg13g2_decap_8
XFILLER_39_585 VPWR VGND sg13g2_decap_8
XFILLER_57_1008 VPWR VGND sg13g2_decap_8
XFILLER_26_224 VPWR VGND sg13g2_decap_8
XFILLER_82_875 VPWR VGND sg13g2_decap_8
XFILLER_81_396 VPWR VGND sg13g2_decap_8
XFILLER_54_599 VPWR VGND sg13g2_decap_8
XFILLER_53_49 VPWR VGND sg13g2_decap_8
XFILLER_42_739 VPWR VGND sg13g2_decap_8
XFILLER_23_931 VPWR VGND sg13g2_decap_8
XFILLER_35_791 VPWR VGND sg13g2_decap_8
XFILLER_41_238 VPWR VGND sg13g2_decap_8
XFILLER_22_452 VPWR VGND sg13g2_decap_8
XFILLER_10_669 VPWR VGND sg13g2_decap_8
XFILLER_2_802 VPWR VGND sg13g2_decap_8
XFILLER_1_301 VPWR VGND sg13g2_decap_8
XFILLER_89_441 VPWR VGND sg13g2_decap_8
XFILLER_78_46 VPWR VGND sg13g2_decap_8
XFILLER_104_763 VPWR VGND sg13g2_decap_8
XFILLER_49_305 VPWR VGND sg13g2_decap_8
XFILLER_2_879 VPWR VGND sg13g2_decap_8
XFILLER_103_273 VPWR VGND sg13g2_decap_8
XFILLER_76_102 VPWR VGND sg13g2_decap_8
XFILLER_1_378 VPWR VGND sg13g2_decap_8
XFILLER_77_658 VPWR VGND sg13g2_decap_8
XFILLER_58_861 VPWR VGND sg13g2_decap_8
XFILLER_40_1001 VPWR VGND sg13g2_decap_8
XFILLER_100_980 VPWR VGND sg13g2_decap_8
XFILLER_94_56 VPWR VGND sg13g2_decap_8
XFILLER_91_105 VPWR VGND sg13g2_decap_8
XFILLER_76_179 VPWR VGND sg13g2_decap_8
XFILLER_64_319 VPWR VGND sg13g2_decap_8
XFILLER_57_371 VPWR VGND sg13g2_decap_8
XFILLER_45_511 VPWR VGND sg13g2_decap_8
XFILLER_18_714 VPWR VGND sg13g2_decap_8
XFILLER_17_235 VPWR VGND sg13g2_decap_8
XFILLER_73_886 VPWR VGND sg13g2_decap_8
XFILLER_45_588 VPWR VGND sg13g2_decap_8
XFILLER_33_728 VPWR VGND sg13g2_decap_8
XFILLER_72_385 VPWR VGND sg13g2_decap_8
XFILLER_60_536 VPWR VGND sg13g2_decap_8
XFILLER_14_931 VPWR VGND sg13g2_decap_8
XFILLER_26_791 VPWR VGND sg13g2_decap_8
XFILLER_13_441 VPWR VGND sg13g2_decap_8
XFILLER_32_249 VPWR VGND sg13g2_decap_8
XFILLER_9_434 VPWR VGND sg13g2_decap_8
XFILLER_5_662 VPWR VGND sg13g2_decap_8
XFILLER_99_238 VPWR VGND sg13g2_decap_8
XFILLER_4_161 VPWR VGND sg13g2_decap_8
XFILLER_4_21 VPWR VGND sg13g2_decap_8
XFILLER_68_614 VPWR VGND sg13g2_decap_8
XFILLER_96_945 VPWR VGND sg13g2_decap_8
XFILLER_4_98 VPWR VGND sg13g2_decap_8
XFILLER_95_466 VPWR VGND sg13g2_decap_8
XFILLER_83_606 VPWR VGND sg13g2_decap_8
XFILLER_56_809 VPWR VGND sg13g2_decap_8
XFILLER_82_105 VPWR VGND sg13g2_decap_8
XFILLER_67_168 VPWR VGND sg13g2_decap_8
XFILLER_55_308 VPWR VGND sg13g2_decap_8
XFILLER_49_872 VPWR VGND sg13g2_decap_8
XFILLER_48_371 VPWR VGND sg13g2_decap_8
XFILLER_36_511 VPWR VGND sg13g2_decap_8
XFILLER_91_672 VPWR VGND sg13g2_decap_8
XFILLER_64_886 VPWR VGND sg13g2_decap_8
XFILLER_36_588 VPWR VGND sg13g2_decap_8
XFILLER_63_385 VPWR VGND sg13g2_decap_8
XFILLER_51_536 VPWR VGND sg13g2_decap_8
XFILLER_23_238 VPWR VGND sg13g2_decap_8
XFILLER_24_739 VPWR VGND sg13g2_decap_8
XFILLER_90_193 VPWR VGND sg13g2_decap_8
XFILLER_20_956 VPWR VGND sg13g2_decap_8
XFILLER_2_109 VPWR VGND sg13g2_decap_8
XFILLER_101_700 VPWR VGND sg13g2_decap_8
XFILLER_63_1001 VPWR VGND sg13g2_decap_8
XFILLER_59_614 VPWR VGND sg13g2_decap_8
XFILLER_100_210 VPWR VGND sg13g2_decap_8
XFILLER_87_945 VPWR VGND sg13g2_decap_8
XFILLER_48_49 VPWR VGND sg13g2_decap_8
XFILLER_86_466 VPWR VGND sg13g2_decap_8
XFILLER_101_777 VPWR VGND sg13g2_decap_8
XFILLER_74_617 VPWR VGND sg13g2_decap_8
XFILLER_73_116 VPWR VGND sg13g2_decap_8
XFILLER_58_168 VPWR VGND sg13g2_decap_8
XFILLER_46_319 VPWR VGND sg13g2_decap_8
XFILLER_104_77 VPWR VGND sg13g2_decap_8
XFILLER_100_287 VPWR VGND sg13g2_decap_8
XFILLER_27_522 VPWR VGND sg13g2_decap_8
XFILLER_39_382 VPWR VGND sg13g2_decap_8
XFILLER_82_672 VPWR VGND sg13g2_decap_8
XFILLER_70_812 VPWR VGND sg13g2_decap_8
XFILLER_55_875 VPWR VGND sg13g2_decap_8
XFILLER_54_396 VPWR VGND sg13g2_decap_8
XFILLER_42_536 VPWR VGND sg13g2_decap_8
XFILLER_14_238 VPWR VGND sg13g2_decap_8
XFILLER_15_739 VPWR VGND sg13g2_decap_8
XFILLER_27_599 VPWR VGND sg13g2_decap_8
XFILLER_81_193 VPWR VGND sg13g2_decap_8
XFILLER_80_14 VPWR VGND sg13g2_decap_8
XFILLER_70_889 VPWR VGND sg13g2_decap_8
XFILLER_11_945 VPWR VGND sg13g2_decap_8
XFILLER_10_466 VPWR VGND sg13g2_decap_8
XFILLER_7_949 VPWR VGND sg13g2_decap_8
XFILLER_13_63 VPWR VGND sg13g2_decap_8
XFILLER_6_448 VPWR VGND sg13g2_decap_8
XFILLER_89_56 VPWR VGND sg13g2_decap_8
XFILLER_2_676 VPWR VGND sg13g2_decap_8
XFILLER_104_560 VPWR VGND sg13g2_decap_8
XFILLER_78_923 VPWR VGND sg13g2_decap_8
XFILLER_49_102 VPWR VGND sg13g2_decap_8
XFILLER_1_175 VPWR VGND sg13g2_decap_8
XFILLER_93_915 VPWR VGND sg13g2_decap_8
XFILLER_77_455 VPWR VGND sg13g2_decap_8
XFILLER_64_116 VPWR VGND sg13g2_decap_8
XFILLER_49_179 VPWR VGND sg13g2_decap_8
XFILLER_18_511 VPWR VGND sg13g2_decap_8
XFILLER_37_319 VPWR VGND sg13g2_decap_8
XFILLER_92_469 VPWR VGND sg13g2_decap_8
XFILLER_80_609 VPWR VGND sg13g2_decap_8
XFILLER_46_886 VPWR VGND sg13g2_decap_8
XFILLER_73_683 VPWR VGND sg13g2_decap_8
XFILLER_72_182 VPWR VGND sg13g2_decap_8
XFILLER_61_823 VPWR VGND sg13g2_decap_8
XFILLER_45_385 VPWR VGND sg13g2_decap_8
XFILLER_18_588 VPWR VGND sg13g2_decap_8
XFILLER_33_525 VPWR VGND sg13g2_decap_8
XFILLER_60_333 VPWR VGND sg13g2_decap_8
XFILLER_54_81 VPWR VGND sg13g2_decap_8
XFILLER_9_231 VPWR VGND sg13g2_decap_8
XFILLER_70_91 VPWR VGND sg13g2_decap_8
XFILLER_86_1012 VPWR VGND sg13g2_decap_8
XFILLER_68_411 VPWR VGND sg13g2_decap_8
XFILLER_96_742 VPWR VGND sg13g2_decap_8
XFILLER_69_967 VPWR VGND sg13g2_decap_8
XFILLER_56_606 VPWR VGND sg13g2_decap_8
XFILLER_29_809 VPWR VGND sg13g2_decap_8
XFILLER_95_263 VPWR VGND sg13g2_decap_8
XFILLER_83_403 VPWR VGND sg13g2_decap_8
XFILLER_68_488 VPWR VGND sg13g2_decap_8
XFILLER_55_105 VPWR VGND sg13g2_decap_8
XFILLER_28_308 VPWR VGND sg13g2_decap_8
XFILLER_84_959 VPWR VGND sg13g2_decap_8
XFILLER_52_812 VPWR VGND sg13g2_decap_8
XFILLER_37_886 VPWR VGND sg13g2_decap_8
XFILLER_93_1027 VPWR VGND sg13g2_fill_2
XFILLER_70_119 VPWR VGND sg13g2_decap_8
XFILLER_64_683 VPWR VGND sg13g2_decap_8
XFILLER_63_182 VPWR VGND sg13g2_decap_8
XFILLER_24_536 VPWR VGND sg13g2_decap_8
XFILLER_34_18 VPWR VGND sg13g2_decap_8
XFILLER_36_385 VPWR VGND sg13g2_decap_8
XFILLER_51_333 VPWR VGND sg13g2_decap_8
XFILLER_52_889 VPWR VGND sg13g2_decap_8
XFILLER_50_28 VPWR VGND sg13g2_decap_8
XFILLER_20_753 VPWR VGND sg13g2_decap_8
XFILLER_30_1022 VPWR VGND sg13g2_decap_8
XFILLER_106_847 VPWR VGND sg13g2_decap_8
XFILLER_105_357 VPWR VGND sg13g2_decap_8
XFILLER_59_411 VPWR VGND sg13g2_decap_8
XFILLER_8_1001 VPWR VGND sg13g2_decap_8
XFILLER_87_742 VPWR VGND sg13g2_decap_8
XFILLER_101_574 VPWR VGND sg13g2_decap_8
XFILLER_86_263 VPWR VGND sg13g2_decap_8
XFILLER_75_14 VPWR VGND sg13g2_decap_8
XFILLER_74_414 VPWR VGND sg13g2_decap_8
XFILLER_59_488 VPWR VGND sg13g2_decap_8
XFILLER_19_308 VPWR VGND sg13g2_decap_8
XFILLER_90_907 VPWR VGND sg13g2_decap_8
XFILLER_75_959 VPWR VGND sg13g2_decap_8
XFILLER_75_58 VPWR VGND sg13g2_fill_1
XFILLER_46_116 VPWR VGND sg13g2_decap_8
XFILLER_83_970 VPWR VGND sg13g2_decap_8
XFILLER_62_609 VPWR VGND sg13g2_decap_8
XFILLER_43_812 VPWR VGND sg13g2_decap_8
XFILLER_28_875 VPWR VGND sg13g2_decap_8
XFILLER_55_672 VPWR VGND sg13g2_decap_8
XFILLER_15_536 VPWR VGND sg13g2_decap_8
XFILLER_27_396 VPWR VGND sg13g2_decap_8
XFILLER_91_35 VPWR VGND sg13g2_decap_8
XFILLER_54_193 VPWR VGND sg13g2_decap_8
XFILLER_42_333 VPWR VGND sg13g2_decap_8
XFILLER_70_686 VPWR VGND sg13g2_decap_8
XFILLER_43_889 VPWR VGND sg13g2_decap_8
XFILLER_11_742 VPWR VGND sg13g2_decap_8
XFILLER_30_539 VPWR VGND sg13g2_decap_8
XFILLER_24_95 VPWR VGND sg13g2_decap_8
XFILLER_10_263 VPWR VGND sg13g2_decap_8
XFILLER_7_746 VPWR VGND sg13g2_decap_8
XFILLER_6_245 VPWR VGND sg13g2_decap_8
XFILLER_3_952 VPWR VGND sg13g2_decap_8
XFILLER_97_539 VPWR VGND sg13g2_decap_8
XFILLER_78_720 VPWR VGND sg13g2_decap_8
XFILLER_2_473 VPWR VGND sg13g2_decap_8
XFILLER_49_81 VPWR VGND sg13g2_decap_8
XFILLER_93_712 VPWR VGND sg13g2_decap_8
XFILLER_78_797 VPWR VGND sg13g2_decap_8
XFILLER_77_252 VPWR VGND sg13g2_decap_8
XFILLER_66_937 VPWR VGND sg13g2_decap_8
XFILLER_37_116 VPWR VGND sg13g2_decap_8
XFILLER_93_789 VPWR VGND sg13g2_decap_8
XFILLER_92_266 VPWR VGND sg13g2_decap_8
XFILLER_81_907 VPWR VGND sg13g2_decap_8
XFILLER_80_406 VPWR VGND sg13g2_decap_8
XFILLER_65_469 VPWR VGND sg13g2_decap_8
XFILLER_53_609 VPWR VGND sg13g2_decap_8
XFILLER_1_77 VPWR VGND sg13g2_decap_8
XFILLER_19_875 VPWR VGND sg13g2_decap_8
XFILLER_74_981 VPWR VGND sg13g2_decap_8
XFILLER_73_480 VPWR VGND sg13g2_decap_8
XFILLER_65_91 VPWR VGND sg13g2_decap_8
XFILLER_61_620 VPWR VGND sg13g2_decap_8
XFILLER_52_119 VPWR VGND sg13g2_decap_8
XFILLER_46_683 VPWR VGND sg13g2_decap_8
XFILLER_18_385 VPWR VGND sg13g2_decap_8
XFILLER_34_823 VPWR VGND sg13g2_decap_8
XFILLER_60_130 VPWR VGND sg13g2_decap_4
XFILLER_45_182 VPWR VGND sg13g2_decap_8
XFILLER_33_322 VPWR VGND sg13g2_decap_8
XFILLER_61_697 VPWR VGND sg13g2_decap_8
XFILLER_53_1022 VPWR VGND sg13g2_decap_8
XFILLER_21_539 VPWR VGND sg13g2_decap_8
XFILLER_33_399 VPWR VGND sg13g2_decap_8
XFILLER_53_0 VPWR VGND sg13g2_decap_8
XFILLER_69_764 VPWR VGND sg13g2_decap_8
XFILLER_29_18 VPWR VGND sg13g2_decap_8
XFILLER_60_1026 VPWR VGND sg13g2_fill_2
XFILLER_56_403 VPWR VGND sg13g2_decap_8
XFILLER_28_105 VPWR VGND sg13g2_decap_8
XFILLER_29_606 VPWR VGND sg13g2_decap_8
XFILLER_84_756 VPWR VGND sg13g2_decap_8
XFILLER_83_200 VPWR VGND sg13g2_decap_8
XFILLER_68_285 VPWR VGND sg13g2_decap_8
XFILLER_57_959 VPWR VGND sg13g2_decap_8
XFILLER_45_28 VPWR VGND sg13g2_decap_8
XFILLER_83_277 VPWR VGND sg13g2_decap_8
XFILLER_71_417 VPWR VGND sg13g2_decap_8
XFILLER_64_480 VPWR VGND sg13g2_decap_8
XFILLER_43_119 VPWR VGND sg13g2_decap_8
XFILLER_25_812 VPWR VGND sg13g2_decap_8
XFILLER_37_683 VPWR VGND sg13g2_decap_8
XFILLER_51_130 VPWR VGND sg13g2_decap_8
XFILLER_24_333 VPWR VGND sg13g2_decap_8
XFILLER_36_182 VPWR VGND sg13g2_decap_8
XFILLER_101_56 VPWR VGND sg13g2_decap_8
XFILLER_80_973 VPWR VGND sg13g2_decap_8
XFILLER_52_686 VPWR VGND sg13g2_decap_8
XFILLER_25_889 VPWR VGND sg13g2_decap_8
XFILLER_40_826 VPWR VGND sg13g2_decap_8
XFILLER_61_27 VPWR VGND sg13g2_decap_4
XFILLER_20_550 VPWR VGND sg13g2_decap_8
XFILLER_4_749 VPWR VGND sg13g2_decap_8
XFILLER_106_644 VPWR VGND sg13g2_decap_8
XFILLER_10_53 VPWR VGND sg13g2_decap_8
XFILLER_3_259 VPWR VGND sg13g2_decap_8
XFILLER_105_154 VPWR VGND sg13g2_decap_8
XFILLER_86_46 VPWR VGND sg13g2_decap_8
XFILLER_0_966 VPWR VGND sg13g2_decap_8
XFILLER_102_861 VPWR VGND sg13g2_decap_8
XFILLER_19_105 VPWR VGND sg13g2_decap_8
XFILLER_101_371 VPWR VGND sg13g2_decap_8
XFILLER_75_756 VPWR VGND sg13g2_decap_8
XFILLER_74_211 VPWR VGND sg13g2_decap_8
XFILLER_59_285 VPWR VGND sg13g2_decap_8
XFILLER_48_959 VPWR VGND sg13g2_decap_8
XFILLER_90_704 VPWR VGND sg13g2_decap_8
XFILLER_62_406 VPWR VGND sg13g2_decap_8
XFILLER_56_970 VPWR VGND sg13g2_decap_8
XFILLER_47_469 VPWR VGND sg13g2_decap_8
XFILLER_19_84 VPWR VGND sg13g2_decap_8
XFILLER_35_609 VPWR VGND sg13g2_decap_8
XFILLER_74_288 VPWR VGND sg13g2_decap_8
XFILLER_16_812 VPWR VGND sg13g2_decap_8
XFILLER_28_672 VPWR VGND sg13g2_decap_8
XFILLER_42_130 VPWR VGND sg13g2_decap_8
XFILLER_15_333 VPWR VGND sg13g2_decap_8
XFILLER_27_193 VPWR VGND sg13g2_decap_8
XFILLER_71_984 VPWR VGND sg13g2_decap_8
XFILLER_43_686 VPWR VGND sg13g2_decap_8
XFILLER_16_889 VPWR VGND sg13g2_decap_8
XFILLER_31_826 VPWR VGND sg13g2_decap_8
XFILLER_37_1028 VPWR VGND sg13g2_fill_1
XFILLER_70_483 VPWR VGND sg13g2_decap_8
XFILLER_30_336 VPWR VGND sg13g2_decap_8
XFILLER_51_60 VPWR VGND sg13g2_decap_8
XFILLER_7_543 VPWR VGND sg13g2_decap_8
XFILLER_83_1026 VPWR VGND sg13g2_fill_2
XFILLER_98_837 VPWR VGND sg13g2_decap_8
XFILLER_97_336 VPWR VGND sg13g2_decap_8
XFILLER_2_270 VPWR VGND sg13g2_decap_8
XFILLER_78_594 VPWR VGND sg13g2_decap_8
XFILLER_66_734 VPWR VGND sg13g2_decap_8
XFILLER_81_704 VPWR VGND sg13g2_decap_8
XFILLER_65_266 VPWR VGND sg13g2_decap_8
XFILLER_54_907 VPWR VGND sg13g2_decap_8
XFILLER_53_406 VPWR VGND sg13g2_decap_8
XFILLER_26_609 VPWR VGND sg13g2_decap_8
XFILLER_38_469 VPWR VGND sg13g2_decap_8
XFILLER_93_586 VPWR VGND sg13g2_decap_8
XFILLER_80_203 VPWR VGND sg13g2_decap_8
XFILLER_19_672 VPWR VGND sg13g2_decap_8
XFILLER_25_119 VPWR VGND sg13g2_decap_8
XFILLER_46_480 VPWR VGND sg13g2_decap_8
XFILLER_18_182 VPWR VGND sg13g2_decap_8
XFILLER_34_620 VPWR VGND sg13g2_decap_8
XFILLER_90_1019 VPWR VGND sg13g2_decap_8
XFILLER_62_973 VPWR VGND sg13g2_decap_8
XFILLER_61_494 VPWR VGND sg13g2_decap_8
XFILLER_21_336 VPWR VGND sg13g2_decap_8
XFILLER_22_837 VPWR VGND sg13g2_decap_8
XFILLER_33_196 VPWR VGND sg13g2_decap_8
XFILLER_34_697 VPWR VGND sg13g2_decap_8
Xoutput19 net19 uo_out[2] VPWR VGND sg13g2_buf_1
XFILLER_89_826 VPWR VGND sg13g2_decap_8
XFILLER_103_658 VPWR VGND sg13g2_decap_8
XFILLER_88_347 VPWR VGND sg13g2_decap_8
XFILLER_102_168 VPWR VGND sg13g2_decap_8
XFILLER_69_561 VPWR VGND sg13g2_decap_8
XFILLER_29_403 VPWR VGND sg13g2_decap_8
XFILLER_99_1022 VPWR VGND sg13g2_decap_8
XFILLER_56_200 VPWR VGND sg13g2_decap_8
XFILLER_5_1026 VPWR VGND sg13g2_fill_2
XFILLER_84_553 VPWR VGND sg13g2_decap_8
XFILLER_57_756 VPWR VGND sg13g2_decap_8
XFILLER_71_214 VPWR VGND sg13g2_decap_8
XFILLER_56_277 VPWR VGND sg13g2_decap_8
XFILLER_44_417 VPWR VGND sg13g2_decap_8
XFILLER_16_119 VPWR VGND sg13g2_decap_8
XFILLER_37_480 VPWR VGND sg13g2_decap_8
XFILLER_80_770 VPWR VGND sg13g2_decap_8
XFILLER_53_973 VPWR VGND sg13g2_decap_8
XFILLER_13_826 VPWR VGND sg13g2_decap_8
XFILLER_24_130 VPWR VGND sg13g2_decap_8
XFILLER_25_686 VPWR VGND sg13g2_decap_8
XFILLER_52_483 VPWR VGND sg13g2_decap_8
XFILLER_40_623 VPWR VGND sg13g2_decap_8
XFILLER_9_819 VPWR VGND sg13g2_decap_8
XFILLER_12_347 VPWR VGND sg13g2_decap_8
XFILLER_8_329 VPWR VGND sg13g2_decap_8
XFILLER_21_63 VPWR VGND sg13g2_decap_8
XFILLER_106_441 VPWR VGND sg13g2_decap_8
XFILLER_4_546 VPWR VGND sg13g2_decap_8
XFILLER_97_56 VPWR VGND sg13g2_decap_8
XFILLER_79_347 VPWR VGND sg13g2_decap_8
XFILLER_0_763 VPWR VGND sg13g2_decap_8
XFILLER_75_553 VPWR VGND sg13g2_decap_8
XFILLER_48_756 VPWR VGND sg13g2_decap_8
XFILLER_90_501 VPWR VGND sg13g2_decap_8
XFILLER_62_203 VPWR VGND sg13g2_decap_8
XFILLER_47_266 VPWR VGND sg13g2_decap_8
XFILLER_46_60 VPWR VGND sg13g2_decap_8
XFILLER_29_970 VPWR VGND sg13g2_decap_8
XFILLER_35_406 VPWR VGND sg13g2_decap_8
XFILLER_90_578 VPWR VGND sg13g2_decap_8
XFILLER_44_984 VPWR VGND sg13g2_decap_8
XFILLER_15_130 VPWR VGND sg13g2_decap_8
XFILLER_16_686 VPWR VGND sg13g2_decap_8
XFILLER_94_7 VPWR VGND sg13g2_decap_8
XFILLER_71_781 VPWR VGND sg13g2_decap_8
XFILLER_70_280 VPWR VGND sg13g2_decap_8
XFILLER_43_483 VPWR VGND sg13g2_decap_8
XFILLER_31_623 VPWR VGND sg13g2_decap_8
XFILLER_30_133 VPWR VGND sg13g2_decap_8
XFILLER_7_340 VPWR VGND sg13g2_decap_8
XFILLER_7_32 VPWR VGND sg13g2_decap_8
XFILLER_8_896 VPWR VGND sg13g2_decap_8
XFILLER_98_634 VPWR VGND sg13g2_decap_8
XFILLER_97_133 VPWR VGND sg13g2_decap_8
XFILLER_94_840 VPWR VGND sg13g2_decap_8
XFILLER_78_391 VPWR VGND sg13g2_decap_8
XFILLER_66_531 VPWR VGND sg13g2_decap_8
XFILLER_54_704 VPWR VGND sg13g2_decap_8
XFILLER_16_0 VPWR VGND sg13g2_decap_8
XFILLER_27_907 VPWR VGND sg13g2_decap_8
XFILLER_39_767 VPWR VGND sg13g2_decap_8
XFILLER_93_383 VPWR VGND sg13g2_decap_8
XFILLER_81_501 VPWR VGND sg13g2_decap_8
XFILLER_53_203 VPWR VGND sg13g2_decap_8
XFILLER_26_406 VPWR VGND sg13g2_decap_8
XFILLER_38_266 VPWR VGND sg13g2_decap_8
XFILLER_81_578 VPWR VGND sg13g2_decap_8
XFILLER_62_770 VPWR VGND sg13g2_decap_8
XFILLER_50_910 VPWR VGND sg13g2_decap_8
XFILLER_35_973 VPWR VGND sg13g2_decap_8
XFILLER_22_634 VPWR VGND sg13g2_decap_8
XFILLER_34_494 VPWR VGND sg13g2_decap_8
XFILLER_61_291 VPWR VGND sg13g2_decap_8
XFILLER_50_987 VPWR VGND sg13g2_decap_8
XFILLER_42_18 VPWR VGND sg13g2_decap_8
XFILLER_21_133 VPWR VGND sg13g2_decap_8
XFILLER_89_623 VPWR VGND sg13g2_decap_8
XFILLER_66_1021 VPWR VGND sg13g2_decap_8
XFILLER_104_945 VPWR VGND sg13g2_decap_8
XFILLER_27_1005 VPWR VGND sg13g2_decap_8
XFILLER_103_455 VPWR VGND sg13g2_decap_8
XFILLER_88_144 VPWR VGND sg13g2_decap_8
XFILLER_29_200 VPWR VGND sg13g2_decap_8
XFILLER_85_840 VPWR VGND sg13g2_decap_8
XFILLER_57_553 VPWR VGND sg13g2_decap_8
XFILLER_84_350 VPWR VGND sg13g2_decap_8
XFILLER_83_25 VPWR VGND sg13g2_decap_8
XFILLER_44_214 VPWR VGND sg13g2_decap_8
XFILLER_17_417 VPWR VGND sg13g2_decap_8
XFILLER_29_277 VPWR VGND sg13g2_decap_8
XFILLER_72_567 VPWR VGND sg13g2_decap_8
XFILLER_60_718 VPWR VGND sg13g2_decap_8
XFILLER_53_770 VPWR VGND sg13g2_decap_8
XFILLER_41_910 VPWR VGND sg13g2_decap_8
XFILLER_26_973 VPWR VGND sg13g2_decap_8
XFILLER_52_280 VPWR VGND sg13g2_decap_8
XFILLER_13_623 VPWR VGND sg13g2_decap_8
XFILLER_16_63 VPWR VGND sg13g2_decap_8
XFILLER_25_483 VPWR VGND sg13g2_decap_8
XFILLER_40_420 VPWR VGND sg13g2_decap_8
XFILLER_9_616 VPWR VGND sg13g2_decap_8
XFILLER_12_144 VPWR VGND sg13g2_decap_8
XFILLER_41_987 VPWR VGND sg13g2_decap_8
XFILLER_8_126 VPWR VGND sg13g2_decap_8
XFILLER_40_497 VPWR VGND sg13g2_decap_8
XFILLER_32_95 VPWR VGND sg13g2_decap_8
XFILLER_5_844 VPWR VGND sg13g2_decap_8
XFILLER_4_343 VPWR VGND sg13g2_decap_8
XFILLER_79_144 VPWR VGND sg13g2_decap_8
XFILLER_95_648 VPWR VGND sg13g2_decap_8
XFILLER_0_560 VPWR VGND sg13g2_decap_8
XFILLER_94_147 VPWR VGND sg13g2_decap_8
XFILLER_76_851 VPWR VGND sg13g2_decap_8
XFILLER_57_70 VPWR VGND sg13g2_decap_8
XFILLER_48_553 VPWR VGND sg13g2_decap_8
XFILLER_75_350 VPWR VGND sg13g2_decap_8
XFILLER_35_203 VPWR VGND sg13g2_decap_8
XFILLER_91_854 VPWR VGND sg13g2_decap_8
XFILLER_90_375 VPWR VGND sg13g2_decap_8
XFILLER_63_567 VPWR VGND sg13g2_decap_8
XFILLER_51_718 VPWR VGND sg13g2_decap_8
XFILLER_17_984 VPWR VGND sg13g2_decap_8
XFILLER_50_217 VPWR VGND sg13g2_decap_8
XFILLER_44_781 VPWR VGND sg13g2_decap_8
XFILLER_16_483 VPWR VGND sg13g2_decap_8
XFILLER_31_420 VPWR VGND sg13g2_decap_8
XFILLER_32_921 VPWR VGND sg13g2_decap_8
XFILLER_43_280 VPWR VGND sg13g2_decap_8
XFILLER_32_998 VPWR VGND sg13g2_decap_8
XFILLER_31_497 VPWR VGND sg13g2_decap_8
XFILLER_8_693 VPWR VGND sg13g2_decap_8
XFILLER_99_910 VPWR VGND sg13g2_decap_8
XFILLER_98_431 VPWR VGND sg13g2_decap_8
XFILLER_99_987 VPWR VGND sg13g2_decap_8
XFILLER_101_959 VPWR VGND sg13g2_decap_8
XFILLER_86_648 VPWR VGND sg13g2_decap_8
XFILLER_100_469 VPWR VGND sg13g2_decap_8
XFILLER_85_147 VPWR VGND sg13g2_decap_8
XFILLER_67_840 VPWR VGND sg13g2_decap_8
XFILLER_37_18 VPWR VGND sg13g2_decap_8
XFILLER_54_501 VPWR VGND sg13g2_decap_8
XFILLER_26_203 VPWR VGND sg13g2_decap_8
XFILLER_27_704 VPWR VGND sg13g2_decap_8
XFILLER_39_564 VPWR VGND sg13g2_decap_8
XFILLER_93_180 VPWR VGND sg13g2_decap_8
XFILLER_82_854 VPWR VGND sg13g2_decap_8
XFILLER_54_578 VPWR VGND sg13g2_decap_8
XFILLER_42_718 VPWR VGND sg13g2_decap_8
XFILLER_81_375 VPWR VGND sg13g2_decap_8
XFILLER_53_28 VPWR VGND sg13g2_decap_8
XFILLER_23_910 VPWR VGND sg13g2_decap_8
XFILLER_35_770 VPWR VGND sg13g2_decap_8
XFILLER_41_217 VPWR VGND sg13g2_decap_8
XFILLER_22_431 VPWR VGND sg13g2_decap_8
XFILLER_34_291 VPWR VGND sg13g2_decap_8
XFILLER_50_784 VPWR VGND sg13g2_decap_8
XFILLER_23_987 VPWR VGND sg13g2_decap_8
XFILLER_10_648 VPWR VGND sg13g2_decap_8
XFILLER_104_742 VPWR VGND sg13g2_decap_8
XFILLER_89_420 VPWR VGND sg13g2_decap_8
XFILLER_78_25 VPWR VGND sg13g2_decap_8
XFILLER_2_858 VPWR VGND sg13g2_decap_8
XFILLER_103_252 VPWR VGND sg13g2_decap_8
XFILLER_78_69 VPWR VGND sg13g2_decap_8
XFILLER_1_357 VPWR VGND sg13g2_decap_8
XFILLER_89_497 VPWR VGND sg13g2_decap_8
XFILLER_77_637 VPWR VGND sg13g2_decap_8
XFILLER_94_35 VPWR VGND sg13g2_decap_8
XFILLER_76_158 VPWR VGND sg13g2_decap_8
XFILLER_58_840 VPWR VGND sg13g2_decap_8
XFILLER_57_350 VPWR VGND sg13g2_decap_8
XFILLER_17_214 VPWR VGND sg13g2_decap_8
XFILLER_73_865 VPWR VGND sg13g2_decap_8
XFILLER_72_364 VPWR VGND sg13g2_decap_8
XFILLER_45_567 VPWR VGND sg13g2_decap_8
XFILLER_27_95 VPWR VGND sg13g2_decap_8
XFILLER_33_707 VPWR VGND sg13g2_decap_8
XFILLER_60_515 VPWR VGND sg13g2_decap_8
XFILLER_14_910 VPWR VGND sg13g2_decap_8
XFILLER_26_770 VPWR VGND sg13g2_decap_8
XFILLER_32_228 VPWR VGND sg13g2_decap_8
XFILLER_13_420 VPWR VGND sg13g2_decap_8
XFILLER_25_280 VPWR VGND sg13g2_decap_8
XFILLER_41_784 VPWR VGND sg13g2_decap_8
XFILLER_9_413 VPWR VGND sg13g2_decap_8
XFILLER_14_987 VPWR VGND sg13g2_decap_8
XFILLER_13_497 VPWR VGND sg13g2_decap_8
XFILLER_40_294 VPWR VGND sg13g2_decap_8
XFILLER_5_641 VPWR VGND sg13g2_decap_8
XFILLER_99_217 VPWR VGND sg13g2_decap_8
XFILLER_57_7 VPWR VGND sg13g2_decap_8
XFILLER_4_140 VPWR VGND sg13g2_decap_8
XFILLER_4_77 VPWR VGND sg13g2_decap_8
XFILLER_96_924 VPWR VGND sg13g2_decap_8
XFILLER_95_445 VPWR VGND sg13g2_decap_8
XFILLER_67_147 VPWR VGND sg13g2_decap_8
XFILLER_49_851 VPWR VGND sg13g2_decap_8
XFILLER_48_350 VPWR VGND sg13g2_decap_8
XFILLER_91_651 VPWR VGND sg13g2_decap_8
XFILLER_64_865 VPWR VGND sg13g2_decap_8
XFILLER_63_364 VPWR VGND sg13g2_decap_8
XFILLER_24_718 VPWR VGND sg13g2_decap_8
XFILLER_36_567 VPWR VGND sg13g2_decap_8
XFILLER_90_172 VPWR VGND sg13g2_decap_8
XFILLER_51_515 VPWR VGND sg13g2_decap_8
XFILLER_17_781 VPWR VGND sg13g2_decap_8
XFILLER_23_217 VPWR VGND sg13g2_decap_8
XFILLER_16_280 VPWR VGND sg13g2_decap_8
XFILLER_17_1026 VPWR VGND sg13g2_fill_2
XFILLER_20_935 VPWR VGND sg13g2_decap_8
XFILLER_31_294 VPWR VGND sg13g2_decap_8
XFILLER_32_795 VPWR VGND sg13g2_decap_8
XFILLER_9_980 VPWR VGND sg13g2_decap_8
XFILLER_8_490 VPWR VGND sg13g2_decap_8
XFILLER_105_539 VPWR VGND sg13g2_decap_8
XFILLER_99_784 VPWR VGND sg13g2_decap_8
XFILLER_87_924 VPWR VGND sg13g2_decap_8
XFILLER_48_28 VPWR VGND sg13g2_decap_8
XFILLER_101_756 VPWR VGND sg13g2_decap_8
XFILLER_86_445 VPWR VGND sg13g2_decap_8
XFILLER_58_147 VPWR VGND sg13g2_decap_8
XFILLER_24_1019 VPWR VGND sg13g2_decap_8
XFILLER_100_266 VPWR VGND sg13g2_decap_8
XFILLER_27_501 VPWR VGND sg13g2_decap_8
XFILLER_39_361 VPWR VGND sg13g2_decap_8
XFILLER_104_56 VPWR VGND sg13g2_decap_8
XFILLER_55_854 VPWR VGND sg13g2_decap_8
XFILLER_82_651 VPWR VGND sg13g2_decap_8
XFILLER_15_718 VPWR VGND sg13g2_decap_8
XFILLER_27_578 VPWR VGND sg13g2_decap_8
XFILLER_81_172 VPWR VGND sg13g2_decap_8
XFILLER_54_375 VPWR VGND sg13g2_decap_8
XFILLER_42_515 VPWR VGND sg13g2_decap_8
XFILLER_14_217 VPWR VGND sg13g2_decap_8
XFILLER_70_868 VPWR VGND sg13g2_decap_8
XFILLER_11_924 VPWR VGND sg13g2_decap_8
XFILLER_23_784 VPWR VGND sg13g2_decap_8
XFILLER_50_581 VPWR VGND sg13g2_decap_8
XFILLER_13_42 VPWR VGND sg13g2_decap_8
XFILLER_10_445 VPWR VGND sg13g2_decap_8
XFILLER_7_928 VPWR VGND sg13g2_decap_8
XFILLER_6_427 VPWR VGND sg13g2_decap_8
XFILLER_89_35 VPWR VGND sg13g2_decap_8
XFILLER_78_902 VPWR VGND sg13g2_decap_8
XFILLER_2_655 VPWR VGND sg13g2_decap_8
XFILLER_1_154 VPWR VGND sg13g2_decap_8
XFILLER_89_294 VPWR VGND sg13g2_decap_8
XFILLER_78_979 VPWR VGND sg13g2_decap_8
XFILLER_77_434 VPWR VGND sg13g2_decap_8
XFILLER_49_158 VPWR VGND sg13g2_decap_8
XFILLER_92_448 VPWR VGND sg13g2_decap_8
XFILLER_73_662 VPWR VGND sg13g2_decap_8
XFILLER_61_802 VPWR VGND sg13g2_decap_8
XFILLER_46_865 VPWR VGND sg13g2_decap_8
XFILLER_18_567 VPWR VGND sg13g2_decap_8
XFILLER_33_504 VPWR VGND sg13g2_decap_8
XFILLER_72_161 VPWR VGND sg13g2_decap_8
XFILLER_60_312 VPWR VGND sg13g2_decap_8
XFILLER_45_364 VPWR VGND sg13g2_decap_8
XFILLER_61_879 VPWR VGND sg13g2_decap_8
XFILLER_54_60 VPWR VGND sg13g2_decap_8
XFILLER_60_389 VPWR VGND sg13g2_decap_8
XFILLER_14_784 VPWR VGND sg13g2_decap_8
XFILLER_9_210 VPWR VGND sg13g2_decap_8
XFILLER_13_294 VPWR VGND sg13g2_decap_8
XFILLER_41_581 VPWR VGND sg13g2_decap_8
XFILLER_70_70 VPWR VGND sg13g2_decap_8
XFILLER_9_287 VPWR VGND sg13g2_decap_8
XFILLER_47_1008 VPWR VGND sg13g2_decap_8
XFILLER_6_994 VPWR VGND sg13g2_decap_8
XFILLER_96_721 VPWR VGND sg13g2_decap_8
XFILLER_69_946 VPWR VGND sg13g2_decap_8
XFILLER_95_242 VPWR VGND sg13g2_decap_8
XFILLER_96_798 VPWR VGND sg13g2_decap_8
XFILLER_84_938 VPWR VGND sg13g2_decap_8
XFILLER_68_467 VPWR VGND sg13g2_decap_8
XFILLER_83_459 VPWR VGND sg13g2_decap_8
XFILLER_64_662 VPWR VGND sg13g2_decap_8
XFILLER_37_865 VPWR VGND sg13g2_decap_8
XFILLER_93_1006 VPWR VGND sg13g2_decap_8
XFILLER_63_161 VPWR VGND sg13g2_decap_8
XFILLER_51_312 VPWR VGND sg13g2_decap_8
XFILLER_24_515 VPWR VGND sg13g2_decap_8
XFILLER_36_364 VPWR VGND sg13g2_decap_8
XFILLER_52_868 VPWR VGND sg13g2_decap_8
XFILLER_51_389 VPWR VGND sg13g2_decap_8
XFILLER_20_732 VPWR VGND sg13g2_decap_8
XFILLER_32_592 VPWR VGND sg13g2_decap_8
XFILLER_30_1001 VPWR VGND sg13g2_decap_8
XFILLER_106_826 VPWR VGND sg13g2_decap_8
XFILLER_105_336 VPWR VGND sg13g2_decap_8
XFILLER_78_209 VPWR VGND sg13g2_decap_8
XFILLER_99_581 VPWR VGND sg13g2_decap_8
XFILLER_87_721 VPWR VGND sg13g2_decap_8
XFILLER_101_553 VPWR VGND sg13g2_decap_8
XFILLER_87_798 VPWR VGND sg13g2_decap_8
XFILLER_86_242 VPWR VGND sg13g2_decap_8
XFILLER_75_938 VPWR VGND sg13g2_decap_8
XFILLER_59_467 VPWR VGND sg13g2_decap_8
XFILLER_55_651 VPWR VGND sg13g2_decap_8
XFILLER_28_854 VPWR VGND sg13g2_decap_8
XFILLER_91_14 VPWR VGND sg13g2_decap_8
XFILLER_61_109 VPWR VGND sg13g2_decap_8
XFILLER_54_172 VPWR VGND sg13g2_decap_8
XFILLER_42_312 VPWR VGND sg13g2_decap_8
XFILLER_15_515 VPWR VGND sg13g2_decap_8
XFILLER_27_375 VPWR VGND sg13g2_decap_8
XFILLER_43_868 VPWR VGND sg13g2_decap_8
XFILLER_70_665 VPWR VGND sg13g2_decap_8
XFILLER_42_389 VPWR VGND sg13g2_decap_8
XFILLER_30_518 VPWR VGND sg13g2_decap_8
XFILLER_11_721 VPWR VGND sg13g2_decap_8
XFILLER_23_581 VPWR VGND sg13g2_decap_8
XFILLER_24_74 VPWR VGND sg13g2_decap_8
XFILLER_10_242 VPWR VGND sg13g2_decap_8
XFILLER_7_725 VPWR VGND sg13g2_decap_8
XFILLER_6_224 VPWR VGND sg13g2_decap_8
XFILLER_11_798 VPWR VGND sg13g2_decap_8
XFILLER_3_931 VPWR VGND sg13g2_decap_8
XFILLER_40_84 VPWR VGND sg13g2_decap_8
XFILLER_97_518 VPWR VGND sg13g2_decap_8
XFILLER_2_452 VPWR VGND sg13g2_decap_8
XFILLER_77_231 VPWR VGND sg13g2_decap_8
XFILLER_49_60 VPWR VGND sg13g2_decap_8
XFILLER_78_776 VPWR VGND sg13g2_decap_8
XFILLER_66_916 VPWR VGND sg13g2_decap_8
XFILLER_65_448 VPWR VGND sg13g2_decap_8
XFILLER_1_56 VPWR VGND sg13g2_decap_8
XFILLER_93_768 VPWR VGND sg13g2_decap_8
XFILLER_92_245 VPWR VGND sg13g2_decap_8
XFILLER_74_960 VPWR VGND sg13g2_decap_8
XFILLER_46_662 VPWR VGND sg13g2_decap_8
XFILLER_19_854 VPWR VGND sg13g2_decap_8
XFILLER_34_802 VPWR VGND sg13g2_decap_8
XFILLER_65_70 VPWR VGND sg13g2_decap_8
XFILLER_45_161 VPWR VGND sg13g2_decap_8
XFILLER_18_364 VPWR VGND sg13g2_decap_8
XFILLER_33_301 VPWR VGND sg13g2_decap_8
XFILLER_61_676 VPWR VGND sg13g2_decap_8
XFILLER_53_1001 VPWR VGND sg13g2_decap_8
XFILLER_21_518 VPWR VGND sg13g2_decap_8
XFILLER_33_378 VPWR VGND sg13g2_decap_8
XFILLER_34_879 VPWR VGND sg13g2_decap_8
XFILLER_60_186 VPWR VGND sg13g2_decap_8
XFILLER_14_581 VPWR VGND sg13g2_decap_8
XFILLER_6_791 VPWR VGND sg13g2_decap_8
XFILLER_88_529 VPWR VGND sg13g2_decap_8
XFILLER_69_743 VPWR VGND sg13g2_decap_8
XFILLER_60_1005 VPWR VGND sg13g2_decap_8
XFILLER_68_264 VPWR VGND sg13g2_decap_8
XFILLER_57_938 VPWR VGND sg13g2_decap_8
XFILLER_96_595 VPWR VGND sg13g2_decap_8
XFILLER_84_735 VPWR VGND sg13g2_decap_8
XFILLER_83_256 VPWR VGND sg13g2_decap_8
XFILLER_56_459 VPWR VGND sg13g2_decap_8
XFILLER_36_161 VPWR VGND sg13g2_decap_8
XFILLER_37_662 VPWR VGND sg13g2_decap_8
XFILLER_80_952 VPWR VGND sg13g2_decap_8
XFILLER_24_312 VPWR VGND sg13g2_decap_8
XFILLER_25_868 VPWR VGND sg13g2_decap_8
XFILLER_101_35 VPWR VGND sg13g2_decap_8
XFILLER_52_665 VPWR VGND sg13g2_decap_8
XFILLER_40_805 VPWR VGND sg13g2_decap_8
XFILLER_51_186 VPWR VGND sg13g2_decap_8
XFILLER_12_529 VPWR VGND sg13g2_decap_8
XFILLER_24_389 VPWR VGND sg13g2_decap_8
XFILLER_106_623 VPWR VGND sg13g2_decap_8
XFILLER_4_728 VPWR VGND sg13g2_decap_8
XFILLER_105_133 VPWR VGND sg13g2_decap_8
XFILLER_10_32 VPWR VGND sg13g2_decap_8
XFILLER_3_238 VPWR VGND sg13g2_decap_8
XFILLER_79_529 VPWR VGND sg13g2_decap_8
XFILLER_102_840 VPWR VGND sg13g2_decap_8
XFILLER_86_25 VPWR VGND sg13g2_decap_8
XFILLER_0_945 VPWR VGND sg13g2_decap_8
XFILLER_101_350 VPWR VGND sg13g2_decap_8
XFILLER_59_264 VPWR VGND sg13g2_decap_8
XFILLER_87_595 VPWR VGND sg13g2_decap_8
XFILLER_75_735 VPWR VGND sg13g2_decap_8
XFILLER_48_938 VPWR VGND sg13g2_decap_8
XFILLER_19_63 VPWR VGND sg13g2_decap_8
XFILLER_47_448 VPWR VGND sg13g2_decap_8
XFILLER_28_651 VPWR VGND sg13g2_decap_8
XFILLER_76_1012 VPWR VGND sg13g2_decap_8
XFILLER_74_267 VPWR VGND sg13g2_decap_8
XFILLER_34_109 VPWR VGND sg13g2_decap_8
XFILLER_71_963 VPWR VGND sg13g2_decap_8
XFILLER_15_312 VPWR VGND sg13g2_decap_8
XFILLER_16_868 VPWR VGND sg13g2_decap_8
XFILLER_27_172 VPWR VGND sg13g2_decap_8
XFILLER_70_462 VPWR VGND sg13g2_decap_8
XFILLER_43_665 VPWR VGND sg13g2_decap_8
XFILLER_31_805 VPWR VGND sg13g2_decap_8
XFILLER_35_84 VPWR VGND sg13g2_decap_8
XFILLER_42_186 VPWR VGND sg13g2_decap_8
XFILLER_15_389 VPWR VGND sg13g2_decap_8
XFILLER_30_315 VPWR VGND sg13g2_decap_8
XFILLER_7_522 VPWR VGND sg13g2_decap_8
XFILLER_11_595 VPWR VGND sg13g2_decap_8
XFILLER_7_599 VPWR VGND sg13g2_decap_8
XFILLER_98_816 VPWR VGND sg13g2_decap_8
XFILLER_83_1005 VPWR VGND sg13g2_decap_8
XFILLER_97_315 VPWR VGND sg13g2_decap_8
XFILLER_78_573 VPWR VGND sg13g2_decap_8
XFILLER_66_713 VPWR VGND sg13g2_decap_8
XFILLER_39_949 VPWR VGND sg13g2_decap_8
XFILLER_93_565 VPWR VGND sg13g2_decap_8
XFILLER_65_245 VPWR VGND sg13g2_decap_8
XFILLER_19_651 VPWR VGND sg13g2_decap_8
XFILLER_38_448 VPWR VGND sg13g2_decap_8
XFILLER_18_161 VPWR VGND sg13g2_decap_8
XFILLER_62_952 VPWR VGND sg13g2_decap_8
XFILLER_80_259 VPWR VGND sg13g2_decap_8
XFILLER_22_816 VPWR VGND sg13g2_decap_8
XFILLER_34_676 VPWR VGND sg13g2_decap_8
XFILLER_61_473 VPWR VGND sg13g2_decap_8
XFILLER_21_315 VPWR VGND sg13g2_decap_8
XFILLER_33_175 VPWR VGND sg13g2_decap_8
XFILLER_30_882 VPWR VGND sg13g2_decap_8
XFILLER_89_805 VPWR VGND sg13g2_decap_8
XFILLER_103_637 VPWR VGND sg13g2_decap_8
XFILLER_88_326 VPWR VGND sg13g2_decap_8
XFILLER_102_147 VPWR VGND sg13g2_decap_8
XFILLER_69_540 VPWR VGND sg13g2_decap_8
XFILLER_5_1005 VPWR VGND sg13g2_decap_8
XFILLER_99_1001 VPWR VGND sg13g2_decap_8
XFILLER_97_882 VPWR VGND sg13g2_decap_8
XFILLER_57_735 VPWR VGND sg13g2_decap_8
XFILLER_96_392 VPWR VGND sg13g2_decap_8
XFILLER_84_532 VPWR VGND sg13g2_decap_8
XFILLER_56_256 VPWR VGND sg13g2_decap_8
XFILLER_56_39 VPWR VGND sg13g2_decap_8
XFILLER_29_459 VPWR VGND sg13g2_decap_8
XFILLER_72_749 VPWR VGND sg13g2_decap_8
XFILLER_53_952 VPWR VGND sg13g2_decap_8
XFILLER_72_49 VPWR VGND sg13g2_decap_8
XFILLER_52_462 VPWR VGND sg13g2_decap_8
XFILLER_13_805 VPWR VGND sg13g2_decap_8
XFILLER_25_665 VPWR VGND sg13g2_decap_8
XFILLER_40_602 VPWR VGND sg13g2_decap_8
XFILLER_12_326 VPWR VGND sg13g2_decap_8
XFILLER_24_186 VPWR VGND sg13g2_decap_8
XFILLER_8_308 VPWR VGND sg13g2_decap_8
XFILLER_40_679 VPWR VGND sg13g2_decap_8
XFILLER_21_882 VPWR VGND sg13g2_decap_8
XFILLER_4_525 VPWR VGND sg13g2_decap_8
XFILLER_21_42 VPWR VGND sg13g2_decap_8
XFILLER_106_420 VPWR VGND sg13g2_decap_8
XFILLER_97_35 VPWR VGND sg13g2_decap_8
XFILLER_106_497 VPWR VGND sg13g2_decap_8
XFILLER_79_326 VPWR VGND sg13g2_decap_8
XFILLER_43_1022 VPWR VGND sg13g2_decap_8
XFILLER_0_742 VPWR VGND sg13g2_decap_8
XFILLER_94_329 VPWR VGND sg13g2_decap_8
XFILLER_88_893 VPWR VGND sg13g2_decap_8
XFILLER_48_735 VPWR VGND sg13g2_decap_8
XFILLER_87_392 VPWR VGND sg13g2_decap_8
XFILLER_75_532 VPWR VGND sg13g2_decap_8
XFILLER_47_245 VPWR VGND sg13g2_decap_8
XFILLER_90_557 VPWR VGND sg13g2_decap_8
XFILLER_63_749 VPWR VGND sg13g2_decap_8
XFILLER_71_760 VPWR VGND sg13g2_decap_8
XFILLER_62_259 VPWR VGND sg13g2_decap_8
XFILLER_44_963 VPWR VGND sg13g2_decap_8
XFILLER_43_462 VPWR VGND sg13g2_decap_8
XFILLER_16_665 VPWR VGND sg13g2_decap_8
XFILLER_31_602 VPWR VGND sg13g2_decap_8
XFILLER_15_186 VPWR VGND sg13g2_decap_8
XFILLER_30_112 VPWR VGND sg13g2_decap_8
XFILLER_87_7 VPWR VGND sg13g2_decap_8
XFILLER_50_1015 VPWR VGND sg13g2_decap_8
XFILLER_7_11 VPWR VGND sg13g2_decap_8
XFILLER_31_679 VPWR VGND sg13g2_decap_8
XFILLER_11_392 VPWR VGND sg13g2_decap_8
XFILLER_12_893 VPWR VGND sg13g2_decap_8
XFILLER_30_189 VPWR VGND sg13g2_decap_8
XFILLER_8_875 VPWR VGND sg13g2_decap_8
XFILLER_7_88 VPWR VGND sg13g2_decap_8
XFILLER_7_396 VPWR VGND sg13g2_decap_8
XFILLER_98_613 VPWR VGND sg13g2_decap_8
XFILLER_97_112 VPWR VGND sg13g2_decap_8
XFILLER_97_189 VPWR VGND sg13g2_decap_8
XFILLER_85_329 VPWR VGND sg13g2_decap_8
XFILLER_79_893 VPWR VGND sg13g2_decap_8
XFILLER_78_370 VPWR VGND sg13g2_decap_8
XFILLER_66_510 VPWR VGND sg13g2_decap_8
XFILLER_38_245 VPWR VGND sg13g2_decap_8
XFILLER_39_746 VPWR VGND sg13g2_decap_8
XFILLER_94_896 VPWR VGND sg13g2_decap_8
XFILLER_93_362 VPWR VGND sg13g2_decap_8
XFILLER_66_587 VPWR VGND sg13g2_decap_8
XFILLER_81_557 VPWR VGND sg13g2_decap_8
XFILLER_53_259 VPWR VGND sg13g2_decap_8
XFILLER_35_952 VPWR VGND sg13g2_decap_8
XFILLER_61_270 VPWR VGND sg13g2_decap_8
XFILLER_21_112 VPWR VGND sg13g2_decap_8
XFILLER_22_613 VPWR VGND sg13g2_decap_8
XFILLER_34_473 VPWR VGND sg13g2_decap_8
XFILLER_50_966 VPWR VGND sg13g2_decap_8
XFILLER_21_189 VPWR VGND sg13g2_decap_8
XFILLER_66_1000 VPWR VGND sg13g2_decap_8
XFILLER_104_924 VPWR VGND sg13g2_decap_8
XFILLER_89_602 VPWR VGND sg13g2_decap_8
XFILLER_103_434 VPWR VGND sg13g2_decap_8
XFILLER_88_123 VPWR VGND sg13g2_decap_8
XFILLER_1_539 VPWR VGND sg13g2_decap_8
XFILLER_27_1028 VPWR VGND sg13g2_fill_1
XFILLER_89_679 VPWR VGND sg13g2_decap_8
XFILLER_77_819 VPWR VGND sg13g2_decap_8
XFILLER_67_38 VPWR VGND sg13g2_decap_8
XFILLER_57_532 VPWR VGND sg13g2_decap_8
XFILLER_85_896 VPWR VGND sg13g2_decap_8
XFILLER_29_256 VPWR VGND sg13g2_decap_8
XFILLER_72_546 VPWR VGND sg13g2_decap_8
XFILLER_45_749 VPWR VGND sg13g2_decap_8
XFILLER_16_42 VPWR VGND sg13g2_decap_8
XFILLER_26_952 VPWR VGND sg13g2_decap_8
XFILLER_73_1026 VPWR VGND sg13g2_fill_2
XFILLER_13_602 VPWR VGND sg13g2_decap_8
XFILLER_25_462 VPWR VGND sg13g2_decap_8
XFILLER_41_966 VPWR VGND sg13g2_decap_8
XFILLER_12_123 VPWR VGND sg13g2_decap_8
XFILLER_8_105 VPWR VGND sg13g2_decap_8
XFILLER_13_679 VPWR VGND sg13g2_decap_8
XFILLER_40_476 VPWR VGND sg13g2_decap_8
XFILLER_32_74 VPWR VGND sg13g2_decap_8
XFILLER_5_823 VPWR VGND sg13g2_decap_8
XFILLER_4_322 VPWR VGND sg13g2_decap_8
XFILLER_106_294 VPWR VGND sg13g2_decap_8
XFILLER_79_123 VPWR VGND sg13g2_decap_8
XFILLER_4_399 VPWR VGND sg13g2_decap_8
XFILLER_80_1008 VPWR VGND sg13g2_decap_8
XFILLER_95_627 VPWR VGND sg13g2_decap_8
XFILLER_94_126 VPWR VGND sg13g2_decap_8
XFILLER_67_329 VPWR VGND sg13g2_decap_8
XFILLER_88_690 VPWR VGND sg13g2_decap_8
XFILLER_76_830 VPWR VGND sg13g2_decap_8
XFILLER_48_532 VPWR VGND sg13g2_decap_8
XFILLER_91_833 VPWR VGND sg13g2_decap_8
XFILLER_63_546 VPWR VGND sg13g2_decap_8
XFILLER_36_749 VPWR VGND sg13g2_decap_8
XFILLER_90_354 VPWR VGND sg13g2_decap_8
XFILLER_44_760 VPWR VGND sg13g2_decap_8
XFILLER_17_963 VPWR VGND sg13g2_decap_8
XFILLER_32_900 VPWR VGND sg13g2_decap_8
XFILLER_35_259 VPWR VGND sg13g2_decap_8
XFILLER_73_81 VPWR VGND sg13g2_decap_8
XFILLER_16_462 VPWR VGND sg13g2_decap_8
XFILLER_32_977 VPWR VGND sg13g2_decap_8
XFILLER_31_476 VPWR VGND sg13g2_decap_8
XFILLER_12_690 VPWR VGND sg13g2_decap_8
XFILLER_89_1022 VPWR VGND sg13g2_decap_8
XFILLER_8_672 VPWR VGND sg13g2_decap_8
XFILLER_7_193 VPWR VGND sg13g2_decap_8
XFILLER_98_410 VPWR VGND sg13g2_decap_8
XFILLER_99_966 VPWR VGND sg13g2_decap_8
XFILLER_101_938 VPWR VGND sg13g2_decap_8
XFILLER_98_487 VPWR VGND sg13g2_decap_8
XFILLER_86_627 VPWR VGND sg13g2_decap_8
XFILLER_58_329 VPWR VGND sg13g2_decap_8
XFILLER_100_448 VPWR VGND sg13g2_decap_8
XFILLER_85_126 VPWR VGND sg13g2_decap_8
XFILLER_79_690 VPWR VGND sg13g2_decap_8
XFILLER_39_543 VPWR VGND sg13g2_decap_8
XFILLER_67_896 VPWR VGND sg13g2_decap_8
XFILLER_2_1019 VPWR VGND sg13g2_decap_8
XFILLER_96_1015 VPWR VGND sg13g2_decap_8
XFILLER_94_693 VPWR VGND sg13g2_decap_8
XFILLER_82_833 VPWR VGND sg13g2_decap_8
XFILLER_66_384 VPWR VGND sg13g2_decap_8
XFILLER_81_354 VPWR VGND sg13g2_decap_8
XFILLER_54_557 VPWR VGND sg13g2_decap_8
XFILLER_26_259 VPWR VGND sg13g2_decap_8
XFILLER_22_410 VPWR VGND sg13g2_decap_8
XFILLER_34_270 VPWR VGND sg13g2_decap_8
XFILLER_23_966 VPWR VGND sg13g2_decap_8
XFILLER_50_763 VPWR VGND sg13g2_decap_8
XFILLER_10_627 VPWR VGND sg13g2_decap_8
XFILLER_6_609 VPWR VGND sg13g2_decap_8
XFILLER_22_487 VPWR VGND sg13g2_decap_8
XFILLER_104_721 VPWR VGND sg13g2_decap_8
XFILLER_2_837 VPWR VGND sg13g2_decap_8
XFILLER_103_231 VPWR VGND sg13g2_decap_8
XFILLER_1_336 VPWR VGND sg13g2_decap_8
XFILLER_104_798 VPWR VGND sg13g2_decap_8
XFILLER_89_476 VPWR VGND sg13g2_decap_8
XFILLER_77_616 VPWR VGND sg13g2_decap_8
XFILLER_94_14 VPWR VGND sg13g2_decap_8
XFILLER_76_137 VPWR VGND sg13g2_decap_8
XFILLER_58_896 VPWR VGND sg13g2_decap_8
XFILLER_85_693 VPWR VGND sg13g2_decap_8
XFILLER_73_844 VPWR VGND sg13g2_decap_8
XFILLER_45_546 VPWR VGND sg13g2_decap_8
XFILLER_18_749 VPWR VGND sg13g2_decap_8
XFILLER_72_343 VPWR VGND sg13g2_decap_8
XFILLER_27_74 VPWR VGND sg13g2_decap_8
XFILLER_32_207 VPWR VGND sg13g2_decap_8
XFILLER_14_966 VPWR VGND sg13g2_decap_8
XFILLER_41_763 VPWR VGND sg13g2_decap_8
XFILLER_13_476 VPWR VGND sg13g2_decap_8
XFILLER_43_84 VPWR VGND sg13g2_decap_8
XFILLER_40_273 VPWR VGND sg13g2_decap_8
XFILLER_9_469 VPWR VGND sg13g2_decap_8
XFILLER_5_620 VPWR VGND sg13g2_decap_8
XFILLER_5_697 VPWR VGND sg13g2_decap_8
XFILLER_96_903 VPWR VGND sg13g2_decap_8
XFILLER_4_196 VPWR VGND sg13g2_decap_8
XFILLER_4_56 VPWR VGND sg13g2_decap_8
XFILLER_95_424 VPWR VGND sg13g2_decap_8
XFILLER_68_649 VPWR VGND sg13g2_decap_8
XFILLER_67_126 VPWR VGND sg13g2_decap_8
XFILLER_49_830 VPWR VGND sg13g2_decap_8
XFILLER_91_630 VPWR VGND sg13g2_decap_8
XFILLER_64_844 VPWR VGND sg13g2_decap_8
XFILLER_84_91 VPWR VGND sg13g2_decap_8
XFILLER_63_343 VPWR VGND sg13g2_decap_8
XFILLER_36_546 VPWR VGND sg13g2_decap_8
XFILLER_90_151 VPWR VGND sg13g2_decap_8
XFILLER_17_760 VPWR VGND sg13g2_decap_8
XFILLER_17_1005 VPWR VGND sg13g2_decap_8
XFILLER_20_914 VPWR VGND sg13g2_decap_8
XFILLER_32_774 VPWR VGND sg13g2_decap_8
XFILLER_104_1008 VPWR VGND sg13g2_decap_8
XFILLER_31_273 VPWR VGND sg13g2_decap_8
XFILLER_105_518 VPWR VGND sg13g2_decap_8
XFILLER_99_763 VPWR VGND sg13g2_decap_8
XFILLER_87_903 VPWR VGND sg13g2_decap_8
XFILLER_86_424 VPWR VGND sg13g2_decap_8
XFILLER_101_735 VPWR VGND sg13g2_decap_8
XFILLER_98_284 VPWR VGND sg13g2_decap_8
XFILLER_59_649 VPWR VGND sg13g2_decap_8
XFILLER_58_137 VPWR VGND sg13g2_fill_2
XFILLER_58_126 VPWR VGND sg13g2_decap_8
XFILLER_104_35 VPWR VGND sg13g2_decap_8
XFILLER_100_245 VPWR VGND sg13g2_decap_8
XFILLER_39_340 VPWR VGND sg13g2_decap_8
XFILLER_95_991 VPWR VGND sg13g2_decap_8
XFILLER_94_490 VPWR VGND sg13g2_decap_8
XFILLER_82_630 VPWR VGND sg13g2_decap_8
XFILLER_67_693 VPWR VGND sg13g2_decap_8
XFILLER_66_181 VPWR VGND sg13g2_decap_8
XFILLER_55_833 VPWR VGND sg13g2_decap_8
XFILLER_64_39 VPWR VGND sg13g2_decap_8
XFILLER_54_354 VPWR VGND sg13g2_decap_8
XFILLER_27_557 VPWR VGND sg13g2_decap_8
XFILLER_81_151 VPWR VGND sg13g2_decap_8
XFILLER_70_847 VPWR VGND sg13g2_decap_8
XFILLER_50_560 VPWR VGND sg13g2_decap_8
XFILLER_11_903 VPWR VGND sg13g2_decap_8
XFILLER_23_763 VPWR VGND sg13g2_decap_8
XFILLER_80_49 VPWR VGND sg13g2_decap_8
XFILLER_10_424 VPWR VGND sg13g2_decap_8
XFILLER_7_907 VPWR VGND sg13g2_decap_8
XFILLER_13_21 VPWR VGND sg13g2_decap_8
XFILLER_22_284 VPWR VGND sg13g2_decap_8
XFILLER_6_406 VPWR VGND sg13g2_decap_8
XFILLER_89_14 VPWR VGND sg13g2_decap_8
XFILLER_13_98 VPWR VGND sg13g2_decap_8
XFILLER_2_634 VPWR VGND sg13g2_decap_8
XFILLER_1_133 VPWR VGND sg13g2_decap_8
XFILLER_89_273 VPWR VGND sg13g2_decap_8
XFILLER_77_413 VPWR VGND sg13g2_decap_8
XFILLER_104_595 VPWR VGND sg13g2_decap_8
XFILLER_78_958 VPWR VGND sg13g2_decap_8
XFILLER_49_137 VPWR VGND sg13g2_decap_8
XFILLER_92_427 VPWR VGND sg13g2_decap_8
XFILLER_86_991 VPWR VGND sg13g2_decap_8
XFILLER_58_693 VPWR VGND sg13g2_decap_8
XFILLER_46_844 VPWR VGND sg13g2_decap_8
XFILLER_38_84 VPWR VGND sg13g2_decap_8
XFILLER_85_490 VPWR VGND sg13g2_decap_8
XFILLER_73_641 VPWR VGND sg13g2_decap_8
XFILLER_72_140 VPWR VGND sg13g2_decap_8
XFILLER_45_343 VPWR VGND sg13g2_decap_8
XFILLER_18_546 VPWR VGND sg13g2_decap_8
XFILLER_61_858 VPWR VGND sg13g2_decap_8
XFILLER_60_368 VPWR VGND sg13g2_decap_8
XFILLER_14_763 VPWR VGND sg13g2_decap_8
XFILLER_41_560 VPWR VGND sg13g2_decap_8
XFILLER_13_273 VPWR VGND sg13g2_decap_8
XFILLER_9_266 VPWR VGND sg13g2_decap_8
XFILLER_10_991 VPWR VGND sg13g2_decap_8
XFILLER_6_973 VPWR VGND sg13g2_decap_8
XFILLER_5_494 VPWR VGND sg13g2_decap_8
XFILLER_96_700 VPWR VGND sg13g2_decap_8
XFILLER_69_925 VPWR VGND sg13g2_decap_8
XFILLER_95_221 VPWR VGND sg13g2_decap_8
XFILLER_68_446 VPWR VGND sg13g2_decap_8
XFILLER_96_777 VPWR VGND sg13g2_decap_8
XFILLER_84_917 VPWR VGND sg13g2_decap_8
XFILLER_95_298 VPWR VGND sg13g2_decap_8
XFILLER_83_438 VPWR VGND sg13g2_decap_8
XFILLER_77_980 VPWR VGND sg13g2_decap_8
XFILLER_37_844 VPWR VGND sg13g2_decap_8
XFILLER_64_641 VPWR VGND sg13g2_decap_8
XFILLER_36_343 VPWR VGND sg13g2_decap_8
XFILLER_92_994 VPWR VGND sg13g2_decap_8
XFILLER_63_140 VPWR VGND sg13g2_decap_8
XFILLER_52_847 VPWR VGND sg13g2_decap_8
XFILLER_51_368 VPWR VGND sg13g2_decap_8
XFILLER_20_711 VPWR VGND sg13g2_decap_8
XFILLER_32_571 VPWR VGND sg13g2_decap_8
XFILLER_20_788 VPWR VGND sg13g2_decap_8
XFILLER_106_805 VPWR VGND sg13g2_decap_8
XFILLER_105_315 VPWR VGND sg13g2_decap_8
XFILLER_59_39 VPWR VGND sg13g2_decap_8
XFILLER_99_560 VPWR VGND sg13g2_decap_8
XFILLER_87_700 VPWR VGND sg13g2_decap_8
XFILLER_101_532 VPWR VGND sg13g2_decap_8
XFILLER_86_221 VPWR VGND sg13g2_decap_8
XFILLER_59_446 VPWR VGND sg13g2_decap_8
XFILLER_87_777 VPWR VGND sg13g2_decap_8
XFILLER_75_917 VPWR VGND sg13g2_decap_8
XFILLER_86_298 VPWR VGND sg13g2_decap_8
XFILLER_75_49 VPWR VGND sg13g2_decap_8
XFILLER_74_449 VPWR VGND sg13g2_decap_8
XFILLER_28_833 VPWR VGND sg13g2_decap_8
XFILLER_67_490 VPWR VGND sg13g2_decap_8
XFILLER_55_630 VPWR VGND sg13g2_decap_8
XFILLER_54_151 VPWR VGND sg13g2_decap_8
XFILLER_27_354 VPWR VGND sg13g2_decap_8
XFILLER_70_644 VPWR VGND sg13g2_decap_8
XFILLER_43_847 VPWR VGND sg13g2_decap_8
XFILLER_42_368 VPWR VGND sg13g2_decap_8
XFILLER_11_700 VPWR VGND sg13g2_decap_8
XFILLER_23_560 VPWR VGND sg13g2_decap_8
XFILLER_24_53 VPWR VGND sg13g2_decap_8
XFILLER_10_221 VPWR VGND sg13g2_decap_8
XFILLER_7_704 VPWR VGND sg13g2_decap_8
XFILLER_6_203 VPWR VGND sg13g2_decap_8
XFILLER_11_777 VPWR VGND sg13g2_decap_8
XFILLER_10_298 VPWR VGND sg13g2_decap_8
XFILLER_40_63 VPWR VGND sg13g2_decap_8
XFILLER_3_910 VPWR VGND sg13g2_decap_8
XFILLER_6_0 VPWR VGND sg13g2_decap_8
XFILLER_2_431 VPWR VGND sg13g2_decap_8
XFILLER_105_882 VPWR VGND sg13g2_decap_8
XFILLER_3_987 VPWR VGND sg13g2_decap_8
XFILLER_104_392 VPWR VGND sg13g2_decap_8
XFILLER_78_755 VPWR VGND sg13g2_decap_8
XFILLER_77_210 VPWR VGND sg13g2_decap_8
XFILLER_93_747 VPWR VGND sg13g2_decap_8
XFILLER_92_224 VPWR VGND sg13g2_decap_8
XFILLER_77_287 VPWR VGND sg13g2_decap_8
XFILLER_65_427 VPWR VGND sg13g2_decap_8
XFILLER_1_35 VPWR VGND sg13g2_decap_8
XFILLER_19_833 VPWR VGND sg13g2_decap_8
XFILLER_58_490 VPWR VGND sg13g2_decap_8
XFILLER_46_641 VPWR VGND sg13g2_decap_8
XFILLER_18_343 VPWR VGND sg13g2_decap_8
XFILLER_45_140 VPWR VGND sg13g2_decap_8
XFILLER_61_655 VPWR VGND sg13g2_decap_8
XFILLER_34_858 VPWR VGND sg13g2_decap_8
XFILLER_60_165 VPWR VGND sg13g2_decap_8
XFILLER_33_357 VPWR VGND sg13g2_decap_8
XFILLER_81_81 VPWR VGND sg13g2_decap_8
XFILLER_14_560 VPWR VGND sg13g2_decap_8
XFILLER_14_1008 VPWR VGND sg13g2_decap_8
XFILLER_6_770 VPWR VGND sg13g2_decap_8
XFILLER_88_508 VPWR VGND sg13g2_decap_8
XFILLER_5_291 VPWR VGND sg13g2_decap_8
XFILLER_103_819 VPWR VGND sg13g2_decap_8
XFILLER_102_329 VPWR VGND sg13g2_decap_8
XFILLER_69_722 VPWR VGND sg13g2_decap_8
XFILLER_96_574 VPWR VGND sg13g2_decap_8
XFILLER_84_714 VPWR VGND sg13g2_decap_8
XFILLER_68_243 VPWR VGND sg13g2_decap_8
XFILLER_60_1028 VPWR VGND sg13g2_fill_1
XFILLER_57_917 VPWR VGND sg13g2_decap_8
XFILLER_69_799 VPWR VGND sg13g2_decap_8
Xinput1 ui_in[0] net1 VPWR VGND sg13g2_buf_1
XFILLER_56_438 VPWR VGND sg13g2_decap_8
XFILLER_83_235 VPWR VGND sg13g2_decap_8
XFILLER_37_641 VPWR VGND sg13g2_decap_8
XFILLER_65_994 VPWR VGND sg13g2_decap_8
XFILLER_36_140 VPWR VGND sg13g2_decap_8
XFILLER_101_14 VPWR VGND sg13g2_decap_8
XFILLER_92_791 VPWR VGND sg13g2_decap_8
XFILLER_80_931 VPWR VGND sg13g2_decap_8
XFILLER_52_644 VPWR VGND sg13g2_decap_8
XFILLER_25_847 VPWR VGND sg13g2_decap_8
XFILLER_12_508 VPWR VGND sg13g2_decap_8
XFILLER_24_368 VPWR VGND sg13g2_decap_8
XFILLER_51_165 VPWR VGND sg13g2_decap_8
XFILLER_20_585 VPWR VGND sg13g2_decap_8
XFILLER_4_707 VPWR VGND sg13g2_decap_8
XFILLER_106_602 VPWR VGND sg13g2_decap_8
XFILLER_10_11 VPWR VGND sg13g2_decap_8
XFILLER_3_217 VPWR VGND sg13g2_decap_8
XFILLER_105_112 VPWR VGND sg13g2_decap_8
XFILLER_106_679 VPWR VGND sg13g2_decap_8
XFILLER_79_508 VPWR VGND sg13g2_decap_8
XFILLER_10_88 VPWR VGND sg13g2_decap_8
XFILLER_105_189 VPWR VGND sg13g2_decap_8
XFILLER_0_924 VPWR VGND sg13g2_decap_8
XFILLER_59_243 VPWR VGND sg13g2_decap_8
XFILLER_48_917 VPWR VGND sg13g2_decap_8
XFILLER_102_896 VPWR VGND sg13g2_decap_8
XFILLER_87_574 VPWR VGND sg13g2_decap_8
XFILLER_75_714 VPWR VGND sg13g2_decap_8
XFILLER_47_427 VPWR VGND sg13g2_decap_8
XFILLER_19_42 VPWR VGND sg13g2_decap_8
XFILLER_74_246 VPWR VGND sg13g2_decap_8
XFILLER_28_630 VPWR VGND sg13g2_decap_8
XFILLER_90_739 VPWR VGND sg13g2_decap_8
XFILLER_27_151 VPWR VGND sg13g2_decap_8
XFILLER_71_942 VPWR VGND sg13g2_decap_8
XFILLER_43_644 VPWR VGND sg13g2_decap_8
XFILLER_16_847 VPWR VGND sg13g2_decap_8
XFILLER_70_441 VPWR VGND sg13g2_decap_8
XFILLER_15_368 VPWR VGND sg13g2_decap_8
XFILLER_35_63 VPWR VGND sg13g2_decap_8
XFILLER_37_1019 VPWR VGND sg13g2_decap_8
XFILLER_42_165 VPWR VGND sg13g2_decap_8
XFILLER_7_501 VPWR VGND sg13g2_decap_8
XFILLER_11_574 VPWR VGND sg13g2_decap_8
XFILLER_51_95 VPWR VGND sg13g2_decap_8
XFILLER_100_1022 VPWR VGND sg13g2_decap_8
XFILLER_7_578 VPWR VGND sg13g2_decap_8
XFILLER_83_1028 VPWR VGND sg13g2_fill_1
XFILLER_3_784 VPWR VGND sg13g2_decap_8
XFILLER_78_552 VPWR VGND sg13g2_decap_8
XFILLER_39_928 VPWR VGND sg13g2_decap_8
XFILLER_38_427 VPWR VGND sg13g2_decap_8
XFILLER_93_544 VPWR VGND sg13g2_decap_8
XFILLER_76_81 VPWR VGND sg13g2_decap_8
XFILLER_66_769 VPWR VGND sg13g2_decap_8
XFILLER_65_224 VPWR VGND sg13g2_decap_8
XFILLER_19_630 VPWR VGND sg13g2_decap_8
XFILLER_20_1012 VPWR VGND sg13g2_decap_8
XFILLER_81_739 VPWR VGND sg13g2_decap_8
XFILLER_47_994 VPWR VGND sg13g2_decap_8
XFILLER_18_140 VPWR VGND sg13g2_decap_8
XFILLER_80_238 VPWR VGND sg13g2_decap_8
XFILLER_62_931 VPWR VGND sg13g2_decap_8
XFILLER_61_452 VPWR VGND sg13g2_decap_8
XFILLER_33_154 VPWR VGND sg13g2_decap_8
XFILLER_34_655 VPWR VGND sg13g2_decap_8
XFILLER_92_91 VPWR VGND sg13g2_decap_8
XFILLER_30_861 VPWR VGND sg13g2_decap_8
XFILLER_103_616 VPWR VGND sg13g2_decap_8
XFILLER_88_305 VPWR VGND sg13g2_decap_8
XFILLER_102_126 VPWR VGND sg13g2_decap_8
XFILLER_97_861 VPWR VGND sg13g2_decap_8
XFILLER_96_371 VPWR VGND sg13g2_decap_8
XFILLER_84_511 VPWR VGND sg13g2_decap_8
XFILLER_69_596 VPWR VGND sg13g2_decap_8
XFILLER_57_714 VPWR VGND sg13g2_decap_8
XFILLER_56_18 VPWR VGND sg13g2_decap_8
XFILLER_5_1028 VPWR VGND sg13g2_fill_1
XFILLER_56_235 VPWR VGND sg13g2_decap_8
XFILLER_29_438 VPWR VGND sg13g2_decap_8
XFILLER_84_588 VPWR VGND sg13g2_decap_8
XFILLER_72_728 VPWR VGND sg13g2_decap_8
XFILLER_71_249 VPWR VGND sg13g2_decap_8
XFILLER_65_791 VPWR VGND sg13g2_decap_8
XFILLER_53_931 VPWR VGND sg13g2_decap_8
XFILLER_25_644 VPWR VGND sg13g2_decap_8
XFILLER_38_994 VPWR VGND sg13g2_decap_8
XFILLER_72_28 VPWR VGND sg13g2_decap_8
XFILLER_52_441 VPWR VGND sg13g2_decap_8
XFILLER_12_305 VPWR VGND sg13g2_decap_8
XFILLER_24_165 VPWR VGND sg13g2_decap_8
XFILLER_40_658 VPWR VGND sg13g2_decap_8
XFILLER_21_861 VPWR VGND sg13g2_decap_8
XFILLER_20_382 VPWR VGND sg13g2_decap_8
XFILLER_21_21 VPWR VGND sg13g2_decap_8
XFILLER_4_504 VPWR VGND sg13g2_decap_8
XFILLER_97_14 VPWR VGND sg13g2_decap_8
XFILLER_21_98 VPWR VGND sg13g2_decap_8
XFILLER_106_476 VPWR VGND sg13g2_decap_8
XFILLER_79_305 VPWR VGND sg13g2_decap_8
XFILLER_0_721 VPWR VGND sg13g2_decap_8
XFILLER_95_809 VPWR VGND sg13g2_decap_8
XFILLER_94_308 VPWR VGND sg13g2_decap_8
XFILLER_88_872 VPWR VGND sg13g2_decap_8
XFILLER_43_1001 VPWR VGND sg13g2_decap_8
XFILLER_87_371 VPWR VGND sg13g2_decap_8
XFILLER_75_511 VPWR VGND sg13g2_decap_8
XFILLER_48_714 VPWR VGND sg13g2_decap_8
XFILLER_0_798 VPWR VGND sg13g2_decap_8
XFILLER_102_693 VPWR VGND sg13g2_decap_8
XFILLER_47_224 VPWR VGND sg13g2_decap_8
XFILLER_75_588 VPWR VGND sg13g2_decap_8
XFILLER_63_728 VPWR VGND sg13g2_decap_8
XFILLER_90_536 VPWR VGND sg13g2_decap_8
XFILLER_62_238 VPWR VGND sg13g2_decap_8
XFILLER_46_95 VPWR VGND sg13g2_decap_8
XFILLER_44_942 VPWR VGND sg13g2_decap_8
XFILLER_43_441 VPWR VGND sg13g2_decap_8
XFILLER_16_644 VPWR VGND sg13g2_decap_8
XFILLER_15_165 VPWR VGND sg13g2_decap_8
XFILLER_31_658 VPWR VGND sg13g2_decap_8
XFILLER_62_83 VPWR VGND sg13g2_decap_8
XFILLER_12_872 VPWR VGND sg13g2_decap_8
XFILLER_30_168 VPWR VGND sg13g2_decap_8
XFILLER_8_854 VPWR VGND sg13g2_decap_8
XFILLER_11_371 VPWR VGND sg13g2_decap_8
XFILLER_7_375 VPWR VGND sg13g2_decap_8
XFILLER_7_67 VPWR VGND sg13g2_decap_8
XFILLER_3_581 VPWR VGND sg13g2_decap_8
XFILLER_98_669 VPWR VGND sg13g2_decap_8
XFILLER_86_809 VPWR VGND sg13g2_decap_8
XFILLER_85_308 VPWR VGND sg13g2_decap_8
XFILLER_97_168 VPWR VGND sg13g2_decap_8
XFILLER_87_91 VPWR VGND sg13g2_decap_8
XFILLER_79_872 VPWR VGND sg13g2_decap_8
XFILLER_39_725 VPWR VGND sg13g2_decap_8
XFILLER_38_224 VPWR VGND sg13g2_decap_8
XFILLER_94_875 VPWR VGND sg13g2_decap_8
XFILLER_93_341 VPWR VGND sg13g2_decap_8
XFILLER_66_566 VPWR VGND sg13g2_decap_8
XFILLER_81_536 VPWR VGND sg13g2_decap_8
XFILLER_54_739 VPWR VGND sg13g2_decap_8
XFILLER_53_238 VPWR VGND sg13g2_decap_8
XFILLER_47_791 VPWR VGND sg13g2_decap_8
XFILLER_35_931 VPWR VGND sg13g2_decap_8
XFILLER_34_452 VPWR VGND sg13g2_decap_8
XFILLER_50_945 VPWR VGND sg13g2_decap_8
XFILLER_10_809 VPWR VGND sg13g2_decap_8
XFILLER_22_669 VPWR VGND sg13g2_decap_8
XFILLER_21_168 VPWR VGND sg13g2_decap_8
XFILLER_104_903 VPWR VGND sg13g2_decap_8
XFILLER_103_413 VPWR VGND sg13g2_decap_8
XFILLER_88_102 VPWR VGND sg13g2_decap_8
XFILLER_1_518 VPWR VGND sg13g2_decap_8
XFILLER_89_658 VPWR VGND sg13g2_decap_8
XFILLER_88_179 VPWR VGND sg13g2_decap_8
XFILLER_76_319 VPWR VGND sg13g2_decap_8
XFILLER_57_511 VPWR VGND sg13g2_decap_8
XFILLER_69_393 VPWR VGND sg13g2_decap_8
XFILLER_29_235 VPWR VGND sg13g2_decap_8
XFILLER_85_875 VPWR VGND sg13g2_decap_8
XFILLER_57_588 VPWR VGND sg13g2_decap_8
XFILLER_45_728 VPWR VGND sg13g2_decap_8
XFILLER_84_385 VPWR VGND sg13g2_decap_8
XFILLER_72_525 VPWR VGND sg13g2_decap_8
XFILLER_26_931 VPWR VGND sg13g2_decap_8
XFILLER_38_791 VPWR VGND sg13g2_decap_8
XFILLER_44_249 VPWR VGND sg13g2_decap_8
XFILLER_16_21 VPWR VGND sg13g2_decap_8
XFILLER_25_441 VPWR VGND sg13g2_decap_8
XFILLER_73_1005 VPWR VGND sg13g2_decap_8
XFILLER_12_102 VPWR VGND sg13g2_decap_8
XFILLER_41_945 VPWR VGND sg13g2_decap_8
XFILLER_13_658 VPWR VGND sg13g2_decap_8
XFILLER_16_98 VPWR VGND sg13g2_decap_8
XFILLER_40_455 VPWR VGND sg13g2_decap_8
XFILLER_12_179 VPWR VGND sg13g2_decap_8
XFILLER_32_53 VPWR VGND sg13g2_decap_8
XFILLER_5_802 VPWR VGND sg13g2_decap_8
XFILLER_4_301 VPWR VGND sg13g2_decap_8
XFILLER_106_0 VPWR VGND sg13g2_decap_8
XFILLER_5_879 VPWR VGND sg13g2_decap_8
XFILLER_106_273 VPWR VGND sg13g2_decap_8
XFILLER_79_102 VPWR VGND sg13g2_decap_8
XFILLER_4_378 VPWR VGND sg13g2_decap_8
XFILLER_95_606 VPWR VGND sg13g2_decap_8
XFILLER_103_980 VPWR VGND sg13g2_decap_8
XFILLER_94_105 VPWR VGND sg13g2_decap_8
XFILLER_79_179 VPWR VGND sg13g2_decap_8
XFILLER_67_308 VPWR VGND sg13g2_decap_8
XFILLER_48_511 VPWR VGND sg13g2_decap_8
XFILLER_102_490 VPWR VGND sg13g2_decap_8
XFILLER_0_595 VPWR VGND sg13g2_decap_8
XFILLER_91_812 VPWR VGND sg13g2_decap_8
XFILLER_76_886 VPWR VGND sg13g2_decap_8
XFILLER_48_588 VPWR VGND sg13g2_decap_8
XFILLER_36_728 VPWR VGND sg13g2_decap_8
XFILLER_75_385 VPWR VGND sg13g2_decap_8
XFILLER_63_525 VPWR VGND sg13g2_decap_8
XFILLER_35_238 VPWR VGND sg13g2_decap_8
XFILLER_91_889 VPWR VGND sg13g2_decap_8
XFILLER_90_333 VPWR VGND sg13g2_decap_8
XFILLER_16_441 VPWR VGND sg13g2_decap_8
XFILLER_17_942 VPWR VGND sg13g2_decap_8
XFILLER_32_956 VPWR VGND sg13g2_decap_8
XFILLER_31_455 VPWR VGND sg13g2_decap_8
XFILLER_89_1001 VPWR VGND sg13g2_decap_8
XFILLER_78_4 VPWR VGND sg13g2_decap_8
XFILLER_8_651 VPWR VGND sg13g2_decap_8
XFILLER_7_172 VPWR VGND sg13g2_decap_8
XFILLER_99_945 VPWR VGND sg13g2_decap_8
XFILLER_98_466 VPWR VGND sg13g2_decap_8
XFILLER_86_606 VPWR VGND sg13g2_decap_8
XFILLER_101_917 VPWR VGND sg13g2_decap_8
XFILLER_85_105 VPWR VGND sg13g2_decap_8
XFILLER_58_308 VPWR VGND sg13g2_decap_8
XFILLER_21_0 VPWR VGND sg13g2_decap_8
XFILLER_100_427 VPWR VGND sg13g2_decap_8
XFILLER_39_522 VPWR VGND sg13g2_decap_8
XFILLER_94_672 VPWR VGND sg13g2_decap_8
XFILLER_82_812 VPWR VGND sg13g2_decap_8
XFILLER_67_875 VPWR VGND sg13g2_decap_8
XFILLER_66_363 VPWR VGND sg13g2_decap_8
XFILLER_54_536 VPWR VGND sg13g2_decap_8
XFILLER_27_739 VPWR VGND sg13g2_decap_8
XFILLER_39_599 VPWR VGND sg13g2_decap_8
XFILLER_82_889 VPWR VGND sg13g2_decap_8
XFILLER_81_333 VPWR VGND sg13g2_decap_8
XFILLER_26_238 VPWR VGND sg13g2_decap_8
XFILLER_50_742 VPWR VGND sg13g2_decap_8
XFILLER_23_945 VPWR VGND sg13g2_decap_8
XFILLER_10_606 VPWR VGND sg13g2_decap_8
XFILLER_22_466 VPWR VGND sg13g2_decap_8
XFILLER_33_1022 VPWR VGND sg13g2_decap_8
XFILLER_5_109 VPWR VGND sg13g2_decap_8
XFILLER_2_816 VPWR VGND sg13g2_decap_8
XFILLER_104_700 VPWR VGND sg13g2_decap_8
XFILLER_1_315 VPWR VGND sg13g2_decap_8
XFILLER_103_210 VPWR VGND sg13g2_decap_8
XFILLER_89_455 VPWR VGND sg13g2_decap_8
XFILLER_104_777 VPWR VGND sg13g2_decap_8
XFILLER_76_116 VPWR VGND sg13g2_decap_8
XFILLER_49_319 VPWR VGND sg13g2_decap_8
XFILLER_103_287 VPWR VGND sg13g2_decap_8
XFILLER_92_609 VPWR VGND sg13g2_decap_8
XFILLER_85_672 VPWR VGND sg13g2_decap_8
XFILLER_69_190 VPWR VGND sg13g2_decap_8
XFILLER_58_875 VPWR VGND sg13g2_decap_8
XFILLER_40_1015 VPWR VGND sg13g2_decap_8
XFILLER_100_994 VPWR VGND sg13g2_decap_8
XFILLER_91_119 VPWR VGND sg13g2_decap_8
XFILLER_84_182 VPWR VGND sg13g2_decap_8
XFILLER_73_823 VPWR VGND sg13g2_decap_8
XFILLER_72_322 VPWR VGND sg13g2_decap_8
XFILLER_57_385 VPWR VGND sg13g2_decap_8
XFILLER_45_525 VPWR VGND sg13g2_decap_8
XFILLER_18_728 VPWR VGND sg13g2_decap_8
XFILLER_27_53 VPWR VGND sg13g2_decap_8
XFILLER_17_249 VPWR VGND sg13g2_decap_8
XFILLER_72_399 VPWR VGND sg13g2_decap_8
XFILLER_41_742 VPWR VGND sg13g2_decap_8
XFILLER_14_945 VPWR VGND sg13g2_decap_8
XFILLER_43_63 VPWR VGND sg13g2_decap_8
XFILLER_13_455 VPWR VGND sg13g2_decap_8
XFILLER_40_252 VPWR VGND sg13g2_decap_8
XFILLER_9_448 VPWR VGND sg13g2_decap_8
XFILLER_5_676 VPWR VGND sg13g2_decap_8
XFILLER_4_175 VPWR VGND sg13g2_decap_8
XFILLER_4_35 VPWR VGND sg13g2_decap_8
XFILLER_95_403 VPWR VGND sg13g2_decap_8
XFILLER_68_628 VPWR VGND sg13g2_decap_8
XFILLER_67_105 VPWR VGND sg13g2_decap_8
XFILLER_96_959 VPWR VGND sg13g2_decap_8
XFILLER_68_82 VPWR VGND sg13g2_decap_8
XFILLER_1_882 VPWR VGND sg13g2_decap_8
XFILLER_49_886 VPWR VGND sg13g2_decap_8
XFILLER_0_392 VPWR VGND sg13g2_decap_8
XFILLER_82_119 VPWR VGND sg13g2_decap_8
XFILLER_76_683 VPWR VGND sg13g2_decap_8
XFILLER_64_823 VPWR VGND sg13g2_decap_8
XFILLER_63_322 VPWR VGND sg13g2_decap_8
XFILLER_48_385 VPWR VGND sg13g2_decap_8
XFILLER_36_525 VPWR VGND sg13g2_decap_8
XFILLER_90_130 VPWR VGND sg13g2_decap_8
XFILLER_84_70 VPWR VGND sg13g2_decap_8
XFILLER_75_182 VPWR VGND sg13g2_decap_8
XFILLER_91_686 VPWR VGND sg13g2_decap_8
XFILLER_63_399 VPWR VGND sg13g2_decap_8
XFILLER_17_1028 VPWR VGND sg13g2_fill_1
XFILLER_31_252 VPWR VGND sg13g2_decap_8
XFILLER_32_753 VPWR VGND sg13g2_decap_8
XFILLER_69_0 VPWR VGND sg13g2_decap_8
XFILLER_99_742 VPWR VGND sg13g2_decap_8
XFILLER_63_1015 VPWR VGND sg13g2_decap_8
XFILLER_101_714 VPWR VGND sg13g2_decap_8
XFILLER_98_263 VPWR VGND sg13g2_decap_8
XFILLER_86_403 VPWR VGND sg13g2_decap_8
XFILLER_59_628 VPWR VGND sg13g2_decap_8
XFILLER_58_105 VPWR VGND sg13g2_decap_8
XFILLER_100_224 VPWR VGND sg13g2_decap_8
XFILLER_87_959 VPWR VGND sg13g2_decap_8
XFILLER_104_14 VPWR VGND sg13g2_decap_8
XFILLER_95_970 VPWR VGND sg13g2_decap_8
XFILLER_67_672 VPWR VGND sg13g2_decap_8
XFILLER_66_160 VPWR VGND sg13g2_decap_8
XFILLER_64_18 VPWR VGND sg13g2_decap_8
XFILLER_55_812 VPWR VGND sg13g2_decap_8
XFILLER_27_536 VPWR VGND sg13g2_decap_8
XFILLER_81_130 VPWR VGND sg13g2_decap_8
XFILLER_54_333 VPWR VGND sg13g2_decap_8
XFILLER_39_396 VPWR VGND sg13g2_decap_8
XFILLER_82_686 VPWR VGND sg13g2_decap_8
XFILLER_70_826 VPWR VGND sg13g2_decap_8
XFILLER_55_889 VPWR VGND sg13g2_decap_8
XFILLER_23_742 VPWR VGND sg13g2_decap_8
XFILLER_80_28 VPWR VGND sg13g2_decap_8
XFILLER_70_1008 VPWR VGND sg13g2_decap_8
XFILLER_10_403 VPWR VGND sg13g2_decap_8
XFILLER_11_959 VPWR VGND sg13g2_decap_8
XFILLER_22_263 VPWR VGND sg13g2_decap_8
XFILLER_13_77 VPWR VGND sg13g2_decap_8
XFILLER_2_613 VPWR VGND sg13g2_decap_8
XFILLER_1_112 VPWR VGND sg13g2_decap_8
XFILLER_104_574 VPWR VGND sg13g2_decap_8
XFILLER_89_252 VPWR VGND sg13g2_decap_8
XFILLER_78_937 VPWR VGND sg13g2_decap_8
XFILLER_49_116 VPWR VGND sg13g2_decap_8
XFILLER_1_189 VPWR VGND sg13g2_decap_8
XFILLER_93_929 VPWR VGND sg13g2_decap_8
XFILLER_92_406 VPWR VGND sg13g2_decap_8
XFILLER_86_970 VPWR VGND sg13g2_decap_8
XFILLER_77_469 VPWR VGND sg13g2_decap_8
XFILLER_65_609 VPWR VGND sg13g2_decap_8
XFILLER_38_63 VPWR VGND sg13g2_decap_8
XFILLER_73_620 VPWR VGND sg13g2_decap_8
XFILLER_58_672 VPWR VGND sg13g2_decap_8
XFILLER_46_823 VPWR VGND sg13g2_decap_8
XFILLER_18_525 VPWR VGND sg13g2_decap_8
XFILLER_100_791 VPWR VGND sg13g2_decap_8
XFILLER_57_182 VPWR VGND sg13g2_decap_8
XFILLER_45_322 VPWR VGND sg13g2_decap_8
XFILLER_73_697 VPWR VGND sg13g2_decap_8
XFILLER_61_837 VPWR VGND sg13g2_decap_8
XFILLER_72_196 VPWR VGND sg13g2_decap_8
XFILLER_60_347 VPWR VGND sg13g2_decap_8
XFILLER_45_399 VPWR VGND sg13g2_decap_8
XFILLER_14_742 VPWR VGND sg13g2_decap_8
XFILLER_33_539 VPWR VGND sg13g2_decap_8
XFILLER_54_95 VPWR VGND sg13g2_decap_8
XFILLER_13_252 VPWR VGND sg13g2_decap_8
XFILLER_9_245 VPWR VGND sg13g2_decap_8
XFILLER_10_970 VPWR VGND sg13g2_decap_8
XFILLER_86_1026 VPWR VGND sg13g2_fill_2
XFILLER_62_7 VPWR VGND sg13g2_decap_8
XFILLER_6_952 VPWR VGND sg13g2_decap_8
XFILLER_5_473 VPWR VGND sg13g2_decap_8
XFILLER_79_81 VPWR VGND sg13g2_decap_8
XFILLER_69_904 VPWR VGND sg13g2_decap_8
XFILLER_96_756 VPWR VGND sg13g2_decap_8
XFILLER_95_200 VPWR VGND sg13g2_decap_8
XFILLER_68_425 VPWR VGND sg13g2_decap_8
XFILLER_95_277 VPWR VGND sg13g2_decap_8
XFILLER_83_417 VPWR VGND sg13g2_decap_8
XFILLER_76_480 VPWR VGND sg13g2_decap_8
XFILLER_64_620 VPWR VGND sg13g2_decap_8
XFILLER_55_119 VPWR VGND sg13g2_decap_8
XFILLER_49_683 VPWR VGND sg13g2_decap_8
XFILLER_37_823 VPWR VGND sg13g2_decap_8
XFILLER_48_182 VPWR VGND sg13g2_decap_8
XFILLER_36_322 VPWR VGND sg13g2_decap_8
XFILLER_92_973 VPWR VGND sg13g2_decap_8
XFILLER_52_826 VPWR VGND sg13g2_decap_8
XFILLER_91_483 VPWR VGND sg13g2_decap_8
XFILLER_64_697 VPWR VGND sg13g2_decap_8
XFILLER_63_196 VPWR VGND sg13g2_decap_8
XFILLER_51_347 VPWR VGND sg13g2_decap_8
XFILLER_36_399 VPWR VGND sg13g2_decap_8
XFILLER_32_550 VPWR VGND sg13g2_decap_8
XFILLER_20_767 VPWR VGND sg13g2_decap_8
XFILLER_59_18 VPWR VGND sg13g2_decap_8
XFILLER_8_1015 VPWR VGND sg13g2_decap_8
XFILLER_101_511 VPWR VGND sg13g2_decap_8
XFILLER_87_756 VPWR VGND sg13g2_decap_8
XFILLER_86_200 VPWR VGND sg13g2_decap_8
XFILLER_59_425 VPWR VGND sg13g2_decap_8
XFILLER_75_28 VPWR VGND sg13g2_decap_8
XFILLER_47_609 VPWR VGND sg13g2_decap_8
XFILLER_101_588 VPWR VGND sg13g2_decap_8
XFILLER_86_277 VPWR VGND sg13g2_decap_8
XFILLER_74_428 VPWR VGND sg13g2_decap_8
XFILLER_68_992 VPWR VGND sg13g2_decap_8
XFILLER_28_812 VPWR VGND sg13g2_decap_8
XFILLER_54_130 VPWR VGND sg13g2_decap_8
XFILLER_27_333 VPWR VGND sg13g2_decap_8
XFILLER_39_193 VPWR VGND sg13g2_decap_8
XFILLER_83_984 VPWR VGND sg13g2_decap_8
XFILLER_55_686 VPWR VGND sg13g2_decap_8
XFILLER_43_826 VPWR VGND sg13g2_decap_8
XFILLER_28_889 VPWR VGND sg13g2_decap_8
XFILLER_91_49 VPWR VGND sg13g2_decap_8
XFILLER_82_483 VPWR VGND sg13g2_decap_8
XFILLER_70_623 VPWR VGND sg13g2_decap_8
XFILLER_42_347 VPWR VGND sg13g2_decap_8
XFILLER_24_32 VPWR VGND sg13g2_decap_8
XFILLER_10_200 VPWR VGND sg13g2_decap_8
XFILLER_11_756 VPWR VGND sg13g2_decap_8
XFILLER_10_277 VPWR VGND sg13g2_decap_8
XFILLER_6_259 VPWR VGND sg13g2_decap_8
XFILLER_40_42 VPWR VGND sg13g2_decap_8
XFILLER_2_410 VPWR VGND sg13g2_decap_8
XFILLER_105_861 VPWR VGND sg13g2_decap_8
XFILLER_3_966 VPWR VGND sg13g2_decap_8
XFILLER_104_371 VPWR VGND sg13g2_decap_8
XFILLER_78_734 VPWR VGND sg13g2_decap_8
XFILLER_2_487 VPWR VGND sg13g2_decap_8
XFILLER_49_95 VPWR VGND sg13g2_decap_8
XFILLER_1_14 VPWR VGND sg13g2_decap_8
XFILLER_38_609 VPWR VGND sg13g2_decap_8
XFILLER_93_726 VPWR VGND sg13g2_decap_8
XFILLER_92_203 VPWR VGND sg13g2_decap_8
XFILLER_77_266 VPWR VGND sg13g2_decap_8
XFILLER_65_406 VPWR VGND sg13g2_decap_8
XFILLER_59_992 VPWR VGND sg13g2_decap_8
XFILLER_19_812 VPWR VGND sg13g2_decap_8
XFILLER_46_620 VPWR VGND sg13g2_decap_8
XFILLER_18_322 VPWR VGND sg13g2_decap_8
XFILLER_74_995 VPWR VGND sg13g2_decap_8
XFILLER_19_889 VPWR VGND sg13g2_decap_8
XFILLER_73_494 VPWR VGND sg13g2_decap_8
XFILLER_61_634 VPWR VGND sg13g2_decap_8
XFILLER_46_697 VPWR VGND sg13g2_decap_8
XFILLER_45_196 VPWR VGND sg13g2_decap_8
XFILLER_18_399 VPWR VGND sg13g2_decap_8
XFILLER_33_336 VPWR VGND sg13g2_decap_8
XFILLER_34_837 VPWR VGND sg13g2_decap_8
XFILLER_60_144 VPWR VGND sg13g2_decap_8
XFILLER_81_60 VPWR VGND sg13g2_decap_8
XFILLER_5_270 VPWR VGND sg13g2_decap_8
XFILLER_102_308 VPWR VGND sg13g2_decap_8
XFILLER_69_701 VPWR VGND sg13g2_decap_8
XFILLER_68_222 VPWR VGND sg13g2_decap_8
XFILLER_96_553 VPWR VGND sg13g2_decap_8
XFILLER_69_778 VPWR VGND sg13g2_decap_8
XFILLER_83_214 VPWR VGND sg13g2_decap_8
Xinput2 ui_in[1] net2 VPWR VGND sg13g2_buf_1
XFILLER_56_417 VPWR VGND sg13g2_decap_8
XFILLER_28_119 VPWR VGND sg13g2_decap_8
XFILLER_68_299 VPWR VGND sg13g2_decap_8
XFILLER_49_480 VPWR VGND sg13g2_decap_8
XFILLER_37_620 VPWR VGND sg13g2_decap_8
XFILLER_92_770 VPWR VGND sg13g2_decap_8
XFILLER_80_910 VPWR VGND sg13g2_decap_8
XFILLER_65_973 VPWR VGND sg13g2_decap_8
XFILLER_25_826 VPWR VGND sg13g2_decap_8
XFILLER_91_280 VPWR VGND sg13g2_decap_8
XFILLER_64_494 VPWR VGND sg13g2_decap_8
XFILLER_52_623 VPWR VGND sg13g2_decap_8
XFILLER_36_196 VPWR VGND sg13g2_decap_8
XFILLER_37_697 VPWR VGND sg13g2_decap_8
XFILLER_80_987 VPWR VGND sg13g2_decap_8
XFILLER_51_144 VPWR VGND sg13g2_decap_8
XFILLER_24_347 VPWR VGND sg13g2_decap_8
XFILLER_20_564 VPWR VGND sg13g2_decap_8
XFILLER_106_658 VPWR VGND sg13g2_decap_8
XFILLER_105_168 VPWR VGND sg13g2_decap_8
XFILLER_10_67 VPWR VGND sg13g2_decap_8
XFILLER_0_903 VPWR VGND sg13g2_decap_8
XFILLER_59_222 VPWR VGND sg13g2_decap_8
XFILLER_87_553 VPWR VGND sg13g2_decap_8
XFILLER_19_21 VPWR VGND sg13g2_decap_8
XFILLER_102_875 VPWR VGND sg13g2_decap_8
XFILLER_47_406 VPWR VGND sg13g2_decap_8
XFILLER_19_119 VPWR VGND sg13g2_decap_8
XFILLER_101_385 VPWR VGND sg13g2_decap_8
XFILLER_74_225 VPWR VGND sg13g2_decap_8
XFILLER_59_299 VPWR VGND sg13g2_decap_8
XFILLER_19_98 VPWR VGND sg13g2_decap_8
XFILLER_90_718 VPWR VGND sg13g2_decap_8
XFILLER_56_984 VPWR VGND sg13g2_decap_8
XFILLER_16_826 VPWR VGND sg13g2_decap_8
XFILLER_27_130 VPWR VGND sg13g2_decap_8
XFILLER_83_781 VPWR VGND sg13g2_decap_8
XFILLER_82_280 VPWR VGND sg13g2_decap_8
XFILLER_71_921 VPWR VGND sg13g2_decap_8
XFILLER_70_420 VPWR VGND sg13g2_decap_8
XFILLER_55_483 VPWR VGND sg13g2_decap_8
XFILLER_43_623 VPWR VGND sg13g2_decap_8
XFILLER_28_686 VPWR VGND sg13g2_decap_8
XFILLER_35_42 VPWR VGND sg13g2_decap_8
XFILLER_42_144 VPWR VGND sg13g2_decap_8
XFILLER_15_347 VPWR VGND sg13g2_decap_8
XFILLER_71_998 VPWR VGND sg13g2_decap_8
XFILLER_70_497 VPWR VGND sg13g2_decap_8
XFILLER_11_553 VPWR VGND sg13g2_decap_8
XFILLER_100_1001 VPWR VGND sg13g2_decap_8
XFILLER_51_74 VPWR VGND sg13g2_decap_8
XFILLER_7_557 VPWR VGND sg13g2_decap_8
XFILLER_3_763 VPWR VGND sg13g2_decap_8
XFILLER_78_531 VPWR VGND sg13g2_decap_8
XFILLER_2_284 VPWR VGND sg13g2_decap_8
XFILLER_25_7 VPWR VGND sg13g2_decap_8
XFILLER_39_907 VPWR VGND sg13g2_decap_8
XFILLER_93_523 VPWR VGND sg13g2_decap_8
XFILLER_76_60 VPWR VGND sg13g2_decap_8
XFILLER_65_203 VPWR VGND sg13g2_decap_8
XFILLER_38_406 VPWR VGND sg13g2_decap_8
XFILLER_66_748 VPWR VGND sg13g2_decap_8
XFILLER_81_718 VPWR VGND sg13g2_decap_8
XFILLER_62_910 VPWR VGND sg13g2_decap_8
XFILLER_47_973 VPWR VGND sg13g2_decap_8
XFILLER_80_217 VPWR VGND sg13g2_decap_8
XFILLER_74_792 VPWR VGND sg13g2_decap_8
XFILLER_46_494 VPWR VGND sg13g2_decap_8
XFILLER_19_686 VPWR VGND sg13g2_decap_8
XFILLER_34_634 VPWR VGND sg13g2_decap_8
XFILLER_92_70 VPWR VGND sg13g2_decap_8
XFILLER_73_291 VPWR VGND sg13g2_decap_8
XFILLER_62_987 VPWR VGND sg13g2_decap_8
XFILLER_61_431 VPWR VGND sg13g2_decap_8
XFILLER_18_196 VPWR VGND sg13g2_decap_8
XFILLER_33_133 VPWR VGND sg13g2_decap_8
XFILLER_30_840 VPWR VGND sg13g2_decap_8
XFILLER_102_105 VPWR VGND sg13g2_decap_8
XFILLER_97_840 VPWR VGND sg13g2_decap_8
XFILLER_96_350 VPWR VGND sg13g2_decap_8
XFILLER_69_575 VPWR VGND sg13g2_decap_8
XFILLER_29_417 VPWR VGND sg13g2_decap_8
XFILLER_56_214 VPWR VGND sg13g2_decap_8
XFILLER_84_567 VPWR VGND sg13g2_decap_8
XFILLER_72_707 VPWR VGND sg13g2_decap_8
XFILLER_65_770 VPWR VGND sg13g2_decap_8
XFILLER_53_910 VPWR VGND sg13g2_decap_8
XFILLER_38_973 VPWR VGND sg13g2_decap_8
XFILLER_71_228 VPWR VGND sg13g2_decap_8
XFILLER_52_420 VPWR VGND sg13g2_decap_8
XFILLER_25_623 VPWR VGND sg13g2_decap_8
XFILLER_37_494 VPWR VGND sg13g2_decap_8
XFILLER_64_291 VPWR VGND sg13g2_decap_8
XFILLER_24_144 VPWR VGND sg13g2_decap_8
XFILLER_80_784 VPWR VGND sg13g2_decap_8
XFILLER_53_987 VPWR VGND sg13g2_decap_8
XFILLER_52_497 VPWR VGND sg13g2_decap_8
XFILLER_21_840 VPWR VGND sg13g2_decap_8
XFILLER_40_637 VPWR VGND sg13g2_decap_8
XFILLER_20_361 VPWR VGND sg13g2_decap_8
XFILLER_21_77 VPWR VGND sg13g2_decap_8
XFILLER_106_455 VPWR VGND sg13g2_decap_8
XFILLER_0_700 VPWR VGND sg13g2_decap_8
XFILLER_88_851 VPWR VGND sg13g2_decap_8
XFILLER_102_672 VPWR VGND sg13g2_decap_8
XFILLER_87_350 VPWR VGND sg13g2_decap_8
XFILLER_47_203 VPWR VGND sg13g2_decap_8
XFILLER_0_777 VPWR VGND sg13g2_decap_8
XFILLER_101_182 VPWR VGND sg13g2_decap_8
XFILLER_90_515 VPWR VGND sg13g2_decap_8
XFILLER_75_567 VPWR VGND sg13g2_decap_8
XFILLER_63_707 VPWR VGND sg13g2_decap_8
XFILLER_29_984 VPWR VGND sg13g2_decap_8
XFILLER_62_217 VPWR VGND sg13g2_decap_8
XFILLER_56_781 VPWR VGND sg13g2_decap_8
XFILLER_46_74 VPWR VGND sg13g2_decap_8
XFILLER_44_921 VPWR VGND sg13g2_decap_8
XFILLER_16_623 VPWR VGND sg13g2_decap_8
XFILLER_28_483 VPWR VGND sg13g2_decap_8
XFILLER_55_280 VPWR VGND sg13g2_decap_8
XFILLER_43_420 VPWR VGND sg13g2_decap_8
XFILLER_15_144 VPWR VGND sg13g2_decap_8
XFILLER_102_91 VPWR VGND sg13g2_decap_8
XFILLER_71_795 VPWR VGND sg13g2_decap_8
XFILLER_44_998 VPWR VGND sg13g2_decap_8
XFILLER_70_294 VPWR VGND sg13g2_decap_8
XFILLER_62_62 VPWR VGND sg13g2_decap_8
XFILLER_43_497 VPWR VGND sg13g2_decap_8
XFILLER_31_637 VPWR VGND sg13g2_decap_8
XFILLER_11_350 VPWR VGND sg13g2_decap_8
XFILLER_12_851 VPWR VGND sg13g2_decap_8
XFILLER_30_147 VPWR VGND sg13g2_decap_8
XFILLER_8_833 VPWR VGND sg13g2_decap_8
XFILLER_7_46 VPWR VGND sg13g2_decap_8
XFILLER_7_354 VPWR VGND sg13g2_decap_8
XFILLER_98_648 VPWR VGND sg13g2_decap_8
XFILLER_3_560 VPWR VGND sg13g2_decap_8
XFILLER_100_609 VPWR VGND sg13g2_decap_8
XFILLER_97_147 VPWR VGND sg13g2_decap_8
XFILLER_87_70 VPWR VGND sg13g2_decap_8
XFILLER_79_851 VPWR VGND sg13g2_decap_8
XFILLER_38_203 VPWR VGND sg13g2_decap_8
XFILLER_39_704 VPWR VGND sg13g2_decap_8
XFILLER_94_854 VPWR VGND sg13g2_decap_8
XFILLER_93_320 VPWR VGND sg13g2_decap_8
XFILLER_66_545 VPWR VGND sg13g2_decap_8
XFILLER_54_718 VPWR VGND sg13g2_decap_8
XFILLER_93_397 VPWR VGND sg13g2_decap_8
XFILLER_81_515 VPWR VGND sg13g2_decap_8
XFILLER_59_1020 VPWR VGND sg13g2_decap_8
XFILLER_53_217 VPWR VGND sg13g2_decap_8
XFILLER_47_770 VPWR VGND sg13g2_decap_8
XFILLER_19_483 VPWR VGND sg13g2_decap_8
XFILLER_35_910 VPWR VGND sg13g2_decap_8
XFILLER_46_291 VPWR VGND sg13g2_decap_8
XFILLER_34_431 VPWR VGND sg13g2_decap_8
XFILLER_62_784 VPWR VGND sg13g2_decap_8
XFILLER_50_924 VPWR VGND sg13g2_decap_8
XFILLER_35_987 VPWR VGND sg13g2_decap_8
XFILLER_99_0 VPWR VGND sg13g2_decap_8
XFILLER_22_648 VPWR VGND sg13g2_decap_8
XFILLER_21_147 VPWR VGND sg13g2_decap_8
XFILLER_89_637 VPWR VGND sg13g2_decap_8
XFILLER_27_1019 VPWR VGND sg13g2_decap_8
XFILLER_104_959 VPWR VGND sg13g2_decap_8
XFILLER_88_158 VPWR VGND sg13g2_decap_8
XFILLER_103_469 VPWR VGND sg13g2_decap_8
XFILLER_69_372 VPWR VGND sg13g2_decap_8
XFILLER_85_854 VPWR VGND sg13g2_decap_8
XFILLER_29_214 VPWR VGND sg13g2_decap_8
XFILLER_84_364 VPWR VGND sg13g2_decap_8
XFILLER_72_504 VPWR VGND sg13g2_decap_8
XFILLER_57_567 VPWR VGND sg13g2_decap_8
XFILLER_45_707 VPWR VGND sg13g2_decap_8
XFILLER_83_39 VPWR VGND sg13g2_decap_8
XFILLER_44_228 VPWR VGND sg13g2_decap_8
XFILLER_26_910 VPWR VGND sg13g2_decap_8
XFILLER_38_770 VPWR VGND sg13g2_decap_8
XFILLER_25_420 VPWR VGND sg13g2_decap_8
XFILLER_37_291 VPWR VGND sg13g2_decap_8
XFILLER_73_1028 VPWR VGND sg13g2_fill_1
XFILLER_53_784 VPWR VGND sg13g2_decap_8
XFILLER_41_924 VPWR VGND sg13g2_decap_8
XFILLER_16_77 VPWR VGND sg13g2_decap_8
XFILLER_26_987 VPWR VGND sg13g2_decap_8
XFILLER_80_581 VPWR VGND sg13g2_decap_8
XFILLER_52_294 VPWR VGND sg13g2_decap_8
XFILLER_13_637 VPWR VGND sg13g2_decap_8
XFILLER_25_497 VPWR VGND sg13g2_decap_8
XFILLER_40_434 VPWR VGND sg13g2_decap_8
XFILLER_12_158 VPWR VGND sg13g2_decap_8
XFILLER_32_32 VPWR VGND sg13g2_decap_8
XFILLER_10_1012 VPWR VGND sg13g2_decap_8
XFILLER_5_858 VPWR VGND sg13g2_decap_8
XFILLER_4_357 VPWR VGND sg13g2_decap_8
XFILLER_106_252 VPWR VGND sg13g2_decap_8
XFILLER_79_158 VPWR VGND sg13g2_decap_8
XFILLER_0_574 VPWR VGND sg13g2_decap_8
XFILLER_76_865 VPWR VGND sg13g2_decap_8
XFILLER_75_364 VPWR VGND sg13g2_decap_8
XFILLER_63_504 VPWR VGND sg13g2_decap_8
XFILLER_57_84 VPWR VGND sg13g2_decap_8
XFILLER_48_567 VPWR VGND sg13g2_decap_8
XFILLER_36_707 VPWR VGND sg13g2_decap_8
XFILLER_90_312 VPWR VGND sg13g2_decap_8
XFILLER_17_921 VPWR VGND sg13g2_decap_8
XFILLER_29_781 VPWR VGND sg13g2_decap_8
XFILLER_35_217 VPWR VGND sg13g2_decap_8
XFILLER_91_868 VPWR VGND sg13g2_decap_8
XFILLER_16_420 VPWR VGND sg13g2_decap_8
XFILLER_28_280 VPWR VGND sg13g2_decap_8
XFILLER_90_389 VPWR VGND sg13g2_decap_8
XFILLER_17_998 VPWR VGND sg13g2_decap_8
XFILLER_92_7 VPWR VGND sg13g2_decap_8
XFILLER_71_592 VPWR VGND sg13g2_decap_8
XFILLER_44_795 VPWR VGND sg13g2_decap_8
XFILLER_43_294 VPWR VGND sg13g2_decap_8
XFILLER_16_497 VPWR VGND sg13g2_decap_8
XFILLER_31_434 VPWR VGND sg13g2_decap_8
XFILLER_32_935 VPWR VGND sg13g2_decap_8
XFILLER_8_630 VPWR VGND sg13g2_decap_8
XFILLER_7_151 VPWR VGND sg13g2_decap_8
XFILLER_99_924 VPWR VGND sg13g2_decap_8
XFILLER_98_445 VPWR VGND sg13g2_decap_8
XFILLER_100_406 VPWR VGND sg13g2_decap_8
XFILLER_39_501 VPWR VGND sg13g2_decap_8
XFILLER_94_651 VPWR VGND sg13g2_decap_8
XFILLER_67_854 VPWR VGND sg13g2_decap_8
XFILLER_66_342 VPWR VGND sg13g2_decap_8
XFILLER_14_0 VPWR VGND sg13g2_decap_8
XFILLER_27_718 VPWR VGND sg13g2_decap_8
XFILLER_39_578 VPWR VGND sg13g2_decap_8
XFILLER_81_312 VPWR VGND sg13g2_decap_8
XFILLER_54_515 VPWR VGND sg13g2_decap_8
XFILLER_26_217 VPWR VGND sg13g2_decap_8
XFILLER_93_194 VPWR VGND sg13g2_decap_8
XFILLER_82_868 VPWR VGND sg13g2_decap_8
XFILLER_19_280 VPWR VGND sg13g2_decap_8
XFILLER_81_389 VPWR VGND sg13g2_decap_8
XFILLER_23_924 VPWR VGND sg13g2_decap_8
XFILLER_35_784 VPWR VGND sg13g2_decap_8
XFILLER_62_581 VPWR VGND sg13g2_decap_8
XFILLER_50_721 VPWR VGND sg13g2_decap_8
XFILLER_22_445 VPWR VGND sg13g2_decap_8
XFILLER_33_1001 VPWR VGND sg13g2_decap_8
XFILLER_50_798 VPWR VGND sg13g2_decap_8
XFILLER_78_39 VPWR VGND sg13g2_decap_8
XFILLER_104_756 VPWR VGND sg13g2_decap_8
XFILLER_89_434 VPWR VGND sg13g2_decap_8
XFILLER_103_266 VPWR VGND sg13g2_decap_8
XFILLER_100_973 VPWR VGND sg13g2_decap_8
XFILLER_94_49 VPWR VGND sg13g2_decap_8
XFILLER_85_651 VPWR VGND sg13g2_decap_8
XFILLER_73_802 VPWR VGND sg13g2_decap_8
XFILLER_58_854 VPWR VGND sg13g2_decap_8
XFILLER_18_707 VPWR VGND sg13g2_decap_8
XFILLER_84_161 VPWR VGND sg13g2_decap_8
XFILLER_72_301 VPWR VGND sg13g2_decap_8
XFILLER_57_364 VPWR VGND sg13g2_decap_8
XFILLER_45_504 VPWR VGND sg13g2_decap_8
XFILLER_17_228 VPWR VGND sg13g2_decap_8
XFILLER_27_32 VPWR VGND sg13g2_decap_8
XFILLER_73_879 VPWR VGND sg13g2_decap_8
XFILLER_72_378 VPWR VGND sg13g2_decap_8
XFILLER_60_529 VPWR VGND sg13g2_decap_8
XFILLER_14_924 VPWR VGND sg13g2_decap_8
XFILLER_26_784 VPWR VGND sg13g2_decap_8
XFILLER_53_581 VPWR VGND sg13g2_decap_8
XFILLER_41_721 VPWR VGND sg13g2_decap_8
XFILLER_13_434 VPWR VGND sg13g2_decap_8
XFILLER_25_294 VPWR VGND sg13g2_decap_8
XFILLER_43_42 VPWR VGND sg13g2_decap_8
XFILLER_40_231 VPWR VGND sg13g2_decap_8
XFILLER_41_798 VPWR VGND sg13g2_decap_8
XFILLER_9_427 VPWR VGND sg13g2_decap_8
XFILLER_5_655 VPWR VGND sg13g2_decap_8
XFILLER_4_154 VPWR VGND sg13g2_decap_8
XFILLER_4_14 VPWR VGND sg13g2_decap_8
XFILLER_96_938 VPWR VGND sg13g2_decap_8
XFILLER_68_607 VPWR VGND sg13g2_decap_8
XFILLER_68_50 VPWR VGND sg13g2_fill_2
XFILLER_1_861 VPWR VGND sg13g2_decap_8
XFILLER_0_371 VPWR VGND sg13g2_decap_8
XFILLER_95_459 VPWR VGND sg13g2_decap_8
XFILLER_76_662 VPWR VGND sg13g2_decap_8
XFILLER_64_802 VPWR VGND sg13g2_decap_8
XFILLER_49_865 VPWR VGND sg13g2_decap_8
XFILLER_75_161 VPWR VGND sg13g2_decap_8
XFILLER_63_301 VPWR VGND sg13g2_decap_8
XFILLER_48_364 VPWR VGND sg13g2_decap_8
XFILLER_36_504 VPWR VGND sg13g2_decap_8
XFILLER_64_879 VPWR VGND sg13g2_decap_8
XFILLER_91_665 VPWR VGND sg13g2_decap_8
XFILLER_63_378 VPWR VGND sg13g2_decap_8
XFILLER_56_1012 VPWR VGND sg13g2_decap_8
XFILLER_51_529 VPWR VGND sg13g2_decap_8
XFILLER_90_186 VPWR VGND sg13g2_decap_8
XFILLER_44_592 VPWR VGND sg13g2_decap_8
XFILLER_17_795 VPWR VGND sg13g2_decap_8
XFILLER_32_732 VPWR VGND sg13g2_decap_8
XFILLER_90_4 VPWR VGND sg13g2_decap_8
XFILLER_16_294 VPWR VGND sg13g2_decap_8
XFILLER_31_231 VPWR VGND sg13g2_decap_8
XFILLER_20_949 VPWR VGND sg13g2_decap_8
XFILLER_9_994 VPWR VGND sg13g2_decap_8
XFILLER_99_721 VPWR VGND sg13g2_decap_8
XFILLER_99_798 VPWR VGND sg13g2_decap_8
XFILLER_98_242 VPWR VGND sg13g2_decap_8
XFILLER_87_938 VPWR VGND sg13g2_decap_8
XFILLER_59_607 VPWR VGND sg13g2_decap_8
XFILLER_100_203 VPWR VGND sg13g2_decap_8
XFILLER_86_459 VPWR VGND sg13g2_decap_8
XFILLER_67_651 VPWR VGND sg13g2_decap_8
XFILLER_73_109 VPWR VGND sg13g2_decap_8
XFILLER_54_312 VPWR VGND sg13g2_decap_8
XFILLER_27_515 VPWR VGND sg13g2_decap_8
XFILLER_39_375 VPWR VGND sg13g2_decap_8
XFILLER_55_868 VPWR VGND sg13g2_decap_8
XFILLER_82_665 VPWR VGND sg13g2_decap_8
XFILLER_70_805 VPWR VGND sg13g2_decap_8
XFILLER_42_529 VPWR VGND sg13g2_decap_8
XFILLER_81_186 VPWR VGND sg13g2_decap_8
XFILLER_54_389 VPWR VGND sg13g2_decap_8
XFILLER_23_721 VPWR VGND sg13g2_decap_8
XFILLER_35_581 VPWR VGND sg13g2_decap_8
XFILLER_22_242 VPWR VGND sg13g2_decap_8
XFILLER_50_595 VPWR VGND sg13g2_decap_8
XFILLER_11_938 VPWR VGND sg13g2_decap_8
XFILLER_23_798 VPWR VGND sg13g2_decap_8
XFILLER_10_459 VPWR VGND sg13g2_decap_8
XFILLER_13_56 VPWR VGND sg13g2_decap_8
XFILLER_89_49 VPWR VGND sg13g2_decap_8
XFILLER_89_231 VPWR VGND sg13g2_decap_8
XFILLER_104_553 VPWR VGND sg13g2_decap_8
XFILLER_78_916 VPWR VGND sg13g2_decap_8
XFILLER_2_669 VPWR VGND sg13g2_decap_8
XFILLER_77_448 VPWR VGND sg13g2_decap_8
XFILLER_1_168 VPWR VGND sg13g2_decap_8
XFILLER_93_908 VPWR VGND sg13g2_decap_8
XFILLER_58_651 VPWR VGND sg13g2_decap_8
XFILLER_46_802 VPWR VGND sg13g2_decap_8
XFILLER_38_42 VPWR VGND sg13g2_decap_8
XFILLER_100_770 VPWR VGND sg13g2_decap_8
XFILLER_79_1012 VPWR VGND sg13g2_decap_8
XFILLER_64_109 VPWR VGND sg13g2_decap_8
XFILLER_57_161 VPWR VGND sg13g2_decap_8
XFILLER_45_301 VPWR VGND sg13g2_decap_8
XFILLER_18_504 VPWR VGND sg13g2_decap_8
XFILLER_73_676 VPWR VGND sg13g2_decap_8
XFILLER_61_816 VPWR VGND sg13g2_decap_8
XFILLER_46_879 VPWR VGND sg13g2_decap_8
XFILLER_45_378 VPWR VGND sg13g2_decap_8
XFILLER_33_518 VPWR VGND sg13g2_decap_8
XFILLER_72_175 VPWR VGND sg13g2_decap_8
XFILLER_60_326 VPWR VGND sg13g2_decap_8
XFILLER_54_74 VPWR VGND sg13g2_decap_8
XFILLER_14_721 VPWR VGND sg13g2_decap_8
XFILLER_26_581 VPWR VGND sg13g2_decap_8
XFILLER_13_231 VPWR VGND sg13g2_decap_8
XFILLER_9_224 VPWR VGND sg13g2_decap_8
XFILLER_14_798 VPWR VGND sg13g2_decap_8
XFILLER_41_595 VPWR VGND sg13g2_decap_8
XFILLER_70_84 VPWR VGND sg13g2_decap_8
XFILLER_6_931 VPWR VGND sg13g2_decap_8
XFILLER_86_1005 VPWR VGND sg13g2_decap_8
XFILLER_55_7 VPWR VGND sg13g2_decap_8
XFILLER_5_452 VPWR VGND sg13g2_decap_8
XFILLER_68_404 VPWR VGND sg13g2_decap_8
XFILLER_96_735 VPWR VGND sg13g2_decap_8
XFILLER_95_256 VPWR VGND sg13g2_decap_8
XFILLER_23_1022 VPWR VGND sg13g2_decap_8
XFILLER_95_81 VPWR VGND sg13g2_decap_8
XFILLER_49_662 VPWR VGND sg13g2_decap_8
XFILLER_48_161 VPWR VGND sg13g2_decap_8
XFILLER_36_301 VPWR VGND sg13g2_decap_8
XFILLER_37_802 VPWR VGND sg13g2_decap_8
XFILLER_92_952 VPWR VGND sg13g2_decap_8
XFILLER_91_462 VPWR VGND sg13g2_decap_8
XFILLER_64_676 VPWR VGND sg13g2_decap_8
XFILLER_52_805 VPWR VGND sg13g2_decap_8
XFILLER_36_378 VPWR VGND sg13g2_decap_8
XFILLER_37_879 VPWR VGND sg13g2_decap_8
XFILLER_63_175 VPWR VGND sg13g2_decap_8
XFILLER_51_326 VPWR VGND sg13g2_decap_8
XFILLER_17_592 VPWR VGND sg13g2_decap_8
XFILLER_24_529 VPWR VGND sg13g2_decap_8
XFILLER_60_893 VPWR VGND sg13g2_decap_8
XFILLER_20_746 VPWR VGND sg13g2_decap_8
XFILLER_30_1015 VPWR VGND sg13g2_decap_8
XFILLER_9_791 VPWR VGND sg13g2_decap_8
XFILLER_59_404 VPWR VGND sg13g2_decap_8
XFILLER_99_595 VPWR VGND sg13g2_decap_8
XFILLER_87_735 VPWR VGND sg13g2_decap_8
XFILLER_101_567 VPWR VGND sg13g2_decap_8
XFILLER_86_256 VPWR VGND sg13g2_decap_8
XFILLER_74_407 VPWR VGND sg13g2_decap_8
XFILLER_68_971 VPWR VGND sg13g2_decap_8
XFILLER_46_109 VPWR VGND sg13g2_decap_8
XFILLER_27_312 VPWR VGND sg13g2_decap_8
XFILLER_28_868 VPWR VGND sg13g2_decap_8
XFILLER_39_172 VPWR VGND sg13g2_decap_8
XFILLER_83_963 VPWR VGND sg13g2_decap_8
XFILLER_82_462 VPWR VGND sg13g2_decap_8
XFILLER_70_602 VPWR VGND sg13g2_decap_8
XFILLER_55_665 VPWR VGND sg13g2_decap_8
XFILLER_43_805 VPWR VGND sg13g2_decap_8
XFILLER_91_28 VPWR VGND sg13g2_decap_8
XFILLER_54_186 VPWR VGND sg13g2_decap_8
XFILLER_42_326 VPWR VGND sg13g2_decap_8
XFILLER_15_529 VPWR VGND sg13g2_decap_8
XFILLER_27_389 VPWR VGND sg13g2_decap_8
XFILLER_70_679 VPWR VGND sg13g2_decap_8
XFILLER_24_11 VPWR VGND sg13g2_decap_8
XFILLER_51_893 VPWR VGND sg13g2_decap_8
XFILLER_50_392 VPWR VGND sg13g2_decap_8
XFILLER_11_735 VPWR VGND sg13g2_decap_8
XFILLER_23_595 VPWR VGND sg13g2_decap_8
XFILLER_24_88 VPWR VGND sg13g2_decap_8
XFILLER_10_256 VPWR VGND sg13g2_decap_8
XFILLER_7_739 VPWR VGND sg13g2_decap_8
XFILLER_6_238 VPWR VGND sg13g2_decap_8
XFILLER_40_21 VPWR VGND sg13g2_decap_8
XFILLER_105_840 VPWR VGND sg13g2_decap_8
XFILLER_3_945 VPWR VGND sg13g2_decap_8
XFILLER_40_98 VPWR VGND sg13g2_decap_8
XFILLER_104_350 VPWR VGND sg13g2_decap_8
XFILLER_78_713 VPWR VGND sg13g2_decap_8
XFILLER_2_466 VPWR VGND sg13g2_decap_8
XFILLER_93_705 VPWR VGND sg13g2_decap_8
XFILLER_77_245 VPWR VGND sg13g2_decap_8
XFILLER_49_74 VPWR VGND sg13g2_decap_8
XFILLER_59_971 VPWR VGND sg13g2_decap_8
XFILLER_18_301 VPWR VGND sg13g2_decap_8
XFILLER_37_109 VPWR VGND sg13g2_decap_8
XFILLER_105_91 VPWR VGND sg13g2_decap_8
XFILLER_92_259 VPWR VGND sg13g2_decap_8
XFILLER_74_974 VPWR VGND sg13g2_decap_8
XFILLER_65_84 VPWR VGND sg13g2_decap_8
XFILLER_46_676 VPWR VGND sg13g2_decap_8
XFILLER_19_868 VPWR VGND sg13g2_decap_8
XFILLER_34_816 VPWR VGND sg13g2_decap_8
XFILLER_73_473 VPWR VGND sg13g2_decap_8
XFILLER_61_613 VPWR VGND sg13g2_decap_8
XFILLER_45_175 VPWR VGND sg13g2_decap_8
XFILLER_18_378 VPWR VGND sg13g2_decap_8
XFILLER_33_315 VPWR VGND sg13g2_decap_8
XFILLER_60_134 VPWR VGND sg13g2_fill_2
XFILLER_60_123 VPWR VGND sg13g2_decap_8
XFILLER_53_1015 VPWR VGND sg13g2_decap_8
XFILLER_42_893 VPWR VGND sg13g2_decap_8
XFILLER_14_595 VPWR VGND sg13g2_decap_8
XFILLER_41_392 VPWR VGND sg13g2_decap_8
XFILLER_68_201 VPWR VGND sg13g2_decap_8
XFILLER_96_532 VPWR VGND sg13g2_decap_8
XFILLER_69_757 VPWR VGND sg13g2_decap_8
XFILLER_60_1019 VPWR VGND sg13g2_decap_8
XFILLER_68_278 VPWR VGND sg13g2_decap_8
XFILLER_84_749 VPWR VGND sg13g2_decap_8
Xinput3 ui_in[2] net3 VPWR VGND sg13g2_buf_1
XFILLER_65_952 VPWR VGND sg13g2_decap_8
XFILLER_52_602 VPWR VGND sg13g2_decap_8
XFILLER_25_805 VPWR VGND sg13g2_decap_8
XFILLER_37_676 VPWR VGND sg13g2_decap_8
XFILLER_64_473 VPWR VGND sg13g2_decap_8
XFILLER_24_326 VPWR VGND sg13g2_decap_8
XFILLER_36_175 VPWR VGND sg13g2_decap_8
XFILLER_101_49 VPWR VGND sg13g2_decap_8
XFILLER_80_966 VPWR VGND sg13g2_decap_8
XFILLER_52_679 VPWR VGND sg13g2_decap_8
XFILLER_51_123 VPWR VGND sg13g2_decap_8
XFILLER_40_819 VPWR VGND sg13g2_decap_8
XFILLER_33_882 VPWR VGND sg13g2_decap_8
XFILLER_60_690 VPWR VGND sg13g2_decap_8
XFILLER_20_543 VPWR VGND sg13g2_decap_8
XFILLER_106_637 VPWR VGND sg13g2_decap_8
XFILLER_10_46 VPWR VGND sg13g2_decap_8
XFILLER_105_147 VPWR VGND sg13g2_decap_8
XFILLER_59_201 VPWR VGND sg13g2_decap_8
XFILLER_102_854 VPWR VGND sg13g2_decap_8
XFILLER_99_392 VPWR VGND sg13g2_decap_8
XFILLER_87_532 VPWR VGND sg13g2_decap_8
XFILLER_86_39 VPWR VGND sg13g2_decap_8
XFILLER_0_959 VPWR VGND sg13g2_decap_8
XFILLER_101_364 VPWR VGND sg13g2_decap_8
XFILLER_74_204 VPWR VGND sg13g2_decap_8
XFILLER_59_278 VPWR VGND sg13g2_decap_8
XFILLER_75_749 VPWR VGND sg13g2_decap_8
XFILLER_19_77 VPWR VGND sg13g2_decap_8
XFILLER_83_760 VPWR VGND sg13g2_decap_8
XFILLER_71_900 VPWR VGND sg13g2_decap_8
XFILLER_56_963 VPWR VGND sg13g2_decap_8
XFILLER_55_462 VPWR VGND sg13g2_decap_8
XFILLER_43_602 VPWR VGND sg13g2_decap_8
XFILLER_16_805 VPWR VGND sg13g2_decap_8
XFILLER_28_665 VPWR VGND sg13g2_decap_8
XFILLER_76_1026 VPWR VGND sg13g2_fill_2
XFILLER_15_326 VPWR VGND sg13g2_decap_8
XFILLER_27_186 VPWR VGND sg13g2_decap_8
XFILLER_35_21 VPWR VGND sg13g2_decap_8
XFILLER_71_977 VPWR VGND sg13g2_decap_8
XFILLER_42_123 VPWR VGND sg13g2_decap_8
XFILLER_70_476 VPWR VGND sg13g2_decap_8
XFILLER_43_679 VPWR VGND sg13g2_decap_8
XFILLER_31_819 VPWR VGND sg13g2_decap_8
XFILLER_35_98 VPWR VGND sg13g2_decap_8
XFILLER_51_690 VPWR VGND sg13g2_decap_8
XFILLER_11_532 VPWR VGND sg13g2_decap_8
XFILLER_23_392 VPWR VGND sg13g2_decap_8
XFILLER_24_893 VPWR VGND sg13g2_decap_8
XFILLER_30_329 VPWR VGND sg13g2_decap_8
XFILLER_51_53 VPWR VGND sg13g2_decap_8
XFILLER_7_536 VPWR VGND sg13g2_decap_8
XFILLER_83_1019 VPWR VGND sg13g2_decap_8
XFILLER_3_742 VPWR VGND sg13g2_decap_8
XFILLER_97_329 VPWR VGND sg13g2_decap_8
XFILLER_78_510 VPWR VGND sg13g2_decap_8
XFILLER_2_263 VPWR VGND sg13g2_decap_8
XFILLER_93_502 VPWR VGND sg13g2_decap_8
XFILLER_78_587 VPWR VGND sg13g2_decap_8
XFILLER_66_727 VPWR VGND sg13g2_decap_8
XFILLER_18_7 VPWR VGND sg13g2_decap_8
XFILLER_93_579 VPWR VGND sg13g2_decap_8
XFILLER_65_259 VPWR VGND sg13g2_decap_8
XFILLER_47_952 VPWR VGND sg13g2_decap_8
XFILLER_19_665 VPWR VGND sg13g2_decap_8
XFILLER_74_771 VPWR VGND sg13g2_decap_8
XFILLER_73_270 VPWR VGND sg13g2_decap_8
XFILLER_61_410 VPWR VGND sg13g2_decap_8
XFILLER_46_473 VPWR VGND sg13g2_decap_8
XFILLER_18_175 VPWR VGND sg13g2_decap_8
XFILLER_34_613 VPWR VGND sg13g2_decap_8
XFILLER_62_966 VPWR VGND sg13g2_decap_8
XFILLER_33_112 VPWR VGND sg13g2_decap_8
XFILLER_61_487 VPWR VGND sg13g2_decap_8
XFILLER_42_690 VPWR VGND sg13g2_decap_8
XFILLER_14_392 VPWR VGND sg13g2_decap_8
XFILLER_15_893 VPWR VGND sg13g2_decap_8
XFILLER_21_329 VPWR VGND sg13g2_decap_8
XFILLER_33_189 VPWR VGND sg13g2_decap_8
XFILLER_30_896 VPWR VGND sg13g2_decap_8
XFILLER_89_819 VPWR VGND sg13g2_decap_8
XFILLER_69_554 VPWR VGND sg13g2_decap_8
XFILLER_99_1015 VPWR VGND sg13g2_decap_8
XFILLER_97_896 VPWR VGND sg13g2_decap_8
XFILLER_5_1019 VPWR VGND sg13g2_decap_8
XFILLER_84_546 VPWR VGND sg13g2_decap_8
XFILLER_57_749 VPWR VGND sg13g2_decap_8
XFILLER_38_952 VPWR VGND sg13g2_decap_8
XFILLER_71_207 VPWR VGND sg13g2_decap_8
XFILLER_64_270 VPWR VGND sg13g2_decap_8
XFILLER_25_602 VPWR VGND sg13g2_decap_8
XFILLER_37_473 VPWR VGND sg13g2_decap_8
XFILLER_53_966 VPWR VGND sg13g2_decap_8
XFILLER_24_123 VPWR VGND sg13g2_decap_8
XFILLER_80_763 VPWR VGND sg13g2_decap_8
XFILLER_52_476 VPWR VGND sg13g2_decap_8
XFILLER_13_819 VPWR VGND sg13g2_decap_8
XFILLER_25_679 VPWR VGND sg13g2_decap_8
XFILLER_40_616 VPWR VGND sg13g2_decap_8
XFILLER_20_340 VPWR VGND sg13g2_decap_8
XFILLER_21_896 VPWR VGND sg13g2_decap_8
XFILLER_4_539 VPWR VGND sg13g2_decap_8
XFILLER_21_56 VPWR VGND sg13g2_decap_8
XFILLER_106_434 VPWR VGND sg13g2_decap_8
XFILLER_97_49 VPWR VGND sg13g2_decap_8
XFILLER_88_830 VPWR VGND sg13g2_decap_8
XFILLER_0_756 VPWR VGND sg13g2_decap_8
XFILLER_102_651 VPWR VGND sg13g2_decap_8
XFILLER_101_161 VPWR VGND sg13g2_decap_8
XFILLER_75_546 VPWR VGND sg13g2_decap_8
XFILLER_48_749 VPWR VGND sg13g2_decap_8
XFILLER_56_760 VPWR VGND sg13g2_decap_8
XFILLER_47_259 VPWR VGND sg13g2_decap_8
XFILLER_44_900 VPWR VGND sg13g2_decap_8
XFILLER_29_963 VPWR VGND sg13g2_decap_8
XFILLER_46_53 VPWR VGND sg13g2_decap_8
XFILLER_16_602 VPWR VGND sg13g2_decap_8
XFILLER_28_462 VPWR VGND sg13g2_decap_8
XFILLER_44_977 VPWR VGND sg13g2_decap_8
XFILLER_15_123 VPWR VGND sg13g2_decap_8
XFILLER_102_70 VPWR VGND sg13g2_decap_8
XFILLER_71_774 VPWR VGND sg13g2_decap_8
XFILLER_43_476 VPWR VGND sg13g2_decap_8
XFILLER_16_679 VPWR VGND sg13g2_decap_8
XFILLER_31_616 VPWR VGND sg13g2_decap_8
XFILLER_70_273 VPWR VGND sg13g2_decap_8
XFILLER_12_830 VPWR VGND sg13g2_decap_8
XFILLER_24_690 VPWR VGND sg13g2_decap_8
XFILLER_30_126 VPWR VGND sg13g2_decap_8
XFILLER_8_812 VPWR VGND sg13g2_decap_8
XFILLER_7_333 VPWR VGND sg13g2_decap_8
XFILLER_7_25 VPWR VGND sg13g2_decap_8
XFILLER_8_889 VPWR VGND sg13g2_decap_8
XFILLER_98_627 VPWR VGND sg13g2_decap_8
XFILLER_97_126 VPWR VGND sg13g2_decap_8
XFILLER_79_830 VPWR VGND sg13g2_decap_8
XFILLER_94_833 VPWR VGND sg13g2_decap_8
XFILLER_78_384 VPWR VGND sg13g2_decap_8
XFILLER_66_524 VPWR VGND sg13g2_decap_8
XFILLER_38_259 VPWR VGND sg13g2_decap_8
XFILLER_93_376 VPWR VGND sg13g2_decap_8
XFILLER_19_462 VPWR VGND sg13g2_decap_8
XFILLER_34_410 VPWR VGND sg13g2_decap_8
XFILLER_46_270 VPWR VGND sg13g2_decap_8
XFILLER_35_966 VPWR VGND sg13g2_decap_8
XFILLER_62_763 VPWR VGND sg13g2_decap_8
XFILLER_50_903 VPWR VGND sg13g2_decap_8
XFILLER_61_284 VPWR VGND sg13g2_decap_8
XFILLER_15_690 VPWR VGND sg13g2_decap_8
XFILLER_21_126 VPWR VGND sg13g2_decap_8
XFILLER_22_627 VPWR VGND sg13g2_decap_8
XFILLER_34_487 VPWR VGND sg13g2_decap_8
XFILLER_30_693 VPWR VGND sg13g2_decap_8
XFILLER_66_1014 VPWR VGND sg13g2_decap_8
XFILLER_104_938 VPWR VGND sg13g2_decap_8
XFILLER_89_616 VPWR VGND sg13g2_decap_8
XFILLER_103_448 VPWR VGND sg13g2_decap_8
XFILLER_88_137 VPWR VGND sg13g2_decap_8
XFILLER_69_351 VPWR VGND sg13g2_decap_8
XFILLER_97_693 VPWR VGND sg13g2_decap_8
XFILLER_85_833 VPWR VGND sg13g2_decap_8
XFILLER_84_343 VPWR VGND sg13g2_decap_8
XFILLER_57_546 VPWR VGND sg13g2_decap_8
XFILLER_83_18 VPWR VGND sg13g2_decap_8
XFILLER_44_207 VPWR VGND sg13g2_decap_8
XFILLER_26_966 VPWR VGND sg13g2_decap_8
XFILLER_37_270 VPWR VGND sg13g2_decap_8
XFILLER_80_560 VPWR VGND sg13g2_decap_8
XFILLER_53_763 VPWR VGND sg13g2_decap_8
XFILLER_41_903 VPWR VGND sg13g2_decap_8
XFILLER_13_616 VPWR VGND sg13g2_decap_8
XFILLER_16_56 VPWR VGND sg13g2_decap_8
XFILLER_25_476 VPWR VGND sg13g2_decap_8
XFILLER_52_273 VPWR VGND sg13g2_decap_8
XFILLER_40_413 VPWR VGND sg13g2_decap_8
XFILLER_9_609 VPWR VGND sg13g2_decap_8
XFILLER_12_137 VPWR VGND sg13g2_decap_8
XFILLER_32_11 VPWR VGND sg13g2_decap_8
XFILLER_8_119 VPWR VGND sg13g2_decap_8
XFILLER_21_693 VPWR VGND sg13g2_decap_8
XFILLER_32_88 VPWR VGND sg13g2_decap_8
XFILLER_5_837 VPWR VGND sg13g2_decap_8
XFILLER_106_231 VPWR VGND sg13g2_decap_8
XFILLER_4_336 VPWR VGND sg13g2_decap_8
XFILLER_79_137 VPWR VGND sg13g2_decap_8
XFILLER_0_553 VPWR VGND sg13g2_decap_8
XFILLER_76_844 VPWR VGND sg13g2_decap_8
XFILLER_75_343 VPWR VGND sg13g2_decap_8
XFILLER_57_63 VPWR VGND sg13g2_decap_8
XFILLER_48_546 VPWR VGND sg13g2_decap_8
XFILLER_91_847 VPWR VGND sg13g2_decap_8
XFILLER_17_900 VPWR VGND sg13g2_decap_8
XFILLER_29_760 VPWR VGND sg13g2_decap_8
XFILLER_90_368 VPWR VGND sg13g2_decap_8
XFILLER_44_774 VPWR VGND sg13g2_decap_8
XFILLER_16_476 VPWR VGND sg13g2_decap_8
XFILLER_17_977 VPWR VGND sg13g2_decap_8
XFILLER_32_914 VPWR VGND sg13g2_decap_8
XFILLER_73_95 VPWR VGND sg13g2_decap_8
XFILLER_71_571 VPWR VGND sg13g2_decap_8
XFILLER_43_273 VPWR VGND sg13g2_decap_8
XFILLER_31_413 VPWR VGND sg13g2_decap_8
XFILLER_85_7 VPWR VGND sg13g2_decap_8
XFILLER_40_980 VPWR VGND sg13g2_decap_8
XFILLER_7_130 VPWR VGND sg13g2_decap_8
XFILLER_8_686 VPWR VGND sg13g2_decap_8
XFILLER_99_903 VPWR VGND sg13g2_decap_8
XFILLER_98_424 VPWR VGND sg13g2_decap_8
XFILLER_98_81 VPWR VGND sg13g2_decap_8
XFILLER_94_630 VPWR VGND sg13g2_decap_8
XFILLER_67_833 VPWR VGND sg13g2_decap_8
XFILLER_66_321 VPWR VGND sg13g2_decap_8
XFILLER_78_181 VPWR VGND sg13g2_decap_8
XFILLER_39_557 VPWR VGND sg13g2_decap_8
XFILLER_93_173 VPWR VGND sg13g2_decap_8
XFILLER_82_847 VPWR VGND sg13g2_decap_8
XFILLER_66_398 VPWR VGND sg13g2_decap_8
XFILLER_81_368 VPWR VGND sg13g2_decap_8
XFILLER_62_560 VPWR VGND sg13g2_decap_8
XFILLER_50_700 VPWR VGND sg13g2_decap_8
XFILLER_23_903 VPWR VGND sg13g2_decap_8
XFILLER_35_763 VPWR VGND sg13g2_decap_8
XFILLER_22_424 VPWR VGND sg13g2_decap_8
XFILLER_34_284 VPWR VGND sg13g2_decap_8
XFILLER_50_777 VPWR VGND sg13g2_decap_8
XFILLER_31_980 VPWR VGND sg13g2_decap_8
XFILLER_30_490 VPWR VGND sg13g2_decap_8
XFILLER_89_413 VPWR VGND sg13g2_decap_8
XFILLER_78_18 VPWR VGND sg13g2_decap_8
XFILLER_104_735 VPWR VGND sg13g2_decap_8
XFILLER_103_245 VPWR VGND sg13g2_decap_8
XFILLER_98_991 VPWR VGND sg13g2_decap_8
XFILLER_58_833 VPWR VGND sg13g2_decap_8
XFILLER_100_952 VPWR VGND sg13g2_decap_8
XFILLER_97_490 VPWR VGND sg13g2_decap_8
XFILLER_94_28 VPWR VGND sg13g2_decap_8
XFILLER_85_630 VPWR VGND sg13g2_decap_8
XFILLER_57_343 VPWR VGND sg13g2_decap_8
XFILLER_27_11 VPWR VGND sg13g2_decap_8
XFILLER_84_140 VPWR VGND sg13g2_decap_8
XFILLER_17_207 VPWR VGND sg13g2_decap_8
XFILLER_73_858 VPWR VGND sg13g2_decap_8
XFILLER_72_357 VPWR VGND sg13g2_decap_8
XFILLER_60_508 VPWR VGND sg13g2_decap_8
XFILLER_53_560 VPWR VGND sg13g2_decap_8
XFILLER_41_700 VPWR VGND sg13g2_decap_8
XFILLER_14_903 VPWR VGND sg13g2_decap_8
XFILLER_26_763 VPWR VGND sg13g2_decap_8
XFILLER_27_88 VPWR VGND sg13g2_decap_8
XFILLER_43_21 VPWR VGND sg13g2_decap_8
XFILLER_13_413 VPWR VGND sg13g2_decap_8
XFILLER_25_273 VPWR VGND sg13g2_decap_8
XFILLER_40_210 VPWR VGND sg13g2_decap_8
XFILLER_41_777 VPWR VGND sg13g2_decap_8
XFILLER_9_406 VPWR VGND sg13g2_decap_8
XFILLER_43_98 VPWR VGND sg13g2_decap_8
XFILLER_40_287 VPWR VGND sg13g2_decap_8
XFILLER_21_490 VPWR VGND sg13g2_decap_8
XFILLER_22_991 VPWR VGND sg13g2_decap_8
XFILLER_5_634 VPWR VGND sg13g2_decap_8
XFILLER_4_133 VPWR VGND sg13g2_decap_8
XFILLER_96_917 VPWR VGND sg13g2_decap_8
XFILLER_1_840 VPWR VGND sg13g2_decap_8
XFILLER_95_438 VPWR VGND sg13g2_decap_8
XFILLER_89_980 VPWR VGND sg13g2_decap_8
XFILLER_0_350 VPWR VGND sg13g2_decap_8
XFILLER_76_641 VPWR VGND sg13g2_decap_8
XFILLER_49_844 VPWR VGND sg13g2_decap_8
XFILLER_48_343 VPWR VGND sg13g2_decap_8
XFILLER_75_140 VPWR VGND sg13g2_decap_8
XFILLER_91_644 VPWR VGND sg13g2_decap_8
XFILLER_64_858 VPWR VGND sg13g2_decap_8
XFILLER_1_1022 VPWR VGND sg13g2_decap_8
XFILLER_90_165 VPWR VGND sg13g2_decap_8
XFILLER_63_357 VPWR VGND sg13g2_decap_8
XFILLER_51_508 VPWR VGND sg13g2_decap_8
XFILLER_17_774 VPWR VGND sg13g2_decap_8
XFILLER_44_571 VPWR VGND sg13g2_decap_8
XFILLER_16_273 VPWR VGND sg13g2_decap_8
XFILLER_31_210 VPWR VGND sg13g2_decap_8
XFILLER_32_711 VPWR VGND sg13g2_decap_8
XFILLER_17_1019 VPWR VGND sg13g2_decap_8
XFILLER_83_4 VPWR VGND sg13g2_decap_8
XFILLER_13_980 VPWR VGND sg13g2_decap_8
XFILLER_20_928 VPWR VGND sg13g2_decap_8
XFILLER_32_788 VPWR VGND sg13g2_decap_8
XFILLER_31_287 VPWR VGND sg13g2_decap_8
XFILLER_9_973 VPWR VGND sg13g2_decap_8
XFILLER_8_483 VPWR VGND sg13g2_decap_8
XFILLER_99_700 VPWR VGND sg13g2_decap_8
XFILLER_98_221 VPWR VGND sg13g2_decap_8
XFILLER_99_777 VPWR VGND sg13g2_decap_8
XFILLER_87_917 VPWR VGND sg13g2_decap_8
XFILLER_101_749 VPWR VGND sg13g2_decap_8
XFILLER_98_298 VPWR VGND sg13g2_decap_8
XFILLER_86_438 VPWR VGND sg13g2_decap_8
XFILLER_100_259 VPWR VGND sg13g2_decap_8
XFILLER_67_630 VPWR VGND sg13g2_decap_8
XFILLER_104_49 VPWR VGND sg13g2_decap_8
XFILLER_39_354 VPWR VGND sg13g2_decap_8
XFILLER_82_644 VPWR VGND sg13g2_decap_8
XFILLER_66_195 VPWR VGND sg13g2_decap_8
XFILLER_55_847 VPWR VGND sg13g2_decap_8
XFILLER_81_165 VPWR VGND sg13g2_decap_8
XFILLER_54_368 VPWR VGND sg13g2_decap_8
XFILLER_42_508 VPWR VGND sg13g2_decap_8
XFILLER_23_700 VPWR VGND sg13g2_decap_8
XFILLER_35_560 VPWR VGND sg13g2_decap_8
XFILLER_22_221 VPWR VGND sg13g2_decap_8
XFILLER_50_574 VPWR VGND sg13g2_decap_8
XFILLER_11_917 VPWR VGND sg13g2_decap_8
XFILLER_23_777 VPWR VGND sg13g2_decap_8
XFILLER_10_438 VPWR VGND sg13g2_decap_8
XFILLER_13_35 VPWR VGND sg13g2_decap_8
XFILLER_22_298 VPWR VGND sg13g2_decap_8
XFILLER_89_28 VPWR VGND sg13g2_decap_8
XFILLER_104_532 VPWR VGND sg13g2_decap_8
XFILLER_89_210 VPWR VGND sg13g2_decap_8
XFILLER_2_648 VPWR VGND sg13g2_decap_8
XFILLER_1_147 VPWR VGND sg13g2_decap_8
XFILLER_89_287 VPWR VGND sg13g2_decap_8
XFILLER_77_427 VPWR VGND sg13g2_decap_8
XFILLER_38_21 VPWR VGND sg13g2_decap_8
XFILLER_58_630 VPWR VGND sg13g2_decap_8
XFILLER_57_140 VPWR VGND sg13g2_decap_8
XFILLER_46_858 VPWR VGND sg13g2_decap_8
XFILLER_38_98 VPWR VGND sg13g2_decap_8
XFILLER_73_655 VPWR VGND sg13g2_decap_8
XFILLER_72_154 VPWR VGND sg13g2_decap_8
XFILLER_45_357 VPWR VGND sg13g2_decap_8
XFILLER_60_305 VPWR VGND sg13g2_decap_8
XFILLER_54_53 VPWR VGND sg13g2_decap_8
XFILLER_14_700 VPWR VGND sg13g2_decap_8
XFILLER_26_560 VPWR VGND sg13g2_decap_8
XFILLER_13_210 VPWR VGND sg13g2_decap_8
XFILLER_9_203 VPWR VGND sg13g2_decap_8
XFILLER_14_777 VPWR VGND sg13g2_decap_8
XFILLER_41_574 VPWR VGND sg13g2_decap_8
XFILLER_13_287 VPWR VGND sg13g2_decap_8
XFILLER_103_1022 VPWR VGND sg13g2_decap_8
XFILLER_70_63 VPWR VGND sg13g2_decap_8
XFILLER_6_910 VPWR VGND sg13g2_decap_8
XFILLER_5_431 VPWR VGND sg13g2_decap_8
XFILLER_86_1028 VPWR VGND sg13g2_fill_1
XFILLER_6_987 VPWR VGND sg13g2_decap_8
XFILLER_48_7 VPWR VGND sg13g2_decap_8
XFILLER_96_714 VPWR VGND sg13g2_decap_8
XFILLER_69_939 VPWR VGND sg13g2_decap_8
XFILLER_95_235 VPWR VGND sg13g2_decap_8
XFILLER_49_641 VPWR VGND sg13g2_decap_8
XFILLER_23_1001 VPWR VGND sg13g2_decap_8
XFILLER_95_60 VPWR VGND sg13g2_decap_8
XFILLER_77_994 VPWR VGND sg13g2_decap_8
XFILLER_48_140 VPWR VGND sg13g2_decap_8
XFILLER_92_931 VPWR VGND sg13g2_decap_8
XFILLER_37_858 VPWR VGND sg13g2_decap_8
XFILLER_91_441 VPWR VGND sg13g2_decap_8
XFILLER_64_655 VPWR VGND sg13g2_decap_8
XFILLER_63_154 VPWR VGND sg13g2_decap_8
XFILLER_24_508 VPWR VGND sg13g2_decap_8
XFILLER_36_357 VPWR VGND sg13g2_decap_8
XFILLER_51_305 VPWR VGND sg13g2_decap_8
XFILLER_17_571 VPWR VGND sg13g2_decap_8
XFILLER_60_872 VPWR VGND sg13g2_decap_8
XFILLER_20_725 VPWR VGND sg13g2_decap_8
XFILLER_32_585 VPWR VGND sg13g2_decap_8
XFILLER_74_0 VPWR VGND sg13g2_decap_8
XFILLER_9_770 VPWR VGND sg13g2_decap_8
XFILLER_8_280 VPWR VGND sg13g2_decap_8
XFILLER_106_819 VPWR VGND sg13g2_decap_8
XFILLER_105_329 VPWR VGND sg13g2_decap_8
XFILLER_99_574 VPWR VGND sg13g2_decap_8
XFILLER_87_714 VPWR VGND sg13g2_decap_8
XFILLER_101_546 VPWR VGND sg13g2_decap_8
XFILLER_86_235 VPWR VGND sg13g2_decap_8
XFILLER_68_950 VPWR VGND sg13g2_decap_8
XFILLER_39_151 VPWR VGND sg13g2_decap_8
XFILLER_83_942 VPWR VGND sg13g2_decap_8
XFILLER_55_644 VPWR VGND sg13g2_decap_8
XFILLER_28_847 VPWR VGND sg13g2_decap_8
XFILLER_82_441 VPWR VGND sg13g2_decap_8
XFILLER_15_508 VPWR VGND sg13g2_decap_8
XFILLER_27_368 VPWR VGND sg13g2_decap_8
XFILLER_54_165 VPWR VGND sg13g2_decap_8
XFILLER_42_305 VPWR VGND sg13g2_decap_8
XFILLER_70_658 VPWR VGND sg13g2_decap_8
XFILLER_51_872 VPWR VGND sg13g2_decap_8
XFILLER_11_714 VPWR VGND sg13g2_decap_8
XFILLER_23_574 VPWR VGND sg13g2_decap_8
XFILLER_24_67 VPWR VGND sg13g2_decap_8
XFILLER_50_371 VPWR VGND sg13g2_decap_8
XFILLER_10_235 VPWR VGND sg13g2_decap_8
XFILLER_7_718 VPWR VGND sg13g2_decap_8
XFILLER_6_217 VPWR VGND sg13g2_decap_8
XFILLER_40_77 VPWR VGND sg13g2_decap_8
XFILLER_3_924 VPWR VGND sg13g2_decap_8
XFILLER_46_1012 VPWR VGND sg13g2_decap_8
XFILLER_2_445 VPWR VGND sg13g2_decap_8
XFILLER_105_896 VPWR VGND sg13g2_decap_8
XFILLER_49_53 VPWR VGND sg13g2_decap_8
XFILLER_78_769 VPWR VGND sg13g2_decap_8
XFILLER_77_224 VPWR VGND sg13g2_decap_8
XFILLER_66_909 VPWR VGND sg13g2_decap_8
XFILLER_59_950 VPWR VGND sg13g2_decap_8
XFILLER_105_70 VPWR VGND sg13g2_decap_8
XFILLER_92_238 VPWR VGND sg13g2_decap_8
XFILLER_74_953 VPWR VGND sg13g2_decap_8
XFILLER_1_49 VPWR VGND sg13g2_decap_8
XFILLER_19_847 VPWR VGND sg13g2_decap_8
XFILLER_73_452 VPWR VGND sg13g2_decap_8
XFILLER_65_63 VPWR VGND sg13g2_decap_8
XFILLER_46_655 VPWR VGND sg13g2_decap_8
XFILLER_45_154 VPWR VGND sg13g2_decap_8
XFILLER_18_357 VPWR VGND sg13g2_decap_8
XFILLER_60_102 VPWR VGND sg13g2_decap_8
XFILLER_61_669 VPWR VGND sg13g2_decap_8
XFILLER_60_179 VPWR VGND sg13g2_decap_8
XFILLER_42_872 VPWR VGND sg13g2_decap_8
XFILLER_14_574 VPWR VGND sg13g2_decap_8
XFILLER_81_95 VPWR VGND sg13g2_decap_8
XFILLER_41_371 VPWR VGND sg13g2_decap_8
XFILLER_6_784 VPWR VGND sg13g2_decap_8
XFILLER_46_4 VPWR VGND sg13g2_decap_8
XFILLER_96_511 VPWR VGND sg13g2_decap_8
XFILLER_69_736 VPWR VGND sg13g2_decap_8
XFILLER_96_588 VPWR VGND sg13g2_decap_8
XFILLER_84_728 VPWR VGND sg13g2_decap_8
XFILLER_68_257 VPWR VGND sg13g2_decap_8
XFILLER_83_249 VPWR VGND sg13g2_decap_8
XFILLER_77_791 VPWR VGND sg13g2_decap_8
Xinput4 ui_in[3] net4 VPWR VGND sg13g2_buf_1
XFILLER_65_931 VPWR VGND sg13g2_decap_8
XFILLER_64_452 VPWR VGND sg13g2_decap_8
XFILLER_37_655 VPWR VGND sg13g2_decap_8
XFILLER_80_945 VPWR VGND sg13g2_decap_8
XFILLER_51_102 VPWR VGND sg13g2_decap_8
XFILLER_24_305 VPWR VGND sg13g2_decap_8
XFILLER_36_154 VPWR VGND sg13g2_decap_8
XFILLER_101_28 VPWR VGND sg13g2_decap_8
XFILLER_52_658 VPWR VGND sg13g2_decap_8
XFILLER_51_179 VPWR VGND sg13g2_decap_8
XFILLER_33_861 VPWR VGND sg13g2_decap_8
XFILLER_20_522 VPWR VGND sg13g2_decap_8
XFILLER_32_382 VPWR VGND sg13g2_decap_8
XFILLER_20_599 VPWR VGND sg13g2_decap_8
XFILLER_106_616 VPWR VGND sg13g2_decap_8
XFILLER_69_1023 VPWR VGND sg13g2_decap_4
XFILLER_105_126 VPWR VGND sg13g2_decap_8
XFILLER_10_25 VPWR VGND sg13g2_decap_8
XFILLER_99_371 VPWR VGND sg13g2_decap_8
XFILLER_87_511 VPWR VGND sg13g2_decap_8
XFILLER_86_18 VPWR VGND sg13g2_decap_8
XFILLER_0_938 VPWR VGND sg13g2_decap_8
XFILLER_102_833 VPWR VGND sg13g2_decap_8
XFILLER_101_343 VPWR VGND sg13g2_decap_8
XFILLER_87_588 VPWR VGND sg13g2_decap_8
XFILLER_75_728 VPWR VGND sg13g2_decap_8
XFILLER_59_257 VPWR VGND sg13g2_decap_8
XFILLER_19_56 VPWR VGND sg13g2_decap_8
XFILLER_56_942 VPWR VGND sg13g2_decap_8
XFILLER_55_441 VPWR VGND sg13g2_decap_8
XFILLER_28_644 VPWR VGND sg13g2_decap_8
XFILLER_76_1005 VPWR VGND sg13g2_decap_8
XFILLER_42_102 VPWR VGND sg13g2_decap_8
XFILLER_15_305 VPWR VGND sg13g2_decap_8
XFILLER_27_165 VPWR VGND sg13g2_decap_8
XFILLER_71_956 VPWR VGND sg13g2_decap_8
XFILLER_43_658 VPWR VGND sg13g2_decap_8
XFILLER_70_455 VPWR VGND sg13g2_decap_8
XFILLER_42_179 VPWR VGND sg13g2_decap_8
XFILLER_24_872 VPWR VGND sg13g2_decap_8
XFILLER_30_308 VPWR VGND sg13g2_decap_8
XFILLER_35_77 VPWR VGND sg13g2_decap_8
XFILLER_11_511 VPWR VGND sg13g2_decap_8
XFILLER_23_371 VPWR VGND sg13g2_decap_8
XFILLER_51_32 VPWR VGND sg13g2_decap_8
XFILLER_7_515 VPWR VGND sg13g2_decap_8
XFILLER_11_588 VPWR VGND sg13g2_decap_8
XFILLER_13_1022 VPWR VGND sg13g2_decap_8
XFILLER_3_721 VPWR VGND sg13g2_decap_8
XFILLER_98_809 VPWR VGND sg13g2_decap_8
XFILLER_4_0 VPWR VGND sg13g2_decap_8
XFILLER_97_308 VPWR VGND sg13g2_decap_8
XFILLER_3_798 VPWR VGND sg13g2_decap_8
XFILLER_2_242 VPWR VGND sg13g2_decap_8
XFILLER_105_693 VPWR VGND sg13g2_decap_8
XFILLER_78_566 VPWR VGND sg13g2_decap_8
XFILLER_66_706 VPWR VGND sg13g2_decap_8
XFILLER_65_238 VPWR VGND sg13g2_decap_8
XFILLER_47_931 VPWR VGND sg13g2_decap_8
XFILLER_93_558 VPWR VGND sg13g2_decap_8
XFILLER_76_95 VPWR VGND sg13g2_decap_8
XFILLER_74_750 VPWR VGND sg13g2_decap_8
XFILLER_46_452 VPWR VGND sg13g2_decap_8
XFILLER_19_644 VPWR VGND sg13g2_decap_8
XFILLER_20_1026 VPWR VGND sg13g2_fill_2
XFILLER_18_154 VPWR VGND sg13g2_decap_8
XFILLER_62_945 VPWR VGND sg13g2_decap_8
XFILLER_22_809 VPWR VGND sg13g2_decap_8
XFILLER_34_669 VPWR VGND sg13g2_decap_8
XFILLER_61_466 VPWR VGND sg13g2_decap_8
XFILLER_15_872 VPWR VGND sg13g2_decap_8
XFILLER_21_308 VPWR VGND sg13g2_decap_8
XFILLER_33_168 VPWR VGND sg13g2_decap_8
XFILLER_14_371 VPWR VGND sg13g2_decap_8
XFILLER_30_875 VPWR VGND sg13g2_decap_8
XFILLER_6_581 VPWR VGND sg13g2_decap_8
XFILLER_88_319 VPWR VGND sg13g2_decap_8
XFILLER_69_533 VPWR VGND sg13g2_decap_8
XFILLER_97_875 VPWR VGND sg13g2_decap_8
XFILLER_57_728 VPWR VGND sg13g2_decap_8
XFILLER_96_385 VPWR VGND sg13g2_decap_8
XFILLER_84_525 VPWR VGND sg13g2_decap_8
XFILLER_38_931 VPWR VGND sg13g2_decap_8
XFILLER_56_249 VPWR VGND sg13g2_decap_8
XFILLER_2_81 VPWR VGND sg13g2_decap_8
XFILLER_37_452 VPWR VGND sg13g2_decap_8
XFILLER_24_102 VPWR VGND sg13g2_decap_8
XFILLER_80_742 VPWR VGND sg13g2_decap_8
XFILLER_53_945 VPWR VGND sg13g2_decap_8
XFILLER_25_658 VPWR VGND sg13g2_decap_8
XFILLER_52_455 VPWR VGND sg13g2_decap_8
XFILLER_12_319 VPWR VGND sg13g2_decap_8
XFILLER_24_179 VPWR VGND sg13g2_decap_8
XFILLER_36_1022 VPWR VGND sg13g2_decap_8
XFILLER_21_875 VPWR VGND sg13g2_decap_8
XFILLER_20_396 VPWR VGND sg13g2_decap_8
XFILLER_21_35 VPWR VGND sg13g2_decap_8
XFILLER_106_413 VPWR VGND sg13g2_decap_8
XFILLER_4_518 VPWR VGND sg13g2_decap_8
XFILLER_97_28 VPWR VGND sg13g2_decap_8
XFILLER_79_319 VPWR VGND sg13g2_decap_8
XFILLER_102_630 VPWR VGND sg13g2_decap_8
XFILLER_43_1015 VPWR VGND sg13g2_decap_8
XFILLER_0_735 VPWR VGND sg13g2_decap_8
XFILLER_101_140 VPWR VGND sg13g2_decap_8
XFILLER_88_886 VPWR VGND sg13g2_decap_8
XFILLER_48_728 VPWR VGND sg13g2_decap_8
XFILLER_87_385 VPWR VGND sg13g2_decap_8
XFILLER_75_525 VPWR VGND sg13g2_decap_8
XFILLER_47_238 VPWR VGND sg13g2_decap_8
XFILLER_46_32 VPWR VGND sg13g2_decap_8
XFILLER_28_441 VPWR VGND sg13g2_decap_8
XFILLER_29_942 VPWR VGND sg13g2_decap_8
XFILLER_71_753 VPWR VGND sg13g2_decap_8
XFILLER_44_956 VPWR VGND sg13g2_decap_8
XFILLER_15_102 VPWR VGND sg13g2_decap_8
XFILLER_16_658 VPWR VGND sg13g2_decap_8
XFILLER_70_252 VPWR VGND sg13g2_decap_8
XFILLER_43_455 VPWR VGND sg13g2_decap_8
XFILLER_62_42 VPWR VGND sg13g2_decap_8
XFILLER_15_179 VPWR VGND sg13g2_decap_8
XFILLER_30_105 VPWR VGND sg13g2_decap_8
XFILLER_50_1008 VPWR VGND sg13g2_decap_8
XFILLER_7_312 VPWR VGND sg13g2_decap_8
XFILLER_12_886 VPWR VGND sg13g2_decap_8
XFILLER_8_868 VPWR VGND sg13g2_decap_8
XFILLER_11_385 VPWR VGND sg13g2_decap_8
XFILLER_7_389 VPWR VGND sg13g2_decap_8
XFILLER_98_606 VPWR VGND sg13g2_decap_8
XFILLER_106_980 VPWR VGND sg13g2_decap_8
XFILLER_97_105 VPWR VGND sg13g2_decap_8
XFILLER_105_490 VPWR VGND sg13g2_decap_8
XFILLER_3_595 VPWR VGND sg13g2_decap_8
XFILLER_30_7 VPWR VGND sg13g2_decap_8
XFILLER_94_812 VPWR VGND sg13g2_decap_8
XFILLER_79_886 VPWR VGND sg13g2_decap_8
XFILLER_78_363 VPWR VGND sg13g2_decap_8
XFILLER_66_503 VPWR VGND sg13g2_decap_8
XFILLER_39_739 VPWR VGND sg13g2_decap_8
XFILLER_94_889 VPWR VGND sg13g2_decap_8
XFILLER_93_355 VPWR VGND sg13g2_decap_8
XFILLER_19_441 VPWR VGND sg13g2_decap_8
XFILLER_38_238 VPWR VGND sg13g2_decap_8
XFILLER_62_742 VPWR VGND sg13g2_decap_8
XFILLER_35_945 VPWR VGND sg13g2_decap_8
XFILLER_22_606 VPWR VGND sg13g2_decap_8
XFILLER_34_466 VPWR VGND sg13g2_decap_8
XFILLER_61_263 VPWR VGND sg13g2_decap_8
XFILLER_50_959 VPWR VGND sg13g2_decap_8
XFILLER_21_105 VPWR VGND sg13g2_decap_8
XFILLER_30_672 VPWR VGND sg13g2_decap_8
XFILLER_104_917 VPWR VGND sg13g2_decap_8
XFILLER_103_427 VPWR VGND sg13g2_decap_8
XFILLER_88_116 VPWR VGND sg13g2_decap_8
XFILLER_85_812 VPWR VGND sg13g2_decap_8
XFILLER_69_330 VPWR VGND sg13g2_decap_8
XFILLER_97_672 VPWR VGND sg13g2_decap_8
XFILLER_84_322 VPWR VGND sg13g2_decap_8
XFILLER_57_525 VPWR VGND sg13g2_decap_8
XFILLER_96_182 VPWR VGND sg13g2_decap_8
XFILLER_29_249 VPWR VGND sg13g2_decap_8
XFILLER_85_889 VPWR VGND sg13g2_decap_8
XFILLER_84_399 VPWR VGND sg13g2_decap_8
XFILLER_72_539 VPWR VGND sg13g2_decap_8
XFILLER_53_742 VPWR VGND sg13g2_decap_8
XFILLER_16_35 VPWR VGND sg13g2_decap_8
XFILLER_26_945 VPWR VGND sg13g2_decap_8
XFILLER_73_1019 VPWR VGND sg13g2_decap_8
XFILLER_52_252 VPWR VGND sg13g2_decap_8
XFILLER_25_455 VPWR VGND sg13g2_decap_8
XFILLER_41_959 VPWR VGND sg13g2_decap_8
XFILLER_12_116 VPWR VGND sg13g2_decap_8
XFILLER_40_469 VPWR VGND sg13g2_decap_8
XFILLER_21_672 VPWR VGND sg13g2_decap_8
XFILLER_20_193 VPWR VGND sg13g2_decap_8
XFILLER_32_67 VPWR VGND sg13g2_decap_8
XFILLER_5_816 VPWR VGND sg13g2_decap_8
XFILLER_4_315 VPWR VGND sg13g2_decap_8
XFILLER_106_210 VPWR VGND sg13g2_decap_8
XFILLER_106_287 VPWR VGND sg13g2_decap_8
XFILLER_79_116 VPWR VGND sg13g2_decap_8
XFILLER_0_532 VPWR VGND sg13g2_decap_8
XFILLER_103_994 VPWR VGND sg13g2_decap_8
XFILLER_94_119 VPWR VGND sg13g2_decap_8
XFILLER_88_683 VPWR VGND sg13g2_decap_8
XFILLER_76_823 VPWR VGND sg13g2_decap_8
XFILLER_57_42 VPWR VGND sg13g2_decap_8
XFILLER_48_525 VPWR VGND sg13g2_decap_8
XFILLER_87_182 VPWR VGND sg13g2_decap_8
XFILLER_75_322 VPWR VGND sg13g2_decap_8
XFILLER_91_826 VPWR VGND sg13g2_decap_8
XFILLER_90_347 VPWR VGND sg13g2_decap_8
XFILLER_75_399 VPWR VGND sg13g2_decap_8
XFILLER_63_539 VPWR VGND sg13g2_decap_8
XFILLER_17_956 VPWR VGND sg13g2_decap_8
XFILLER_73_74 VPWR VGND sg13g2_decap_8
XFILLER_71_550 VPWR VGND sg13g2_decap_8
XFILLER_44_753 VPWR VGND sg13g2_decap_8
XFILLER_43_252 VPWR VGND sg13g2_decap_8
XFILLER_16_455 VPWR VGND sg13g2_decap_8
XFILLER_31_469 VPWR VGND sg13g2_decap_8
XFILLER_89_1015 VPWR VGND sg13g2_decap_8
XFILLER_8_665 VPWR VGND sg13g2_decap_8
XFILLER_11_182 VPWR VGND sg13g2_decap_8
XFILLER_12_683 VPWR VGND sg13g2_decap_8
XFILLER_7_186 VPWR VGND sg13g2_decap_8
XFILLER_98_403 VPWR VGND sg13g2_decap_8
XFILLER_98_60 VPWR VGND sg13g2_decap_8
XFILLER_99_959 VPWR VGND sg13g2_decap_8
XFILLER_4_882 VPWR VGND sg13g2_decap_8
XFILLER_3_392 VPWR VGND sg13g2_decap_8
XFILLER_85_119 VPWR VGND sg13g2_decap_8
XFILLER_79_683 VPWR VGND sg13g2_decap_8
XFILLER_78_160 VPWR VGND sg13g2_decap_8
XFILLER_67_812 VPWR VGND sg13g2_decap_8
XFILLER_66_300 VPWR VGND sg13g2_decap_8
XFILLER_39_536 VPWR VGND sg13g2_decap_8
XFILLER_96_1008 VPWR VGND sg13g2_decap_8
XFILLER_94_686 VPWR VGND sg13g2_decap_8
XFILLER_93_152 VPWR VGND sg13g2_decap_8
XFILLER_82_826 VPWR VGND sg13g2_decap_8
XFILLER_67_889 VPWR VGND sg13g2_decap_8
XFILLER_66_377 VPWR VGND sg13g2_decap_8
XFILLER_81_347 VPWR VGND sg13g2_decap_8
XFILLER_35_742 VPWR VGND sg13g2_decap_8
XFILLER_22_403 VPWR VGND sg13g2_decap_8
XFILLER_34_263 VPWR VGND sg13g2_decap_8
XFILLER_50_756 VPWR VGND sg13g2_decap_8
XFILLER_23_959 VPWR VGND sg13g2_decap_8
XFILLER_8_91 VPWR VGND sg13g2_decap_8
XFILLER_104_714 VPWR VGND sg13g2_decap_8
XFILLER_103_224 VPWR VGND sg13g2_decap_8
XFILLER_1_329 VPWR VGND sg13g2_decap_8
XFILLER_98_970 VPWR VGND sg13g2_decap_8
XFILLER_89_469 VPWR VGND sg13g2_decap_8
XFILLER_77_609 VPWR VGND sg13g2_decap_8
XFILLER_58_812 VPWR VGND sg13g2_decap_8
XFILLER_100_931 VPWR VGND sg13g2_decap_8
XFILLER_57_322 VPWR VGND sg13g2_decap_8
XFILLER_85_686 VPWR VGND sg13g2_decap_8
XFILLER_73_837 VPWR VGND sg13g2_decap_8
XFILLER_58_889 VPWR VGND sg13g2_decap_8
XFILLER_84_196 VPWR VGND sg13g2_decap_8
XFILLER_72_336 VPWR VGND sg13g2_decap_8
XFILLER_57_399 VPWR VGND sg13g2_decap_8
XFILLER_45_539 VPWR VGND sg13g2_decap_8
XFILLER_27_67 VPWR VGND sg13g2_decap_8
XFILLER_26_742 VPWR VGND sg13g2_decap_8
XFILLER_25_252 VPWR VGND sg13g2_decap_8
XFILLER_41_756 VPWR VGND sg13g2_decap_8
XFILLER_14_959 VPWR VGND sg13g2_decap_8
XFILLER_43_77 VPWR VGND sg13g2_decap_8
XFILLER_13_469 VPWR VGND sg13g2_decap_8
XFILLER_22_970 VPWR VGND sg13g2_decap_8
XFILLER_40_266 VPWR VGND sg13g2_decap_8
XFILLER_5_613 VPWR VGND sg13g2_decap_8
XFILLER_4_112 VPWR VGND sg13g2_decap_8
XFILLER_104_0 VPWR VGND sg13g2_decap_8
XFILLER_4_189 VPWR VGND sg13g2_decap_8
XFILLER_4_49 VPWR VGND sg13g2_decap_8
XFILLER_95_417 VPWR VGND sg13g2_decap_8
XFILLER_76_620 VPWR VGND sg13g2_decap_8
XFILLER_68_96 VPWR VGND sg13g2_decap_8
XFILLER_67_119 VPWR VGND sg13g2_decap_8
XFILLER_49_823 VPWR VGND sg13g2_decap_8
XFILLER_1_896 VPWR VGND sg13g2_decap_8
XFILLER_103_791 VPWR VGND sg13g2_decap_8
XFILLER_88_480 VPWR VGND sg13g2_decap_8
XFILLER_48_322 VPWR VGND sg13g2_decap_8
XFILLER_91_623 VPWR VGND sg13g2_decap_8
XFILLER_76_697 VPWR VGND sg13g2_decap_8
XFILLER_75_196 VPWR VGND sg13g2_decap_8
XFILLER_64_837 VPWR VGND sg13g2_decap_8
XFILLER_63_336 VPWR VGND sg13g2_decap_8
XFILLER_48_399 VPWR VGND sg13g2_decap_8
XFILLER_1_1001 VPWR VGND sg13g2_decap_8
XFILLER_36_539 VPWR VGND sg13g2_decap_8
XFILLER_90_144 VPWR VGND sg13g2_decap_8
XFILLER_84_84 VPWR VGND sg13g2_decap_8
XFILLER_44_550 VPWR VGND sg13g2_decap_8
XFILLER_17_753 VPWR VGND sg13g2_decap_8
XFILLER_16_252 VPWR VGND sg13g2_decap_8
XFILLER_20_907 VPWR VGND sg13g2_decap_8
XFILLER_32_767 VPWR VGND sg13g2_decap_8
XFILLER_31_266 VPWR VGND sg13g2_decap_8
XFILLER_9_952 VPWR VGND sg13g2_decap_8
XFILLER_12_480 VPWR VGND sg13g2_decap_8
XFILLER_76_4 VPWR VGND sg13g2_decap_8
XFILLER_8_462 VPWR VGND sg13g2_decap_8
XFILLER_98_200 VPWR VGND sg13g2_decap_8
XFILLER_99_756 VPWR VGND sg13g2_decap_8
XFILLER_101_728 VPWR VGND sg13g2_decap_8
XFILLER_98_277 VPWR VGND sg13g2_decap_8
XFILLER_86_417 VPWR VGND sg13g2_decap_8
XFILLER_58_119 VPWR VGND sg13g2_decap_8
XFILLER_100_238 VPWR VGND sg13g2_decap_8
XFILLER_79_480 VPWR VGND sg13g2_decap_8
XFILLER_39_333 VPWR VGND sg13g2_decap_8
XFILLER_104_28 VPWR VGND sg13g2_decap_8
XFILLER_95_984 VPWR VGND sg13g2_decap_8
XFILLER_67_686 VPWR VGND sg13g2_decap_8
XFILLER_55_826 VPWR VGND sg13g2_decap_8
XFILLER_94_483 VPWR VGND sg13g2_decap_8
XFILLER_82_623 VPWR VGND sg13g2_decap_8
XFILLER_66_174 VPWR VGND sg13g2_decap_8
XFILLER_81_144 VPWR VGND sg13g2_decap_8
XFILLER_54_347 VPWR VGND sg13g2_decap_8
XFILLER_22_200 VPWR VGND sg13g2_decap_8
XFILLER_23_756 VPWR VGND sg13g2_decap_8
XFILLER_50_553 VPWR VGND sg13g2_decap_8
XFILLER_10_417 VPWR VGND sg13g2_decap_8
XFILLER_13_14 VPWR VGND sg13g2_decap_8
XFILLER_22_277 VPWR VGND sg13g2_decap_8
XFILLER_104_511 VPWR VGND sg13g2_decap_8
XFILLER_8_7 VPWR VGND sg13g2_decap_8
XFILLER_2_627 VPWR VGND sg13g2_decap_8
XFILLER_1_126 VPWR VGND sg13g2_decap_8
XFILLER_104_588 VPWR VGND sg13g2_decap_8
XFILLER_89_266 VPWR VGND sg13g2_decap_8
XFILLER_77_406 VPWR VGND sg13g2_decap_8
XFILLER_86_984 VPWR VGND sg13g2_decap_8
XFILLER_58_686 VPWR VGND sg13g2_decap_8
XFILLER_38_77 VPWR VGND sg13g2_decap_8
XFILLER_85_483 VPWR VGND sg13g2_decap_8
XFILLER_73_634 VPWR VGND sg13g2_decap_8
XFILLER_57_196 VPWR VGND sg13g2_decap_8
XFILLER_46_837 VPWR VGND sg13g2_decap_8
XFILLER_45_336 VPWR VGND sg13g2_decap_8
XFILLER_18_539 VPWR VGND sg13g2_decap_8
XFILLER_72_133 VPWR VGND sg13g2_decap_8
XFILLER_54_32 VPWR VGND sg13g2_decap_8
XFILLER_14_756 VPWR VGND sg13g2_decap_8
XFILLER_13_266 VPWR VGND sg13g2_decap_8
XFILLER_41_553 VPWR VGND sg13g2_decap_8
XFILLER_103_1001 VPWR VGND sg13g2_decap_8
XFILLER_70_42 VPWR VGND sg13g2_decap_8
XFILLER_9_259 VPWR VGND sg13g2_decap_8
XFILLER_5_410 VPWR VGND sg13g2_decap_8
XFILLER_10_984 VPWR VGND sg13g2_decap_8
XFILLER_6_966 VPWR VGND sg13g2_decap_8
XFILLER_5_487 VPWR VGND sg13g2_decap_8
XFILLER_79_95 VPWR VGND sg13g2_decap_8
XFILLER_69_918 VPWR VGND sg13g2_decap_8
XFILLER_95_214 VPWR VGND sg13g2_decap_8
XFILLER_68_439 VPWR VGND sg13g2_decap_8
XFILLER_49_620 VPWR VGND sg13g2_decap_8
XFILLER_1_693 VPWR VGND sg13g2_decap_8
XFILLER_92_910 VPWR VGND sg13g2_decap_8
XFILLER_77_973 VPWR VGND sg13g2_decap_8
XFILLER_91_420 VPWR VGND sg13g2_decap_8
XFILLER_76_494 VPWR VGND sg13g2_decap_8
XFILLER_64_634 VPWR VGND sg13g2_decap_8
XFILLER_49_697 VPWR VGND sg13g2_decap_8
XFILLER_36_336 VPWR VGND sg13g2_decap_8
XFILLER_37_837 VPWR VGND sg13g2_decap_8
XFILLER_92_987 VPWR VGND sg13g2_decap_8
XFILLER_63_133 VPWR VGND sg13g2_decap_8
XFILLER_48_196 VPWR VGND sg13g2_decap_8
XFILLER_91_497 VPWR VGND sg13g2_decap_8
XFILLER_17_550 VPWR VGND sg13g2_decap_8
XFILLER_60_851 VPWR VGND sg13g2_decap_8
XFILLER_20_704 VPWR VGND sg13g2_decap_8
XFILLER_32_564 VPWR VGND sg13g2_decap_8
XFILLER_67_0 VPWR VGND sg13g2_decap_8
XFILLER_105_308 VPWR VGND sg13g2_decap_8
XFILLER_99_553 VPWR VGND sg13g2_decap_8
XFILLER_5_81 VPWR VGND sg13g2_decap_8
XFILLER_86_214 VPWR VGND sg13g2_decap_8
XFILLER_101_525 VPWR VGND sg13g2_decap_8
XFILLER_59_439 VPWR VGND sg13g2_decap_8
XFILLER_39_130 VPWR VGND sg13g2_decap_8
XFILLER_95_781 VPWR VGND sg13g2_decap_8
XFILLER_94_280 VPWR VGND sg13g2_decap_8
XFILLER_83_921 VPWR VGND sg13g2_decap_8
XFILLER_82_420 VPWR VGND sg13g2_decap_8
XFILLER_67_483 VPWR VGND sg13g2_decap_8
XFILLER_55_623 VPWR VGND sg13g2_decap_8
XFILLER_28_826 VPWR VGND sg13g2_decap_8
XFILLER_54_144 VPWR VGND sg13g2_decap_8
XFILLER_27_347 VPWR VGND sg13g2_decap_8
XFILLER_83_998 VPWR VGND sg13g2_decap_8
XFILLER_82_497 VPWR VGND sg13g2_decap_8
XFILLER_70_637 VPWR VGND sg13g2_decap_8
XFILLER_51_851 VPWR VGND sg13g2_decap_8
XFILLER_50_350 VPWR VGND sg13g2_decap_8
XFILLER_23_553 VPWR VGND sg13g2_decap_8
XFILLER_24_46 VPWR VGND sg13g2_decap_8
XFILLER_10_214 VPWR VGND sg13g2_decap_8
XFILLER_3_903 VPWR VGND sg13g2_decap_8
XFILLER_40_56 VPWR VGND sg13g2_decap_8
XFILLER_2_424 VPWR VGND sg13g2_decap_8
XFILLER_105_875 VPWR VGND sg13g2_decap_8
XFILLER_77_203 VPWR VGND sg13g2_decap_8
XFILLER_49_32 VPWR VGND sg13g2_decap_8
XFILLER_104_385 VPWR VGND sg13g2_decap_8
XFILLER_78_748 VPWR VGND sg13g2_decap_8
XFILLER_1_28 VPWR VGND sg13g2_decap_8
XFILLER_92_217 VPWR VGND sg13g2_decap_8
XFILLER_86_781 VPWR VGND sg13g2_decap_8
XFILLER_85_280 VPWR VGND sg13g2_decap_8
XFILLER_74_932 VPWR VGND sg13g2_decap_8
XFILLER_65_42 VPWR VGND sg13g2_decap_8
XFILLER_58_483 VPWR VGND sg13g2_decap_8
XFILLER_46_634 VPWR VGND sg13g2_decap_8
XFILLER_19_826 VPWR VGND sg13g2_decap_8
XFILLER_73_431 VPWR VGND sg13g2_decap_8
XFILLER_45_133 VPWR VGND sg13g2_decap_8
XFILLER_18_336 VPWR VGND sg13g2_decap_8
XFILLER_92_1022 VPWR VGND sg13g2_decap_8
XFILLER_61_648 VPWR VGND sg13g2_decap_8
XFILLER_60_158 VPWR VGND sg13g2_decap_8
XFILLER_42_851 VPWR VGND sg13g2_decap_8
XFILLER_14_553 VPWR VGND sg13g2_decap_8
XFILLER_41_350 VPWR VGND sg13g2_decap_8
XFILLER_81_74 VPWR VGND sg13g2_decap_8
XFILLER_10_781 VPWR VGND sg13g2_decap_8
XFILLER_60_7 VPWR VGND sg13g2_decap_8
XFILLER_6_763 VPWR VGND sg13g2_decap_8
XFILLER_5_284 VPWR VGND sg13g2_decap_8
XFILLER_69_715 VPWR VGND sg13g2_decap_8
XFILLER_39_4 VPWR VGND sg13g2_decap_8
XFILLER_68_236 VPWR VGND sg13g2_decap_8
XFILLER_2_991 VPWR VGND sg13g2_decap_8
XFILLER_96_567 VPWR VGND sg13g2_decap_8
XFILLER_84_707 VPWR VGND sg13g2_decap_8
XFILLER_65_910 VPWR VGND sg13g2_decap_8
XFILLER_1_490 VPWR VGND sg13g2_decap_8
XFILLER_83_228 VPWR VGND sg13g2_decap_8
XFILLER_77_770 VPWR VGND sg13g2_decap_8
Xinput5 ui_in[4] net5 VPWR VGND sg13g2_buf_1
XFILLER_49_494 VPWR VGND sg13g2_decap_8
XFILLER_37_634 VPWR VGND sg13g2_decap_8
XFILLER_76_291 VPWR VGND sg13g2_decap_8
XFILLER_64_431 VPWR VGND sg13g2_decap_8
XFILLER_36_133 VPWR VGND sg13g2_decap_8
XFILLER_92_784 VPWR VGND sg13g2_decap_8
XFILLER_80_924 VPWR VGND sg13g2_decap_8
XFILLER_65_987 VPWR VGND sg13g2_decap_8
XFILLER_91_294 VPWR VGND sg13g2_decap_8
XFILLER_52_637 VPWR VGND sg13g2_decap_8
XFILLER_33_840 VPWR VGND sg13g2_decap_8
XFILLER_51_158 VPWR VGND sg13g2_decap_8
XFILLER_20_501 VPWR VGND sg13g2_decap_8
XFILLER_32_361 VPWR VGND sg13g2_decap_8
XFILLER_20_578 VPWR VGND sg13g2_decap_8
XFILLER_69_1002 VPWR VGND sg13g2_decap_8
XFILLER_105_105 VPWR VGND sg13g2_decap_8
XFILLER_102_812 VPWR VGND sg13g2_decap_8
XFILLER_99_350 VPWR VGND sg13g2_decap_8
XFILLER_0_917 VPWR VGND sg13g2_decap_8
XFILLER_101_322 VPWR VGND sg13g2_decap_8
XFILLER_59_236 VPWR VGND sg13g2_decap_8
XFILLER_102_889 VPWR VGND sg13g2_decap_8
XFILLER_87_567 VPWR VGND sg13g2_decap_8
XFILLER_75_707 VPWR VGND sg13g2_decap_8
XFILLER_19_35 VPWR VGND sg13g2_decap_8
XFILLER_101_399 VPWR VGND sg13g2_decap_8
XFILLER_74_239 VPWR VGND sg13g2_decap_8
XFILLER_56_921 VPWR VGND sg13g2_decap_8
XFILLER_28_623 VPWR VGND sg13g2_decap_8
XFILLER_67_280 VPWR VGND sg13g2_decap_8
XFILLER_55_420 VPWR VGND sg13g2_decap_8
XFILLER_27_144 VPWR VGND sg13g2_decap_8
XFILLER_83_795 VPWR VGND sg13g2_decap_8
XFILLER_76_1028 VPWR VGND sg13g2_fill_1
XFILLER_71_935 VPWR VGND sg13g2_decap_8
XFILLER_56_998 VPWR VGND sg13g2_decap_8
XFILLER_82_294 VPWR VGND sg13g2_decap_8
XFILLER_70_434 VPWR VGND sg13g2_decap_8
XFILLER_55_497 VPWR VGND sg13g2_decap_8
XFILLER_43_637 VPWR VGND sg13g2_decap_8
XFILLER_35_56 VPWR VGND sg13g2_decap_8
XFILLER_42_158 VPWR VGND sg13g2_decap_8
XFILLER_23_350 VPWR VGND sg13g2_decap_8
XFILLER_24_851 VPWR VGND sg13g2_decap_8
XFILLER_51_11 VPWR VGND sg13g2_decap_8
XFILLER_11_567 VPWR VGND sg13g2_decap_8
XFILLER_13_1001 VPWR VGND sg13g2_decap_8
XFILLER_51_88 VPWR VGND sg13g2_decap_8
XFILLER_100_1015 VPWR VGND sg13g2_decap_8
XFILLER_3_700 VPWR VGND sg13g2_decap_8
XFILLER_2_221 VPWR VGND sg13g2_decap_8
XFILLER_105_672 VPWR VGND sg13g2_decap_8
XFILLER_3_777 VPWR VGND sg13g2_decap_8
XFILLER_104_182 VPWR VGND sg13g2_decap_8
XFILLER_78_545 VPWR VGND sg13g2_decap_8
XFILLER_2_298 VPWR VGND sg13g2_decap_8
XFILLER_93_537 VPWR VGND sg13g2_decap_8
XFILLER_76_74 VPWR VGND sg13g2_decap_8
XFILLER_65_217 VPWR VGND sg13g2_decap_8
XFILLER_47_910 VPWR VGND sg13g2_decap_8
XFILLER_19_623 VPWR VGND sg13g2_decap_8
XFILLER_58_280 VPWR VGND sg13g2_decap_8
XFILLER_46_431 VPWR VGND sg13g2_decap_8
XFILLER_18_133 VPWR VGND sg13g2_decap_8
XFILLER_20_1005 VPWR VGND sg13g2_decap_8
XFILLER_62_924 VPWR VGND sg13g2_decap_8
XFILLER_47_987 VPWR VGND sg13g2_decap_8
XFILLER_61_445 VPWR VGND sg13g2_decap_8
XFILLER_34_648 VPWR VGND sg13g2_decap_8
XFILLER_92_84 VPWR VGND sg13g2_decap_8
XFILLER_14_350 VPWR VGND sg13g2_decap_8
XFILLER_15_851 VPWR VGND sg13g2_decap_8
XFILLER_33_147 VPWR VGND sg13g2_decap_8
XFILLER_30_854 VPWR VGND sg13g2_decap_8
XFILLER_6_560 VPWR VGND sg13g2_decap_8
XFILLER_103_609 VPWR VGND sg13g2_decap_8
XFILLER_102_119 VPWR VGND sg13g2_decap_8
XFILLER_97_854 VPWR VGND sg13g2_decap_8
XFILLER_69_512 VPWR VGND sg13g2_decap_8
XFILLER_96_364 VPWR VGND sg13g2_decap_8
XFILLER_84_504 VPWR VGND sg13g2_decap_8
XFILLER_57_707 VPWR VGND sg13g2_decap_8
XFILLER_69_589 VPWR VGND sg13g2_decap_8
XFILLER_56_228 VPWR VGND sg13g2_decap_8
XFILLER_2_60 VPWR VGND sg13g2_decap_8
XFILLER_38_910 VPWR VGND sg13g2_decap_8
XFILLER_49_291 VPWR VGND sg13g2_decap_8
XFILLER_37_431 VPWR VGND sg13g2_decap_8
X_59_ net7 net15 _25_ VPWR VGND sg13g2_nor2_1
XFILLER_65_784 VPWR VGND sg13g2_decap_8
XFILLER_53_924 VPWR VGND sg13g2_decap_8
XFILLER_38_987 VPWR VGND sg13g2_decap_8
XFILLER_92_581 VPWR VGND sg13g2_decap_8
XFILLER_80_721 VPWR VGND sg13g2_decap_8
XFILLER_52_434 VPWR VGND sg13g2_decap_8
XFILLER_25_637 VPWR VGND sg13g2_decap_8
XFILLER_24_158 VPWR VGND sg13g2_decap_8
XFILLER_36_1001 VPWR VGND sg13g2_decap_8
XFILLER_80_798 VPWR VGND sg13g2_decap_8
XFILLER_21_854 VPWR VGND sg13g2_decap_8
XFILLER_20_375 VPWR VGND sg13g2_decap_8
XFILLER_21_14 VPWR VGND sg13g2_decap_8
XFILLER_106_469 VPWR VGND sg13g2_decap_8
XFILLER_0_714 VPWR VGND sg13g2_decap_8
XFILLER_88_865 VPWR VGND sg13g2_decap_8
XFILLER_87_364 VPWR VGND sg13g2_decap_8
XFILLER_75_504 VPWR VGND sg13g2_decap_8
XFILLER_48_707 VPWR VGND sg13g2_decap_8
XFILLER_102_686 VPWR VGND sg13g2_decap_8
XFILLER_47_217 VPWR VGND sg13g2_decap_8
XFILLER_29_921 VPWR VGND sg13g2_decap_8
XFILLER_101_196 VPWR VGND sg13g2_decap_8
XFILLER_46_11 VPWR VGND sg13g2_decap_8
XFILLER_28_420 VPWR VGND sg13g2_decap_8
XFILLER_90_529 VPWR VGND sg13g2_decap_8
XFILLER_29_998 VPWR VGND sg13g2_decap_8
XFILLER_83_592 VPWR VGND sg13g2_decap_8
XFILLER_71_732 VPWR VGND sg13g2_decap_8
XFILLER_56_795 VPWR VGND sg13g2_decap_8
XFILLER_55_294 VPWR VGND sg13g2_decap_8
XFILLER_46_88 VPWR VGND sg13g2_decap_8
XFILLER_44_935 VPWR VGND sg13g2_decap_8
XFILLER_43_434 VPWR VGND sg13g2_decap_8
XFILLER_16_637 VPWR VGND sg13g2_decap_8
XFILLER_28_497 VPWR VGND sg13g2_decap_8
XFILLER_70_231 VPWR VGND sg13g2_decap_8
XFILLER_62_21 VPWR VGND sg13g2_decap_8
XFILLER_15_158 VPWR VGND sg13g2_decap_8
XFILLER_62_98 VPWR VGND sg13g2_decap_8
XFILLER_62_76 VPWR VGND sg13g2_decap_8
XFILLER_12_865 VPWR VGND sg13g2_decap_8
XFILLER_8_847 VPWR VGND sg13g2_decap_8
XFILLER_11_364 VPWR VGND sg13g2_decap_8
XFILLER_7_368 VPWR VGND sg13g2_decap_8
XFILLER_11_91 VPWR VGND sg13g2_decap_8
XFILLER_3_574 VPWR VGND sg13g2_decap_8
XFILLER_87_84 VPWR VGND sg13g2_decap_8
XFILLER_79_865 VPWR VGND sg13g2_decap_8
XFILLER_78_342 VPWR VGND sg13g2_decap_8
XFILLER_23_7 VPWR VGND sg13g2_decap_8
XFILLER_39_718 VPWR VGND sg13g2_decap_8
XFILLER_38_217 VPWR VGND sg13g2_decap_8
XFILLER_94_868 VPWR VGND sg13g2_decap_8
XFILLER_93_334 VPWR VGND sg13g2_decap_8
XFILLER_66_559 VPWR VGND sg13g2_decap_8
XFILLER_19_420 VPWR VGND sg13g2_decap_8
XFILLER_81_529 VPWR VGND sg13g2_decap_8
XFILLER_47_784 VPWR VGND sg13g2_decap_8
XFILLER_35_924 VPWR VGND sg13g2_decap_8
XFILLER_62_721 VPWR VGND sg13g2_decap_8
XFILLER_19_497 VPWR VGND sg13g2_decap_8
XFILLER_61_242 VPWR VGND sg13g2_decap_8
XFILLER_34_445 VPWR VGND sg13g2_decap_8
XFILLER_62_798 VPWR VGND sg13g2_decap_8
XFILLER_50_938 VPWR VGND sg13g2_decap_8
XFILLER_30_651 VPWR VGND sg13g2_decap_8
XFILLER_103_406 VPWR VGND sg13g2_decap_8
XFILLER_97_651 VPWR VGND sg13g2_decap_8
XFILLER_96_161 VPWR VGND sg13g2_decap_8
XFILLER_84_301 VPWR VGND sg13g2_decap_8
XFILLER_69_386 VPWR VGND sg13g2_decap_8
XFILLER_57_504 VPWR VGND sg13g2_decap_8
XFILLER_85_868 VPWR VGND sg13g2_decap_8
XFILLER_29_228 VPWR VGND sg13g2_decap_8
XFILLER_84_378 VPWR VGND sg13g2_decap_8
XFILLER_72_518 VPWR VGND sg13g2_decap_8
XFILLER_26_924 VPWR VGND sg13g2_decap_8
XFILLER_38_784 VPWR VGND sg13g2_decap_8
XFILLER_65_581 VPWR VGND sg13g2_decap_8
XFILLER_53_721 VPWR VGND sg13g2_decap_8
XFILLER_16_14 VPWR VGND sg13g2_decap_8
XFILLER_25_434 VPWR VGND sg13g2_decap_8
XFILLER_52_231 VPWR VGND sg13g2_decap_8
XFILLER_80_595 VPWR VGND sg13g2_decap_8
XFILLER_53_798 VPWR VGND sg13g2_decap_8
XFILLER_41_938 VPWR VGND sg13g2_decap_8
XFILLER_40_448 VPWR VGND sg13g2_decap_8
XFILLER_21_651 VPWR VGND sg13g2_decap_8
XFILLER_32_46 VPWR VGND sg13g2_decap_8
XFILLER_20_172 VPWR VGND sg13g2_decap_8
XFILLER_10_1026 VPWR VGND sg13g2_fill_2
XFILLER_106_266 VPWR VGND sg13g2_decap_8
XFILLER_0_511 VPWR VGND sg13g2_decap_8
XFILLER_88_662 VPWR VGND sg13g2_decap_8
XFILLER_76_802 VPWR VGND sg13g2_decap_8
XFILLER_103_973 VPWR VGND sg13g2_decap_8
XFILLER_87_161 VPWR VGND sg13g2_decap_8
XFILLER_75_301 VPWR VGND sg13g2_decap_8
XFILLER_57_21 VPWR VGND sg13g2_decap_8
XFILLER_48_504 VPWR VGND sg13g2_decap_8
XFILLER_0_588 VPWR VGND sg13g2_decap_8
XFILLER_102_483 VPWR VGND sg13g2_decap_8
XFILLER_91_805 VPWR VGND sg13g2_decap_8
XFILLER_76_879 VPWR VGND sg13g2_decap_8
XFILLER_75_378 VPWR VGND sg13g2_decap_8
XFILLER_63_518 VPWR VGND sg13g2_decap_8
XFILLER_57_98 VPWR VGND sg13g2_decap_8
XFILLER_90_326 VPWR VGND sg13g2_decap_8
XFILLER_56_592 VPWR VGND sg13g2_decap_8
XFILLER_44_732 VPWR VGND sg13g2_decap_8
XFILLER_17_935 VPWR VGND sg13g2_decap_8
XFILLER_29_795 VPWR VGND sg13g2_decap_8
XFILLER_73_53 VPWR VGND sg13g2_decap_4
XFILLER_43_231 VPWR VGND sg13g2_decap_8
XFILLER_16_434 VPWR VGND sg13g2_decap_8
XFILLER_28_294 VPWR VGND sg13g2_decap_8
XFILLER_32_949 VPWR VGND sg13g2_decap_8
XFILLER_31_448 VPWR VGND sg13g2_decap_8
XFILLER_12_662 VPWR VGND sg13g2_decap_8
XFILLER_8_644 VPWR VGND sg13g2_decap_8
XFILLER_11_161 VPWR VGND sg13g2_decap_8
XFILLER_7_165 VPWR VGND sg13g2_decap_8
XFILLER_99_938 VPWR VGND sg13g2_decap_8
XFILLER_4_861 VPWR VGND sg13g2_decap_8
XFILLER_3_371 VPWR VGND sg13g2_decap_8
XFILLER_98_459 VPWR VGND sg13g2_decap_8
XFILLER_26_1022 VPWR VGND sg13g2_decap_8
XFILLER_79_662 VPWR VGND sg13g2_decap_8
XFILLER_39_515 VPWR VGND sg13g2_decap_8
XFILLER_93_131 VPWR VGND sg13g2_decap_8
XFILLER_67_868 VPWR VGND sg13g2_decap_8
XFILLER_94_665 VPWR VGND sg13g2_decap_8
XFILLER_82_805 VPWR VGND sg13g2_decap_8
XFILLER_66_356 VPWR VGND sg13g2_decap_8
XFILLER_81_326 VPWR VGND sg13g2_decap_8
XFILLER_54_529 VPWR VGND sg13g2_decap_8
XFILLER_47_581 VPWR VGND sg13g2_decap_8
XFILLER_35_721 VPWR VGND sg13g2_decap_8
XFILLER_19_294 VPWR VGND sg13g2_decap_8
XFILLER_34_242 VPWR VGND sg13g2_decap_8
XFILLER_90_893 VPWR VGND sg13g2_decap_8
XFILLER_50_735 VPWR VGND sg13g2_decap_8
XFILLER_23_938 VPWR VGND sg13g2_decap_8
XFILLER_35_798 VPWR VGND sg13g2_decap_8
XFILLER_97_0 VPWR VGND sg13g2_decap_8
XFILLER_62_595 VPWR VGND sg13g2_decap_8
XFILLER_22_459 VPWR VGND sg13g2_decap_8
XFILLER_33_1015 VPWR VGND sg13g2_decap_8
XFILLER_8_70 VPWR VGND sg13g2_decap_8
XFILLER_2_809 VPWR VGND sg13g2_decap_8
XFILLER_103_203 VPWR VGND sg13g2_decap_8
XFILLER_1_308 VPWR VGND sg13g2_decap_8
XFILLER_89_448 VPWR VGND sg13g2_decap_8
XFILLER_100_910 VPWR VGND sg13g2_decap_8
XFILLER_76_109 VPWR VGND sg13g2_decap_8
XFILLER_57_301 VPWR VGND sg13g2_decap_8
XFILLER_69_183 VPWR VGND sg13g2_decap_8
XFILLER_58_868 VPWR VGND sg13g2_decap_8
XFILLER_40_1008 VPWR VGND sg13g2_decap_8
XFILLER_100_987 VPWR VGND sg13g2_decap_8
XFILLER_85_665 VPWR VGND sg13g2_decap_8
XFILLER_73_816 VPWR VGND sg13g2_decap_8
XFILLER_57_378 VPWR VGND sg13g2_decap_8
XFILLER_45_518 VPWR VGND sg13g2_decap_8
XFILLER_84_175 VPWR VGND sg13g2_decap_8
XFILLER_72_315 VPWR VGND sg13g2_decap_8
XFILLER_26_721 VPWR VGND sg13g2_decap_8
XFILLER_27_46 VPWR VGND sg13g2_decap_8
XFILLER_38_581 VPWR VGND sg13g2_decap_8
XFILLER_25_231 VPWR VGND sg13g2_decap_8
XFILLER_81_893 VPWR VGND sg13g2_decap_8
XFILLER_14_938 VPWR VGND sg13g2_decap_8
XFILLER_26_798 VPWR VGND sg13g2_decap_8
XFILLER_80_392 VPWR VGND sg13g2_decap_8
XFILLER_53_595 VPWR VGND sg13g2_decap_8
XFILLER_43_56 VPWR VGND sg13g2_decap_8
XFILLER_41_735 VPWR VGND sg13g2_decap_8
XFILLER_13_448 VPWR VGND sg13g2_decap_8
XFILLER_40_245 VPWR VGND sg13g2_decap_8
XFILLER_5_669 VPWR VGND sg13g2_decap_8
XFILLER_4_168 VPWR VGND sg13g2_decap_8
XFILLER_4_28 VPWR VGND sg13g2_decap_8
XFILLER_103_770 VPWR VGND sg13g2_decap_8
XFILLER_68_75 VPWR VGND sg13g2_decap_8
XFILLER_49_802 VPWR VGND sg13g2_decap_8
XFILLER_48_301 VPWR VGND sg13g2_decap_8
XFILLER_1_875 VPWR VGND sg13g2_decap_8
XFILLER_102_280 VPWR VGND sg13g2_decap_8
XFILLER_0_385 VPWR VGND sg13g2_decap_8
XFILLER_91_602 VPWR VGND sg13g2_decap_8
XFILLER_76_676 VPWR VGND sg13g2_decap_8
XFILLER_64_816 VPWR VGND sg13g2_decap_8
XFILLER_49_879 VPWR VGND sg13g2_decap_8
XFILLER_48_378 VPWR VGND sg13g2_decap_8
XFILLER_36_518 VPWR VGND sg13g2_decap_8
XFILLER_90_123 VPWR VGND sg13g2_decap_8
XFILLER_84_63 VPWR VGND sg13g2_decap_8
XFILLER_75_175 VPWR VGND sg13g2_decap_8
XFILLER_63_315 VPWR VGND sg13g2_decap_8
XFILLER_17_732 VPWR VGND sg13g2_decap_8
XFILLER_91_679 VPWR VGND sg13g2_decap_8
XFILLER_16_231 VPWR VGND sg13g2_decap_8
XFILLER_29_592 VPWR VGND sg13g2_decap_8
XFILLER_72_882 VPWR VGND sg13g2_decap_8
XFILLER_56_1026 VPWR VGND sg13g2_fill_2
XFILLER_32_746 VPWR VGND sg13g2_decap_8
XFILLER_31_245 VPWR VGND sg13g2_decap_8
XFILLER_9_931 VPWR VGND sg13g2_decap_8
XFILLER_8_441 VPWR VGND sg13g2_decap_8
XFILLER_99_735 VPWR VGND sg13g2_decap_8
XFILLER_101_707 VPWR VGND sg13g2_decap_8
XFILLER_98_256 VPWR VGND sg13g2_decap_8
XFILLER_63_1008 VPWR VGND sg13g2_decap_8
XFILLER_100_217 VPWR VGND sg13g2_decap_8
XFILLER_39_312 VPWR VGND sg13g2_decap_8
XFILLER_95_963 VPWR VGND sg13g2_decap_8
XFILLER_94_462 VPWR VGND sg13g2_decap_8
XFILLER_82_602 VPWR VGND sg13g2_decap_8
XFILLER_67_665 VPWR VGND sg13g2_decap_8
XFILLER_66_153 VPWR VGND sg13g2_decap_8
XFILLER_55_805 VPWR VGND sg13g2_decap_8
XFILLER_54_326 VPWR VGND sg13g2_decap_8
XFILLER_27_529 VPWR VGND sg13g2_decap_8
XFILLER_39_389 VPWR VGND sg13g2_decap_8
XFILLER_82_679 VPWR VGND sg13g2_decap_8
XFILLER_81_123 VPWR VGND sg13g2_decap_8
XFILLER_70_819 VPWR VGND sg13g2_decap_8
XFILLER_63_882 VPWR VGND sg13g2_decap_8
XFILLER_90_690 VPWR VGND sg13g2_decap_8
XFILLER_62_392 VPWR VGND sg13g2_decap_8
XFILLER_50_532 VPWR VGND sg13g2_decap_8
XFILLER_23_735 VPWR VGND sg13g2_decap_8
XFILLER_35_595 VPWR VGND sg13g2_decap_8
XFILLER_22_256 VPWR VGND sg13g2_decap_8
XFILLER_2_606 VPWR VGND sg13g2_decap_8
XFILLER_1_105 VPWR VGND sg13g2_decap_8
XFILLER_89_245 VPWR VGND sg13g2_decap_8
XFILLER_104_567 VPWR VGND sg13g2_decap_8
XFILLER_49_109 VPWR VGND sg13g2_decap_8
XFILLER_86_963 VPWR VGND sg13g2_decap_8
XFILLER_85_462 VPWR VGND sg13g2_decap_8
XFILLER_58_665 VPWR VGND sg13g2_decap_8
XFILLER_46_816 VPWR VGND sg13g2_decap_8
XFILLER_38_56 VPWR VGND sg13g2_decap_8
XFILLER_100_784 VPWR VGND sg13g2_decap_8
XFILLER_79_1026 VPWR VGND sg13g2_fill_2
XFILLER_73_613 VPWR VGND sg13g2_decap_8
XFILLER_72_112 VPWR VGND sg13g2_decap_8
XFILLER_57_175 VPWR VGND sg13g2_decap_8
XFILLER_45_315 VPWR VGND sg13g2_decap_8
XFILLER_18_518 VPWR VGND sg13g2_decap_8
XFILLER_54_11 VPWR VGND sg13g2_decap_8
XFILLER_72_189 VPWR VGND sg13g2_decap_8
XFILLER_81_690 VPWR VGND sg13g2_decap_8
XFILLER_54_893 VPWR VGND sg13g2_decap_8
XFILLER_54_88 VPWR VGND sg13g2_decap_8
XFILLER_53_392 VPWR VGND sg13g2_decap_8
XFILLER_14_735 VPWR VGND sg13g2_decap_8
XFILLER_26_595 VPWR VGND sg13g2_decap_8
XFILLER_41_532 VPWR VGND sg13g2_decap_8
XFILLER_13_245 VPWR VGND sg13g2_decap_8
XFILLER_70_21 VPWR VGND sg13g2_decap_8
XFILLER_9_238 VPWR VGND sg13g2_decap_8
XFILLER_10_963 VPWR VGND sg13g2_decap_8
XFILLER_70_98 VPWR VGND sg13g2_decap_8
XFILLER_6_945 VPWR VGND sg13g2_decap_8
XFILLER_86_1019 VPWR VGND sg13g2_decap_8
XFILLER_5_466 VPWR VGND sg13g2_decap_8
XFILLER_79_74 VPWR VGND sg13g2_decap_8
XFILLER_68_418 VPWR VGND sg13g2_decap_8
XFILLER_96_749 VPWR VGND sg13g2_decap_8
XFILLER_77_952 VPWR VGND sg13g2_decap_8
XFILLER_1_672 VPWR VGND sg13g2_decap_8
XFILLER_49_676 VPWR VGND sg13g2_decap_8
XFILLER_0_182 VPWR VGND sg13g2_decap_8
XFILLER_37_816 VPWR VGND sg13g2_decap_8
XFILLER_95_95 VPWR VGND sg13g2_decap_8
XFILLER_76_473 VPWR VGND sg13g2_decap_8
XFILLER_64_613 VPWR VGND sg13g2_decap_8
XFILLER_63_112 VPWR VGND sg13g2_decap_8
XFILLER_48_175 VPWR VGND sg13g2_decap_8
XFILLER_36_315 VPWR VGND sg13g2_decap_8
XFILLER_92_966 VPWR VGND sg13g2_decap_8
XFILLER_52_819 VPWR VGND sg13g2_decap_8
XFILLER_91_476 VPWR VGND sg13g2_decap_8
XFILLER_45_882 VPWR VGND sg13g2_decap_8
XFILLER_63_189 VPWR VGND sg13g2_decap_8
XFILLER_60_830 VPWR VGND sg13g2_decap_8
XFILLER_32_543 VPWR VGND sg13g2_decap_8
XFILLER_99_532 VPWR VGND sg13g2_decap_8
XFILLER_5_60 VPWR VGND sg13g2_decap_8
XFILLER_101_504 VPWR VGND sg13g2_decap_8
XFILLER_59_418 VPWR VGND sg13g2_decap_8
XFILLER_8_1008 VPWR VGND sg13g2_decap_8
XFILLER_87_749 VPWR VGND sg13g2_decap_8
XFILLER_95_760 VPWR VGND sg13g2_decap_8
XFILLER_83_900 VPWR VGND sg13g2_decap_8
XFILLER_68_985 VPWR VGND sg13g2_decap_8
XFILLER_55_602 VPWR VGND sg13g2_decap_8
XFILLER_28_805 VPWR VGND sg13g2_decap_8
XFILLER_67_462 VPWR VGND sg13g2_decap_8
XFILLER_27_326 VPWR VGND sg13g2_decap_8
XFILLER_39_186 VPWR VGND sg13g2_decap_8
XFILLER_83_977 VPWR VGND sg13g2_decap_8
XFILLER_54_123 VPWR VGND sg13g2_decap_8
XFILLER_82_476 VPWR VGND sg13g2_decap_8
XFILLER_70_616 VPWR VGND sg13g2_decap_8
XFILLER_55_679 VPWR VGND sg13g2_decap_8
XFILLER_43_819 VPWR VGND sg13g2_decap_8
XFILLER_36_882 VPWR VGND sg13g2_decap_8
XFILLER_51_830 VPWR VGND sg13g2_decap_8
XFILLER_23_532 VPWR VGND sg13g2_decap_8
XFILLER_35_392 VPWR VGND sg13g2_decap_8
XFILLER_24_25 VPWR VGND sg13g2_decap_8
XFILLER_11_749 VPWR VGND sg13g2_decap_8
XFILLER_40_35 VPWR VGND sg13g2_decap_8
XFILLER_2_403 VPWR VGND sg13g2_decap_8
XFILLER_105_854 VPWR VGND sg13g2_decap_8
XFILLER_49_11 VPWR VGND sg13g2_decap_8
XFILLER_3_959 VPWR VGND sg13g2_decap_8
XFILLER_104_364 VPWR VGND sg13g2_decap_8
XFILLER_78_727 VPWR VGND sg13g2_decap_8
XFILLER_49_88 VPWR VGND sg13g2_decap_8
XFILLER_93_719 VPWR VGND sg13g2_decap_8
XFILLER_86_760 VPWR VGND sg13g2_decap_8
XFILLER_77_259 VPWR VGND sg13g2_decap_8
XFILLER_19_805 VPWR VGND sg13g2_decap_8
XFILLER_100_581 VPWR VGND sg13g2_decap_8
XFILLER_74_911 VPWR VGND sg13g2_decap_8
XFILLER_73_410 VPWR VGND sg13g2_decap_8
XFILLER_65_21 VPWR VGND sg13g2_decap_8
XFILLER_59_985 VPWR VGND sg13g2_decap_8
XFILLER_58_462 VPWR VGND sg13g2_decap_8
XFILLER_46_613 VPWR VGND sg13g2_decap_8
XFILLER_18_315 VPWR VGND sg13g2_decap_8
XFILLER_45_112 VPWR VGND sg13g2_decap_8
XFILLER_74_988 VPWR VGND sg13g2_decap_8
XFILLER_73_487 VPWR VGND sg13g2_decap_8
XFILLER_65_98 VPWR VGND sg13g2_decap_8
XFILLER_61_627 VPWR VGND sg13g2_decap_8
XFILLER_92_1001 VPWR VGND sg13g2_decap_8
XFILLER_54_690 VPWR VGND sg13g2_decap_8
XFILLER_45_189 VPWR VGND sg13g2_decap_8
XFILLER_42_830 VPWR VGND sg13g2_decap_8
XFILLER_14_532 VPWR VGND sg13g2_decap_8
XFILLER_26_392 VPWR VGND sg13g2_decap_8
XFILLER_27_893 VPWR VGND sg13g2_decap_8
XFILLER_33_329 VPWR VGND sg13g2_decap_8
XFILLER_81_53 VPWR VGND sg13g2_decap_8
XFILLER_10_760 VPWR VGND sg13g2_decap_8
XFILLER_14_91 VPWR VGND sg13g2_decap_8
XFILLER_6_742 VPWR VGND sg13g2_decap_8
XFILLER_53_7 VPWR VGND sg13g2_decap_8
XFILLER_5_263 VPWR VGND sg13g2_decap_8
XFILLER_2_970 VPWR VGND sg13g2_decap_8
XFILLER_96_546 VPWR VGND sg13g2_decap_8
XFILLER_68_215 VPWR VGND sg13g2_decap_8
XFILLER_83_207 VPWR VGND sg13g2_decap_8
XFILLER_76_270 VPWR VGND sg13g2_decap_8
Xinput6 ui_in[5] net6 VPWR VGND sg13g2_buf_1
XFILLER_64_410 VPWR VGND sg13g2_decap_8
XFILLER_49_473 VPWR VGND sg13g2_decap_8
XFILLER_37_613 VPWR VGND sg13g2_decap_8
XFILLER_65_966 VPWR VGND sg13g2_decap_8
XFILLER_36_112 VPWR VGND sg13g2_decap_8
XFILLER_92_763 VPWR VGND sg13g2_decap_8
XFILLER_80_903 VPWR VGND sg13g2_decap_8
XFILLER_64_487 VPWR VGND sg13g2_decap_8
XFILLER_52_616 VPWR VGND sg13g2_decap_8
XFILLER_25_819 VPWR VGND sg13g2_decap_8
XFILLER_91_273 VPWR VGND sg13g2_decap_8
XFILLER_51_137 VPWR VGND sg13g2_decap_8
XFILLER_18_882 VPWR VGND sg13g2_decap_8
XFILLER_36_189 VPWR VGND sg13g2_decap_8
XFILLER_32_340 VPWR VGND sg13g2_decap_8
XFILLER_33_896 VPWR VGND sg13g2_decap_8
XFILLER_20_557 VPWR VGND sg13g2_decap_8
XFILLER_101_301 VPWR VGND sg13g2_decap_8
XFILLER_87_546 VPWR VGND sg13g2_decap_8
XFILLER_59_215 VPWR VGND sg13g2_decap_8
XFILLER_102_868 VPWR VGND sg13g2_decap_8
XFILLER_56_900 VPWR VGND sg13g2_decap_8
XFILLER_19_14 VPWR VGND sg13g2_decap_8
XFILLER_101_378 VPWR VGND sg13g2_decap_8
XFILLER_74_218 VPWR VGND sg13g2_decap_8
XFILLER_68_782 VPWR VGND sg13g2_decap_8
XFILLER_28_602 VPWR VGND sg13g2_decap_8
XFILLER_27_123 VPWR VGND sg13g2_decap_8
XFILLER_83_774 VPWR VGND sg13g2_decap_8
XFILLER_71_914 VPWR VGND sg13g2_decap_8
XFILLER_56_977 VPWR VGND sg13g2_decap_8
XFILLER_55_476 VPWR VGND sg13g2_decap_8
XFILLER_43_616 VPWR VGND sg13g2_decap_8
XFILLER_16_819 VPWR VGND sg13g2_decap_8
XFILLER_28_679 VPWR VGND sg13g2_decap_8
XFILLER_82_273 VPWR VGND sg13g2_decap_8
XFILLER_70_413 VPWR VGND sg13g2_decap_8
XFILLER_24_830 VPWR VGND sg13g2_decap_8
XFILLER_35_35 VPWR VGND sg13g2_decap_8
XFILLER_42_137 VPWR VGND sg13g2_decap_8
XFILLER_11_546 VPWR VGND sg13g2_decap_8
XFILLER_51_67 VPWR VGND sg13g2_decap_8
XFILLER_2_200 VPWR VGND sg13g2_decap_8
XFILLER_105_651 VPWR VGND sg13g2_decap_8
XFILLER_3_756 VPWR VGND sg13g2_decap_8
XFILLER_104_161 VPWR VGND sg13g2_decap_8
XFILLER_78_524 VPWR VGND sg13g2_decap_8
XFILLER_2_277 VPWR VGND sg13g2_decap_8
XFILLER_93_516 VPWR VGND sg13g2_decap_8
XFILLER_76_53 VPWR VGND sg13g2_decap_8
XFILLER_59_782 VPWR VGND sg13g2_decap_8
XFILLER_19_602 VPWR VGND sg13g2_decap_8
XFILLER_47_966 VPWR VGND sg13g2_decap_8
XFILLER_46_410 VPWR VGND sg13g2_decap_8
XFILLER_18_112 VPWR VGND sg13g2_decap_8
XFILLER_20_1028 VPWR VGND sg13g2_fill_1
XFILLER_74_785 VPWR VGND sg13g2_decap_8
XFILLER_62_903 VPWR VGND sg13g2_decap_8
XFILLER_19_679 VPWR VGND sg13g2_decap_8
XFILLER_92_63 VPWR VGND sg13g2_decap_8
XFILLER_73_284 VPWR VGND sg13g2_decap_8
XFILLER_61_424 VPWR VGND sg13g2_decap_8
XFILLER_46_487 VPWR VGND sg13g2_decap_8
XFILLER_15_830 VPWR VGND sg13g2_decap_8
XFILLER_18_189 VPWR VGND sg13g2_decap_8
XFILLER_27_690 VPWR VGND sg13g2_decap_8
XFILLER_33_126 VPWR VGND sg13g2_decap_8
XFILLER_34_627 VPWR VGND sg13g2_decap_8
XFILLER_70_980 VPWR VGND sg13g2_decap_8
XFILLER_30_833 VPWR VGND sg13g2_decap_8
XFILLER_51_4 VPWR VGND sg13g2_decap_8
XFILLER_97_833 VPWR VGND sg13g2_decap_8
XFILLER_96_343 VPWR VGND sg13g2_decap_8
XFILLER_69_568 VPWR VGND sg13g2_decap_8
XFILLER_56_207 VPWR VGND sg13g2_decap_8
XFILLER_49_270 VPWR VGND sg13g2_decap_8
XFILLER_37_410 VPWR VGND sg13g2_decap_8
XFILLER_38_966 VPWR VGND sg13g2_decap_8
XFILLER_92_560 VPWR VGND sg13g2_decap_8
XFILLER_80_700 VPWR VGND sg13g2_decap_8
X_58_ _24_ net7 net15 VPWR VGND sg13g2_nand2_1
XFILLER_65_763 VPWR VGND sg13g2_decap_8
XFILLER_53_903 VPWR VGND sg13g2_decap_8
XFILLER_25_616 VPWR VGND sg13g2_decap_8
XFILLER_64_284 VPWR VGND sg13g2_decap_8
XFILLER_52_413 VPWR VGND sg13g2_decap_8
XFILLER_37_487 VPWR VGND sg13g2_decap_8
XFILLER_80_777 VPWR VGND sg13g2_decap_8
XFILLER_24_137 VPWR VGND sg13g2_decap_8
XFILLER_61_991 VPWR VGND sg13g2_decap_8
XFILLER_21_833 VPWR VGND sg13g2_decap_8
XFILLER_33_693 VPWR VGND sg13g2_decap_8
XFILLER_20_354 VPWR VGND sg13g2_decap_8
XFILLER_106_448 VPWR VGND sg13g2_decap_8
XFILLER_88_844 VPWR VGND sg13g2_decap_8
XFILLER_82_1022 VPWR VGND sg13g2_decap_8
XFILLER_87_343 VPWR VGND sg13g2_decap_8
XFILLER_102_665 VPWR VGND sg13g2_decap_8
XFILLER_29_900 VPWR VGND sg13g2_decap_8
XFILLER_101_175 VPWR VGND sg13g2_decap_8
XFILLER_90_508 VPWR VGND sg13g2_decap_8
XFILLER_56_774 VPWR VGND sg13g2_decap_8
XFILLER_46_67 VPWR VGND sg13g2_decap_8
XFILLER_44_914 VPWR VGND sg13g2_decap_8
XFILLER_16_616 VPWR VGND sg13g2_decap_8
XFILLER_28_476 VPWR VGND sg13g2_decap_8
XFILLER_29_977 VPWR VGND sg13g2_decap_8
XFILLER_83_571 VPWR VGND sg13g2_decap_8
XFILLER_71_711 VPWR VGND sg13g2_decap_8
XFILLER_70_210 VPWR VGND sg13g2_decap_8
XFILLER_55_273 VPWR VGND sg13g2_decap_8
XFILLER_43_413 VPWR VGND sg13g2_decap_8
XFILLER_15_137 VPWR VGND sg13g2_decap_8
XFILLER_102_84 VPWR VGND sg13g2_decap_8
XFILLER_71_788 VPWR VGND sg13g2_decap_8
XFILLER_70_287 VPWR VGND sg13g2_decap_8
XFILLER_52_980 VPWR VGND sg13g2_decap_8
XFILLER_12_844 VPWR VGND sg13g2_decap_8
XFILLER_8_826 VPWR VGND sg13g2_decap_8
XFILLER_11_343 VPWR VGND sg13g2_decap_8
XFILLER_7_347 VPWR VGND sg13g2_decap_8
XFILLER_7_39 VPWR VGND sg13g2_decap_8
XFILLER_3_553 VPWR VGND sg13g2_decap_8
XFILLER_11_70 VPWR VGND sg13g2_decap_8
XFILLER_79_844 VPWR VGND sg13g2_decap_8
XFILLER_87_63 VPWR VGND sg13g2_decap_8
XFILLER_78_321 VPWR VGND sg13g2_decap_8
XFILLER_93_313 VPWR VGND sg13g2_decap_8
XFILLER_94_847 VPWR VGND sg13g2_decap_8
XFILLER_78_398 VPWR VGND sg13g2_decap_8
XFILLER_66_538 VPWR VGND sg13g2_decap_8
XFILLER_4_1022 VPWR VGND sg13g2_decap_8
XFILLER_16_7 VPWR VGND sg13g2_decap_8
XFILLER_81_508 VPWR VGND sg13g2_decap_8
XFILLER_62_700 VPWR VGND sg13g2_decap_8
XFILLER_59_1013 VPWR VGND sg13g2_decap_8
XFILLER_47_763 VPWR VGND sg13g2_decap_8
XFILLER_35_903 VPWR VGND sg13g2_decap_8
XFILLER_74_582 VPWR VGND sg13g2_decap_8
XFILLER_46_284 VPWR VGND sg13g2_decap_8
XFILLER_19_476 VPWR VGND sg13g2_decap_8
XFILLER_34_424 VPWR VGND sg13g2_decap_8
XFILLER_62_777 VPWR VGND sg13g2_decap_8
XFILLER_61_221 VPWR VGND sg13g2_decap_8
XFILLER_50_917 VPWR VGND sg13g2_decap_8
XFILLER_43_980 VPWR VGND sg13g2_decap_8
XFILLER_61_298 VPWR VGND sg13g2_decap_8
XFILLER_30_630 VPWR VGND sg13g2_decap_8
XFILLER_66_1028 VPWR VGND sg13g2_fill_1
XFILLER_97_630 VPWR VGND sg13g2_decap_8
XFILLER_96_140 VPWR VGND sg13g2_decap_8
XFILLER_69_365 VPWR VGND sg13g2_decap_8
XFILLER_29_207 VPWR VGND sg13g2_decap_8
XFILLER_85_847 VPWR VGND sg13g2_decap_8
XFILLER_84_357 VPWR VGND sg13g2_decap_8
XFILLER_65_560 VPWR VGND sg13g2_decap_8
XFILLER_53_700 VPWR VGND sg13g2_decap_8
XFILLER_26_903 VPWR VGND sg13g2_decap_8
XFILLER_38_763 VPWR VGND sg13g2_decap_8
XFILLER_93_880 VPWR VGND sg13g2_decap_8
XFILLER_52_210 VPWR VGND sg13g2_decap_8
XFILLER_25_413 VPWR VGND sg13g2_decap_8
XFILLER_37_284 VPWR VGND sg13g2_decap_8
XFILLER_41_917 VPWR VGND sg13g2_decap_8
XFILLER_80_574 VPWR VGND sg13g2_decap_8
XFILLER_53_777 VPWR VGND sg13g2_decap_8
XFILLER_40_427 VPWR VGND sg13g2_decap_8
XFILLER_52_287 VPWR VGND sg13g2_decap_8
XFILLER_21_630 VPWR VGND sg13g2_decap_8
XFILLER_33_490 VPWR VGND sg13g2_decap_8
XFILLER_34_991 VPWR VGND sg13g2_decap_8
XFILLER_32_25 VPWR VGND sg13g2_decap_8
XFILLER_20_151 VPWR VGND sg13g2_decap_8
XFILLER_10_1005 VPWR VGND sg13g2_decap_8
XFILLER_106_245 VPWR VGND sg13g2_decap_8
XFILLER_103_952 VPWR VGND sg13g2_decap_8
XFILLER_88_641 VPWR VGND sg13g2_decap_8
XFILLER_102_462 VPWR VGND sg13g2_decap_8
XFILLER_87_140 VPWR VGND sg13g2_decap_8
XFILLER_0_567 VPWR VGND sg13g2_decap_8
XFILLER_76_858 VPWR VGND sg13g2_decap_8
XFILLER_57_77 VPWR VGND sg13g2_decap_8
XFILLER_90_305 VPWR VGND sg13g2_decap_8
XFILLER_75_357 VPWR VGND sg13g2_decap_8
XFILLER_17_914 VPWR VGND sg13g2_decap_8
XFILLER_29_774 VPWR VGND sg13g2_decap_8
XFILLER_56_571 VPWR VGND sg13g2_decap_8
XFILLER_44_711 VPWR VGND sg13g2_decap_8
XFILLER_43_210 VPWR VGND sg13g2_decap_8
XFILLER_16_413 VPWR VGND sg13g2_decap_8
XFILLER_28_273 VPWR VGND sg13g2_decap_8
XFILLER_73_32 VPWR VGND sg13g2_decap_8
XFILLER_71_585 VPWR VGND sg13g2_decap_8
XFILLER_44_788 VPWR VGND sg13g2_decap_8
XFILLER_25_980 VPWR VGND sg13g2_decap_8
XFILLER_32_928 VPWR VGND sg13g2_decap_8
XFILLER_43_287 VPWR VGND sg13g2_decap_8
XFILLER_31_427 VPWR VGND sg13g2_decap_8
XFILLER_106_1022 VPWR VGND sg13g2_decap_8
XFILLER_11_140 VPWR VGND sg13g2_decap_8
XFILLER_12_641 VPWR VGND sg13g2_decap_8
XFILLER_8_623 VPWR VGND sg13g2_decap_8
XFILLER_40_994 VPWR VGND sg13g2_decap_8
XFILLER_7_144 VPWR VGND sg13g2_decap_8
XFILLER_99_917 VPWR VGND sg13g2_decap_8
XFILLER_4_840 VPWR VGND sg13g2_decap_8
XFILLER_98_438 VPWR VGND sg13g2_decap_8
XFILLER_98_95 VPWR VGND sg13g2_decap_8
XFILLER_3_350 VPWR VGND sg13g2_decap_8
XFILLER_79_641 VPWR VGND sg13g2_decap_8
XFILLER_26_1001 VPWR VGND sg13g2_decap_8
XFILLER_94_644 VPWR VGND sg13g2_decap_8
XFILLER_93_110 VPWR VGND sg13g2_decap_8
XFILLER_78_195 VPWR VGND sg13g2_decap_8
XFILLER_67_847 VPWR VGND sg13g2_decap_8
XFILLER_66_335 VPWR VGND sg13g2_decap_8
XFILLER_81_305 VPWR VGND sg13g2_decap_8
XFILLER_54_508 VPWR VGND sg13g2_decap_8
XFILLER_93_187 VPWR VGND sg13g2_decap_8
XFILLER_47_560 VPWR VGND sg13g2_decap_8
XFILLER_19_273 VPWR VGND sg13g2_decap_8
XFILLER_35_700 VPWR VGND sg13g2_decap_8
XFILLER_34_221 VPWR VGND sg13g2_decap_8
XFILLER_90_872 VPWR VGND sg13g2_decap_8
XFILLER_62_574 VPWR VGND sg13g2_decap_8
XFILLER_50_714 VPWR VGND sg13g2_decap_8
XFILLER_16_980 VPWR VGND sg13g2_decap_8
XFILLER_23_917 VPWR VGND sg13g2_decap_8
XFILLER_35_777 VPWR VGND sg13g2_decap_8
XFILLER_22_438 VPWR VGND sg13g2_decap_8
XFILLER_34_298 VPWR VGND sg13g2_decap_8
XFILLER_31_994 VPWR VGND sg13g2_decap_8
XFILLER_89_427 VPWR VGND sg13g2_decap_8
XFILLER_104_749 VPWR VGND sg13g2_decap_8
XFILLER_103_259 VPWR VGND sg13g2_decap_8
XFILLER_69_162 VPWR VGND sg13g2_decap_8
XFILLER_85_644 VPWR VGND sg13g2_decap_8
XFILLER_58_847 VPWR VGND sg13g2_decap_8
XFILLER_100_966 VPWR VGND sg13g2_decap_8
XFILLER_84_154 VPWR VGND sg13g2_decap_8
XFILLER_57_357 VPWR VGND sg13g2_decap_8
XFILLER_27_25 VPWR VGND sg13g2_decap_8
XFILLER_26_700 VPWR VGND sg13g2_decap_8
XFILLER_38_560 VPWR VGND sg13g2_decap_8
XFILLER_25_210 VPWR VGND sg13g2_decap_8
XFILLER_81_872 VPWR VGND sg13g2_decap_8
XFILLER_53_574 VPWR VGND sg13g2_decap_8
XFILLER_41_714 VPWR VGND sg13g2_decap_8
XFILLER_14_917 VPWR VGND sg13g2_decap_8
XFILLER_26_777 VPWR VGND sg13g2_decap_8
XFILLER_80_371 VPWR VGND sg13g2_decap_8
XFILLER_43_35 VPWR VGND sg13g2_decap_8
XFILLER_13_427 VPWR VGND sg13g2_decap_8
XFILLER_25_287 VPWR VGND sg13g2_decap_8
XFILLER_40_224 VPWR VGND sg13g2_decap_8
XFILLER_5_648 VPWR VGND sg13g2_decap_8
XFILLER_49_1012 VPWR VGND sg13g2_decap_8
XFILLER_4_147 VPWR VGND sg13g2_decap_8
XFILLER_68_32 VPWR VGND sg13g2_decap_8
XFILLER_1_854 VPWR VGND sg13g2_decap_8
XFILLER_89_994 VPWR VGND sg13g2_decap_8
XFILLER_0_364 VPWR VGND sg13g2_decap_8
XFILLER_49_858 VPWR VGND sg13g2_decap_8
XFILLER_76_655 VPWR VGND sg13g2_decap_8
XFILLER_75_154 VPWR VGND sg13g2_decap_8
XFILLER_48_357 VPWR VGND sg13g2_decap_8
XFILLER_90_102 VPWR VGND sg13g2_decap_8
XFILLER_84_42 VPWR VGND sg13g2_decap_8
XFILLER_17_711 VPWR VGND sg13g2_decap_8
XFILLER_29_571 VPWR VGND sg13g2_decap_8
XFILLER_91_658 VPWR VGND sg13g2_decap_8
XFILLER_16_210 VPWR VGND sg13g2_decap_8
XFILLER_90_179 VPWR VGND sg13g2_decap_8
XFILLER_72_861 VPWR VGND sg13g2_decap_8
XFILLER_56_1005 VPWR VGND sg13g2_decap_8
XFILLER_17_788 VPWR VGND sg13g2_decap_8
XFILLER_32_725 VPWR VGND sg13g2_decap_8
XFILLER_71_382 VPWR VGND sg13g2_decap_8
XFILLER_44_585 VPWR VGND sg13g2_decap_8
XFILLER_16_287 VPWR VGND sg13g2_decap_8
XFILLER_31_224 VPWR VGND sg13g2_decap_8
XFILLER_9_910 VPWR VGND sg13g2_decap_8
XFILLER_8_420 VPWR VGND sg13g2_decap_8
XFILLER_13_994 VPWR VGND sg13g2_decap_8
XFILLER_40_791 VPWR VGND sg13g2_decap_8
XFILLER_9_987 VPWR VGND sg13g2_decap_8
XFILLER_8_497 VPWR VGND sg13g2_decap_8
XFILLER_99_714 VPWR VGND sg13g2_decap_8
XFILLER_98_235 VPWR VGND sg13g2_decap_8
XFILLER_95_942 VPWR VGND sg13g2_decap_8
XFILLER_67_644 VPWR VGND sg13g2_decap_8
XFILLER_94_441 VPWR VGND sg13g2_decap_8
XFILLER_66_132 VPWR VGND sg13g2_decap_8
XFILLER_27_508 VPWR VGND sg13g2_decap_8
XFILLER_39_368 VPWR VGND sg13g2_decap_8
XFILLER_81_102 VPWR VGND sg13g2_decap_8
XFILLER_54_305 VPWR VGND sg13g2_decap_8
XFILLER_82_658 VPWR VGND sg13g2_decap_8
XFILLER_81_179 VPWR VGND sg13g2_decap_8
XFILLER_63_861 VPWR VGND sg13g2_decap_8
XFILLER_23_714 VPWR VGND sg13g2_decap_8
XFILLER_35_574 VPWR VGND sg13g2_decap_8
XFILLER_62_371 VPWR VGND sg13g2_decap_8
XFILLER_50_511 VPWR VGND sg13g2_decap_8
XFILLER_22_235 VPWR VGND sg13g2_decap_8
XFILLER_50_588 VPWR VGND sg13g2_decap_8
XFILLER_13_49 VPWR VGND sg13g2_decap_8
XFILLER_31_791 VPWR VGND sg13g2_decap_8
XFILLER_104_546 VPWR VGND sg13g2_decap_8
XFILLER_89_224 VPWR VGND sg13g2_decap_8
XFILLER_78_909 VPWR VGND sg13g2_decap_8
XFILLER_86_942 VPWR VGND sg13g2_decap_8
XFILLER_38_35 VPWR VGND sg13g2_decap_8
XFILLER_100_763 VPWR VGND sg13g2_decap_8
XFILLER_85_441 VPWR VGND sg13g2_decap_8
XFILLER_79_1005 VPWR VGND sg13g2_decap_8
XFILLER_58_644 VPWR VGND sg13g2_decap_8
XFILLER_57_154 VPWR VGND sg13g2_decap_8
XFILLER_73_669 VPWR VGND sg13g2_decap_8
XFILLER_61_809 VPWR VGND sg13g2_decap_8
XFILLER_72_168 VPWR VGND sg13g2_decap_8
XFILLER_60_319 VPWR VGND sg13g2_decap_8
XFILLER_54_872 VPWR VGND sg13g2_decap_8
XFILLER_14_714 VPWR VGND sg13g2_decap_8
XFILLER_26_574 VPWR VGND sg13g2_decap_8
XFILLER_54_67 VPWR VGND sg13g2_decap_8
XFILLER_53_371 VPWR VGND sg13g2_decap_8
XFILLER_13_224 VPWR VGND sg13g2_decap_8
XFILLER_41_511 VPWR VGND sg13g2_decap_8
XFILLER_9_217 VPWR VGND sg13g2_decap_8
XFILLER_16_1022 VPWR VGND sg13g2_decap_8
XFILLER_41_588 VPWR VGND sg13g2_decap_8
XFILLER_70_77 VPWR VGND sg13g2_decap_8
XFILLER_10_942 VPWR VGND sg13g2_decap_8
XFILLER_6_924 VPWR VGND sg13g2_decap_8
XFILLER_5_445 VPWR VGND sg13g2_decap_8
XFILLER_79_42 VPWR VGND sg13g2_decap_8
XFILLER_96_728 VPWR VGND sg13g2_decap_8
XFILLER_1_651 VPWR VGND sg13g2_decap_8
XFILLER_89_791 VPWR VGND sg13g2_decap_8
XFILLER_77_931 VPWR VGND sg13g2_decap_8
XFILLER_0_161 VPWR VGND sg13g2_decap_8
XFILLER_95_249 VPWR VGND sg13g2_decap_8
XFILLER_95_74 VPWR VGND sg13g2_decap_8
XFILLER_76_452 VPWR VGND sg13g2_decap_8
XFILLER_49_655 VPWR VGND sg13g2_decap_8
XFILLER_23_1015 VPWR VGND sg13g2_decap_8
XFILLER_92_945 VPWR VGND sg13g2_decap_8
XFILLER_48_154 VPWR VGND sg13g2_decap_8
XFILLER_91_455 VPWR VGND sg13g2_decap_8
XFILLER_64_669 VPWR VGND sg13g2_decap_8
XFILLER_63_168 VPWR VGND sg13g2_decap_8
XFILLER_51_319 VPWR VGND sg13g2_decap_8
XFILLER_45_861 VPWR VGND sg13g2_decap_8
XFILLER_44_382 VPWR VGND sg13g2_decap_8
XFILLER_17_585 VPWR VGND sg13g2_decap_8
XFILLER_32_522 VPWR VGND sg13g2_decap_8
XFILLER_81_4 VPWR VGND sg13g2_decap_8
XFILLER_60_886 VPWR VGND sg13g2_decap_8
XFILLER_20_739 VPWR VGND sg13g2_decap_8
XFILLER_32_599 VPWR VGND sg13g2_decap_8
XFILLER_13_791 VPWR VGND sg13g2_decap_8
XFILLER_30_1008 VPWR VGND sg13g2_decap_8
XFILLER_9_784 VPWR VGND sg13g2_decap_8
XFILLER_8_294 VPWR VGND sg13g2_decap_8
XFILLER_99_511 VPWR VGND sg13g2_decap_8
XFILLER_99_588 VPWR VGND sg13g2_decap_8
XFILLER_87_728 VPWR VGND sg13g2_decap_8
XFILLER_86_249 VPWR VGND sg13g2_decap_8
XFILLER_68_964 VPWR VGND sg13g2_decap_8
XFILLER_67_441 VPWR VGND sg13g2_decap_8
XFILLER_54_102 VPWR VGND sg13g2_decap_8
XFILLER_27_305 VPWR VGND sg13g2_decap_8
XFILLER_39_165 VPWR VGND sg13g2_decap_8
XFILLER_83_956 VPWR VGND sg13g2_decap_8
XFILLER_55_658 VPWR VGND sg13g2_decap_8
XFILLER_82_455 VPWR VGND sg13g2_decap_8
XFILLER_54_179 VPWR VGND sg13g2_decap_8
XFILLER_42_319 VPWR VGND sg13g2_decap_8
XFILLER_36_861 VPWR VGND sg13g2_decap_8
XFILLER_23_511 VPWR VGND sg13g2_decap_8
XFILLER_35_371 VPWR VGND sg13g2_decap_8
XFILLER_51_886 VPWR VGND sg13g2_decap_8
XFILLER_50_385 VPWR VGND sg13g2_decap_8
XFILLER_11_728 VPWR VGND sg13g2_decap_8
XFILLER_23_588 VPWR VGND sg13g2_decap_8
XFILLER_10_249 VPWR VGND sg13g2_decap_8
XFILLER_40_14 VPWR VGND sg13g2_decap_8
XFILLER_3_938 VPWR VGND sg13g2_decap_8
XFILLER_105_833 VPWR VGND sg13g2_decap_8
XFILLER_104_343 VPWR VGND sg13g2_decap_8
XFILLER_78_706 VPWR VGND sg13g2_decap_8
XFILLER_46_1026 VPWR VGND sg13g2_fill_2
XFILLER_2_459 VPWR VGND sg13g2_decap_8
XFILLER_77_238 VPWR VGND sg13g2_decap_8
XFILLER_49_67 VPWR VGND sg13g2_decap_8
XFILLER_59_964 VPWR VGND sg13g2_decap_8
XFILLER_58_441 VPWR VGND sg13g2_decap_8
XFILLER_105_84 VPWR VGND sg13g2_decap_8
XFILLER_100_560 VPWR VGND sg13g2_decap_8
XFILLER_74_967 VPWR VGND sg13g2_decap_8
XFILLER_34_809 VPWR VGND sg13g2_decap_8
XFILLER_73_466 VPWR VGND sg13g2_decap_8
XFILLER_65_77 VPWR VGND sg13g2_decap_8
XFILLER_61_606 VPWR VGND sg13g2_decap_8
XFILLER_46_669 VPWR VGND sg13g2_decap_8
XFILLER_45_168 VPWR VGND sg13g2_decap_8
XFILLER_27_872 VPWR VGND sg13g2_decap_8
XFILLER_33_308 VPWR VGND sg13g2_decap_8
XFILLER_60_116 VPWR VGND sg13g2_decap_8
XFILLER_14_511 VPWR VGND sg13g2_decap_8
XFILLER_26_371 VPWR VGND sg13g2_decap_8
XFILLER_81_32 VPWR VGND sg13g2_decap_8
XFILLER_53_1008 VPWR VGND sg13g2_decap_8
XFILLER_42_886 VPWR VGND sg13g2_decap_8
XFILLER_14_588 VPWR VGND sg13g2_decap_8
XFILLER_41_385 VPWR VGND sg13g2_decap_8
XFILLER_14_70 VPWR VGND sg13g2_decap_8
XFILLER_6_721 VPWR VGND sg13g2_decap_8
XFILLER_5_242 VPWR VGND sg13g2_decap_8
XFILLER_6_798 VPWR VGND sg13g2_decap_8
XFILLER_30_91 VPWR VGND sg13g2_decap_8
XFILLER_96_525 VPWR VGND sg13g2_decap_8
Xinput7 ui_in[6] net7 VPWR VGND sg13g2_buf_1
XFILLER_49_452 VPWR VGND sg13g2_decap_8
XFILLER_92_742 VPWR VGND sg13g2_decap_8
XFILLER_65_945 VPWR VGND sg13g2_decap_8
XFILLER_91_252 VPWR VGND sg13g2_decap_8
XFILLER_64_466 VPWR VGND sg13g2_decap_8
XFILLER_18_861 VPWR VGND sg13g2_decap_8
XFILLER_36_168 VPWR VGND sg13g2_decap_8
XFILLER_37_669 VPWR VGND sg13g2_decap_8
XFILLER_80_959 VPWR VGND sg13g2_decap_8
XFILLER_51_116 VPWR VGND sg13g2_decap_8
XFILLER_17_382 VPWR VGND sg13g2_decap_8
XFILLER_24_319 VPWR VGND sg13g2_decap_8
XFILLER_60_683 VPWR VGND sg13g2_decap_8
XFILLER_33_875 VPWR VGND sg13g2_decap_8
XFILLER_20_536 VPWR VGND sg13g2_decap_8
XFILLER_32_396 VPWR VGND sg13g2_decap_8
XFILLER_72_0 VPWR VGND sg13g2_decap_8
XFILLER_9_581 VPWR VGND sg13g2_decap_8
XFILLER_10_39 VPWR VGND sg13g2_decap_8
XFILLER_102_847 VPWR VGND sg13g2_decap_8
XFILLER_99_385 VPWR VGND sg13g2_decap_8
XFILLER_87_525 VPWR VGND sg13g2_decap_8
XFILLER_101_357 VPWR VGND sg13g2_decap_8
XFILLER_68_761 VPWR VGND sg13g2_decap_8
XFILLER_83_753 VPWR VGND sg13g2_decap_8
XFILLER_56_956 VPWR VGND sg13g2_decap_8
XFILLER_27_102 VPWR VGND sg13g2_decap_8
XFILLER_28_658 VPWR VGND sg13g2_decap_8
XFILLER_82_252 VPWR VGND sg13g2_decap_8
XFILLER_76_1019 VPWR VGND sg13g2_decap_8
XFILLER_55_455 VPWR VGND sg13g2_decap_8
XFILLER_35_14 VPWR VGND sg13g2_decap_8
XFILLER_42_116 VPWR VGND sg13g2_decap_8
XFILLER_15_319 VPWR VGND sg13g2_decap_8
XFILLER_27_179 VPWR VGND sg13g2_decap_8
XFILLER_70_469 VPWR VGND sg13g2_decap_8
XFILLER_51_683 VPWR VGND sg13g2_decap_8
XFILLER_24_886 VPWR VGND sg13g2_decap_8
XFILLER_50_182 VPWR VGND sg13g2_decap_8
XFILLER_11_525 VPWR VGND sg13g2_decap_8
XFILLER_23_385 VPWR VGND sg13g2_decap_8
XFILLER_51_46 VPWR VGND sg13g2_decap_8
XFILLER_7_529 VPWR VGND sg13g2_decap_8
XFILLER_105_630 VPWR VGND sg13g2_decap_8
XFILLER_3_735 VPWR VGND sg13g2_decap_8
XFILLER_104_140 VPWR VGND sg13g2_decap_8
XFILLER_78_503 VPWR VGND sg13g2_decap_8
XFILLER_2_256 VPWR VGND sg13g2_decap_8
XFILLER_76_32 VPWR VGND sg13g2_decap_8
XFILLER_59_761 VPWR VGND sg13g2_decap_8
XFILLER_47_945 VPWR VGND sg13g2_decap_8
XFILLER_19_658 VPWR VGND sg13g2_decap_8
XFILLER_74_764 VPWR VGND sg13g2_decap_8
XFILLER_46_466 VPWR VGND sg13g2_decap_8
XFILLER_18_168 VPWR VGND sg13g2_decap_8
XFILLER_34_606 VPWR VGND sg13g2_decap_8
XFILLER_92_42 VPWR VGND sg13g2_decap_8
XFILLER_73_263 VPWR VGND sg13g2_decap_8
XFILLER_62_959 VPWR VGND sg13g2_decap_8
XFILLER_61_403 VPWR VGND sg13g2_decap_8
XFILLER_33_105 VPWR VGND sg13g2_decap_8
XFILLER_42_683 VPWR VGND sg13g2_decap_8
XFILLER_15_886 VPWR VGND sg13g2_decap_8
XFILLER_30_812 VPWR VGND sg13g2_decap_8
XFILLER_14_385 VPWR VGND sg13g2_decap_8
XFILLER_25_91 VPWR VGND sg13g2_decap_8
XFILLER_41_182 VPWR VGND sg13g2_decap_8
XFILLER_30_889 VPWR VGND sg13g2_decap_8
XFILLER_6_595 VPWR VGND sg13g2_decap_8
XFILLER_44_4 VPWR VGND sg13g2_decap_8
XFILLER_97_812 VPWR VGND sg13g2_decap_8
XFILLER_96_322 VPWR VGND sg13g2_decap_8
XFILLER_69_547 VPWR VGND sg13g2_decap_8
XFILLER_99_1008 VPWR VGND sg13g2_decap_8
XFILLER_97_889 VPWR VGND sg13g2_decap_8
XFILLER_96_399 VPWR VGND sg13g2_decap_8
XFILLER_84_539 VPWR VGND sg13g2_decap_8
XFILLER_65_742 VPWR VGND sg13g2_decap_8
XFILLER_2_95 VPWR VGND sg13g2_decap_8
XFILLER_38_945 VPWR VGND sg13g2_decap_8
X_57_ VPWR VGND _21_ _22_ _13_ net6 _23_ net14 sg13g2_a221oi_1
XFILLER_37_466 VPWR VGND sg13g2_decap_8
XFILLER_64_263 VPWR VGND sg13g2_decap_8
XFILLER_53_959 VPWR VGND sg13g2_decap_8
XFILLER_24_116 VPWR VGND sg13g2_decap_8
XFILLER_80_756 VPWR VGND sg13g2_decap_8
XFILLER_52_469 VPWR VGND sg13g2_decap_8
XFILLER_40_609 VPWR VGND sg13g2_decap_8
XFILLER_61_970 VPWR VGND sg13g2_decap_8
XFILLER_21_812 VPWR VGND sg13g2_decap_8
XFILLER_33_672 VPWR VGND sg13g2_decap_8
XFILLER_60_480 VPWR VGND sg13g2_decap_8
XFILLER_20_333 VPWR VGND sg13g2_decap_8
XFILLER_32_193 VPWR VGND sg13g2_decap_8
XFILLER_21_889 VPWR VGND sg13g2_decap_8
XFILLER_21_49 VPWR VGND sg13g2_decap_8
XFILLER_106_427 VPWR VGND sg13g2_decap_8
XFILLER_82_1001 VPWR VGND sg13g2_decap_8
XFILLER_88_823 VPWR VGND sg13g2_decap_8
XFILLER_102_644 VPWR VGND sg13g2_decap_8
XFILLER_99_182 VPWR VGND sg13g2_decap_8
XFILLER_87_322 VPWR VGND sg13g2_decap_8
XFILLER_0_749 VPWR VGND sg13g2_decap_8
XFILLER_101_154 VPWR VGND sg13g2_decap_8
XFILLER_87_399 VPWR VGND sg13g2_decap_8
XFILLER_75_539 VPWR VGND sg13g2_decap_8
XFILLER_29_956 VPWR VGND sg13g2_decap_8
XFILLER_83_550 VPWR VGND sg13g2_decap_8
XFILLER_56_753 VPWR VGND sg13g2_decap_8
XFILLER_55_252 VPWR VGND sg13g2_decap_8
XFILLER_46_46 VPWR VGND sg13g2_decap_8
XFILLER_28_455 VPWR VGND sg13g2_decap_8
XFILLER_15_116 VPWR VGND sg13g2_decap_8
XFILLER_102_63 VPWR VGND sg13g2_decap_8
XFILLER_71_767 VPWR VGND sg13g2_decap_8
XFILLER_31_609 VPWR VGND sg13g2_decap_8
XFILLER_70_266 VPWR VGND sg13g2_decap_8
XFILLER_43_469 VPWR VGND sg13g2_decap_8
XFILLER_30_119 VPWR VGND sg13g2_decap_8
XFILLER_62_56 VPWR VGND sg13g2_fill_1
XFILLER_51_480 VPWR VGND sg13g2_decap_8
XFILLER_8_805 VPWR VGND sg13g2_decap_8
XFILLER_11_322 VPWR VGND sg13g2_decap_8
XFILLER_12_823 VPWR VGND sg13g2_decap_8
XFILLER_23_182 VPWR VGND sg13g2_decap_8
XFILLER_24_683 VPWR VGND sg13g2_decap_8
XFILLER_7_18 VPWR VGND sg13g2_decap_8
XFILLER_7_326 VPWR VGND sg13g2_decap_8
XFILLER_11_399 VPWR VGND sg13g2_decap_8
XFILLER_3_532 VPWR VGND sg13g2_decap_8
XFILLER_106_994 VPWR VGND sg13g2_decap_8
XFILLER_97_119 VPWR VGND sg13g2_decap_8
XFILLER_87_42 VPWR VGND sg13g2_decap_8
XFILLER_79_823 VPWR VGND sg13g2_decap_8
XFILLER_78_300 VPWR VGND sg13g2_decap_8
XFILLER_94_826 VPWR VGND sg13g2_decap_8
XFILLER_78_377 VPWR VGND sg13g2_decap_8
XFILLER_66_517 VPWR VGND sg13g2_decap_8
XFILLER_4_1001 VPWR VGND sg13g2_decap_8
XFILLER_93_369 VPWR VGND sg13g2_decap_8
XFILLER_47_742 VPWR VGND sg13g2_decap_8
XFILLER_19_455 VPWR VGND sg13g2_decap_8
XFILLER_74_561 VPWR VGND sg13g2_decap_8
XFILLER_61_200 VPWR VGND sg13g2_decap_8
XFILLER_46_263 VPWR VGND sg13g2_decap_8
XFILLER_34_403 VPWR VGND sg13g2_decap_8
XFILLER_62_756 VPWR VGND sg13g2_decap_8
XFILLER_35_959 VPWR VGND sg13g2_decap_8
XFILLER_61_277 VPWR VGND sg13g2_decap_8
XFILLER_42_480 VPWR VGND sg13g2_decap_8
XFILLER_14_182 VPWR VGND sg13g2_decap_8
XFILLER_15_683 VPWR VGND sg13g2_decap_8
XFILLER_21_119 VPWR VGND sg13g2_decap_8
Xinput10 uio_in[1] net10 VPWR VGND sg13g2_buf_1
XFILLER_30_686 VPWR VGND sg13g2_decap_8
XFILLER_66_1007 VPWR VGND sg13g2_decap_8
XFILLER_7_893 VPWR VGND sg13g2_decap_8
XFILLER_89_609 VPWR VGND sg13g2_decap_8
XFILLER_6_392 VPWR VGND sg13g2_decap_8
XFILLER_69_344 VPWR VGND sg13g2_decap_8
XFILLER_35_0 VPWR VGND sg13g2_decap_8
XFILLER_97_686 VPWR VGND sg13g2_decap_8
XFILLER_85_826 VPWR VGND sg13g2_decap_8
XFILLER_96_196 VPWR VGND sg13g2_decap_8
XFILLER_84_336 VPWR VGND sg13g2_decap_8
XFILLER_57_539 VPWR VGND sg13g2_decap_8
XFILLER_38_742 VPWR VGND sg13g2_decap_8
XFILLER_37_263 VPWR VGND sg13g2_decap_8
XFILLER_80_553 VPWR VGND sg13g2_decap_8
XFILLER_53_756 VPWR VGND sg13g2_decap_8
XFILLER_16_49 VPWR VGND sg13g2_decap_8
XFILLER_26_959 VPWR VGND sg13g2_decap_8
XFILLER_52_266 VPWR VGND sg13g2_decap_8
XFILLER_13_609 VPWR VGND sg13g2_decap_8
XFILLER_25_469 VPWR VGND sg13g2_decap_8
XFILLER_34_970 VPWR VGND sg13g2_decap_8
XFILLER_40_406 VPWR VGND sg13g2_decap_8
XFILLER_20_130 VPWR VGND sg13g2_decap_8
XFILLER_21_686 VPWR VGND sg13g2_decap_8
XFILLER_106_224 VPWR VGND sg13g2_decap_8
XFILLER_4_329 VPWR VGND sg13g2_decap_8
XFILLER_10_1028 VPWR VGND sg13g2_fill_1
XFILLER_103_931 VPWR VGND sg13g2_decap_8
XFILLER_88_620 VPWR VGND sg13g2_decap_8
XFILLER_0_546 VPWR VGND sg13g2_decap_8
XFILLER_102_441 VPWR VGND sg13g2_decap_8
XFILLER_88_697 VPWR VGND sg13g2_decap_8
XFILLER_87_196 VPWR VGND sg13g2_decap_8
XFILLER_76_837 VPWR VGND sg13g2_decap_8
XFILLER_75_336 VPWR VGND sg13g2_decap_8
XFILLER_57_56 VPWR VGND sg13g2_decap_8
XFILLER_48_539 VPWR VGND sg13g2_decap_8
XFILLER_56_550 VPWR VGND sg13g2_decap_8
XFILLER_29_753 VPWR VGND sg13g2_decap_8
XFILLER_73_11 VPWR VGND sg13g2_decap_8
XFILLER_28_252 VPWR VGND sg13g2_decap_8
XFILLER_44_767 VPWR VGND sg13g2_decap_8
XFILLER_32_907 VPWR VGND sg13g2_decap_8
XFILLER_73_88 VPWR VGND sg13g2_decap_8
XFILLER_71_564 VPWR VGND sg13g2_decap_8
XFILLER_43_266 VPWR VGND sg13g2_decap_8
XFILLER_16_469 VPWR VGND sg13g2_decap_8
XFILLER_31_406 VPWR VGND sg13g2_decap_8
XFILLER_106_1001 VPWR VGND sg13g2_decap_8
XFILLER_12_620 VPWR VGND sg13g2_decap_8
XFILLER_24_480 VPWR VGND sg13g2_decap_8
XFILLER_8_602 VPWR VGND sg13g2_decap_8
XFILLER_40_973 VPWR VGND sg13g2_decap_8
XFILLER_7_123 VPWR VGND sg13g2_decap_8
XFILLER_12_697 VPWR VGND sg13g2_decap_8
XFILLER_8_679 VPWR VGND sg13g2_decap_8
XFILLER_11_196 VPWR VGND sg13g2_decap_8
XFILLER_22_81 VPWR VGND sg13g2_decap_8
XFILLER_98_417 VPWR VGND sg13g2_decap_8
XFILLER_98_74 VPWR VGND sg13g2_decap_8
XFILLER_4_896 VPWR VGND sg13g2_decap_8
XFILLER_106_791 VPWR VGND sg13g2_decap_8
XFILLER_79_620 VPWR VGND sg13g2_decap_8
XFILLER_67_826 VPWR VGND sg13g2_decap_8
XFILLER_94_623 VPWR VGND sg13g2_decap_8
XFILLER_79_697 VPWR VGND sg13g2_decap_8
XFILLER_78_174 VPWR VGND sg13g2_decap_8
XFILLER_66_314 VPWR VGND sg13g2_decap_8
XFILLER_93_166 VPWR VGND sg13g2_decap_8
XFILLER_19_252 VPWR VGND sg13g2_decap_8
XFILLER_34_200 VPWR VGND sg13g2_decap_8
XFILLER_90_851 VPWR VGND sg13g2_decap_8
XFILLER_35_756 VPWR VGND sg13g2_decap_8
XFILLER_62_553 VPWR VGND sg13g2_decap_8
XFILLER_22_417 VPWR VGND sg13g2_decap_8
XFILLER_72_1022 VPWR VGND sg13g2_decap_8
XFILLER_15_480 VPWR VGND sg13g2_decap_8
XFILLER_34_277 VPWR VGND sg13g2_decap_8
XFILLER_31_973 VPWR VGND sg13g2_decap_8
XFILLER_30_483 VPWR VGND sg13g2_decap_8
XFILLER_7_690 VPWR VGND sg13g2_decap_8
XFILLER_104_728 VPWR VGND sg13g2_decap_8
XFILLER_89_406 VPWR VGND sg13g2_decap_8
XFILLER_103_238 VPWR VGND sg13g2_decap_8
XFILLER_98_984 VPWR VGND sg13g2_decap_8
XFILLER_69_141 VPWR VGND sg13g2_decap_8
XFILLER_58_826 VPWR VGND sg13g2_decap_8
XFILLER_100_945 VPWR VGND sg13g2_decap_8
XFILLER_97_483 VPWR VGND sg13g2_decap_8
XFILLER_85_623 VPWR VGND sg13g2_decap_8
XFILLER_57_336 VPWR VGND sg13g2_decap_8
XFILLER_84_133 VPWR VGND sg13g2_decap_8
XFILLER_66_881 VPWR VGND sg13g2_decap_8
XFILLER_81_851 VPWR VGND sg13g2_decap_8
XFILLER_26_756 VPWR VGND sg13g2_decap_8
XFILLER_80_350 VPWR VGND sg13g2_decap_8
XFILLER_53_553 VPWR VGND sg13g2_decap_8
XFILLER_43_14 VPWR VGND sg13g2_decap_8
XFILLER_13_406 VPWR VGND sg13g2_decap_8
XFILLER_25_266 VPWR VGND sg13g2_decap_8
XFILLER_40_203 VPWR VGND sg13g2_decap_8
XFILLER_22_984 VPWR VGND sg13g2_decap_8
XFILLER_21_483 VPWR VGND sg13g2_decap_8
XFILLER_5_627 VPWR VGND sg13g2_decap_8
XFILLER_4_126 VPWR VGND sg13g2_decap_8
XFILLER_68_11 VPWR VGND sg13g2_decap_8
XFILLER_1_833 VPWR VGND sg13g2_decap_8
XFILLER_89_973 VPWR VGND sg13g2_decap_8
XFILLER_0_343 VPWR VGND sg13g2_decap_8
XFILLER_88_494 VPWR VGND sg13g2_decap_8
XFILLER_76_634 VPWR VGND sg13g2_decap_8
XFILLER_49_837 VPWR VGND sg13g2_decap_8
XFILLER_84_21 VPWR VGND sg13g2_decap_8
XFILLER_75_133 VPWR VGND sg13g2_decap_8
XFILLER_48_336 VPWR VGND sg13g2_decap_8
XFILLER_91_637 VPWR VGND sg13g2_decap_8
XFILLER_1_1015 VPWR VGND sg13g2_decap_8
XFILLER_29_550 VPWR VGND sg13g2_decap_8
XFILLER_84_98 VPWR VGND sg13g2_decap_8
XFILLER_72_840 VPWR VGND sg13g2_decap_8
XFILLER_90_158 VPWR VGND sg13g2_decap_8
XFILLER_71_361 VPWR VGND sg13g2_decap_8
XFILLER_56_1028 VPWR VGND sg13g2_fill_1
XFILLER_44_564 VPWR VGND sg13g2_decap_8
XFILLER_16_266 VPWR VGND sg13g2_decap_8
XFILLER_17_81 VPWR VGND sg13g2_decap_8
XFILLER_17_767 VPWR VGND sg13g2_decap_8
XFILLER_32_704 VPWR VGND sg13g2_decap_8
XFILLER_31_203 VPWR VGND sg13g2_decap_8
XFILLER_13_973 VPWR VGND sg13g2_decap_8
XFILLER_40_770 VPWR VGND sg13g2_decap_8
XFILLER_9_966 VPWR VGND sg13g2_decap_8
XFILLER_12_494 VPWR VGND sg13g2_decap_8
XFILLER_33_91 VPWR VGND sg13g2_decap_8
XFILLER_8_476 VPWR VGND sg13g2_decap_8
XFILLER_98_214 VPWR VGND sg13g2_decap_8
XFILLER_4_693 VPWR VGND sg13g2_decap_8
XFILLER_95_921 VPWR VGND sg13g2_decap_8
XFILLER_94_420 VPWR VGND sg13g2_decap_8
XFILLER_79_494 VPWR VGND sg13g2_decap_8
XFILLER_67_623 VPWR VGND sg13g2_decap_8
XFILLER_66_111 VPWR VGND sg13g2_decap_8
XFILLER_39_347 VPWR VGND sg13g2_decap_8
XFILLER_95_998 VPWR VGND sg13g2_decap_8
XFILLER_82_637 VPWR VGND sg13g2_decap_8
XFILLER_94_497 VPWR VGND sg13g2_decap_8
XFILLER_66_188 VPWR VGND sg13g2_decap_8
XFILLER_63_840 VPWR VGND sg13g2_decap_8
XFILLER_81_158 VPWR VGND sg13g2_decap_8
XFILLER_62_350 VPWR VGND sg13g2_decap_8
XFILLER_35_553 VPWR VGND sg13g2_decap_8
XFILLER_22_214 VPWR VGND sg13g2_decap_8
XFILLER_50_567 VPWR VGND sg13g2_decap_8
XFILLER_13_28 VPWR VGND sg13g2_decap_8
XFILLER_31_770 VPWR VGND sg13g2_decap_8
XFILLER_30_280 VPWR VGND sg13g2_decap_8
XFILLER_89_203 VPWR VGND sg13g2_decap_8
XFILLER_104_525 VPWR VGND sg13g2_decap_8
XFILLER_98_781 VPWR VGND sg13g2_decap_8
XFILLER_86_921 VPWR VGND sg13g2_decap_8
XFILLER_85_420 VPWR VGND sg13g2_decap_8
XFILLER_58_623 VPWR VGND sg13g2_decap_8
XFILLER_38_14 VPWR VGND sg13g2_decap_8
XFILLER_100_742 VPWR VGND sg13g2_decap_8
XFILLER_97_280 VPWR VGND sg13g2_decap_8
XFILLER_57_133 VPWR VGND sg13g2_decap_8
XFILLER_86_998 VPWR VGND sg13g2_decap_8
XFILLER_79_1028 VPWR VGND sg13g2_fill_1
XFILLER_85_497 VPWR VGND sg13g2_decap_8
XFILLER_73_648 VPWR VGND sg13g2_decap_8
XFILLER_72_147 VPWR VGND sg13g2_decap_8
XFILLER_54_851 VPWR VGND sg13g2_decap_8
XFILLER_54_46 VPWR VGND sg13g2_decap_8
XFILLER_53_350 VPWR VGND sg13g2_decap_8
XFILLER_26_553 VPWR VGND sg13g2_decap_8
XFILLER_13_203 VPWR VGND sg13g2_decap_8
XFILLER_16_1001 VPWR VGND sg13g2_decap_8
XFILLER_41_567 VPWR VGND sg13g2_decap_8
XFILLER_10_921 VPWR VGND sg13g2_decap_8
XFILLER_22_781 VPWR VGND sg13g2_decap_8
XFILLER_103_1015 VPWR VGND sg13g2_decap_8
XFILLER_70_56 VPWR VGND sg13g2_decap_8
XFILLER_6_903 VPWR VGND sg13g2_decap_8
XFILLER_21_280 VPWR VGND sg13g2_decap_8
XFILLER_5_424 VPWR VGND sg13g2_decap_8
XFILLER_10_998 VPWR VGND sg13g2_decap_8
XFILLER_102_0 VPWR VGND sg13g2_decap_8
XFILLER_79_21 VPWR VGND sg13g2_decap_8
XFILLER_96_707 VPWR VGND sg13g2_decap_8
XFILLER_1_630 VPWR VGND sg13g2_decap_8
XFILLER_95_228 VPWR VGND sg13g2_decap_8
XFILLER_89_770 VPWR VGND sg13g2_decap_8
XFILLER_77_910 VPWR VGND sg13g2_decap_8
XFILLER_49_634 VPWR VGND sg13g2_decap_8
XFILLER_0_140 VPWR VGND sg13g2_decap_8
XFILLER_95_53 VPWR VGND sg13g2_decap_8
XFILLER_88_291 VPWR VGND sg13g2_decap_8
XFILLER_76_431 VPWR VGND sg13g2_decap_8
XFILLER_48_133 VPWR VGND sg13g2_decap_8
XFILLER_92_924 VPWR VGND sg13g2_decap_8
XFILLER_77_987 VPWR VGND sg13g2_decap_8
XFILLER_91_434 VPWR VGND sg13g2_decap_8
XFILLER_64_648 VPWR VGND sg13g2_decap_8
XFILLER_45_840 VPWR VGND sg13g2_decap_8
XFILLER_28_91 VPWR VGND sg13g2_decap_8
XFILLER_63_147 VPWR VGND sg13g2_decap_8
XFILLER_17_564 VPWR VGND sg13g2_decap_8
XFILLER_44_361 VPWR VGND sg13g2_decap_8
XFILLER_32_501 VPWR VGND sg13g2_decap_8
XFILLER_60_865 VPWR VGND sg13g2_decap_8
XFILLER_13_770 VPWR VGND sg13g2_decap_8
XFILLER_20_718 VPWR VGND sg13g2_decap_8
XFILLER_32_578 VPWR VGND sg13g2_decap_8
XFILLER_9_763 VPWR VGND sg13g2_decap_8
XFILLER_8_273 VPWR VGND sg13g2_decap_8
XFILLER_12_291 VPWR VGND sg13g2_decap_8
XFILLER_5_991 VPWR VGND sg13g2_decap_8
XFILLER_99_567 VPWR VGND sg13g2_decap_8
XFILLER_87_707 VPWR VGND sg13g2_decap_8
XFILLER_5_95 VPWR VGND sg13g2_decap_8
XFILLER_4_490 VPWR VGND sg13g2_decap_8
XFILLER_101_539 VPWR VGND sg13g2_decap_8
XFILLER_86_228 VPWR VGND sg13g2_decap_8
XFILLER_79_291 VPWR VGND sg13g2_decap_8
XFILLER_68_943 VPWR VGND sg13g2_decap_8
XFILLER_67_420 VPWR VGND sg13g2_decap_8
XFILLER_95_795 VPWR VGND sg13g2_decap_8
XFILLER_83_935 VPWR VGND sg13g2_decap_8
XFILLER_39_144 VPWR VGND sg13g2_decap_8
XFILLER_94_294 VPWR VGND sg13g2_decap_8
XFILLER_82_434 VPWR VGND sg13g2_decap_8
XFILLER_67_497 VPWR VGND sg13g2_decap_8
XFILLER_55_637 VPWR VGND sg13g2_decap_8
XFILLER_36_840 VPWR VGND sg13g2_decap_8
XFILLER_54_158 VPWR VGND sg13g2_decap_8
XFILLER_35_350 VPWR VGND sg13g2_decap_8
XFILLER_39_1012 VPWR VGND sg13g2_decap_8
XFILLER_51_865 VPWR VGND sg13g2_decap_8
XFILLER_11_707 VPWR VGND sg13g2_decap_8
XFILLER_50_364 VPWR VGND sg13g2_decap_8
XFILLER_23_567 VPWR VGND sg13g2_decap_8
XFILLER_10_228 VPWR VGND sg13g2_decap_8
XFILLER_105_812 VPWR VGND sg13g2_decap_8
XFILLER_3_917 VPWR VGND sg13g2_decap_8
XFILLER_104_322 VPWR VGND sg13g2_decap_8
XFILLER_46_1005 VPWR VGND sg13g2_decap_8
XFILLER_6_7 VPWR VGND sg13g2_decap_8
XFILLER_2_438 VPWR VGND sg13g2_decap_8
XFILLER_105_889 VPWR VGND sg13g2_decap_8
XFILLER_49_46 VPWR VGND sg13g2_decap_8
XFILLER_104_399 VPWR VGND sg13g2_decap_8
XFILLER_77_217 VPWR VGND sg13g2_decap_8
XFILLER_59_943 VPWR VGND sg13g2_decap_8
XFILLER_58_420 VPWR VGND sg13g2_decap_8
XFILLER_105_63 VPWR VGND sg13g2_decap_8
XFILLER_86_795 VPWR VGND sg13g2_decap_8
XFILLER_85_294 VPWR VGND sg13g2_decap_8
XFILLER_74_946 VPWR VGND sg13g2_decap_8
XFILLER_73_445 VPWR VGND sg13g2_decap_8
XFILLER_65_56 VPWR VGND sg13g2_decap_8
XFILLER_58_497 VPWR VGND sg13g2_decap_8
XFILLER_46_648 VPWR VGND sg13g2_decap_8
XFILLER_45_147 VPWR VGND sg13g2_decap_8
XFILLER_27_851 VPWR VGND sg13g2_decap_8
XFILLER_81_11 VPWR VGND sg13g2_decap_8
XFILLER_26_350 VPWR VGND sg13g2_decap_8
XFILLER_42_865 VPWR VGND sg13g2_decap_8
XFILLER_14_567 VPWR VGND sg13g2_decap_8
XFILLER_41_364 VPWR VGND sg13g2_decap_8
XFILLER_81_88 VPWR VGND sg13g2_decap_8
XFILLER_6_700 VPWR VGND sg13g2_decap_8
XFILLER_5_221 VPWR VGND sg13g2_decap_8
XFILLER_10_795 VPWR VGND sg13g2_decap_8
XFILLER_6_777 VPWR VGND sg13g2_decap_8
XFILLER_5_298 VPWR VGND sg13g2_decap_8
XFILLER_30_70 VPWR VGND sg13g2_decap_8
XFILLER_96_504 VPWR VGND sg13g2_decap_8
XFILLER_69_729 VPWR VGND sg13g2_decap_8
XFILLER_49_431 VPWR VGND sg13g2_decap_8
Xinput8 ui_in[7] net8 VPWR VGND sg13g2_buf_1
XFILLER_77_784 VPWR VGND sg13g2_decap_8
XFILLER_65_924 VPWR VGND sg13g2_decap_8
XFILLER_92_721 VPWR VGND sg13g2_decap_8
XFILLER_37_648 VPWR VGND sg13g2_decap_8
XFILLER_91_231 VPWR VGND sg13g2_decap_8
XFILLER_64_445 VPWR VGND sg13g2_decap_8
XFILLER_18_840 VPWR VGND sg13g2_decap_8
XFILLER_36_147 VPWR VGND sg13g2_decap_8
XFILLER_92_798 VPWR VGND sg13g2_decap_8
XFILLER_80_938 VPWR VGND sg13g2_decap_8
XFILLER_17_361 VPWR VGND sg13g2_decap_8
XFILLER_33_854 VPWR VGND sg13g2_decap_8
XFILLER_60_662 VPWR VGND sg13g2_decap_8
XFILLER_20_515 VPWR VGND sg13g2_decap_8
XFILLER_32_375 VPWR VGND sg13g2_decap_8
XFILLER_9_560 VPWR VGND sg13g2_decap_8
XFILLER_69_1016 VPWR VGND sg13g2_decap_8
XFILLER_65_0 VPWR VGND sg13g2_decap_8
XFILLER_106_609 VPWR VGND sg13g2_decap_8
XFILLER_69_1027 VPWR VGND sg13g2_fill_2
XFILLER_10_18 VPWR VGND sg13g2_decap_8
XFILLER_105_119 VPWR VGND sg13g2_decap_8
XFILLER_102_826 VPWR VGND sg13g2_decap_8
XFILLER_99_364 VPWR VGND sg13g2_decap_8
XFILLER_87_504 VPWR VGND sg13g2_decap_8
XFILLER_101_336 VPWR VGND sg13g2_decap_8
XFILLER_68_740 VPWR VGND sg13g2_decap_8
XFILLER_19_49 VPWR VGND sg13g2_decap_8
XFILLER_95_592 VPWR VGND sg13g2_decap_8
XFILLER_83_732 VPWR VGND sg13g2_decap_8
XFILLER_67_294 VPWR VGND sg13g2_decap_8
XFILLER_56_935 VPWR VGND sg13g2_decap_8
XFILLER_55_434 VPWR VGND sg13g2_decap_8
XFILLER_28_637 VPWR VGND sg13g2_decap_8
XFILLER_82_231 VPWR VGND sg13g2_decap_8
XFILLER_27_158 VPWR VGND sg13g2_decap_8
XFILLER_71_949 VPWR VGND sg13g2_decap_8
XFILLER_70_448 VPWR VGND sg13g2_decap_8
XFILLER_24_865 VPWR VGND sg13g2_decap_8
XFILLER_51_662 VPWR VGND sg13g2_decap_8
XFILLER_11_504 VPWR VGND sg13g2_decap_8
XFILLER_23_364 VPWR VGND sg13g2_decap_8
XFILLER_51_25 VPWR VGND sg13g2_decap_8
XFILLER_50_161 VPWR VGND sg13g2_decap_8
XFILLER_7_508 VPWR VGND sg13g2_decap_8
XFILLER_13_1015 VPWR VGND sg13g2_decap_8
XFILLER_3_714 VPWR VGND sg13g2_decap_8
XFILLER_2_235 VPWR VGND sg13g2_decap_8
XFILLER_105_686 VPWR VGND sg13g2_decap_8
XFILLER_104_196 VPWR VGND sg13g2_decap_8
XFILLER_78_559 VPWR VGND sg13g2_decap_8
XFILLER_76_11 VPWR VGND sg13g2_decap_8
XFILLER_59_740 VPWR VGND sg13g2_decap_8
XFILLER_47_924 VPWR VGND sg13g2_decap_8
XFILLER_86_592 VPWR VGND sg13g2_decap_8
XFILLER_76_88 VPWR VGND sg13g2_decap_8
XFILLER_74_743 VPWR VGND sg13g2_decap_8
XFILLER_58_294 VPWR VGND sg13g2_decap_8
XFILLER_19_637 VPWR VGND sg13g2_decap_8
XFILLER_20_1019 VPWR VGND sg13g2_decap_8
XFILLER_92_21 VPWR VGND sg13g2_decap_8
XFILLER_73_242 VPWR VGND sg13g2_decap_8
XFILLER_46_445 VPWR VGND sg13g2_decap_8
XFILLER_18_147 VPWR VGND sg13g2_decap_8
XFILLER_62_938 VPWR VGND sg13g2_decap_8
XFILLER_61_459 VPWR VGND sg13g2_decap_8
XFILLER_92_98 VPWR VGND sg13g2_decap_8
XFILLER_42_662 VPWR VGND sg13g2_decap_8
XFILLER_14_364 VPWR VGND sg13g2_decap_8
XFILLER_15_865 VPWR VGND sg13g2_decap_8
XFILLER_25_70 VPWR VGND sg13g2_decap_8
XFILLER_41_161 VPWR VGND sg13g2_decap_8
XFILLER_30_868 VPWR VGND sg13g2_decap_8
XFILLER_10_592 VPWR VGND sg13g2_decap_8
XFILLER_41_91 VPWR VGND sg13g2_decap_8
XFILLER_6_574 VPWR VGND sg13g2_decap_8
XFILLER_96_301 VPWR VGND sg13g2_decap_8
XFILLER_69_526 VPWR VGND sg13g2_decap_8
XFILLER_37_4 VPWR VGND sg13g2_decap_8
XFILLER_97_868 VPWR VGND sg13g2_decap_8
XFILLER_96_378 VPWR VGND sg13g2_decap_8
XFILLER_84_518 VPWR VGND sg13g2_decap_8
XFILLER_38_924 VPWR VGND sg13g2_decap_8
XFILLER_77_581 VPWR VGND sg13g2_decap_8
XFILLER_65_721 VPWR VGND sg13g2_decap_8
XFILLER_2_74 VPWR VGND sg13g2_decap_8
X_56_ _14_ _18_ _22_ VPWR VGND sg13g2_nor2_1
XFILLER_64_242 VPWR VGND sg13g2_decap_8
XFILLER_37_445 VPWR VGND sg13g2_decap_8
XFILLER_92_595 VPWR VGND sg13g2_decap_8
XFILLER_80_735 VPWR VGND sg13g2_decap_8
XFILLER_65_798 VPWR VGND sg13g2_decap_8
XFILLER_53_938 VPWR VGND sg13g2_decap_8
XFILLER_52_448 VPWR VGND sg13g2_decap_8
XFILLER_33_651 VPWR VGND sg13g2_decap_8
XFILLER_36_1015 VPWR VGND sg13g2_decap_8
XFILLER_20_312 VPWR VGND sg13g2_decap_8
XFILLER_32_172 VPWR VGND sg13g2_decap_8
XFILLER_21_868 VPWR VGND sg13g2_decap_8
XFILLER_20_389 VPWR VGND sg13g2_decap_8
XFILLER_21_28 VPWR VGND sg13g2_decap_8
XFILLER_106_406 VPWR VGND sg13g2_decap_8
XFILLER_88_802 VPWR VGND sg13g2_decap_8
XFILLER_99_161 VPWR VGND sg13g2_decap_8
XFILLER_87_301 VPWR VGND sg13g2_decap_8
XFILLER_0_728 VPWR VGND sg13g2_decap_8
XFILLER_102_623 VPWR VGND sg13g2_decap_8
XFILLER_43_1008 VPWR VGND sg13g2_decap_8
XFILLER_101_133 VPWR VGND sg13g2_decap_8
XFILLER_88_879 VPWR VGND sg13g2_decap_8
XFILLER_87_378 VPWR VGND sg13g2_decap_8
XFILLER_75_518 VPWR VGND sg13g2_decap_8
XFILLER_56_732 VPWR VGND sg13g2_decap_8
XFILLER_46_25 VPWR VGND sg13g2_decap_8
XFILLER_29_935 VPWR VGND sg13g2_decap_8
XFILLER_55_231 VPWR VGND sg13g2_decap_8
XFILLER_28_434 VPWR VGND sg13g2_decap_8
XFILLER_44_949 VPWR VGND sg13g2_decap_8
XFILLER_102_42 VPWR VGND sg13g2_decap_8
XFILLER_71_746 VPWR VGND sg13g2_decap_8
XFILLER_70_245 VPWR VGND sg13g2_decap_8
XFILLER_43_448 VPWR VGND sg13g2_decap_8
XFILLER_62_35 VPWR VGND sg13g2_decap_8
XFILLER_12_802 VPWR VGND sg13g2_decap_8
XFILLER_24_662 VPWR VGND sg13g2_decap_8
XFILLER_11_301 VPWR VGND sg13g2_decap_8
XFILLER_23_161 VPWR VGND sg13g2_decap_8
XFILLER_7_305 VPWR VGND sg13g2_decap_8
XFILLER_12_879 VPWR VGND sg13g2_decap_8
XFILLER_11_378 VPWR VGND sg13g2_decap_8
XFILLER_3_511 VPWR VGND sg13g2_decap_8
XFILLER_106_973 VPWR VGND sg13g2_decap_8
XFILLER_87_21 VPWR VGND sg13g2_decap_8
XFILLER_79_802 VPWR VGND sg13g2_decap_8
XFILLER_3_588 VPWR VGND sg13g2_decap_8
XFILLER_105_483 VPWR VGND sg13g2_decap_8
XFILLER_94_805 VPWR VGND sg13g2_decap_8
XFILLER_87_98 VPWR VGND sg13g2_decap_8
XFILLER_79_879 VPWR VGND sg13g2_decap_8
XFILLER_78_356 VPWR VGND sg13g2_decap_8
XFILLER_47_721 VPWR VGND sg13g2_decap_8
XFILLER_93_348 VPWR VGND sg13g2_decap_8
XFILLER_74_540 VPWR VGND sg13g2_decap_8
XFILLER_46_242 VPWR VGND sg13g2_decap_8
XFILLER_19_434 VPWR VGND sg13g2_decap_8
XFILLER_47_798 VPWR VGND sg13g2_decap_8
XFILLER_35_938 VPWR VGND sg13g2_decap_8
XFILLER_62_735 VPWR VGND sg13g2_decap_8
XFILLER_34_459 VPWR VGND sg13g2_decap_8
XFILLER_36_91 VPWR VGND sg13g2_decap_8
XFILLER_61_256 VPWR VGND sg13g2_decap_8
XFILLER_15_662 VPWR VGND sg13g2_decap_8
XFILLER_14_161 VPWR VGND sg13g2_decap_8
XFILLER_30_665 VPWR VGND sg13g2_decap_8
Xinput11 uio_in[2] net11 VPWR VGND sg13g2_buf_1
XFILLER_7_872 VPWR VGND sg13g2_decap_8
XFILLER_6_371 VPWR VGND sg13g2_decap_8
XFILLER_88_109 VPWR VGND sg13g2_decap_8
XFILLER_69_323 VPWR VGND sg13g2_decap_8
XFILLER_97_665 VPWR VGND sg13g2_decap_8
XFILLER_85_805 VPWR VGND sg13g2_decap_8
XFILLER_57_518 VPWR VGND sg13g2_decap_8
XFILLER_28_0 VPWR VGND sg13g2_decap_8
XFILLER_96_175 VPWR VGND sg13g2_decap_8
XFILLER_84_315 VPWR VGND sg13g2_decap_8
XFILLER_38_721 VPWR VGND sg13g2_decap_8
XFILLER_37_242 VPWR VGND sg13g2_decap_8
X_39_ net4 net12 _08_ VPWR VGND sg13g2_and2_1
XFILLER_26_938 VPWR VGND sg13g2_decap_8
XFILLER_38_798 VPWR VGND sg13g2_decap_8
XFILLER_92_392 VPWR VGND sg13g2_decap_8
XFILLER_80_532 VPWR VGND sg13g2_decap_8
XFILLER_65_595 VPWR VGND sg13g2_decap_8
XFILLER_53_735 VPWR VGND sg13g2_decap_8
XFILLER_16_28 VPWR VGND sg13g2_decap_8
XFILLER_25_448 VPWR VGND sg13g2_decap_8
XFILLER_52_245 VPWR VGND sg13g2_decap_8
XFILLER_12_109 VPWR VGND sg13g2_decap_8
Xheichips25_example_large_40 VPWR VGND uio_out[7] sg13g2_tielo
XFILLER_21_665 VPWR VGND sg13g2_decap_8
XFILLER_5_809 VPWR VGND sg13g2_decap_8
XFILLER_20_186 VPWR VGND sg13g2_decap_8
XFILLER_106_203 VPWR VGND sg13g2_decap_8
XFILLER_4_308 VPWR VGND sg13g2_decap_8
XFILLER_106_7 VPWR VGND sg13g2_decap_8
XFILLER_103_910 VPWR VGND sg13g2_decap_8
XFILLER_79_109 VPWR VGND sg13g2_decap_8
XFILLER_102_420 VPWR VGND sg13g2_decap_8
XFILLER_0_525 VPWR VGND sg13g2_decap_8
XFILLER_103_987 VPWR VGND sg13g2_decap_8
XFILLER_88_676 VPWR VGND sg13g2_decap_8
XFILLER_76_816 VPWR VGND sg13g2_decap_8
XFILLER_57_35 VPWR VGND sg13g2_decap_8
XFILLER_48_518 VPWR VGND sg13g2_decap_8
XFILLER_102_497 VPWR VGND sg13g2_decap_8
XFILLER_87_175 VPWR VGND sg13g2_decap_8
XFILLER_75_315 VPWR VGND sg13g2_decap_8
XFILLER_69_890 VPWR VGND sg13g2_decap_8
XFILLER_91_819 VPWR VGND sg13g2_decap_8
XFILLER_28_231 VPWR VGND sg13g2_decap_8
XFILLER_29_732 VPWR VGND sg13g2_decap_8
XFILLER_84_882 VPWR VGND sg13g2_decap_8
XFILLER_71_543 VPWR VGND sg13g2_decap_8
XFILLER_44_746 VPWR VGND sg13g2_decap_8
XFILLER_16_448 VPWR VGND sg13g2_decap_8
XFILLER_17_949 VPWR VGND sg13g2_decap_8
XFILLER_73_67 VPWR VGND sg13g2_decap_8
XFILLER_43_245 VPWR VGND sg13g2_decap_8
XFILLER_40_952 VPWR VGND sg13g2_decap_8
XFILLER_89_1008 VPWR VGND sg13g2_decap_8
XFILLER_7_102 VPWR VGND sg13g2_decap_8
XFILLER_12_676 VPWR VGND sg13g2_decap_8
XFILLER_8_658 VPWR VGND sg13g2_decap_8
XFILLER_11_175 VPWR VGND sg13g2_decap_8
XFILLER_22_60 VPWR VGND sg13g2_decap_8
XFILLER_7_179 VPWR VGND sg13g2_decap_8
XFILLER_98_53 VPWR VGND sg13g2_decap_8
XFILLER_106_770 VPWR VGND sg13g2_decap_8
XFILLER_4_875 VPWR VGND sg13g2_decap_8
XFILLER_105_280 VPWR VGND sg13g2_decap_8
XFILLER_3_385 VPWR VGND sg13g2_decap_8
XFILLER_94_602 VPWR VGND sg13g2_decap_8
XFILLER_79_676 VPWR VGND sg13g2_decap_8
XFILLER_78_153 VPWR VGND sg13g2_decap_8
XFILLER_67_805 VPWR VGND sg13g2_decap_8
XFILLER_21_7 VPWR VGND sg13g2_decap_8
XFILLER_39_529 VPWR VGND sg13g2_decap_8
XFILLER_94_679 VPWR VGND sg13g2_decap_8
XFILLER_93_145 VPWR VGND sg13g2_decap_8
XFILLER_82_819 VPWR VGND sg13g2_decap_8
XFILLER_19_231 VPWR VGND sg13g2_decap_8
XFILLER_75_882 VPWR VGND sg13g2_decap_8
XFILLER_90_830 VPWR VGND sg13g2_decap_8
XFILLER_62_532 VPWR VGND sg13g2_decap_8
XFILLER_47_595 VPWR VGND sg13g2_decap_8
XFILLER_35_735 VPWR VGND sg13g2_decap_8
XFILLER_34_256 VPWR VGND sg13g2_decap_8
XFILLER_72_1001 VPWR VGND sg13g2_decap_8
XFILLER_50_749 VPWR VGND sg13g2_decap_8
XFILLER_31_952 VPWR VGND sg13g2_decap_8
XFILLER_30_462 VPWR VGND sg13g2_decap_8
XFILLER_8_84 VPWR VGND sg13g2_decap_8
XFILLER_104_707 VPWR VGND sg13g2_decap_8
XFILLER_103_217 VPWR VGND sg13g2_decap_8
XFILLER_98_963 VPWR VGND sg13g2_decap_8
XFILLER_97_462 VPWR VGND sg13g2_decap_8
XFILLER_85_602 VPWR VGND sg13g2_decap_8
XFILLER_69_120 VPWR VGND sg13g2_decap_8
XFILLER_58_805 VPWR VGND sg13g2_decap_8
XFILLER_100_924 VPWR VGND sg13g2_decap_8
XFILLER_84_112 VPWR VGND sg13g2_decap_8
XFILLER_57_315 VPWR VGND sg13g2_decap_8
XFILLER_69_197 VPWR VGND sg13g2_decap_8
XFILLER_85_679 VPWR VGND sg13g2_decap_8
XFILLER_72_329 VPWR VGND sg13g2_decap_8
XFILLER_66_860 VPWR VGND sg13g2_decap_8
XFILLER_84_189 VPWR VGND sg13g2_decap_8
XFILLER_81_830 VPWR VGND sg13g2_decap_8
XFILLER_65_392 VPWR VGND sg13g2_decap_8
XFILLER_53_532 VPWR VGND sg13g2_decap_8
XFILLER_26_735 VPWR VGND sg13g2_decap_8
XFILLER_38_595 VPWR VGND sg13g2_decap_8
XFILLER_25_245 VPWR VGND sg13g2_decap_8
XFILLER_41_749 VPWR VGND sg13g2_decap_8
XFILLER_22_963 VPWR VGND sg13g2_decap_8
XFILLER_40_259 VPWR VGND sg13g2_decap_8
XFILLER_21_462 VPWR VGND sg13g2_decap_8
XFILLER_5_606 VPWR VGND sg13g2_decap_8
XFILLER_4_105 VPWR VGND sg13g2_decap_8
XFILLER_1_812 VPWR VGND sg13g2_decap_8
XFILLER_89_952 VPWR VGND sg13g2_decap_8
XFILLER_49_816 VPWR VGND sg13g2_decap_8
XFILLER_0_322 VPWR VGND sg13g2_decap_8
XFILLER_103_784 VPWR VGND sg13g2_decap_8
XFILLER_88_473 VPWR VGND sg13g2_decap_8
XFILLER_76_613 VPWR VGND sg13g2_decap_8
XFILLER_75_112 VPWR VGND sg13g2_decap_8
XFILLER_68_89 VPWR VGND sg13g2_decap_8
XFILLER_48_315 VPWR VGND sg13g2_decap_8
XFILLER_1_889 VPWR VGND sg13g2_decap_8
XFILLER_102_294 VPWR VGND sg13g2_decap_8
XFILLER_0_399 VPWR VGND sg13g2_decap_8
XFILLER_91_616 VPWR VGND sg13g2_decap_8
XFILLER_57_882 VPWR VGND sg13g2_decap_8
XFILLER_95_1012 VPWR VGND sg13g2_decap_8
XFILLER_90_137 VPWR VGND sg13g2_decap_8
XFILLER_84_77 VPWR VGND sg13g2_decap_8
XFILLER_75_189 VPWR VGND sg13g2_decap_8
XFILLER_63_329 VPWR VGND sg13g2_decap_8
XFILLER_17_746 VPWR VGND sg13g2_decap_8
XFILLER_71_340 VPWR VGND sg13g2_decap_8
XFILLER_44_543 VPWR VGND sg13g2_decap_8
XFILLER_16_245 VPWR VGND sg13g2_decap_8
XFILLER_17_60 VPWR VGND sg13g2_decap_8
XFILLER_72_896 VPWR VGND sg13g2_decap_8
XFILLER_13_952 VPWR VGND sg13g2_decap_8
XFILLER_31_259 VPWR VGND sg13g2_decap_8
XFILLER_9_945 VPWR VGND sg13g2_decap_8
XFILLER_12_473 VPWR VGND sg13g2_decap_8
XFILLER_33_70 VPWR VGND sg13g2_decap_8
XFILLER_8_455 VPWR VGND sg13g2_decap_8
XFILLER_69_7 VPWR VGND sg13g2_decap_8
XFILLER_99_749 VPWR VGND sg13g2_decap_8
XFILLER_4_672 VPWR VGND sg13g2_decap_8
XFILLER_95_900 VPWR VGND sg13g2_decap_8
XFILLER_3_182 VPWR VGND sg13g2_decap_8
XFILLER_79_473 VPWR VGND sg13g2_decap_8
XFILLER_67_602 VPWR VGND sg13g2_decap_8
XFILLER_39_326 VPWR VGND sg13g2_decap_8
XFILLER_95_977 VPWR VGND sg13g2_decap_8
XFILLER_94_476 VPWR VGND sg13g2_decap_8
XFILLER_82_616 VPWR VGND sg13g2_decap_8
XFILLER_67_679 VPWR VGND sg13g2_decap_8
XFILLER_66_167 VPWR VGND sg13g2_decap_8
XFILLER_55_819 VPWR VGND sg13g2_decap_8
XFILLER_48_882 VPWR VGND sg13g2_decap_8
XFILLER_81_137 VPWR VGND sg13g2_decap_8
XFILLER_47_392 VPWR VGND sg13g2_decap_8
XFILLER_35_532 VPWR VGND sg13g2_decap_8
XFILLER_63_896 VPWR VGND sg13g2_decap_8
XFILLER_23_749 VPWR VGND sg13g2_decap_8
XFILLER_50_546 VPWR VGND sg13g2_decap_8
XFILLER_104_504 VPWR VGND sg13g2_decap_8
XFILLER_1_119 VPWR VGND sg13g2_decap_8
XFILLER_98_760 VPWR VGND sg13g2_decap_8
XFILLER_89_259 VPWR VGND sg13g2_decap_8
XFILLER_86_900 VPWR VGND sg13g2_decap_8
XFILLER_100_721 VPWR VGND sg13g2_decap_8
XFILLER_58_602 VPWR VGND sg13g2_decap_8
XFILLER_86_977 VPWR VGND sg13g2_decap_8
XFILLER_57_112 VPWR VGND sg13g2_decap_8
XFILLER_85_476 VPWR VGND sg13g2_decap_8
XFILLER_73_627 VPWR VGND sg13g2_decap_8
XFILLER_58_679 VPWR VGND sg13g2_decap_8
XFILLER_100_798 VPWR VGND sg13g2_decap_8
XFILLER_72_126 VPWR VGND sg13g2_decap_8
XFILLER_57_189 VPWR VGND sg13g2_decap_8
XFILLER_54_830 VPWR VGND sg13g2_decap_8
XFILLER_45_329 VPWR VGND sg13g2_decap_8
XFILLER_26_532 VPWR VGND sg13g2_decap_8
XFILLER_39_893 VPWR VGND sg13g2_decap_8
XFILLER_54_25 VPWR VGND sg13g2_decap_8
XFILLER_38_392 VPWR VGND sg13g2_decap_8
XFILLER_14_749 VPWR VGND sg13g2_decap_8
XFILLER_41_546 VPWR VGND sg13g2_decap_8
XFILLER_70_35 VPWR VGND sg13g2_decap_8
XFILLER_10_900 VPWR VGND sg13g2_decap_8
XFILLER_13_259 VPWR VGND sg13g2_decap_8
XFILLER_22_760 VPWR VGND sg13g2_decap_8
XFILLER_5_403 VPWR VGND sg13g2_decap_8
XFILLER_10_977 VPWR VGND sg13g2_decap_8
XFILLER_6_959 VPWR VGND sg13g2_decap_8
XFILLER_79_88 VPWR VGND sg13g2_decap_8
XFILLER_95_207 VPWR VGND sg13g2_decap_8
XFILLER_95_32 VPWR VGND sg13g2_decap_8
XFILLER_88_270 VPWR VGND sg13g2_decap_8
XFILLER_76_410 VPWR VGND sg13g2_decap_8
XFILLER_62_1022 VPWR VGND sg13g2_decap_8
XFILLER_49_613 VPWR VGND sg13g2_decap_8
XFILLER_1_686 VPWR VGND sg13g2_decap_8
XFILLER_103_581 VPWR VGND sg13g2_decap_8
XFILLER_77_966 VPWR VGND sg13g2_decap_8
XFILLER_48_112 VPWR VGND sg13g2_decap_8
XFILLER_0_196 VPWR VGND sg13g2_decap_8
XFILLER_92_903 VPWR VGND sg13g2_decap_8
XFILLER_64_627 VPWR VGND sg13g2_decap_8
XFILLER_91_413 VPWR VGND sg13g2_decap_8
XFILLER_76_487 VPWR VGND sg13g2_decap_8
XFILLER_63_126 VPWR VGND sg13g2_decap_8
XFILLER_48_189 VPWR VGND sg13g2_decap_8
XFILLER_28_70 VPWR VGND sg13g2_decap_8
XFILLER_36_329 VPWR VGND sg13g2_decap_8
XFILLER_44_340 VPWR VGND sg13g2_decap_8
XFILLER_17_543 VPWR VGND sg13g2_decap_8
XFILLER_72_693 VPWR VGND sg13g2_decap_8
XFILLER_45_896 VPWR VGND sg13g2_decap_8
XFILLER_60_844 VPWR VGND sg13g2_decap_8
XFILLER_32_557 VPWR VGND sg13g2_decap_8
XFILLER_9_742 VPWR VGND sg13g2_decap_8
XFILLER_12_270 VPWR VGND sg13g2_decap_8
XFILLER_8_252 VPWR VGND sg13g2_decap_8
XFILLER_99_546 VPWR VGND sg13g2_decap_8
XFILLER_5_970 VPWR VGND sg13g2_decap_8
XFILLER_5_74 VPWR VGND sg13g2_decap_8
XFILLER_101_518 VPWR VGND sg13g2_decap_8
XFILLER_86_207 VPWR VGND sg13g2_decap_8
XFILLER_68_922 VPWR VGND sg13g2_decap_8
XFILLER_79_270 VPWR VGND sg13g2_decap_8
XFILLER_39_123 VPWR VGND sg13g2_decap_8
XFILLER_95_774 VPWR VGND sg13g2_decap_8
XFILLER_83_914 VPWR VGND sg13g2_decap_8
XFILLER_68_999 VPWR VGND sg13g2_decap_8
XFILLER_67_476 VPWR VGND sg13g2_decap_8
XFILLER_55_616 VPWR VGND sg13g2_decap_8
XFILLER_28_819 VPWR VGND sg13g2_decap_8
XFILLER_94_273 VPWR VGND sg13g2_decap_8
XFILLER_82_413 VPWR VGND sg13g2_decap_8
XFILLER_54_137 VPWR VGND sg13g2_decap_8
XFILLER_91_980 VPWR VGND sg13g2_decap_8
XFILLER_36_896 VPWR VGND sg13g2_decap_8
XFILLER_63_693 VPWR VGND sg13g2_decap_8
XFILLER_51_844 VPWR VGND sg13g2_decap_8
XFILLER_50_343 VPWR VGND sg13g2_decap_8
XFILLER_23_546 VPWR VGND sg13g2_decap_8
XFILLER_24_39 VPWR VGND sg13g2_decap_8
XFILLER_10_207 VPWR VGND sg13g2_decap_8
XFILLER_40_49 VPWR VGND sg13g2_decap_8
XFILLER_85_1022 VPWR VGND sg13g2_decap_8
XFILLER_104_301 VPWR VGND sg13g2_decap_8
XFILLER_2_417 VPWR VGND sg13g2_decap_8
XFILLER_105_868 VPWR VGND sg13g2_decap_8
XFILLER_49_25 VPWR VGND sg13g2_decap_8
XFILLER_46_1028 VPWR VGND sg13g2_fill_1
XFILLER_104_378 VPWR VGND sg13g2_decap_8
XFILLER_59_922 VPWR VGND sg13g2_decap_8
XFILLER_105_42 VPWR VGND sg13g2_decap_8
XFILLER_86_774 VPWR VGND sg13g2_decap_8
XFILLER_74_925 VPWR VGND sg13g2_decap_8
XFILLER_59_999 VPWR VGND sg13g2_decap_8
XFILLER_58_476 VPWR VGND sg13g2_decap_8
XFILLER_19_819 VPWR VGND sg13g2_decap_8
XFILLER_100_595 VPWR VGND sg13g2_decap_8
XFILLER_85_273 VPWR VGND sg13g2_decap_8
XFILLER_73_424 VPWR VGND sg13g2_decap_8
XFILLER_65_35 VPWR VGND sg13g2_decap_8
XFILLER_46_627 VPWR VGND sg13g2_decap_8
XFILLER_45_126 VPWR VGND sg13g2_decap_8
XFILLER_18_329 VPWR VGND sg13g2_decap_8
XFILLER_27_830 VPWR VGND sg13g2_decap_8
XFILLER_39_690 VPWR VGND sg13g2_decap_8
XFILLER_92_1015 VPWR VGND sg13g2_decap_8
XFILLER_82_980 VPWR VGND sg13g2_decap_8
XFILLER_42_844 VPWR VGND sg13g2_decap_8
XFILLER_14_546 VPWR VGND sg13g2_decap_8
XFILLER_81_67 VPWR VGND sg13g2_decap_8
XFILLER_41_343 VPWR VGND sg13g2_decap_8
XFILLER_5_200 VPWR VGND sg13g2_decap_8
XFILLER_10_774 VPWR VGND sg13g2_decap_8
XFILLER_6_756 VPWR VGND sg13g2_decap_8
XFILLER_5_277 VPWR VGND sg13g2_decap_8
XFILLER_69_708 VPWR VGND sg13g2_decap_8
XFILLER_68_229 VPWR VGND sg13g2_decap_8
XFILLER_2_984 VPWR VGND sg13g2_decap_8
XFILLER_49_410 VPWR VGND sg13g2_decap_8
XFILLER_1_483 VPWR VGND sg13g2_decap_8
XFILLER_92_700 VPWR VGND sg13g2_decap_8
XFILLER_77_763 VPWR VGND sg13g2_decap_8
XFILLER_65_903 VPWR VGND sg13g2_decap_8
XFILLER_91_210 VPWR VGND sg13g2_decap_8
Xinput9 uio_in[0] net9 VPWR VGND sg13g2_buf_1
XFILLER_76_284 VPWR VGND sg13g2_decap_8
XFILLER_64_424 VPWR VGND sg13g2_decap_8
XFILLER_49_487 VPWR VGND sg13g2_decap_8
XFILLER_36_126 VPWR VGND sg13g2_decap_8
XFILLER_37_627 VPWR VGND sg13g2_decap_8
XFILLER_92_777 VPWR VGND sg13g2_decap_8
XFILLER_80_917 VPWR VGND sg13g2_decap_8
XFILLER_17_340 VPWR VGND sg13g2_decap_8
XFILLER_91_287 VPWR VGND sg13g2_decap_8
XFILLER_73_991 VPWR VGND sg13g2_decap_8
XFILLER_18_896 VPWR VGND sg13g2_decap_8
XFILLER_72_490 VPWR VGND sg13g2_decap_8
XFILLER_60_641 VPWR VGND sg13g2_decap_8
XFILLER_45_693 VPWR VGND sg13g2_decap_8
XFILLER_33_833 VPWR VGND sg13g2_decap_8
XFILLER_32_354 VPWR VGND sg13g2_decap_8
XFILLER_58_0 VPWR VGND sg13g2_decap_8
XFILLER_99_343 VPWR VGND sg13g2_decap_8
XFILLER_102_805 VPWR VGND sg13g2_decap_8
XFILLER_101_315 VPWR VGND sg13g2_decap_8
XFILLER_59_229 VPWR VGND sg13g2_decap_8
XFILLER_19_28 VPWR VGND sg13g2_decap_8
XFILLER_56_914 VPWR VGND sg13g2_decap_8
XFILLER_28_616 VPWR VGND sg13g2_decap_8
XFILLER_95_571 VPWR VGND sg13g2_decap_8
XFILLER_83_711 VPWR VGND sg13g2_decap_8
XFILLER_82_210 VPWR VGND sg13g2_decap_8
XFILLER_68_796 VPWR VGND sg13g2_decap_8
XFILLER_67_273 VPWR VGND sg13g2_decap_8
XFILLER_55_413 VPWR VGND sg13g2_decap_8
XFILLER_27_137 VPWR VGND sg13g2_decap_8
XFILLER_83_788 VPWR VGND sg13g2_decap_8
XFILLER_82_287 VPWR VGND sg13g2_decap_8
XFILLER_71_928 VPWR VGND sg13g2_decap_8
XFILLER_70_427 VPWR VGND sg13g2_decap_8
XFILLER_64_991 VPWR VGND sg13g2_decap_8
XFILLER_35_49 VPWR VGND sg13g2_decap_8
XFILLER_63_490 VPWR VGND sg13g2_decap_8
XFILLER_51_641 VPWR VGND sg13g2_decap_8
XFILLER_24_844 VPWR VGND sg13g2_decap_8
XFILLER_36_693 VPWR VGND sg13g2_decap_8
XFILLER_50_140 VPWR VGND sg13g2_decap_8
XFILLER_23_343 VPWR VGND sg13g2_decap_8
XFILLER_100_1008 VPWR VGND sg13g2_decap_8
XFILLER_2_214 VPWR VGND sg13g2_decap_8
XFILLER_105_665 VPWR VGND sg13g2_decap_8
XFILLER_104_175 VPWR VGND sg13g2_decap_8
XFILLER_78_538 VPWR VGND sg13g2_decap_8
XFILLER_76_67 VPWR VGND sg13g2_decap_8
XFILLER_47_903 VPWR VGND sg13g2_decap_8
XFILLER_101_882 VPWR VGND sg13g2_decap_8
XFILLER_86_571 VPWR VGND sg13g2_decap_8
XFILLER_74_722 VPWR VGND sg13g2_decap_8
XFILLER_59_796 VPWR VGND sg13g2_decap_8
XFILLER_58_273 VPWR VGND sg13g2_decap_8
XFILLER_46_424 VPWR VGND sg13g2_decap_8
XFILLER_19_616 VPWR VGND sg13g2_decap_8
XFILLER_100_392 VPWR VGND sg13g2_decap_8
XFILLER_73_221 VPWR VGND sg13g2_decap_8
XFILLER_62_917 VPWR VGND sg13g2_decap_8
XFILLER_18_126 VPWR VGND sg13g2_decap_8
XFILLER_74_799 VPWR VGND sg13g2_decap_8
XFILLER_55_980 VPWR VGND sg13g2_decap_8
XFILLER_92_77 VPWR VGND sg13g2_decap_8
XFILLER_73_298 VPWR VGND sg13g2_decap_8
XFILLER_61_438 VPWR VGND sg13g2_decap_8
XFILLER_15_844 VPWR VGND sg13g2_decap_8
XFILLER_42_641 VPWR VGND sg13g2_decap_8
XFILLER_14_343 VPWR VGND sg13g2_decap_8
XFILLER_41_140 VPWR VGND sg13g2_decap_8
XFILLER_70_994 VPWR VGND sg13g2_decap_8
XFILLER_30_847 VPWR VGND sg13g2_decap_8
XFILLER_10_571 VPWR VGND sg13g2_decap_8
XFILLER_6_553 VPWR VGND sg13g2_decap_8
XFILLER_41_70 VPWR VGND sg13g2_decap_8
XFILLER_29_1012 VPWR VGND sg13g2_decap_8
XFILLER_69_505 VPWR VGND sg13g2_decap_8
XFILLER_97_847 VPWR VGND sg13g2_decap_8
XFILLER_2_781 VPWR VGND sg13g2_decap_8
XFILLER_96_357 VPWR VGND sg13g2_decap_8
XFILLER_77_560 VPWR VGND sg13g2_decap_8
XFILLER_65_700 VPWR VGND sg13g2_decap_8
XFILLER_1_280 VPWR VGND sg13g2_decap_8
XFILLER_2_53 VPWR VGND sg13g2_decap_8
XFILLER_38_903 VPWR VGND sg13g2_decap_8
XFILLER_49_284 VPWR VGND sg13g2_decap_8
XFILLER_37_424 VPWR VGND sg13g2_decap_8
X_55_ _16_ _19_ _21_ VPWR VGND sg13g2_nor2_1
XFILLER_64_221 VPWR VGND sg13g2_decap_8
XFILLER_92_574 VPWR VGND sg13g2_decap_8
XFILLER_80_714 VPWR VGND sg13g2_decap_8
XFILLER_65_777 VPWR VGND sg13g2_decap_8
XFILLER_53_917 VPWR VGND sg13g2_decap_8
XFILLER_64_298 VPWR VGND sg13g2_decap_8
XFILLER_52_427 VPWR VGND sg13g2_decap_8
XFILLER_46_991 VPWR VGND sg13g2_decap_8
XFILLER_45_490 VPWR VGND sg13g2_decap_8
XFILLER_18_693 VPWR VGND sg13g2_decap_8
XFILLER_33_630 VPWR VGND sg13g2_decap_8
XFILLER_21_847 VPWR VGND sg13g2_decap_8
XFILLER_32_151 VPWR VGND sg13g2_decap_8
XFILLER_20_368 VPWR VGND sg13g2_decap_8
XFILLER_102_602 VPWR VGND sg13g2_decap_8
XFILLER_99_140 VPWR VGND sg13g2_decap_8
XFILLER_0_707 VPWR VGND sg13g2_decap_8
XFILLER_101_112 VPWR VGND sg13g2_decap_8
XFILLER_88_858 VPWR VGND sg13g2_decap_8
XFILLER_102_679 VPWR VGND sg13g2_decap_8
XFILLER_87_357 VPWR VGND sg13g2_decap_8
XFILLER_29_914 VPWR VGND sg13g2_decap_8
XFILLER_101_189 VPWR VGND sg13g2_decap_8
XFILLER_68_593 VPWR VGND sg13g2_decap_8
XFILLER_56_711 VPWR VGND sg13g2_decap_8
XFILLER_28_413 VPWR VGND sg13g2_decap_8
XFILLER_55_210 VPWR VGND sg13g2_decap_8
XFILLER_102_21 VPWR VGND sg13g2_decap_8
XFILLER_83_585 VPWR VGND sg13g2_decap_8
XFILLER_71_725 VPWR VGND sg13g2_decap_8
XFILLER_56_788 VPWR VGND sg13g2_decap_8
XFILLER_44_928 VPWR VGND sg13g2_decap_8
XFILLER_70_224 VPWR VGND sg13g2_decap_8
XFILLER_55_287 VPWR VGND sg13g2_decap_8
XFILLER_43_427 VPWR VGND sg13g2_decap_8
XFILLER_36_490 VPWR VGND sg13g2_decap_8
XFILLER_37_991 VPWR VGND sg13g2_decap_8
XFILLER_62_14 VPWR VGND sg13g2_decap_8
XFILLER_23_140 VPWR VGND sg13g2_decap_8
XFILLER_24_641 VPWR VGND sg13g2_decap_8
XFILLER_102_98 VPWR VGND sg13g2_decap_8
XFILLER_62_69 VPWR VGND sg13g2_decap_8
XFILLER_52_994 VPWR VGND sg13g2_decap_8
XFILLER_11_357 VPWR VGND sg13g2_decap_8
XFILLER_12_858 VPWR VGND sg13g2_decap_8
XFILLER_106_952 VPWR VGND sg13g2_decap_8
XFILLER_11_84 VPWR VGND sg13g2_decap_8
XFILLER_105_462 VPWR VGND sg13g2_decap_8
XFILLER_3_567 VPWR VGND sg13g2_decap_8
XFILLER_87_77 VPWR VGND sg13g2_decap_8
XFILLER_79_858 VPWR VGND sg13g2_decap_8
XFILLER_78_335 VPWR VGND sg13g2_decap_8
XFILLER_93_327 VPWR VGND sg13g2_decap_8
XFILLER_47_700 VPWR VGND sg13g2_decap_8
XFILLER_19_413 VPWR VGND sg13g2_decap_8
XFILLER_59_593 VPWR VGND sg13g2_decap_8
XFILLER_46_221 VPWR VGND sg13g2_decap_8
XFILLER_62_714 VPWR VGND sg13g2_decap_8
XFILLER_59_1027 VPWR VGND sg13g2_fill_2
XFILLER_47_777 VPWR VGND sg13g2_decap_8
XFILLER_28_980 VPWR VGND sg13g2_decap_8
XFILLER_35_917 VPWR VGND sg13g2_decap_8
XFILLER_74_596 VPWR VGND sg13g2_decap_8
XFILLER_61_235 VPWR VGND sg13g2_decap_8
XFILLER_46_298 VPWR VGND sg13g2_decap_8
XFILLER_34_438 VPWR VGND sg13g2_decap_8
XFILLER_36_70 VPWR VGND sg13g2_decap_8
XFILLER_14_140 VPWR VGND sg13g2_decap_8
XFILLER_15_641 VPWR VGND sg13g2_decap_8
XFILLER_99_7 VPWR VGND sg13g2_decap_8
XFILLER_70_791 VPWR VGND sg13g2_decap_8
XFILLER_43_994 VPWR VGND sg13g2_decap_8
XFILLER_30_644 VPWR VGND sg13g2_decap_8
Xinput12 uio_in[3] net12 VPWR VGND sg13g2_buf_1
XFILLER_52_91 VPWR VGND sg13g2_decap_8
XFILLER_7_851 VPWR VGND sg13g2_decap_8
XFILLER_6_350 VPWR VGND sg13g2_decap_8
XFILLER_69_302 VPWR VGND sg13g2_decap_8
XFILLER_97_644 VPWR VGND sg13g2_decap_8
XFILLER_96_154 VPWR VGND sg13g2_decap_8
XFILLER_69_379 VPWR VGND sg13g2_decap_8
XFILLER_38_700 VPWR VGND sg13g2_decap_8
XFILLER_37_221 VPWR VGND sg13g2_decap_8
XFILLER_65_574 VPWR VGND sg13g2_decap_8
X_38_ VGND VPWR _07_ net12 net4 sg13g2_or2_1
XFILLER_53_714 VPWR VGND sg13g2_decap_8
XFILLER_26_917 VPWR VGND sg13g2_decap_8
XFILLER_38_777 VPWR VGND sg13g2_decap_8
XFILLER_93_894 VPWR VGND sg13g2_decap_8
XFILLER_92_371 VPWR VGND sg13g2_decap_8
XFILLER_80_511 VPWR VGND sg13g2_decap_8
XFILLER_52_224 VPWR VGND sg13g2_decap_8
XFILLER_19_980 VPWR VGND sg13g2_decap_8
XFILLER_25_427 VPWR VGND sg13g2_decap_8
XFILLER_37_298 VPWR VGND sg13g2_decap_8
Xheichips25_example_large_30 VPWR VGND uio_oe[5] sg13g2_tielo
XFILLER_18_490 VPWR VGND sg13g2_decap_8
XFILLER_80_588 VPWR VGND sg13g2_decap_8
XFILLER_21_644 VPWR VGND sg13g2_decap_8
XFILLER_20_165 VPWR VGND sg13g2_decap_8
XFILLER_32_39 VPWR VGND sg13g2_decap_8
XFILLER_10_1019 VPWR VGND sg13g2_decap_8
XFILLER_106_259 VPWR VGND sg13g2_decap_8
XFILLER_0_504 VPWR VGND sg13g2_decap_8
XFILLER_103_966 VPWR VGND sg13g2_decap_8
XFILLER_88_655 VPWR VGND sg13g2_decap_8
XFILLER_87_154 VPWR VGND sg13g2_decap_8
XFILLER_57_14 VPWR VGND sg13g2_decap_8
XFILLER_102_476 VPWR VGND sg13g2_decap_8
XFILLER_29_711 VPWR VGND sg13g2_decap_8
XFILLER_68_390 VPWR VGND sg13g2_decap_8
XFILLER_28_210 VPWR VGND sg13g2_decap_8
XFILLER_90_319 VPWR VGND sg13g2_decap_8
XFILLER_84_861 VPWR VGND sg13g2_decap_8
XFILLER_17_928 VPWR VGND sg13g2_decap_8
XFILLER_29_788 VPWR VGND sg13g2_decap_8
XFILLER_83_382 VPWR VGND sg13g2_decap_8
XFILLER_73_46 VPWR VGND sg13g2_decap_8
XFILLER_71_522 VPWR VGND sg13g2_decap_8
XFILLER_56_585 VPWR VGND sg13g2_decap_8
XFILLER_44_725 VPWR VGND sg13g2_decap_8
XFILLER_43_224 VPWR VGND sg13g2_decap_8
XFILLER_16_427 VPWR VGND sg13g2_decap_8
XFILLER_28_287 VPWR VGND sg13g2_decap_8
XFILLER_73_57 VPWR VGND sg13g2_fill_2
XFILLER_71_599 VPWR VGND sg13g2_decap_8
XFILLER_19_1022 VPWR VGND sg13g2_decap_8
XFILLER_25_994 VPWR VGND sg13g2_decap_8
XFILLER_40_931 VPWR VGND sg13g2_decap_8
XFILLER_52_791 VPWR VGND sg13g2_decap_8
XFILLER_12_655 VPWR VGND sg13g2_decap_8
XFILLER_8_637 VPWR VGND sg13g2_decap_8
XFILLER_11_154 VPWR VGND sg13g2_decap_8
XFILLER_7_158 VPWR VGND sg13g2_decap_8
XFILLER_98_32 VPWR VGND sg13g2_decap_8
XFILLER_4_854 VPWR VGND sg13g2_decap_8
XFILLER_3_364 VPWR VGND sg13g2_decap_8
XFILLER_79_655 VPWR VGND sg13g2_decap_8
XFILLER_78_132 VPWR VGND sg13g2_decap_8
XFILLER_26_1015 VPWR VGND sg13g2_decap_8
XFILLER_39_508 VPWR VGND sg13g2_decap_8
XFILLER_94_658 VPWR VGND sg13g2_decap_8
XFILLER_93_124 VPWR VGND sg13g2_decap_8
XFILLER_66_349 VPWR VGND sg13g2_decap_8
XFILLER_59_390 VPWR VGND sg13g2_decap_8
XFILLER_14_7 VPWR VGND sg13g2_decap_8
XFILLER_19_210 VPWR VGND sg13g2_decap_8
XFILLER_81_319 VPWR VGND sg13g2_decap_8
XFILLER_75_861 VPWR VGND sg13g2_decap_8
XFILLER_47_574 VPWR VGND sg13g2_decap_8
XFILLER_47_91 VPWR VGND sg13g2_decap_8
XFILLER_35_714 VPWR VGND sg13g2_decap_8
XFILLER_74_393 VPWR VGND sg13g2_decap_8
XFILLER_62_511 VPWR VGND sg13g2_decap_8
XFILLER_19_287 VPWR VGND sg13g2_decap_8
XFILLER_34_235 VPWR VGND sg13g2_decap_8
XFILLER_90_886 VPWR VGND sg13g2_decap_8
XFILLER_62_588 VPWR VGND sg13g2_decap_8
XFILLER_50_728 VPWR VGND sg13g2_decap_8
XFILLER_16_994 VPWR VGND sg13g2_decap_8
XFILLER_43_791 VPWR VGND sg13g2_decap_8
XFILLER_31_931 VPWR VGND sg13g2_decap_8
XFILLER_33_1008 VPWR VGND sg13g2_decap_8
XFILLER_30_441 VPWR VGND sg13g2_decap_8
XFILLER_8_63 VPWR VGND sg13g2_decap_8
XFILLER_98_942 VPWR VGND sg13g2_decap_8
XFILLER_40_0 VPWR VGND sg13g2_decap_8
XFILLER_100_903 VPWR VGND sg13g2_decap_8
XFILLER_97_441 VPWR VGND sg13g2_decap_8
XFILLER_69_176 VPWR VGND sg13g2_decap_8
XFILLER_85_658 VPWR VGND sg13g2_decap_8
XFILLER_73_809 VPWR VGND sg13g2_decap_8
XFILLER_84_168 VPWR VGND sg13g2_decap_8
XFILLER_72_308 VPWR VGND sg13g2_decap_8
XFILLER_26_714 VPWR VGND sg13g2_decap_8
XFILLER_27_39 VPWR VGND sg13g2_decap_8
XFILLER_38_574 VPWR VGND sg13g2_decap_8
XFILLER_93_691 VPWR VGND sg13g2_decap_8
XFILLER_65_371 VPWR VGND sg13g2_decap_8
XFILLER_53_511 VPWR VGND sg13g2_decap_8
XFILLER_25_224 VPWR VGND sg13g2_decap_8
XFILLER_81_886 VPWR VGND sg13g2_decap_8
XFILLER_80_385 VPWR VGND sg13g2_decap_8
XFILLER_53_588 VPWR VGND sg13g2_decap_8
XFILLER_41_728 VPWR VGND sg13g2_decap_8
XFILLER_43_49 VPWR VGND sg13g2_decap_8
XFILLER_22_942 VPWR VGND sg13g2_decap_8
XFILLER_40_238 VPWR VGND sg13g2_decap_8
XFILLER_21_441 VPWR VGND sg13g2_decap_8
XFILLER_49_1026 VPWR VGND sg13g2_fill_2
XFILLER_89_931 VPWR VGND sg13g2_decap_8
XFILLER_0_301 VPWR VGND sg13g2_decap_8
XFILLER_88_452 VPWR VGND sg13g2_decap_8
XFILLER_68_68 VPWR VGND sg13g2_decap_8
XFILLER_68_46 VPWR VGND sg13g2_decap_4
XFILLER_1_868 VPWR VGND sg13g2_decap_8
XFILLER_103_763 VPWR VGND sg13g2_decap_8
XFILLER_0_378 VPWR VGND sg13g2_decap_8
XFILLER_102_273 VPWR VGND sg13g2_decap_8
XFILLER_76_669 VPWR VGND sg13g2_decap_8
XFILLER_64_809 VPWR VGND sg13g2_decap_8
XFILLER_84_56 VPWR VGND sg13g2_decap_8
XFILLER_75_168 VPWR VGND sg13g2_decap_8
XFILLER_63_308 VPWR VGND sg13g2_decap_8
XFILLER_57_861 VPWR VGND sg13g2_decap_8
XFILLER_90_116 VPWR VGND sg13g2_decap_8
XFILLER_56_382 VPWR VGND sg13g2_decap_8
XFILLER_44_522 VPWR VGND sg13g2_decap_8
XFILLER_16_224 VPWR VGND sg13g2_decap_8
XFILLER_17_725 VPWR VGND sg13g2_decap_8
XFILLER_29_585 VPWR VGND sg13g2_decap_8
XFILLER_72_875 VPWR VGND sg13g2_decap_8
XFILLER_56_1019 VPWR VGND sg13g2_decap_8
XFILLER_44_599 VPWR VGND sg13g2_decap_8
XFILLER_32_739 VPWR VGND sg13g2_decap_8
XFILLER_71_396 VPWR VGND sg13g2_decap_8
XFILLER_13_931 VPWR VGND sg13g2_decap_8
XFILLER_25_791 VPWR VGND sg13g2_decap_8
XFILLER_31_238 VPWR VGND sg13g2_decap_8
XFILLER_9_924 VPWR VGND sg13g2_decap_8
XFILLER_12_452 VPWR VGND sg13g2_decap_8
XFILLER_8_434 VPWR VGND sg13g2_decap_8
XFILLER_99_728 VPWR VGND sg13g2_decap_8
XFILLER_4_651 VPWR VGND sg13g2_decap_8
XFILLER_3_161 VPWR VGND sg13g2_decap_8
XFILLER_98_249 VPWR VGND sg13g2_decap_8
XFILLER_79_452 VPWR VGND sg13g2_decap_8
XFILLER_39_305 VPWR VGND sg13g2_decap_8
XFILLER_95_956 VPWR VGND sg13g2_decap_8
XFILLER_67_658 VPWR VGND sg13g2_decap_8
XFILLER_12_4 VPWR VGND sg13g2_decap_8
XFILLER_94_455 VPWR VGND sg13g2_decap_8
XFILLER_66_146 VPWR VGND sg13g2_decap_8
XFILLER_54_319 VPWR VGND sg13g2_decap_8
XFILLER_48_861 VPWR VGND sg13g2_decap_8
XFILLER_81_116 VPWR VGND sg13g2_decap_8
XFILLER_47_371 VPWR VGND sg13g2_decap_8
XFILLER_35_511 VPWR VGND sg13g2_decap_8
XFILLER_74_190 VPWR VGND sg13g2_decap_8
XFILLER_63_875 VPWR VGND sg13g2_decap_8
XFILLER_90_683 VPWR VGND sg13g2_decap_8
XFILLER_62_385 VPWR VGND sg13g2_decap_8
XFILLER_50_525 VPWR VGND sg13g2_decap_8
XFILLER_23_728 VPWR VGND sg13g2_decap_8
XFILLER_35_588 VPWR VGND sg13g2_decap_8
XFILLER_16_791 VPWR VGND sg13g2_decap_8
XFILLER_22_249 VPWR VGND sg13g2_decap_8
XFILLER_89_238 VPWR VGND sg13g2_decap_8
XFILLER_100_700 VPWR VGND sg13g2_decap_8
XFILLER_86_956 VPWR VGND sg13g2_decap_8
XFILLER_58_658 VPWR VGND sg13g2_decap_8
XFILLER_38_49 VPWR VGND sg13g2_decap_8
XFILLER_100_777 VPWR VGND sg13g2_decap_8
XFILLER_85_455 VPWR VGND sg13g2_decap_8
XFILLER_79_1019 VPWR VGND sg13g2_decap_8
XFILLER_73_606 VPWR VGND sg13g2_decap_8
XFILLER_57_168 VPWR VGND sg13g2_decap_8
XFILLER_46_809 VPWR VGND sg13g2_decap_8
XFILLER_45_308 VPWR VGND sg13g2_decap_8
XFILLER_39_872 VPWR VGND sg13g2_decap_8
XFILLER_72_105 VPWR VGND sg13g2_decap_8
XFILLER_26_511 VPWR VGND sg13g2_decap_8
XFILLER_38_371 VPWR VGND sg13g2_decap_8
XFILLER_81_683 VPWR VGND sg13g2_decap_8
XFILLER_54_886 VPWR VGND sg13g2_decap_8
XFILLER_14_728 VPWR VGND sg13g2_decap_8
XFILLER_26_588 VPWR VGND sg13g2_decap_8
XFILLER_41_525 VPWR VGND sg13g2_decap_8
XFILLER_80_182 VPWR VGND sg13g2_decap_8
XFILLER_53_385 VPWR VGND sg13g2_decap_8
XFILLER_13_238 VPWR VGND sg13g2_decap_8
XFILLER_70_14 VPWR VGND sg13g2_decap_8
XFILLER_10_956 VPWR VGND sg13g2_decap_8
XFILLER_6_938 VPWR VGND sg13g2_decap_8
XFILLER_5_459 VPWR VGND sg13g2_decap_8
XFILLER_79_67 VPWR VGND sg13g2_decap_8
XFILLER_79_56 VPWR VGND sg13g2_fill_2
XFILLER_62_1001 VPWR VGND sg13g2_decap_8
XFILLER_103_560 VPWR VGND sg13g2_decap_8
XFILLER_95_11 VPWR VGND sg13g2_decap_8
XFILLER_1_665 VPWR VGND sg13g2_decap_8
XFILLER_77_945 VPWR VGND sg13g2_decap_8
XFILLER_0_175 VPWR VGND sg13g2_decap_8
XFILLER_95_88 VPWR VGND sg13g2_decap_8
XFILLER_76_466 VPWR VGND sg13g2_decap_8
XFILLER_64_606 VPWR VGND sg13g2_decap_8
XFILLER_49_669 VPWR VGND sg13g2_decap_8
XFILLER_48_168 VPWR VGND sg13g2_decap_8
XFILLER_36_308 VPWR VGND sg13g2_decap_8
XFILLER_37_809 VPWR VGND sg13g2_decap_8
XFILLER_92_959 VPWR VGND sg13g2_decap_8
XFILLER_63_105 VPWR VGND sg13g2_decap_8
XFILLER_17_522 VPWR VGND sg13g2_decap_8
XFILLER_29_382 VPWR VGND sg13g2_decap_8
XFILLER_91_469 VPWR VGND sg13g2_decap_8
XFILLER_72_672 VPWR VGND sg13g2_decap_8
XFILLER_60_823 VPWR VGND sg13g2_decap_8
XFILLER_45_875 VPWR VGND sg13g2_decap_8
XFILLER_71_193 VPWR VGND sg13g2_decap_8
XFILLER_44_396 VPWR VGND sg13g2_decap_8
XFILLER_17_599 VPWR VGND sg13g2_decap_8
XFILLER_32_536 VPWR VGND sg13g2_decap_8
XFILLER_44_81 VPWR VGND sg13g2_decap_8
XFILLER_9_721 VPWR VGND sg13g2_decap_8
XFILLER_8_231 VPWR VGND sg13g2_decap_8
XFILLER_9_798 VPWR VGND sg13g2_decap_8
XFILLER_99_525 VPWR VGND sg13g2_decap_8
XFILLER_5_53 VPWR VGND sg13g2_decap_8
XFILLER_68_901 VPWR VGND sg13g2_decap_8
XFILLER_39_102 VPWR VGND sg13g2_decap_8
XFILLER_95_753 VPWR VGND sg13g2_decap_8
XFILLER_94_252 VPWR VGND sg13g2_decap_8
XFILLER_68_978 VPWR VGND sg13g2_decap_8
XFILLER_67_455 VPWR VGND sg13g2_decap_8
XFILLER_54_116 VPWR VGND sg13g2_decap_8
XFILLER_27_319 VPWR VGND sg13g2_decap_8
XFILLER_39_179 VPWR VGND sg13g2_decap_8
XFILLER_82_469 VPWR VGND sg13g2_decap_8
XFILLER_70_609 VPWR VGND sg13g2_decap_8
XFILLER_63_672 VPWR VGND sg13g2_decap_8
XFILLER_51_823 VPWR VGND sg13g2_decap_8
XFILLER_36_875 VPWR VGND sg13g2_decap_8
XFILLER_90_480 VPWR VGND sg13g2_decap_8
XFILLER_62_182 VPWR VGND sg13g2_decap_8
XFILLER_50_322 VPWR VGND sg13g2_decap_8
XFILLER_23_525 VPWR VGND sg13g2_decap_8
XFILLER_24_18 VPWR VGND sg13g2_decap_8
XFILLER_35_385 VPWR VGND sg13g2_decap_8
XFILLER_50_399 VPWR VGND sg13g2_decap_8
XFILLER_40_28 VPWR VGND sg13g2_decap_8
XFILLER_85_1001 VPWR VGND sg13g2_decap_8
XFILLER_105_847 VPWR VGND sg13g2_decap_8
XFILLER_104_357 VPWR VGND sg13g2_decap_8
XFILLER_59_901 VPWR VGND sg13g2_decap_8
XFILLER_105_21 VPWR VGND sg13g2_decap_8
XFILLER_86_753 VPWR VGND sg13g2_decap_8
XFILLER_85_252 VPWR VGND sg13g2_decap_8
XFILLER_74_904 VPWR VGND sg13g2_decap_8
XFILLER_65_14 VPWR VGND sg13g2_decap_8
XFILLER_59_978 VPWR VGND sg13g2_decap_8
XFILLER_58_455 VPWR VGND sg13g2_decap_8
XFILLER_46_606 VPWR VGND sg13g2_decap_8
XFILLER_18_308 VPWR VGND sg13g2_decap_8
XFILLER_105_98 VPWR VGND sg13g2_decap_8
XFILLER_100_574 VPWR VGND sg13g2_decap_8
XFILLER_73_403 VPWR VGND sg13g2_decap_8
XFILLER_45_105 VPWR VGND sg13g2_decap_8
XFILLER_54_683 VPWR VGND sg13g2_decap_8
XFILLER_42_823 VPWR VGND sg13g2_decap_8
XFILLER_27_886 VPWR VGND sg13g2_decap_8
XFILLER_81_480 VPWR VGND sg13g2_decap_8
XFILLER_53_182 VPWR VGND sg13g2_decap_8
XFILLER_14_525 VPWR VGND sg13g2_decap_8
XFILLER_26_385 VPWR VGND sg13g2_decap_8
XFILLER_41_322 VPWR VGND sg13g2_decap_8
XFILLER_81_46 VPWR VGND sg13g2_decap_8
XFILLER_41_399 VPWR VGND sg13g2_decap_8
XFILLER_10_753 VPWR VGND sg13g2_decap_8
XFILLER_14_84 VPWR VGND sg13g2_decap_8
XFILLER_6_735 VPWR VGND sg13g2_decap_8
XFILLER_5_256 VPWR VGND sg13g2_decap_8
XFILLER_68_208 VPWR VGND sg13g2_decap_8
XFILLER_2_963 VPWR VGND sg13g2_decap_8
XFILLER_1_462 VPWR VGND sg13g2_decap_8
XFILLER_96_539 VPWR VGND sg13g2_decap_8
XFILLER_77_742 VPWR VGND sg13g2_decap_8
XFILLER_7_1012 VPWR VGND sg13g2_decap_8
XFILLER_49_466 VPWR VGND sg13g2_decap_8
XFILLER_37_606 VPWR VGND sg13g2_decap_8
XFILLER_39_81 VPWR VGND sg13g2_decap_8
XFILLER_76_263 VPWR VGND sg13g2_decap_8
XFILLER_65_959 VPWR VGND sg13g2_decap_8
XFILLER_64_403 VPWR VGND sg13g2_decap_8
XFILLER_36_105 VPWR VGND sg13g2_decap_8
XFILLER_92_756 VPWR VGND sg13g2_decap_8
XFILLER_52_609 VPWR VGND sg13g2_decap_8
XFILLER_91_266 VPWR VGND sg13g2_decap_8
XFILLER_73_970 VPWR VGND sg13g2_decap_8
XFILLER_45_672 VPWR VGND sg13g2_decap_8
XFILLER_18_875 VPWR VGND sg13g2_decap_8
XFILLER_33_812 VPWR VGND sg13g2_decap_8
XFILLER_60_620 VPWR VGND sg13g2_decap_8
XFILLER_55_91 VPWR VGND sg13g2_decap_8
XFILLER_17_396 VPWR VGND sg13g2_decap_8
XFILLER_44_193 VPWR VGND sg13g2_decap_8
XFILLER_32_333 VPWR VGND sg13g2_decap_8
XFILLER_33_889 VPWR VGND sg13g2_decap_8
XFILLER_60_697 VPWR VGND sg13g2_decap_8
XFILLER_9_595 VPWR VGND sg13g2_decap_8
XFILLER_99_322 VPWR VGND sg13g2_decap_8
XFILLER_59_208 VPWR VGND sg13g2_decap_8
XFILLER_99_399 VPWR VGND sg13g2_decap_8
XFILLER_87_539 VPWR VGND sg13g2_decap_8
XFILLER_95_550 VPWR VGND sg13g2_decap_8
XFILLER_68_775 VPWR VGND sg13g2_decap_8
XFILLER_67_252 VPWR VGND sg13g2_decap_8
XFILLER_27_116 VPWR VGND sg13g2_decap_8
XFILLER_83_767 VPWR VGND sg13g2_decap_8
XFILLER_71_907 VPWR VGND sg13g2_decap_8
XFILLER_82_266 VPWR VGND sg13g2_decap_8
XFILLER_70_406 VPWR VGND sg13g2_decap_8
XFILLER_64_970 VPWR VGND sg13g2_decap_8
XFILLER_55_469 VPWR VGND sg13g2_decap_8
XFILLER_43_609 VPWR VGND sg13g2_decap_8
XFILLER_35_28 VPWR VGND sg13g2_decap_8
XFILLER_36_672 VPWR VGND sg13g2_decap_8
XFILLER_51_620 VPWR VGND sg13g2_decap_8
XFILLER_23_322 VPWR VGND sg13g2_decap_8
XFILLER_24_823 VPWR VGND sg13g2_decap_8
XFILLER_35_182 VPWR VGND sg13g2_decap_8
XFILLER_52_1022 VPWR VGND sg13g2_decap_8
XFILLER_51_697 VPWR VGND sg13g2_decap_8
XFILLER_11_539 VPWR VGND sg13g2_decap_8
XFILLER_23_399 VPWR VGND sg13g2_decap_8
XFILLER_50_196 VPWR VGND sg13g2_decap_8
XFILLER_105_644 VPWR VGND sg13g2_decap_8
XFILLER_3_749 VPWR VGND sg13g2_decap_8
XFILLER_104_154 VPWR VGND sg13g2_decap_8
XFILLER_78_517 VPWR VGND sg13g2_decap_8
XFILLER_101_861 VPWR VGND sg13g2_decap_8
XFILLER_93_509 VPWR VGND sg13g2_decap_8
XFILLER_86_550 VPWR VGND sg13g2_decap_8
XFILLER_76_46 VPWR VGND sg13g2_decap_8
XFILLER_59_775 VPWR VGND sg13g2_decap_8
XFILLER_100_371 VPWR VGND sg13g2_decap_8
XFILLER_74_701 VPWR VGND sg13g2_decap_8
XFILLER_73_200 VPWR VGND sg13g2_decap_8
XFILLER_58_252 VPWR VGND sg13g2_decap_8
XFILLER_46_403 VPWR VGND sg13g2_decap_8
XFILLER_18_105 VPWR VGND sg13g2_decap_8
XFILLER_47_959 VPWR VGND sg13g2_decap_8
XFILLER_74_778 VPWR VGND sg13g2_decap_8
XFILLER_73_277 VPWR VGND sg13g2_decap_8
XFILLER_61_417 VPWR VGND sg13g2_decap_8
XFILLER_92_56 VPWR VGND sg13g2_decap_8
XFILLER_54_480 VPWR VGND sg13g2_decap_8
XFILLER_42_620 VPWR VGND sg13g2_decap_8
XFILLER_14_322 VPWR VGND sg13g2_decap_8
XFILLER_15_823 VPWR VGND sg13g2_decap_8
XFILLER_26_182 VPWR VGND sg13g2_decap_8
XFILLER_27_683 VPWR VGND sg13g2_decap_8
XFILLER_33_119 VPWR VGND sg13g2_decap_8
XFILLER_70_973 VPWR VGND sg13g2_decap_8
XFILLER_42_697 VPWR VGND sg13g2_decap_8
XFILLER_14_399 VPWR VGND sg13g2_decap_8
XFILLER_30_826 VPWR VGND sg13g2_decap_8
XFILLER_41_196 VPWR VGND sg13g2_decap_8
XFILLER_10_550 VPWR VGND sg13g2_decap_8
XFILLER_6_532 VPWR VGND sg13g2_decap_8
XFILLER_97_826 VPWR VGND sg13g2_decap_8
XFILLER_2_760 VPWR VGND sg13g2_decap_8
XFILLER_96_336 VPWR VGND sg13g2_decap_8
XFILLER_2_32 VPWR VGND sg13g2_decap_8
XFILLER_64_200 VPWR VGND sg13g2_decap_8
XFILLER_49_263 VPWR VGND sg13g2_decap_8
XFILLER_37_403 VPWR VGND sg13g2_decap_8
XFILLER_66_90 VPWR VGND sg13g2_decap_8
X_54_ net22 _19_ _20_ VPWR VGND sg13g2_xnor2_1
XFILLER_65_756 VPWR VGND sg13g2_decap_8
XFILLER_38_959 VPWR VGND sg13g2_decap_8
XFILLER_92_553 VPWR VGND sg13g2_decap_8
XFILLER_64_277 VPWR VGND sg13g2_decap_8
XFILLER_52_406 VPWR VGND sg13g2_decap_8
XFILLER_46_970 VPWR VGND sg13g2_decap_8
XFILLER_18_672 VPWR VGND sg13g2_decap_8
XFILLER_25_609 VPWR VGND sg13g2_decap_8
XFILLER_75_1022 VPWR VGND sg13g2_decap_8
XFILLER_17_193 VPWR VGND sg13g2_decap_8
XFILLER_32_130 VPWR VGND sg13g2_decap_8
XFILLER_61_984 VPWR VGND sg13g2_decap_8
XFILLER_21_826 VPWR VGND sg13g2_decap_8
XFILLER_33_686 VPWR VGND sg13g2_decap_8
XFILLER_60_494 VPWR VGND sg13g2_decap_8
XFILLER_20_347 VPWR VGND sg13g2_decap_8
XFILLER_70_0 VPWR VGND sg13g2_decap_8
XFILLER_9_392 VPWR VGND sg13g2_decap_8
XFILLER_82_1015 VPWR VGND sg13g2_decap_8
XFILLER_99_196 VPWR VGND sg13g2_decap_8
XFILLER_88_837 VPWR VGND sg13g2_decap_8
XFILLER_87_336 VPWR VGND sg13g2_decap_8
XFILLER_102_658 VPWR VGND sg13g2_decap_8
XFILLER_101_168 VPWR VGND sg13g2_decap_8
XFILLER_68_572 VPWR VGND sg13g2_decap_8
XFILLER_56_767 VPWR VGND sg13g2_decap_8
XFILLER_44_907 VPWR VGND sg13g2_decap_8
XFILLER_83_564 VPWR VGND sg13g2_decap_8
XFILLER_71_704 VPWR VGND sg13g2_decap_8
XFILLER_55_266 VPWR VGND sg13g2_decap_8
XFILLER_43_406 VPWR VGND sg13g2_decap_8
XFILLER_16_609 VPWR VGND sg13g2_decap_8
XFILLER_28_469 VPWR VGND sg13g2_decap_8
XFILLER_37_970 VPWR VGND sg13g2_decap_8
XFILLER_70_203 VPWR VGND sg13g2_decap_8
XFILLER_24_620 VPWR VGND sg13g2_decap_8
XFILLER_102_77 VPWR VGND sg13g2_decap_8
XFILLER_52_973 VPWR VGND sg13g2_decap_8
XFILLER_12_837 VPWR VGND sg13g2_decap_8
XFILLER_24_697 VPWR VGND sg13g2_decap_8
XFILLER_51_494 VPWR VGND sg13g2_decap_8
XFILLER_8_819 VPWR VGND sg13g2_decap_8
XFILLER_11_336 VPWR VGND sg13g2_decap_8
XFILLER_23_196 VPWR VGND sg13g2_decap_8
XFILLER_106_931 VPWR VGND sg13g2_decap_8
XFILLER_3_546 VPWR VGND sg13g2_decap_8
XFILLER_11_63 VPWR VGND sg13g2_decap_8
XFILLER_105_441 VPWR VGND sg13g2_decap_8
XFILLER_87_56 VPWR VGND sg13g2_decap_8
XFILLER_79_837 VPWR VGND sg13g2_decap_8
XFILLER_78_314 VPWR VGND sg13g2_decap_8
XFILLER_93_306 VPWR VGND sg13g2_decap_8
XFILLER_59_572 VPWR VGND sg13g2_decap_8
XFILLER_46_200 VPWR VGND sg13g2_decap_8
XFILLER_4_1015 VPWR VGND sg13g2_decap_8
XFILLER_47_756 VPWR VGND sg13g2_decap_8
XFILLER_74_575 VPWR VGND sg13g2_decap_8
XFILLER_59_1006 VPWR VGND sg13g2_decap_8
XFILLER_19_469 VPWR VGND sg13g2_decap_8
XFILLER_61_214 VPWR VGND sg13g2_decap_8
XFILLER_46_277 VPWR VGND sg13g2_decap_8
XFILLER_15_620 VPWR VGND sg13g2_decap_8
XFILLER_27_480 VPWR VGND sg13g2_decap_8
XFILLER_34_417 VPWR VGND sg13g2_decap_8
XFILLER_43_973 VPWR VGND sg13g2_decap_8
XFILLER_70_770 VPWR VGND sg13g2_decap_8
XFILLER_15_697 VPWR VGND sg13g2_decap_8
XFILLER_30_623 VPWR VGND sg13g2_decap_8
XFILLER_42_494 VPWR VGND sg13g2_decap_8
XFILLER_14_196 VPWR VGND sg13g2_decap_8
Xinput13 uio_in[4] net13 VPWR VGND sg13g2_buf_1
XFILLER_52_70 VPWR VGND sg13g2_decap_8
XFILLER_7_830 VPWR VGND sg13g2_decap_8
XFILLER_42_4 VPWR VGND sg13g2_decap_8
XFILLER_97_623 VPWR VGND sg13g2_decap_8
XFILLER_96_133 VPWR VGND sg13g2_decap_8
XFILLER_69_358 VPWR VGND sg13g2_decap_8
XFILLER_78_881 VPWR VGND sg13g2_decap_8
XFILLER_37_200 VPWR VGND sg13g2_decap_8
XFILLER_38_756 VPWR VGND sg13g2_decap_8
XFILLER_93_873 VPWR VGND sg13g2_decap_8
XFILLER_92_350 VPWR VGND sg13g2_decap_8
XFILLER_65_553 VPWR VGND sg13g2_decap_8
X_37_ _05_ _03_ net19 VPWR VGND sg13g2_xor2_1
XFILLER_25_406 VPWR VGND sg13g2_decap_8
XFILLER_52_203 VPWR VGND sg13g2_decap_8
XFILLER_37_277 VPWR VGND sg13g2_decap_8
XFILLER_80_567 VPWR VGND sg13g2_decap_8
Xheichips25_example_large_31 VPWR VGND uio_oe[6] sg13g2_tielo
XFILLER_61_781 VPWR VGND sg13g2_decap_8
XFILLER_34_984 VPWR VGND sg13g2_decap_8
XFILLER_60_291 VPWR VGND sg13g2_decap_8
XFILLER_21_623 VPWR VGND sg13g2_decap_8
XFILLER_32_18 VPWR VGND sg13g2_decap_8
XFILLER_33_483 VPWR VGND sg13g2_decap_8
XFILLER_20_144 VPWR VGND sg13g2_decap_8
XFILLER_106_238 VPWR VGND sg13g2_decap_8
XFILLER_103_945 VPWR VGND sg13g2_decap_8
XFILLER_88_634 VPWR VGND sg13g2_decap_8
XFILLER_102_455 VPWR VGND sg13g2_decap_8
XFILLER_87_133 VPWR VGND sg13g2_decap_8
XFILLER_84_840 VPWR VGND sg13g2_decap_8
XFILLER_71_501 VPWR VGND sg13g2_decap_8
XFILLER_56_564 VPWR VGND sg13g2_decap_8
XFILLER_44_704 VPWR VGND sg13g2_decap_8
XFILLER_16_406 VPWR VGND sg13g2_decap_8
XFILLER_17_907 VPWR VGND sg13g2_decap_8
XFILLER_28_266 VPWR VGND sg13g2_decap_8
XFILLER_29_767 VPWR VGND sg13g2_decap_8
XFILLER_83_361 VPWR VGND sg13g2_decap_8
XFILLER_73_25 VPWR VGND sg13g2_decap_8
XFILLER_43_203 VPWR VGND sg13g2_decap_8
XFILLER_19_1001 VPWR VGND sg13g2_decap_8
XFILLER_71_578 VPWR VGND sg13g2_decap_8
XFILLER_52_770 VPWR VGND sg13g2_decap_8
XFILLER_25_973 VPWR VGND sg13g2_decap_8
XFILLER_40_910 VPWR VGND sg13g2_decap_8
XFILLER_106_1015 VPWR VGND sg13g2_decap_8
XFILLER_51_291 VPWR VGND sg13g2_decap_8
XFILLER_12_634 VPWR VGND sg13g2_decap_8
XFILLER_24_494 VPWR VGND sg13g2_decap_8
XFILLER_8_616 VPWR VGND sg13g2_decap_8
XFILLER_11_133 VPWR VGND sg13g2_decap_8
XFILLER_40_987 VPWR VGND sg13g2_decap_8
XFILLER_7_137 VPWR VGND sg13g2_decap_8
XFILLER_98_11 VPWR VGND sg13g2_decap_8
XFILLER_4_833 VPWR VGND sg13g2_decap_8
XFILLER_22_95 VPWR VGND sg13g2_decap_8
XFILLER_3_343 VPWR VGND sg13g2_decap_8
XFILLER_98_88 VPWR VGND sg13g2_decap_8
XFILLER_79_634 VPWR VGND sg13g2_decap_8
XFILLER_78_111 VPWR VGND sg13g2_decap_8
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_93_103 VPWR VGND sg13g2_decap_8
XFILLER_94_637 VPWR VGND sg13g2_decap_8
XFILLER_78_188 VPWR VGND sg13g2_decap_8
XFILLER_75_840 VPWR VGND sg13g2_decap_8
XFILLER_66_328 VPWR VGND sg13g2_decap_8
XFILLER_47_553 VPWR VGND sg13g2_decap_8
XFILLER_47_70 VPWR VGND sg13g2_decap_8
XFILLER_74_372 VPWR VGND sg13g2_decap_8
XFILLER_19_266 VPWR VGND sg13g2_decap_8
XFILLER_34_214 VPWR VGND sg13g2_decap_8
XFILLER_90_865 VPWR VGND sg13g2_decap_8
XFILLER_62_567 VPWR VGND sg13g2_decap_8
XFILLER_50_707 VPWR VGND sg13g2_decap_8
XFILLER_43_770 VPWR VGND sg13g2_decap_8
XFILLER_16_973 VPWR VGND sg13g2_decap_8
XFILLER_31_910 VPWR VGND sg13g2_decap_8
XFILLER_63_91 VPWR VGND sg13g2_decap_8
XFILLER_42_291 VPWR VGND sg13g2_decap_8
XFILLER_15_494 VPWR VGND sg13g2_decap_8
XFILLER_30_420 VPWR VGND sg13g2_decap_8
XFILLER_8_42 VPWR VGND sg13g2_decap_8
XFILLER_31_987 VPWR VGND sg13g2_decap_8
XFILLER_30_497 VPWR VGND sg13g2_decap_8
XFILLER_98_921 VPWR VGND sg13g2_decap_8
XFILLER_97_420 VPWR VGND sg13g2_decap_8
XFILLER_33_0 VPWR VGND sg13g2_decap_8
XFILLER_98_998 VPWR VGND sg13g2_decap_8
XFILLER_69_155 VPWR VGND sg13g2_decap_8
XFILLER_100_959 VPWR VGND sg13g2_decap_8
XFILLER_97_497 VPWR VGND sg13g2_decap_8
XFILLER_85_637 VPWR VGND sg13g2_decap_8
XFILLER_27_18 VPWR VGND sg13g2_decap_8
XFILLER_84_147 VPWR VGND sg13g2_decap_8
XFILLER_65_350 VPWR VGND sg13g2_decap_8
XFILLER_38_553 VPWR VGND sg13g2_decap_8
XFILLER_93_670 VPWR VGND sg13g2_decap_8
XFILLER_66_895 VPWR VGND sg13g2_decap_8
XFILLER_25_203 VPWR VGND sg13g2_decap_8
XFILLER_81_865 VPWR VGND sg13g2_decap_8
XFILLER_53_567 VPWR VGND sg13g2_decap_8
XFILLER_41_707 VPWR VGND sg13g2_decap_8
XFILLER_80_364 VPWR VGND sg13g2_decap_8
XFILLER_43_28 VPWR VGND sg13g2_decap_8
XFILLER_22_921 VPWR VGND sg13g2_decap_8
XFILLER_40_217 VPWR VGND sg13g2_decap_8
XFILLER_21_420 VPWR VGND sg13g2_decap_8
XFILLER_33_280 VPWR VGND sg13g2_decap_8
XFILLER_34_781 VPWR VGND sg13g2_decap_8
XFILLER_21_497 VPWR VGND sg13g2_decap_8
XFILLER_22_998 VPWR VGND sg13g2_decap_8
XFILLER_49_1005 VPWR VGND sg13g2_decap_8
XFILLER_89_910 VPWR VGND sg13g2_decap_8
XFILLER_68_25 VPWR VGND sg13g2_decap_8
XFILLER_103_742 VPWR VGND sg13g2_decap_8
XFILLER_88_431 VPWR VGND sg13g2_decap_8
XFILLER_1_847 VPWR VGND sg13g2_decap_8
XFILLER_102_252 VPWR VGND sg13g2_decap_8
XFILLER_89_987 VPWR VGND sg13g2_decap_8
XFILLER_0_357 VPWR VGND sg13g2_decap_8
XFILLER_76_648 VPWR VGND sg13g2_decap_8
XFILLER_57_840 VPWR VGND sg13g2_decap_8
XFILLER_84_35 VPWR VGND sg13g2_decap_8
XFILLER_75_147 VPWR VGND sg13g2_decap_8
XFILLER_17_704 VPWR VGND sg13g2_decap_8
XFILLER_29_564 VPWR VGND sg13g2_decap_8
XFILLER_56_361 VPWR VGND sg13g2_decap_8
XFILLER_44_501 VPWR VGND sg13g2_decap_8
XFILLER_16_203 VPWR VGND sg13g2_decap_8
XFILLER_72_854 VPWR VGND sg13g2_decap_8
XFILLER_71_375 VPWR VGND sg13g2_decap_8
XFILLER_44_578 VPWR VGND sg13g2_decap_8
XFILLER_13_910 VPWR VGND sg13g2_decap_8
XFILLER_17_95 VPWR VGND sg13g2_decap_8
XFILLER_25_770 VPWR VGND sg13g2_decap_8
XFILLER_31_217 VPWR VGND sg13g2_decap_8
XFILLER_32_718 VPWR VGND sg13g2_decap_8
XFILLER_9_903 VPWR VGND sg13g2_decap_8
XFILLER_8_413 VPWR VGND sg13g2_decap_8
XFILLER_12_431 VPWR VGND sg13g2_decap_8
XFILLER_13_987 VPWR VGND sg13g2_decap_8
XFILLER_24_291 VPWR VGND sg13g2_decap_8
XFILLER_40_784 VPWR VGND sg13g2_decap_8
XFILLER_99_707 VPWR VGND sg13g2_decap_8
XFILLER_4_630 VPWR VGND sg13g2_decap_8
XFILLER_98_228 VPWR VGND sg13g2_decap_8
XFILLER_3_140 VPWR VGND sg13g2_decap_8
XFILLER_79_431 VPWR VGND sg13g2_decap_8
XFILLER_95_935 VPWR VGND sg13g2_decap_8
XFILLER_94_434 VPWR VGND sg13g2_decap_8
XFILLER_67_637 VPWR VGND sg13g2_decap_8
XFILLER_66_125 VPWR VGND sg13g2_decap_8
XFILLER_58_91 VPWR VGND sg13g2_decap_8
XFILLER_48_840 VPWR VGND sg13g2_decap_8
XFILLER_47_350 VPWR VGND sg13g2_decap_8
XFILLER_63_854 VPWR VGND sg13g2_decap_8
XFILLER_90_662 VPWR VGND sg13g2_decap_8
XFILLER_62_364 VPWR VGND sg13g2_decap_8
XFILLER_50_504 VPWR VGND sg13g2_decap_8
XFILLER_16_770 VPWR VGND sg13g2_decap_8
XFILLER_23_707 VPWR VGND sg13g2_decap_8
XFILLER_35_567 VPWR VGND sg13g2_decap_8
XFILLER_22_228 VPWR VGND sg13g2_decap_8
XFILLER_15_291 VPWR VGND sg13g2_decap_8
XFILLER_31_784 VPWR VGND sg13g2_decap_8
XFILLER_30_294 VPWR VGND sg13g2_decap_8
XFILLER_8_980 VPWR VGND sg13g2_decap_8
XFILLER_104_539 VPWR VGND sg13g2_decap_8
XFILLER_89_217 VPWR VGND sg13g2_decap_8
XFILLER_98_795 VPWR VGND sg13g2_decap_8
XFILLER_97_294 VPWR VGND sg13g2_decap_8
XFILLER_86_935 VPWR VGND sg13g2_decap_8
XFILLER_85_434 VPWR VGND sg13g2_decap_8
XFILLER_58_637 VPWR VGND sg13g2_decap_8
XFILLER_38_28 VPWR VGND sg13g2_decap_8
XFILLER_100_756 VPWR VGND sg13g2_decap_8
XFILLER_57_147 VPWR VGND sg13g2_decap_8
XFILLER_39_851 VPWR VGND sg13g2_decap_8
XFILLER_38_350 VPWR VGND sg13g2_decap_8
XFILLER_66_692 VPWR VGND sg13g2_decap_8
XFILLER_54_865 VPWR VGND sg13g2_decap_8
XFILLER_81_662 VPWR VGND sg13g2_decap_8
XFILLER_80_161 VPWR VGND sg13g2_decap_8
XFILLER_53_364 VPWR VGND sg13g2_decap_8
XFILLER_14_707 VPWR VGND sg13g2_decap_8
XFILLER_26_567 VPWR VGND sg13g2_decap_8
XFILLER_41_504 VPWR VGND sg13g2_decap_8
XFILLER_13_217 VPWR VGND sg13g2_decap_8
XFILLER_16_1015 VPWR VGND sg13g2_decap_8
XFILLER_10_935 VPWR VGND sg13g2_decap_8
XFILLER_22_795 VPWR VGND sg13g2_decap_8
XFILLER_6_917 VPWR VGND sg13g2_decap_8
XFILLER_21_294 VPWR VGND sg13g2_decap_8
XFILLER_5_438 VPWR VGND sg13g2_decap_8
XFILLER_79_35 VPWR VGND sg13g2_decap_8
XFILLER_1_644 VPWR VGND sg13g2_decap_8
XFILLER_89_784 VPWR VGND sg13g2_decap_8
XFILLER_77_924 VPWR VGND sg13g2_decap_8
XFILLER_0_154 VPWR VGND sg13g2_decap_8
XFILLER_49_648 VPWR VGND sg13g2_decap_8
XFILLER_23_1008 VPWR VGND sg13g2_decap_8
XFILLER_95_67 VPWR VGND sg13g2_decap_8
XFILLER_76_445 VPWR VGND sg13g2_decap_8
XFILLER_48_147 VPWR VGND sg13g2_decap_8
XFILLER_92_938 VPWR VGND sg13g2_decap_8
XFILLER_17_501 VPWR VGND sg13g2_decap_8
XFILLER_29_361 VPWR VGND sg13g2_decap_8
XFILLER_91_448 VPWR VGND sg13g2_decap_8
XFILLER_45_854 VPWR VGND sg13g2_decap_8
XFILLER_72_651 VPWR VGND sg13g2_decap_8
XFILLER_60_802 VPWR VGND sg13g2_decap_8
XFILLER_44_375 VPWR VGND sg13g2_decap_8
XFILLER_17_578 VPWR VGND sg13g2_decap_8
XFILLER_32_515 VPWR VGND sg13g2_decap_8
XFILLER_71_172 VPWR VGND sg13g2_decap_8
XFILLER_44_60 VPWR VGND sg13g2_decap_8
XFILLER_60_879 VPWR VGND sg13g2_decap_8
XFILLER_9_700 VPWR VGND sg13g2_decap_8
XFILLER_8_210 VPWR VGND sg13g2_decap_8
XFILLER_13_784 VPWR VGND sg13g2_decap_8
XFILLER_40_581 VPWR VGND sg13g2_decap_8
XFILLER_74_7 VPWR VGND sg13g2_decap_8
XFILLER_9_777 VPWR VGND sg13g2_decap_8
XFILLER_60_81 VPWR VGND sg13g2_decap_8
XFILLER_8_287 VPWR VGND sg13g2_decap_8
XFILLER_99_504 VPWR VGND sg13g2_decap_8
XFILLER_5_32 VPWR VGND sg13g2_decap_8
XFILLER_95_732 VPWR VGND sg13g2_decap_8
XFILLER_68_957 VPWR VGND sg13g2_decap_8
XFILLER_67_434 VPWR VGND sg13g2_decap_8
XFILLER_94_231 VPWR VGND sg13g2_decap_8
XFILLER_39_158 VPWR VGND sg13g2_decap_8
XFILLER_83_949 VPWR VGND sg13g2_decap_8
XFILLER_82_448 VPWR VGND sg13g2_decap_8
XFILLER_36_854 VPWR VGND sg13g2_decap_8
XFILLER_63_651 VPWR VGND sg13g2_decap_8
XFILLER_51_802 VPWR VGND sg13g2_decap_8
XFILLER_23_504 VPWR VGND sg13g2_decap_8
XFILLER_35_364 VPWR VGND sg13g2_decap_8
XFILLER_39_1026 VPWR VGND sg13g2_fill_2
XFILLER_62_161 VPWR VGND sg13g2_decap_8
XFILLER_50_301 VPWR VGND sg13g2_decap_8
XFILLER_51_879 VPWR VGND sg13g2_decap_8
XFILLER_50_378 VPWR VGND sg13g2_decap_8
XFILLER_31_581 VPWR VGND sg13g2_decap_8
XFILLER_105_826 VPWR VGND sg13g2_decap_8
XFILLER_104_336 VPWR VGND sg13g2_decap_8
XFILLER_46_1019 VPWR VGND sg13g2_decap_8
XFILLER_98_592 VPWR VGND sg13g2_decap_8
XFILLER_86_732 VPWR VGND sg13g2_decap_8
XFILLER_59_957 VPWR VGND sg13g2_decap_8
XFILLER_58_434 VPWR VGND sg13g2_decap_8
XFILLER_100_553 VPWR VGND sg13g2_decap_8
XFILLER_85_231 VPWR VGND sg13g2_decap_8
XFILLER_105_77 VPWR VGND sg13g2_decap_8
XFILLER_73_459 VPWR VGND sg13g2_decap_8
XFILLER_60_109 VPWR VGND sg13g2_decap_8
XFILLER_54_662 VPWR VGND sg13g2_decap_8
XFILLER_42_802 VPWR VGND sg13g2_decap_8
XFILLER_14_504 VPWR VGND sg13g2_decap_8
XFILLER_26_364 VPWR VGND sg13g2_decap_8
XFILLER_27_865 VPWR VGND sg13g2_decap_8
XFILLER_81_25 VPWR VGND sg13g2_decap_8
XFILLER_53_161 VPWR VGND sg13g2_decap_8
XFILLER_41_301 VPWR VGND sg13g2_decap_8
XFILLER_42_879 VPWR VGND sg13g2_decap_8
XFILLER_14_63 VPWR VGND sg13g2_decap_8
XFILLER_41_378 VPWR VGND sg13g2_decap_8
XFILLER_10_732 VPWR VGND sg13g2_decap_8
XFILLER_22_592 VPWR VGND sg13g2_decap_8
XFILLER_6_714 VPWR VGND sg13g2_decap_8
XFILLER_5_235 VPWR VGND sg13g2_decap_8
XFILLER_100_0 VPWR VGND sg13g2_decap_8
XFILLER_2_942 VPWR VGND sg13g2_decap_8
XFILLER_30_84 VPWR VGND sg13g2_decap_8
XFILLER_96_518 VPWR VGND sg13g2_decap_8
XFILLER_1_441 VPWR VGND sg13g2_decap_8
XFILLER_89_581 VPWR VGND sg13g2_decap_8
XFILLER_77_721 VPWR VGND sg13g2_decap_8
XFILLER_39_60 VPWR VGND sg13g2_decap_8
XFILLER_76_242 VPWR VGND sg13g2_decap_8
XFILLER_49_445 VPWR VGND sg13g2_decap_8
XFILLER_92_735 VPWR VGND sg13g2_decap_8
XFILLER_77_798 VPWR VGND sg13g2_decap_8
XFILLER_65_938 VPWR VGND sg13g2_decap_8
XFILLER_91_245 VPWR VGND sg13g2_decap_8
XFILLER_64_459 VPWR VGND sg13g2_decap_8
XFILLER_18_854 VPWR VGND sg13g2_decap_8
XFILLER_55_70 VPWR VGND sg13g2_decap_8
XFILLER_51_109 VPWR VGND sg13g2_decap_8
XFILLER_45_651 VPWR VGND sg13g2_decap_8
XFILLER_44_172 VPWR VGND sg13g2_decap_8
XFILLER_17_375 VPWR VGND sg13g2_decap_8
XFILLER_32_312 VPWR VGND sg13g2_decap_8
XFILLER_33_868 VPWR VGND sg13g2_decap_8
XFILLER_60_676 VPWR VGND sg13g2_decap_8
XFILLER_20_529 VPWR VGND sg13g2_decap_8
XFILLER_32_389 VPWR VGND sg13g2_decap_8
XFILLER_13_581 VPWR VGND sg13g2_decap_8
XFILLER_9_574 VPWR VGND sg13g2_decap_8
XFILLER_99_301 VPWR VGND sg13g2_decap_8
XFILLER_99_378 VPWR VGND sg13g2_decap_8
XFILLER_87_518 VPWR VGND sg13g2_decap_8
XFILLER_68_754 VPWR VGND sg13g2_decap_8
XFILLER_67_231 VPWR VGND sg13g2_decap_8
XFILLER_56_949 VPWR VGND sg13g2_decap_8
XFILLER_83_746 VPWR VGND sg13g2_decap_8
XFILLER_55_448 VPWR VGND sg13g2_decap_8
XFILLER_82_245 VPWR VGND sg13g2_decap_8
XFILLER_42_109 VPWR VGND sg13g2_decap_8
XFILLER_24_802 VPWR VGND sg13g2_decap_8
XFILLER_36_651 VPWR VGND sg13g2_decap_8
XFILLER_23_301 VPWR VGND sg13g2_decap_8
XFILLER_35_161 VPWR VGND sg13g2_decap_8
XFILLER_24_879 VPWR VGND sg13g2_decap_8
XFILLER_52_1001 VPWR VGND sg13g2_decap_8
XFILLER_51_676 VPWR VGND sg13g2_decap_8
XFILLER_50_175 VPWR VGND sg13g2_decap_8
XFILLER_11_518 VPWR VGND sg13g2_decap_8
XFILLER_23_378 VPWR VGND sg13g2_decap_8
XFILLER_51_39 VPWR VGND sg13g2_decap_8
XFILLER_3_728 VPWR VGND sg13g2_decap_8
XFILLER_105_623 VPWR VGND sg13g2_decap_8
XFILLER_4_7 VPWR VGND sg13g2_decap_8
XFILLER_104_133 VPWR VGND sg13g2_decap_8
XFILLER_2_249 VPWR VGND sg13g2_decap_8
XFILLER_101_840 VPWR VGND sg13g2_decap_8
XFILLER_76_25 VPWR VGND sg13g2_decap_8
XFILLER_59_754 VPWR VGND sg13g2_decap_8
XFILLER_58_231 VPWR VGND sg13g2_decap_8
XFILLER_100_350 VPWR VGND sg13g2_decap_8
XFILLER_47_938 VPWR VGND sg13g2_decap_8
XFILLER_74_757 VPWR VGND sg13g2_decap_8
XFILLER_46_459 VPWR VGND sg13g2_decap_8
XFILLER_92_35 VPWR VGND sg13g2_decap_8
XFILLER_73_256 VPWR VGND sg13g2_decap_8
XFILLER_15_802 VPWR VGND sg13g2_decap_8
XFILLER_27_662 VPWR VGND sg13g2_decap_8
XFILLER_14_301 VPWR VGND sg13g2_decap_8
XFILLER_26_161 VPWR VGND sg13g2_decap_8
XFILLER_70_952 VPWR VGND sg13g2_decap_8
XFILLER_15_879 VPWR VGND sg13g2_decap_8
XFILLER_30_805 VPWR VGND sg13g2_decap_8
XFILLER_42_676 VPWR VGND sg13g2_decap_8
XFILLER_14_378 VPWR VGND sg13g2_decap_8
XFILLER_25_84 VPWR VGND sg13g2_decap_8
XFILLER_41_175 VPWR VGND sg13g2_decap_8
XFILLER_6_511 VPWR VGND sg13g2_decap_8
XFILLER_6_588 VPWR VGND sg13g2_decap_8
XFILLER_97_805 VPWR VGND sg13g2_decap_8
XFILLER_96_315 VPWR VGND sg13g2_decap_8
XFILLER_49_242 VPWR VGND sg13g2_decap_8
XFILLER_2_11 VPWR VGND sg13g2_decap_8
X_53_ _20_ _14_ _17_ VPWR VGND sg13g2_nand2_1
XFILLER_38_938 VPWR VGND sg13g2_decap_8
XFILLER_92_532 VPWR VGND sg13g2_decap_8
XFILLER_77_595 VPWR VGND sg13g2_decap_8
XFILLER_65_735 VPWR VGND sg13g2_decap_8
XFILLER_2_88 VPWR VGND sg13g2_decap_8
XFILLER_64_256 VPWR VGND sg13g2_decap_8
XFILLER_18_651 VPWR VGND sg13g2_decap_8
XFILLER_37_459 VPWR VGND sg13g2_decap_8
XFILLER_80_749 VPWR VGND sg13g2_decap_8
XFILLER_75_1001 VPWR VGND sg13g2_decap_8
XFILLER_17_172 VPWR VGND sg13g2_decap_8
XFILLER_24_109 VPWR VGND sg13g2_decap_8
XFILLER_61_963 VPWR VGND sg13g2_decap_8
XFILLER_21_805 VPWR VGND sg13g2_decap_8
XFILLER_33_665 VPWR VGND sg13g2_decap_8
XFILLER_60_473 VPWR VGND sg13g2_decap_8
XFILLER_20_326 VPWR VGND sg13g2_decap_8
XFILLER_32_186 VPWR VGND sg13g2_decap_8
XFILLER_9_371 VPWR VGND sg13g2_decap_8
XFILLER_63_0 VPWR VGND sg13g2_decap_8
XFILLER_88_816 VPWR VGND sg13g2_decap_8
XFILLER_102_637 VPWR VGND sg13g2_decap_8
XFILLER_99_175 VPWR VGND sg13g2_decap_8
XFILLER_87_315 VPWR VGND sg13g2_decap_8
XFILLER_101_147 VPWR VGND sg13g2_decap_8
XFILLER_96_882 VPWR VGND sg13g2_decap_8
XFILLER_68_551 VPWR VGND sg13g2_decap_8
XFILLER_83_543 VPWR VGND sg13g2_decap_8
XFILLER_56_746 VPWR VGND sg13g2_decap_8
XFILLER_46_39 VPWR VGND sg13g2_decap_8
XFILLER_28_448 VPWR VGND sg13g2_decap_8
XFILLER_29_949 VPWR VGND sg13g2_decap_8
XFILLER_55_245 VPWR VGND sg13g2_decap_8
XFILLER_15_109 VPWR VGND sg13g2_decap_8
XFILLER_102_56 VPWR VGND sg13g2_decap_8
XFILLER_70_259 VPWR VGND sg13g2_decap_8
XFILLER_52_952 VPWR VGND sg13g2_decap_8
XFILLER_62_49 VPWR VGND sg13g2_decap_8
XFILLER_51_473 VPWR VGND sg13g2_decap_8
XFILLER_12_816 VPWR VGND sg13g2_decap_8
XFILLER_24_676 VPWR VGND sg13g2_decap_8
XFILLER_11_315 VPWR VGND sg13g2_decap_8
XFILLER_23_175 VPWR VGND sg13g2_decap_8
XFILLER_7_319 VPWR VGND sg13g2_decap_8
XFILLER_20_893 VPWR VGND sg13g2_decap_8
XFILLER_106_910 VPWR VGND sg13g2_decap_8
XFILLER_11_42 VPWR VGND sg13g2_decap_8
XFILLER_105_420 VPWR VGND sg13g2_decap_8
XFILLER_3_525 VPWR VGND sg13g2_decap_8
XFILLER_106_987 VPWR VGND sg13g2_decap_8
XFILLER_79_816 VPWR VGND sg13g2_decap_8
XFILLER_2_4 VPWR VGND sg13g2_decap_8
XFILLER_105_497 VPWR VGND sg13g2_decap_8
XFILLER_87_35 VPWR VGND sg13g2_decap_8
XFILLER_94_819 VPWR VGND sg13g2_decap_8
XFILLER_87_882 VPWR VGND sg13g2_decap_8
XFILLER_59_551 VPWR VGND sg13g2_decap_8
XFILLER_98_1012 VPWR VGND sg13g2_decap_8
XFILLER_47_735 VPWR VGND sg13g2_decap_8
XFILLER_19_448 VPWR VGND sg13g2_decap_8
XFILLER_74_554 VPWR VGND sg13g2_decap_8
XFILLER_46_256 VPWR VGND sg13g2_decap_8
XFILLER_62_749 VPWR VGND sg13g2_decap_8
XFILLER_43_952 VPWR VGND sg13g2_decap_8
XFILLER_42_473 VPWR VGND sg13g2_decap_8
XFILLER_15_676 VPWR VGND sg13g2_decap_8
XFILLER_30_602 VPWR VGND sg13g2_decap_8
XFILLER_14_175 VPWR VGND sg13g2_decap_8
XFILLER_30_679 VPWR VGND sg13g2_decap_8
Xinput14 uio_in[5] net14 VPWR VGND sg13g2_buf_2
XFILLER_11_882 VPWR VGND sg13g2_decap_8
XFILLER_7_886 VPWR VGND sg13g2_decap_8
XFILLER_6_385 VPWR VGND sg13g2_decap_8
XFILLER_97_602 VPWR VGND sg13g2_decap_8
XFILLER_96_112 VPWR VGND sg13g2_decap_8
XFILLER_69_337 VPWR VGND sg13g2_decap_8
XFILLER_97_679 VPWR VGND sg13g2_decap_8
XFILLER_85_819 VPWR VGND sg13g2_decap_8
XFILLER_78_860 VPWR VGND sg13g2_decap_8
XFILLER_96_189 VPWR VGND sg13g2_decap_8
XFILLER_84_329 VPWR VGND sg13g2_decap_8
XFILLER_77_392 VPWR VGND sg13g2_decap_8
XFILLER_65_532 VPWR VGND sg13g2_decap_8
XFILLER_38_735 VPWR VGND sg13g2_decap_8
XFILLER_93_852 VPWR VGND sg13g2_decap_8
X_36_ _03_ _05_ _06_ VPWR VGND sg13g2_nor2_1
XFILLER_37_256 VPWR VGND sg13g2_decap_8
XFILLER_53_749 VPWR VGND sg13g2_decap_8
XFILLER_80_546 VPWR VGND sg13g2_decap_8
Xheichips25_example_large_32 VPWR VGND uio_oe[7] sg13g2_tielo
XFILLER_52_259 VPWR VGND sg13g2_decap_8
XFILLER_34_963 VPWR VGND sg13g2_decap_8
XFILLER_61_760 VPWR VGND sg13g2_decap_8
XFILLER_21_602 VPWR VGND sg13g2_decap_8
XFILLER_33_462 VPWR VGND sg13g2_decap_8
XFILLER_60_270 VPWR VGND sg13g2_decap_8
XFILLER_20_123 VPWR VGND sg13g2_decap_8
XFILLER_21_679 VPWR VGND sg13g2_decap_8
XFILLER_106_217 VPWR VGND sg13g2_decap_8
XFILLER_103_924 VPWR VGND sg13g2_decap_8
XFILLER_88_613 VPWR VGND sg13g2_decap_8
XFILLER_102_434 VPWR VGND sg13g2_decap_8
XFILLER_87_112 VPWR VGND sg13g2_decap_8
XFILLER_0_539 VPWR VGND sg13g2_decap_8
XFILLER_57_49 VPWR VGND sg13g2_decap_8
XFILLER_87_189 VPWR VGND sg13g2_decap_8
XFILLER_75_329 VPWR VGND sg13g2_decap_8
XFILLER_29_746 VPWR VGND sg13g2_decap_8
XFILLER_83_340 VPWR VGND sg13g2_decap_8
XFILLER_56_543 VPWR VGND sg13g2_decap_8
XFILLER_28_245 VPWR VGND sg13g2_decap_8
XFILLER_84_896 VPWR VGND sg13g2_decap_8
XFILLER_71_557 VPWR VGND sg13g2_decap_8
XFILLER_43_259 VPWR VGND sg13g2_decap_8
XFILLER_25_952 VPWR VGND sg13g2_decap_8
XFILLER_12_613 VPWR VGND sg13g2_decap_8
XFILLER_51_270 VPWR VGND sg13g2_decap_8
XFILLER_11_112 VPWR VGND sg13g2_decap_8
XFILLER_24_473 VPWR VGND sg13g2_decap_8
XFILLER_40_966 VPWR VGND sg13g2_decap_8
XFILLER_7_116 VPWR VGND sg13g2_decap_8
XFILLER_11_189 VPWR VGND sg13g2_decap_8
XFILLER_20_690 VPWR VGND sg13g2_decap_8
XFILLER_22_74 VPWR VGND sg13g2_decap_8
XFILLER_4_812 VPWR VGND sg13g2_decap_8
XFILLER_98_67 VPWR VGND sg13g2_decap_8
XFILLER_3_322 VPWR VGND sg13g2_decap_8
XFILLER_106_784 VPWR VGND sg13g2_decap_8
XFILLER_79_613 VPWR VGND sg13g2_decap_8
XFILLER_65_1022 VPWR VGND sg13g2_decap_8
XFILLER_4_889 VPWR VGND sg13g2_decap_8
XFILLER_105_294 VPWR VGND sg13g2_decap_8
XFILLER_3_399 VPWR VGND sg13g2_decap_8
XFILLER_94_616 VPWR VGND sg13g2_decap_8
XFILLER_78_167 VPWR VGND sg13g2_decap_8
XFILLER_67_819 VPWR VGND sg13g2_decap_8
XFILLER_66_307 VPWR VGND sg13g2_decap_8
XFILLER_47_532 VPWR VGND sg13g2_decap_8
XFILLER_93_159 VPWR VGND sg13g2_decap_8
XFILLER_74_351 VPWR VGND sg13g2_decap_8
XFILLER_19_245 VPWR VGND sg13g2_decap_8
XFILLER_75_896 VPWR VGND sg13g2_decap_8
XFILLER_90_844 VPWR VGND sg13g2_decap_8
XFILLER_62_546 VPWR VGND sg13g2_decap_8
XFILLER_16_952 VPWR VGND sg13g2_decap_8
XFILLER_35_749 VPWR VGND sg13g2_decap_8
XFILLER_72_1015 VPWR VGND sg13g2_decap_8
XFILLER_63_70 VPWR VGND sg13g2_decap_8
XFILLER_42_270 VPWR VGND sg13g2_decap_8
XFILLER_15_473 VPWR VGND sg13g2_decap_8
XFILLER_8_21 VPWR VGND sg13g2_decap_8
XFILLER_31_966 VPWR VGND sg13g2_decap_8
XFILLER_30_476 VPWR VGND sg13g2_decap_8
XFILLER_8_98 VPWR VGND sg13g2_decap_8
XFILLER_7_683 VPWR VGND sg13g2_decap_8
XFILLER_98_900 VPWR VGND sg13g2_decap_8
XFILLER_6_182 VPWR VGND sg13g2_decap_8
XFILLER_69_134 VPWR VGND sg13g2_decap_8
XFILLER_98_977 VPWR VGND sg13g2_decap_8
XFILLER_97_476 VPWR VGND sg13g2_decap_8
XFILLER_85_616 VPWR VGND sg13g2_decap_8
XFILLER_58_819 VPWR VGND sg13g2_decap_8
XFILLER_26_0 VPWR VGND sg13g2_decap_8
XFILLER_100_938 VPWR VGND sg13g2_decap_8
XFILLER_84_126 VPWR VGND sg13g2_decap_8
XFILLER_57_329 VPWR VGND sg13g2_decap_8
XFILLER_66_874 VPWR VGND sg13g2_decap_8
XFILLER_38_532 VPWR VGND sg13g2_decap_8
XFILLER_81_844 VPWR VGND sg13g2_decap_8
XFILLER_80_343 VPWR VGND sg13g2_decap_8
XFILLER_53_546 VPWR VGND sg13g2_decap_8
XFILLER_26_749 VPWR VGND sg13g2_decap_8
XFILLER_22_900 VPWR VGND sg13g2_decap_8
XFILLER_25_259 VPWR VGND sg13g2_decap_8
XFILLER_34_760 VPWR VGND sg13g2_decap_8
XFILLER_22_977 VPWR VGND sg13g2_decap_8
XFILLER_21_476 VPWR VGND sg13g2_decap_8
XFILLER_4_119 VPWR VGND sg13g2_decap_8
XFILLER_104_7 VPWR VGND sg13g2_decap_8
XFILLER_49_1028 VPWR VGND sg13g2_fill_1
XFILLER_88_410 VPWR VGND sg13g2_decap_8
XFILLER_1_826 VPWR VGND sg13g2_decap_8
XFILLER_103_721 VPWR VGND sg13g2_decap_8
XFILLER_89_966 VPWR VGND sg13g2_decap_8
XFILLER_0_336 VPWR VGND sg13g2_decap_8
XFILLER_102_231 VPWR VGND sg13g2_decap_8
XFILLER_103_798 VPWR VGND sg13g2_decap_8
XFILLER_88_487 VPWR VGND sg13g2_decap_8
XFILLER_76_627 VPWR VGND sg13g2_decap_8
XFILLER_75_126 VPWR VGND sg13g2_decap_8
XFILLER_48_329 VPWR VGND sg13g2_decap_8
XFILLER_84_14 VPWR VGND sg13g2_decap_8
XFILLER_56_340 VPWR VGND sg13g2_decap_8
XFILLER_29_543 VPWR VGND sg13g2_decap_8
XFILLER_72_833 VPWR VGND sg13g2_decap_8
XFILLER_57_896 VPWR VGND sg13g2_decap_8
XFILLER_1_1008 VPWR VGND sg13g2_decap_8
XFILLER_95_1026 VPWR VGND sg13g2_fill_2
XFILLER_84_693 VPWR VGND sg13g2_decap_8
XFILLER_44_557 VPWR VGND sg13g2_decap_8
XFILLER_17_74 VPWR VGND sg13g2_decap_8
XFILLER_71_354 VPWR VGND sg13g2_decap_8
XFILLER_16_259 VPWR VGND sg13g2_decap_8
XFILLER_12_410 VPWR VGND sg13g2_decap_8
XFILLER_24_270 VPWR VGND sg13g2_decap_8
XFILLER_13_966 VPWR VGND sg13g2_decap_8
XFILLER_40_763 VPWR VGND sg13g2_decap_8
XFILLER_9_959 VPWR VGND sg13g2_decap_8
XFILLER_12_487 VPWR VGND sg13g2_decap_8
XFILLER_33_84 VPWR VGND sg13g2_decap_8
XFILLER_8_469 VPWR VGND sg13g2_decap_8
XFILLER_98_207 VPWR VGND sg13g2_decap_8
XFILLER_4_686 VPWR VGND sg13g2_decap_8
XFILLER_106_581 VPWR VGND sg13g2_decap_8
XFILLER_79_410 VPWR VGND sg13g2_decap_8
XFILLER_3_196 VPWR VGND sg13g2_decap_8
XFILLER_95_914 VPWR VGND sg13g2_decap_8
XFILLER_67_616 VPWR VGND sg13g2_decap_8
XFILLER_94_413 VPWR VGND sg13g2_decap_8
XFILLER_79_487 VPWR VGND sg13g2_decap_8
XFILLER_66_104 VPWR VGND sg13g2_decap_8
XFILLER_58_70 VPWR VGND sg13g2_decap_8
XFILLER_48_896 VPWR VGND sg13g2_decap_8
XFILLER_90_641 VPWR VGND sg13g2_decap_8
XFILLER_75_693 VPWR VGND sg13g2_decap_8
XFILLER_63_833 VPWR VGND sg13g2_decap_8
XFILLER_35_546 VPWR VGND sg13g2_decap_8
XFILLER_62_343 VPWR VGND sg13g2_decap_8
XFILLER_22_207 VPWR VGND sg13g2_decap_8
XFILLER_15_270 VPWR VGND sg13g2_decap_8
XFILLER_31_763 VPWR VGND sg13g2_decap_8
XFILLER_30_273 VPWR VGND sg13g2_decap_8
XFILLER_7_480 VPWR VGND sg13g2_decap_8
XFILLER_104_518 VPWR VGND sg13g2_decap_8
XFILLER_98_774 VPWR VGND sg13g2_decap_8
XFILLER_86_914 VPWR VGND sg13g2_decap_8
XFILLER_58_616 VPWR VGND sg13g2_decap_8
XFILLER_100_735 VPWR VGND sg13g2_decap_8
XFILLER_97_273 VPWR VGND sg13g2_decap_8
XFILLER_85_413 VPWR VGND sg13g2_decap_8
XFILLER_57_126 VPWR VGND sg13g2_decap_8
XFILLER_39_830 VPWR VGND sg13g2_decap_8
XFILLER_94_980 VPWR VGND sg13g2_decap_8
XFILLER_66_671 VPWR VGND sg13g2_decap_8
XFILLER_81_641 VPWR VGND sg13g2_decap_8
XFILLER_54_844 VPWR VGND sg13g2_decap_8
XFILLER_54_39 VPWR VGND sg13g2_decap_8
XFILLER_26_546 VPWR VGND sg13g2_decap_8
XFILLER_80_140 VPWR VGND sg13g2_decap_8
XFILLER_53_343 VPWR VGND sg13g2_decap_8
XFILLER_103_1008 VPWR VGND sg13g2_decap_8
XFILLER_70_49 VPWR VGND sg13g2_decap_8
XFILLER_10_914 VPWR VGND sg13g2_decap_8
XFILLER_21_273 VPWR VGND sg13g2_decap_8
XFILLER_22_774 VPWR VGND sg13g2_decap_8
XFILLER_5_417 VPWR VGND sg13g2_decap_8
XFILLER_79_14 VPWR VGND sg13g2_decap_8
XFILLER_79_58 VPWR VGND sg13g2_fill_1
XFILLER_1_623 VPWR VGND sg13g2_decap_8
XFILLER_89_763 VPWR VGND sg13g2_decap_8
XFILLER_77_903 VPWR VGND sg13g2_decap_8
XFILLER_0_133 VPWR VGND sg13g2_decap_8
XFILLER_103_595 VPWR VGND sg13g2_decap_8
XFILLER_95_46 VPWR VGND sg13g2_decap_8
XFILLER_88_284 VPWR VGND sg13g2_decap_8
XFILLER_76_424 VPWR VGND sg13g2_decap_8
XFILLER_49_627 VPWR VGND sg13g2_decap_8
XFILLER_48_126 VPWR VGND sg13g2_decap_8
XFILLER_92_917 VPWR VGND sg13g2_decap_8
XFILLER_91_427 VPWR VGND sg13g2_decap_8
XFILLER_85_980 VPWR VGND sg13g2_decap_8
XFILLER_28_84 VPWR VGND sg13g2_decap_8
XFILLER_29_340 VPWR VGND sg13g2_decap_8
XFILLER_84_490 VPWR VGND sg13g2_decap_8
XFILLER_72_630 VPWR VGND sg13g2_decap_8
XFILLER_57_693 VPWR VGND sg13g2_decap_8
XFILLER_45_833 VPWR VGND sg13g2_decap_8
XFILLER_71_151 VPWR VGND sg13g2_decap_8
XFILLER_44_354 VPWR VGND sg13g2_decap_8
XFILLER_17_557 VPWR VGND sg13g2_decap_8
XFILLER_60_858 VPWR VGND sg13g2_decap_8
XFILLER_13_763 VPWR VGND sg13g2_decap_8
XFILLER_40_560 VPWR VGND sg13g2_decap_8
XFILLER_9_756 VPWR VGND sg13g2_decap_8
XFILLER_12_284 VPWR VGND sg13g2_decap_8
XFILLER_67_7 VPWR VGND sg13g2_decap_8
XFILLER_60_60 VPWR VGND sg13g2_decap_8
XFILLER_8_266 VPWR VGND sg13g2_decap_8
XFILLER_5_11 VPWR VGND sg13g2_decap_8
XFILLER_5_984 VPWR VGND sg13g2_decap_8
XFILLER_5_88 VPWR VGND sg13g2_decap_8
XFILLER_4_483 VPWR VGND sg13g2_decap_8
XFILLER_95_711 VPWR VGND sg13g2_decap_8
XFILLER_94_210 VPWR VGND sg13g2_decap_8
XFILLER_79_284 VPWR VGND sg13g2_decap_8
XFILLER_68_936 VPWR VGND sg13g2_decap_8
XFILLER_67_413 VPWR VGND sg13g2_decap_8
XFILLER_39_137 VPWR VGND sg13g2_decap_8
XFILLER_95_788 VPWR VGND sg13g2_decap_8
XFILLER_94_287 VPWR VGND sg13g2_decap_8
XFILLER_83_928 VPWR VGND sg13g2_decap_8
XFILLER_82_427 VPWR VGND sg13g2_decap_8
XFILLER_78_1021 VPWR VGND sg13g2_decap_8
XFILLER_76_991 VPWR VGND sg13g2_decap_8
XFILLER_75_490 VPWR VGND sg13g2_decap_8
XFILLER_63_630 VPWR VGND sg13g2_decap_8
XFILLER_48_693 VPWR VGND sg13g2_decap_8
XFILLER_36_833 VPWR VGND sg13g2_decap_8
XFILLER_62_140 VPWR VGND sg13g2_decap_8
XFILLER_35_343 VPWR VGND sg13g2_decap_8
XFILLER_39_1005 VPWR VGND sg13g2_decap_8
XFILLER_91_994 VPWR VGND sg13g2_decap_8
XFILLER_51_858 VPWR VGND sg13g2_decap_8
XFILLER_50_357 VPWR VGND sg13g2_decap_8
XFILLER_31_560 VPWR VGND sg13g2_decap_8
XFILLER_105_805 VPWR VGND sg13g2_decap_8
XFILLER_104_315 VPWR VGND sg13g2_decap_8
XFILLER_49_39 VPWR VGND sg13g2_decap_8
XFILLER_98_571 VPWR VGND sg13g2_decap_8
XFILLER_86_711 VPWR VGND sg13g2_decap_8
XFILLER_85_210 VPWR VGND sg13g2_decap_8
XFILLER_59_936 VPWR VGND sg13g2_decap_8
XFILLER_58_413 VPWR VGND sg13g2_decap_8
XFILLER_105_56 VPWR VGND sg13g2_decap_8
XFILLER_100_532 VPWR VGND sg13g2_decap_8
XFILLER_86_788 VPWR VGND sg13g2_decap_8
XFILLER_74_939 VPWR VGND sg13g2_decap_8
XFILLER_67_980 VPWR VGND sg13g2_decap_8
XFILLER_65_49 VPWR VGND sg13g2_decap_8
XFILLER_85_287 VPWR VGND sg13g2_decap_8
XFILLER_73_438 VPWR VGND sg13g2_decap_8
XFILLER_27_844 VPWR VGND sg13g2_decap_8
XFILLER_54_641 VPWR VGND sg13g2_decap_8
XFILLER_53_140 VPWR VGND sg13g2_decap_8
XFILLER_26_343 VPWR VGND sg13g2_decap_8
XFILLER_82_994 VPWR VGND sg13g2_decap_8
XFILLER_42_858 VPWR VGND sg13g2_decap_8
XFILLER_41_357 VPWR VGND sg13g2_decap_8
XFILLER_10_711 VPWR VGND sg13g2_decap_8
XFILLER_14_42 VPWR VGND sg13g2_decap_8
XFILLER_22_571 VPWR VGND sg13g2_decap_8
XFILLER_10_788 VPWR VGND sg13g2_decap_8
XFILLER_5_214 VPWR VGND sg13g2_decap_8
XFILLER_30_63 VPWR VGND sg13g2_decap_8
XFILLER_2_921 VPWR VGND sg13g2_decap_8
XFILLER_77_700 VPWR VGND sg13g2_decap_8
XFILLER_1_420 VPWR VGND sg13g2_decap_8
XFILLER_104_882 VPWR VGND sg13g2_decap_8
XFILLER_89_560 VPWR VGND sg13g2_decap_8
XFILLER_49_424 VPWR VGND sg13g2_decap_8
XFILLER_2_998 VPWR VGND sg13g2_decap_8
XFILLER_103_392 VPWR VGND sg13g2_decap_8
XFILLER_76_221 VPWR VGND sg13g2_decap_8
XFILLER_1_497 VPWR VGND sg13g2_decap_8
XFILLER_92_714 VPWR VGND sg13g2_decap_8
XFILLER_77_777 VPWR VGND sg13g2_decap_8
XFILLER_65_917 VPWR VGND sg13g2_decap_8
XFILLER_58_980 VPWR VGND sg13g2_decap_8
XFILLER_91_224 VPWR VGND sg13g2_decap_8
XFILLER_76_298 VPWR VGND sg13g2_decap_8
XFILLER_64_438 VPWR VGND sg13g2_decap_8
XFILLER_57_490 VPWR VGND sg13g2_decap_8
XFILLER_45_630 VPWR VGND sg13g2_decap_8
XFILLER_18_833 VPWR VGND sg13g2_decap_8
XFILLER_17_354 VPWR VGND sg13g2_decap_8
XFILLER_44_151 VPWR VGND sg13g2_decap_8
XFILLER_33_847 VPWR VGND sg13g2_decap_8
XFILLER_60_655 VPWR VGND sg13g2_decap_8
XFILLER_13_560 VPWR VGND sg13g2_decap_8
XFILLER_20_508 VPWR VGND sg13g2_decap_8
XFILLER_32_368 VPWR VGND sg13g2_decap_8
XFILLER_71_81 VPWR VGND sg13g2_decap_8
XFILLER_9_553 VPWR VGND sg13g2_decap_8
XFILLER_69_1009 VPWR VGND sg13g2_decap_8
XFILLER_5_781 VPWR VGND sg13g2_decap_8
XFILLER_102_819 VPWR VGND sg13g2_decap_8
XFILLER_99_357 VPWR VGND sg13g2_decap_8
XFILLER_4_280 VPWR VGND sg13g2_decap_8
XFILLER_101_329 VPWR VGND sg13g2_decap_8
XFILLER_68_733 VPWR VGND sg13g2_decap_8
XFILLER_67_210 VPWR VGND sg13g2_decap_8
XFILLER_95_585 VPWR VGND sg13g2_decap_8
XFILLER_83_725 VPWR VGND sg13g2_decap_8
XFILLER_56_928 VPWR VGND sg13g2_decap_8
XFILLER_82_224 VPWR VGND sg13g2_decap_8
XFILLER_67_287 VPWR VGND sg13g2_decap_8
XFILLER_55_427 VPWR VGND sg13g2_decap_8
XFILLER_49_991 VPWR VGND sg13g2_decap_8
XFILLER_48_490 VPWR VGND sg13g2_decap_8
XFILLER_36_630 VPWR VGND sg13g2_decap_8
XFILLER_35_140 VPWR VGND sg13g2_decap_8
XFILLER_91_791 VPWR VGND sg13g2_decap_8
XFILLER_51_655 VPWR VGND sg13g2_decap_8
XFILLER_23_357 VPWR VGND sg13g2_decap_8
XFILLER_24_858 VPWR VGND sg13g2_decap_8
XFILLER_51_18 VPWR VGND sg13g2_decap_8
XFILLER_50_154 VPWR VGND sg13g2_decap_8
XFILLER_13_1008 VPWR VGND sg13g2_decap_8
XFILLER_105_602 VPWR VGND sg13g2_decap_8
XFILLER_3_707 VPWR VGND sg13g2_decap_8
XFILLER_104_112 VPWR VGND sg13g2_decap_8
XFILLER_2_228 VPWR VGND sg13g2_decap_8
XFILLER_105_679 VPWR VGND sg13g2_decap_8
XFILLER_104_189 VPWR VGND sg13g2_decap_8
XFILLER_59_733 VPWR VGND sg13g2_decap_8
XFILLER_58_210 VPWR VGND sg13g2_decap_8
XFILLER_86_585 VPWR VGND sg13g2_decap_8
XFILLER_47_917 VPWR VGND sg13g2_decap_8
XFILLER_101_896 VPWR VGND sg13g2_decap_8
XFILLER_74_736 VPWR VGND sg13g2_decap_8
XFILLER_73_235 VPWR VGND sg13g2_decap_8
XFILLER_58_287 VPWR VGND sg13g2_decap_8
XFILLER_46_438 VPWR VGND sg13g2_decap_8
XFILLER_92_14 VPWR VGND sg13g2_decap_8
XFILLER_26_140 VPWR VGND sg13g2_decap_8
XFILLER_27_641 VPWR VGND sg13g2_decap_8
XFILLER_82_791 VPWR VGND sg13g2_decap_8
XFILLER_70_931 VPWR VGND sg13g2_decap_8
XFILLER_55_994 VPWR VGND sg13g2_decap_8
XFILLER_42_655 VPWR VGND sg13g2_decap_8
XFILLER_15_858 VPWR VGND sg13g2_decap_8
XFILLER_25_63 VPWR VGND sg13g2_decap_8
XFILLER_14_357 VPWR VGND sg13g2_decap_8
XFILLER_41_154 VPWR VGND sg13g2_decap_8
XFILLER_10_585 VPWR VGND sg13g2_decap_8
XFILLER_41_84 VPWR VGND sg13g2_decap_8
XFILLER_68_1020 VPWR VGND sg13g2_decap_8
XFILLER_6_567 VPWR VGND sg13g2_decap_8
XFILLER_29_1026 VPWR VGND sg13g2_fill_2
XFILLER_69_519 VPWR VGND sg13g2_decap_8
XFILLER_49_221 VPWR VGND sg13g2_decap_8
XFILLER_2_795 VPWR VGND sg13g2_decap_8
XFILLER_1_294 VPWR VGND sg13g2_decap_8
XFILLER_77_574 VPWR VGND sg13g2_decap_8
X_52_ _19_ net6 net14 VPWR VGND sg13g2_xnor2_1
XFILLER_65_714 VPWR VGND sg13g2_decap_8
XFILLER_2_67 VPWR VGND sg13g2_decap_8
XFILLER_38_917 VPWR VGND sg13g2_decap_8
XFILLER_92_511 VPWR VGND sg13g2_decap_8
XFILLER_49_298 VPWR VGND sg13g2_decap_8
XFILLER_37_438 VPWR VGND sg13g2_decap_8
XFILLER_64_235 VPWR VGND sg13g2_decap_8
XFILLER_18_630 VPWR VGND sg13g2_decap_8
XFILLER_92_588 VPWR VGND sg13g2_decap_8
XFILLER_80_728 VPWR VGND sg13g2_decap_8
XFILLER_17_151 VPWR VGND sg13g2_decap_8
XFILLER_61_942 VPWR VGND sg13g2_decap_8
XFILLER_33_644 VPWR VGND sg13g2_decap_8
XFILLER_36_1008 VPWR VGND sg13g2_decap_8
XFILLER_82_91 VPWR VGND sg13g2_decap_8
XFILLER_60_452 VPWR VGND sg13g2_decap_8
XFILLER_20_305 VPWR VGND sg13g2_decap_8
XFILLER_32_165 VPWR VGND sg13g2_decap_8
XFILLER_9_350 VPWR VGND sg13g2_decap_8
XFILLER_99_154 VPWR VGND sg13g2_decap_8
XFILLER_102_616 VPWR VGND sg13g2_decap_8
XFILLER_101_126 VPWR VGND sg13g2_decap_8
XFILLER_68_530 VPWR VGND sg13g2_decap_8
XFILLER_96_861 VPWR VGND sg13g2_decap_8
XFILLER_29_928 VPWR VGND sg13g2_decap_8
XFILLER_95_382 VPWR VGND sg13g2_decap_8
XFILLER_83_522 VPWR VGND sg13g2_decap_8
XFILLER_56_725 VPWR VGND sg13g2_decap_8
XFILLER_55_224 VPWR VGND sg13g2_decap_8
XFILLER_46_18 VPWR VGND sg13g2_decap_8
XFILLER_28_427 VPWR VGND sg13g2_decap_8
XFILLER_102_35 VPWR VGND sg13g2_decap_8
XFILLER_83_599 VPWR VGND sg13g2_decap_8
XFILLER_71_739 VPWR VGND sg13g2_decap_8
XFILLER_70_238 VPWR VGND sg13g2_decap_8
XFILLER_62_28 VPWR VGND sg13g2_decap_8
XFILLER_52_931 VPWR VGND sg13g2_decap_8
XFILLER_24_655 VPWR VGND sg13g2_decap_8
XFILLER_51_452 VPWR VGND sg13g2_decap_8
XFILLER_23_154 VPWR VGND sg13g2_decap_8
XFILLER_20_872 VPWR VGND sg13g2_decap_8
XFILLER_11_21 VPWR VGND sg13g2_decap_8
XFILLER_3_504 VPWR VGND sg13g2_decap_8
XFILLER_106_966 VPWR VGND sg13g2_decap_8
XFILLER_87_14 VPWR VGND sg13g2_decap_8
XFILLER_11_98 VPWR VGND sg13g2_decap_8
XFILLER_105_476 VPWR VGND sg13g2_decap_8
XFILLER_78_349 VPWR VGND sg13g2_decap_8
XFILLER_59_530 VPWR VGND sg13g2_decap_8
XFILLER_87_861 VPWR VGND sg13g2_decap_8
XFILLER_47_714 VPWR VGND sg13g2_decap_8
XFILLER_101_693 VPWR VGND sg13g2_decap_8
XFILLER_86_382 VPWR VGND sg13g2_decap_8
XFILLER_74_533 VPWR VGND sg13g2_decap_8
XFILLER_19_427 VPWR VGND sg13g2_decap_8
XFILLER_46_235 VPWR VGND sg13g2_decap_8
XFILLER_62_728 VPWR VGND sg13g2_decap_8
XFILLER_28_994 VPWR VGND sg13g2_decap_8
XFILLER_61_249 VPWR VGND sg13g2_decap_8
XFILLER_55_791 VPWR VGND sg13g2_decap_8
XFILLER_43_931 VPWR VGND sg13g2_decap_8
XFILLER_36_84 VPWR VGND sg13g2_decap_8
XFILLER_42_452 VPWR VGND sg13g2_decap_8
XFILLER_14_154 VPWR VGND sg13g2_decap_8
XFILLER_15_655 VPWR VGND sg13g2_decap_8
XFILLER_11_861 VPWR VGND sg13g2_decap_8
XFILLER_30_658 VPWR VGND sg13g2_decap_8
Xinput15 uio_in[6] net15 VPWR VGND sg13g2_buf_1
XFILLER_10_382 VPWR VGND sg13g2_decap_8
XFILLER_7_865 VPWR VGND sg13g2_decap_8
XFILLER_6_364 VPWR VGND sg13g2_decap_8
XFILLER_69_316 VPWR VGND sg13g2_decap_8
XFILLER_97_658 VPWR VGND sg13g2_decap_8
XFILLER_2_592 VPWR VGND sg13g2_decap_8
XFILLER_96_168 VPWR VGND sg13g2_decap_8
XFILLER_84_308 VPWR VGND sg13g2_decap_8
XFILLER_77_91 VPWR VGND sg13g2_decap_8
XFILLER_42_1012 VPWR VGND sg13g2_decap_8
XFILLER_38_714 VPWR VGND sg13g2_decap_8
XFILLER_93_831 VPWR VGND sg13g2_decap_8
XFILLER_77_371 VPWR VGND sg13g2_decap_8
XFILLER_65_511 VPWR VGND sg13g2_decap_8
X_35_ _05_ net3 net11 VPWR VGND sg13g2_xnor2_1
XFILLER_37_235 VPWR VGND sg13g2_decap_8
XFILLER_92_385 VPWR VGND sg13g2_decap_8
XFILLER_80_525 VPWR VGND sg13g2_decap_8
XFILLER_65_588 VPWR VGND sg13g2_decap_8
XFILLER_53_728 VPWR VGND sg13g2_decap_8
XFILLER_19_994 VPWR VGND sg13g2_decap_8
XFILLER_52_238 VPWR VGND sg13g2_decap_8
Xheichips25_example_large_33 VPWR VGND uio_out[0] sg13g2_tielo
XFILLER_34_942 VPWR VGND sg13g2_decap_8
XFILLER_33_441 VPWR VGND sg13g2_decap_8
XFILLER_20_102 VPWR VGND sg13g2_decap_8
XFILLER_21_658 VPWR VGND sg13g2_decap_8
XFILLER_20_179 VPWR VGND sg13g2_decap_8
XFILLER_103_903 VPWR VGND sg13g2_decap_8
XFILLER_0_518 VPWR VGND sg13g2_decap_8
XFILLER_102_413 VPWR VGND sg13g2_decap_8
XFILLER_76_809 VPWR VGND sg13g2_decap_8
XFILLER_88_669 VPWR VGND sg13g2_decap_8
XFILLER_87_168 VPWR VGND sg13g2_decap_8
XFILLER_75_308 VPWR VGND sg13g2_decap_8
XFILLER_57_28 VPWR VGND sg13g2_decap_8
XFILLER_69_883 VPWR VGND sg13g2_decap_8
XFILLER_56_522 VPWR VGND sg13g2_decap_8
XFILLER_29_725 VPWR VGND sg13g2_decap_8
XFILLER_84_875 VPWR VGND sg13g2_decap_8
XFILLER_28_224 VPWR VGND sg13g2_decap_8
XFILLER_56_599 VPWR VGND sg13g2_decap_8
XFILLER_44_739 VPWR VGND sg13g2_decap_8
XFILLER_83_396 VPWR VGND sg13g2_decap_8
XFILLER_71_536 VPWR VGND sg13g2_decap_8
XFILLER_43_238 VPWR VGND sg13g2_decap_8
XFILLER_25_931 VPWR VGND sg13g2_decap_8
XFILLER_24_452 VPWR VGND sg13g2_decap_8
XFILLER_40_945 VPWR VGND sg13g2_decap_8
XFILLER_12_669 VPWR VGND sg13g2_decap_8
XFILLER_11_168 VPWR VGND sg13g2_decap_8
XFILLER_22_53 VPWR VGND sg13g2_decap_8
XFILLER_3_301 VPWR VGND sg13g2_decap_8
XFILLER_98_46 VPWR VGND sg13g2_decap_8
XFILLER_65_1001 VPWR VGND sg13g2_decap_8
XFILLER_4_868 VPWR VGND sg13g2_decap_8
XFILLER_106_763 VPWR VGND sg13g2_decap_8
XFILLER_3_378 VPWR VGND sg13g2_decap_8
XFILLER_105_273 VPWR VGND sg13g2_decap_8
XFILLER_79_669 VPWR VGND sg13g2_decap_8
XFILLER_78_146 VPWR VGND sg13g2_decap_8
XFILLER_102_980 VPWR VGND sg13g2_decap_8
XFILLER_47_511 VPWR VGND sg13g2_decap_8
XFILLER_101_490 VPWR VGND sg13g2_decap_8
XFILLER_93_138 VPWR VGND sg13g2_decap_8
XFILLER_74_330 VPWR VGND sg13g2_decap_8
XFILLER_19_224 VPWR VGND sg13g2_decap_8
XFILLER_90_823 VPWR VGND sg13g2_decap_8
XFILLER_75_875 VPWR VGND sg13g2_decap_8
XFILLER_62_525 VPWR VGND sg13g2_decap_8
XFILLER_47_588 VPWR VGND sg13g2_decap_8
XFILLER_35_728 VPWR VGND sg13g2_decap_8
XFILLER_16_931 VPWR VGND sg13g2_decap_8
XFILLER_28_791 VPWR VGND sg13g2_decap_8
XFILLER_34_249 VPWR VGND sg13g2_decap_8
XFILLER_15_452 VPWR VGND sg13g2_decap_8
XFILLER_97_7 VPWR VGND sg13g2_decap_8
XFILLER_31_945 VPWR VGND sg13g2_decap_8
XFILLER_30_455 VPWR VGND sg13g2_decap_8
XFILLER_8_77 VPWR VGND sg13g2_decap_8
XFILLER_7_662 VPWR VGND sg13g2_decap_8
XFILLER_6_161 VPWR VGND sg13g2_decap_8
XFILLER_98_956 VPWR VGND sg13g2_decap_8
XFILLER_69_113 VPWR VGND sg13g2_decap_8
XFILLER_100_917 VPWR VGND sg13g2_decap_8
XFILLER_97_455 VPWR VGND sg13g2_decap_8
XFILLER_57_308 VPWR VGND sg13g2_decap_8
XFILLER_84_105 VPWR VGND sg13g2_decap_8
XFILLER_38_511 VPWR VGND sg13g2_decap_8
XFILLER_66_853 VPWR VGND sg13g2_decap_8
XFILLER_19_0 VPWR VGND sg13g2_decap_8
XFILLER_81_823 VPWR VGND sg13g2_decap_8
XFILLER_26_728 VPWR VGND sg13g2_decap_8
XFILLER_38_588 VPWR VGND sg13g2_decap_8
XFILLER_92_182 VPWR VGND sg13g2_decap_8
XFILLER_80_322 VPWR VGND sg13g2_decap_8
XFILLER_65_385 VPWR VGND sg13g2_decap_8
XFILLER_53_525 VPWR VGND sg13g2_decap_8
XFILLER_19_791 VPWR VGND sg13g2_decap_8
XFILLER_25_238 VPWR VGND sg13g2_decap_8
XFILLER_80_399 VPWR VGND sg13g2_decap_8
XFILLER_21_455 VPWR VGND sg13g2_decap_8
XFILLER_22_956 VPWR VGND sg13g2_decap_8
XFILLER_88_1012 VPWR VGND sg13g2_decap_8
XFILLER_103_700 VPWR VGND sg13g2_decap_8
XFILLER_1_805 VPWR VGND sg13g2_decap_8
XFILLER_102_210 VPWR VGND sg13g2_decap_8
XFILLER_89_945 VPWR VGND sg13g2_decap_8
XFILLER_0_315 VPWR VGND sg13g2_decap_8
XFILLER_103_777 VPWR VGND sg13g2_decap_8
XFILLER_88_466 VPWR VGND sg13g2_decap_8
XFILLER_76_606 VPWR VGND sg13g2_decap_8
XFILLER_49_809 VPWR VGND sg13g2_decap_8
XFILLER_48_308 VPWR VGND sg13g2_decap_8
XFILLER_102_287 VPWR VGND sg13g2_decap_8
XFILLER_75_105 VPWR VGND sg13g2_decap_8
XFILLER_69_680 VPWR VGND sg13g2_decap_8
XFILLER_29_522 VPWR VGND sg13g2_decap_8
XFILLER_91_609 VPWR VGND sg13g2_decap_8
XFILLER_95_1005 VPWR VGND sg13g2_decap_8
XFILLER_84_672 VPWR VGND sg13g2_decap_8
XFILLER_72_812 VPWR VGND sg13g2_decap_8
XFILLER_57_875 VPWR VGND sg13g2_decap_8
XFILLER_83_193 VPWR VGND sg13g2_decap_8
XFILLER_71_333 VPWR VGND sg13g2_decap_8
XFILLER_56_396 VPWR VGND sg13g2_decap_8
XFILLER_44_536 VPWR VGND sg13g2_decap_8
XFILLER_16_238 VPWR VGND sg13g2_decap_8
XFILLER_17_53 VPWR VGND sg13g2_decap_8
XFILLER_17_739 VPWR VGND sg13g2_decap_8
XFILLER_29_599 VPWR VGND sg13g2_decap_8
XFILLER_72_889 VPWR VGND sg13g2_decap_8
XFILLER_13_945 VPWR VGND sg13g2_decap_8
XFILLER_40_742 VPWR VGND sg13g2_decap_8
XFILLER_9_938 VPWR VGND sg13g2_decap_8
XFILLER_12_466 VPWR VGND sg13g2_decap_8
XFILLER_33_63 VPWR VGND sg13g2_decap_8
XFILLER_8_448 VPWR VGND sg13g2_decap_8
XFILLER_106_560 VPWR VGND sg13g2_decap_8
XFILLER_4_665 VPWR VGND sg13g2_decap_8
XFILLER_3_175 VPWR VGND sg13g2_decap_8
XFILLER_79_466 VPWR VGND sg13g2_decap_8
XFILLER_0_882 VPWR VGND sg13g2_decap_8
XFILLER_39_319 VPWR VGND sg13g2_decap_8
XFILLER_94_469 VPWR VGND sg13g2_decap_8
XFILLER_82_609 VPWR VGND sg13g2_decap_8
XFILLER_75_672 VPWR VGND sg13g2_decap_8
XFILLER_63_812 VPWR VGND sg13g2_decap_8
XFILLER_48_875 VPWR VGND sg13g2_decap_8
XFILLER_90_620 VPWR VGND sg13g2_decap_8
XFILLER_62_322 VPWR VGND sg13g2_decap_8
XFILLER_47_385 VPWR VGND sg13g2_decap_8
XFILLER_35_525 VPWR VGND sg13g2_decap_8
XFILLER_74_92 VPWR VGND sg13g2_decap_8
XFILLER_63_889 VPWR VGND sg13g2_decap_8
XFILLER_90_697 VPWR VGND sg13g2_decap_8
XFILLER_62_399 VPWR VGND sg13g2_decap_8
XFILLER_50_539 VPWR VGND sg13g2_decap_8
XFILLER_95_4 VPWR VGND sg13g2_decap_8
XFILLER_31_742 VPWR VGND sg13g2_decap_8
XFILLER_30_252 VPWR VGND sg13g2_decap_8
XFILLER_98_753 VPWR VGND sg13g2_decap_8
XFILLER_97_252 VPWR VGND sg13g2_decap_8
XFILLER_100_714 VPWR VGND sg13g2_decap_8
XFILLER_57_105 VPWR VGND sg13g2_decap_8
XFILLER_85_469 VPWR VGND sg13g2_decap_8
XFILLER_72_119 VPWR VGND sg13g2_decap_8
XFILLER_66_650 VPWR VGND sg13g2_decap_8
XFILLER_54_823 VPWR VGND sg13g2_decap_8
XFILLER_39_886 VPWR VGND sg13g2_decap_8
XFILLER_81_620 VPWR VGND sg13g2_decap_8
XFILLER_65_182 VPWR VGND sg13g2_decap_8
XFILLER_54_18 VPWR VGND sg13g2_decap_8
XFILLER_53_322 VPWR VGND sg13g2_decap_8
XFILLER_26_525 VPWR VGND sg13g2_decap_8
XFILLER_38_385 VPWR VGND sg13g2_decap_8
XFILLER_81_697 VPWR VGND sg13g2_decap_8
XFILLER_55_1022 VPWR VGND sg13g2_decap_8
XFILLER_53_399 VPWR VGND sg13g2_decap_8
XFILLER_41_539 VPWR VGND sg13g2_decap_8
XFILLER_80_196 VPWR VGND sg13g2_decap_8
XFILLER_22_753 VPWR VGND sg13g2_decap_8
XFILLER_70_28 VPWR VGND sg13g2_decap_8
XFILLER_21_252 VPWR VGND sg13g2_decap_8
XFILLER_1_602 VPWR VGND sg13g2_decap_8
XFILLER_89_742 VPWR VGND sg13g2_decap_8
XFILLER_0_112 VPWR VGND sg13g2_decap_8
XFILLER_62_1015 VPWR VGND sg13g2_decap_8
XFILLER_49_606 VPWR VGND sg13g2_decap_8
XFILLER_103_574 VPWR VGND sg13g2_decap_8
XFILLER_95_25 VPWR VGND sg13g2_decap_8
XFILLER_88_263 VPWR VGND sg13g2_decap_8
XFILLER_76_403 VPWR VGND sg13g2_decap_8
XFILLER_48_105 VPWR VGND sg13g2_decap_8
XFILLER_1_679 VPWR VGND sg13g2_decap_8
XFILLER_77_959 VPWR VGND sg13g2_decap_8
XFILLER_0_189 VPWR VGND sg13g2_decap_8
XFILLER_91_406 VPWR VGND sg13g2_decap_8
XFILLER_63_119 VPWR VGND sg13g2_decap_8
XFILLER_57_672 VPWR VGND sg13g2_decap_8
XFILLER_45_812 VPWR VGND sg13g2_decap_8
XFILLER_28_63 VPWR VGND sg13g2_decap_8
XFILLER_17_536 VPWR VGND sg13g2_decap_8
XFILLER_29_396 VPWR VGND sg13g2_decap_8
XFILLER_71_130 VPWR VGND sg13g2_decap_8
XFILLER_56_193 VPWR VGND sg13g2_decap_8
XFILLER_45_889 VPWR VGND sg13g2_decap_8
XFILLER_44_333 VPWR VGND sg13g2_decap_8
XFILLER_72_686 VPWR VGND sg13g2_decap_8
XFILLER_60_837 VPWR VGND sg13g2_decap_8
XFILLER_44_95 VPWR VGND sg13g2_decap_8
XFILLER_13_742 VPWR VGND sg13g2_decap_8
XFILLER_9_735 VPWR VGND sg13g2_decap_8
XFILLER_12_263 VPWR VGND sg13g2_decap_8
XFILLER_8_245 VPWR VGND sg13g2_decap_8
XFILLER_5_963 VPWR VGND sg13g2_decap_8
XFILLER_99_539 VPWR VGND sg13g2_decap_8
XFILLER_5_67 VPWR VGND sg13g2_decap_8
XFILLER_4_462 VPWR VGND sg13g2_decap_8
XFILLER_69_92 VPWR VGND sg13g2_decap_8
XFILLER_68_915 VPWR VGND sg13g2_decap_8
XFILLER_79_263 VPWR VGND sg13g2_decap_8
XFILLER_39_116 VPWR VGND sg13g2_decap_8
XFILLER_95_767 VPWR VGND sg13g2_decap_8
XFILLER_83_907 VPWR VGND sg13g2_decap_8
XFILLER_94_266 VPWR VGND sg13g2_decap_8
XFILLER_82_406 VPWR VGND sg13g2_decap_8
XFILLER_78_1000 VPWR VGND sg13g2_decap_8
XFILLER_76_970 VPWR VGND sg13g2_decap_8
XFILLER_67_469 VPWR VGND sg13g2_decap_8
XFILLER_55_609 VPWR VGND sg13g2_decap_8
XFILLER_48_672 VPWR VGND sg13g2_decap_8
XFILLER_10_4 VPWR VGND sg13g2_decap_8
XFILLER_36_812 VPWR VGND sg13g2_decap_8
XFILLER_85_91 VPWR VGND sg13g2_decap_8
XFILLER_47_182 VPWR VGND sg13g2_decap_8
XFILLER_35_322 VPWR VGND sg13g2_decap_8
XFILLER_91_973 VPWR VGND sg13g2_decap_8
XFILLER_36_889 VPWR VGND sg13g2_decap_8
XFILLER_39_1028 VPWR VGND sg13g2_fill_1
XFILLER_63_686 VPWR VGND sg13g2_decap_8
XFILLER_51_837 VPWR VGND sg13g2_decap_8
XFILLER_23_539 VPWR VGND sg13g2_decap_8
XFILLER_35_399 VPWR VGND sg13g2_decap_8
XFILLER_90_494 VPWR VGND sg13g2_decap_8
XFILLER_62_196 VPWR VGND sg13g2_decap_8
XFILLER_50_336 VPWR VGND sg13g2_decap_8
XFILLER_85_1015 VPWR VGND sg13g2_decap_8
XFILLER_49_18 VPWR VGND sg13g2_decap_8
XFILLER_98_550 VPWR VGND sg13g2_decap_8
XFILLER_59_915 VPWR VGND sg13g2_decap_8
XFILLER_100_511 VPWR VGND sg13g2_decap_8
XFILLER_105_35 VPWR VGND sg13g2_decap_8
XFILLER_86_767 VPWR VGND sg13g2_decap_8
XFILLER_85_266 VPWR VGND sg13g2_decap_8
XFILLER_74_918 VPWR VGND sg13g2_decap_8
XFILLER_73_417 VPWR VGND sg13g2_decap_8
XFILLER_65_28 VPWR VGND sg13g2_decap_8
XFILLER_58_469 VPWR VGND sg13g2_decap_8
XFILLER_100_588 VPWR VGND sg13g2_decap_8
XFILLER_54_620 VPWR VGND sg13g2_decap_8
XFILLER_45_119 VPWR VGND sg13g2_decap_8
XFILLER_26_322 VPWR VGND sg13g2_decap_8
XFILLER_27_823 VPWR VGND sg13g2_decap_8
XFILLER_38_182 VPWR VGND sg13g2_decap_8
XFILLER_39_683 VPWR VGND sg13g2_decap_8
XFILLER_82_973 VPWR VGND sg13g2_decap_8
XFILLER_92_1008 VPWR VGND sg13g2_decap_8
XFILLER_54_697 VPWR VGND sg13g2_decap_8
XFILLER_42_837 VPWR VGND sg13g2_decap_8
XFILLER_14_539 VPWR VGND sg13g2_decap_8
XFILLER_81_494 VPWR VGND sg13g2_decap_8
XFILLER_53_196 VPWR VGND sg13g2_decap_8
XFILLER_26_399 VPWR VGND sg13g2_decap_8
XFILLER_41_336 VPWR VGND sg13g2_decap_8
XFILLER_14_21 VPWR VGND sg13g2_decap_8
XFILLER_22_550 VPWR VGND sg13g2_decap_8
XFILLER_10_767 VPWR VGND sg13g2_decap_8
XFILLER_14_98 VPWR VGND sg13g2_decap_8
XFILLER_6_749 VPWR VGND sg13g2_decap_8
XFILLER_2_900 VPWR VGND sg13g2_decap_8
XFILLER_30_42 VPWR VGND sg13g2_decap_8
XFILLER_104_861 VPWR VGND sg13g2_decap_8
XFILLER_76_200 VPWR VGND sg13g2_decap_8
XFILLER_49_403 VPWR VGND sg13g2_decap_8
XFILLER_7_1026 VPWR VGND sg13g2_fill_2
XFILLER_2_977 VPWR VGND sg13g2_decap_8
XFILLER_1_476 VPWR VGND sg13g2_decap_8
XFILLER_103_371 VPWR VGND sg13g2_decap_8
XFILLER_77_756 VPWR VGND sg13g2_decap_8
XFILLER_76_277 VPWR VGND sg13g2_decap_8
XFILLER_64_417 VPWR VGND sg13g2_decap_8
XFILLER_18_812 VPWR VGND sg13g2_decap_8
XFILLER_39_95 VPWR VGND sg13g2_decap_8
XFILLER_91_203 VPWR VGND sg13g2_decap_8
XFILLER_36_119 VPWR VGND sg13g2_decap_8
XFILLER_44_130 VPWR VGND sg13g2_decap_8
XFILLER_17_333 VPWR VGND sg13g2_decap_8
XFILLER_29_193 VPWR VGND sg13g2_decap_8
XFILLER_73_984 VPWR VGND sg13g2_decap_8
XFILLER_72_483 VPWR VGND sg13g2_decap_8
XFILLER_45_686 VPWR VGND sg13g2_decap_8
XFILLER_18_889 VPWR VGND sg13g2_decap_8
XFILLER_33_826 VPWR VGND sg13g2_decap_8
XFILLER_60_634 VPWR VGND sg13g2_decap_8
XFILLER_32_347 VPWR VGND sg13g2_decap_8
XFILLER_71_60 VPWR VGND sg13g2_decap_8
XFILLER_9_532 VPWR VGND sg13g2_decap_8
XFILLER_99_336 VPWR VGND sg13g2_decap_8
XFILLER_5_760 VPWR VGND sg13g2_decap_8
XFILLER_101_308 VPWR VGND sg13g2_decap_8
XFILLER_68_712 VPWR VGND sg13g2_decap_8
XFILLER_56_907 VPWR VGND sg13g2_decap_8
XFILLER_95_564 VPWR VGND sg13g2_decap_8
XFILLER_83_704 VPWR VGND sg13g2_decap_8
XFILLER_68_789 VPWR VGND sg13g2_decap_8
XFILLER_67_266 VPWR VGND sg13g2_decap_8
XFILLER_55_406 VPWR VGND sg13g2_decap_8
XFILLER_49_970 VPWR VGND sg13g2_decap_8
XFILLER_28_609 VPWR VGND sg13g2_decap_8
XFILLER_82_203 VPWR VGND sg13g2_decap_8
XFILLER_91_770 VPWR VGND sg13g2_decap_8
XFILLER_64_984 VPWR VGND sg13g2_decap_8
XFILLER_63_483 VPWR VGND sg13g2_decap_8
XFILLER_24_837 VPWR VGND sg13g2_decap_8
XFILLER_36_686 VPWR VGND sg13g2_decap_8
XFILLER_90_291 VPWR VGND sg13g2_decap_8
XFILLER_51_634 VPWR VGND sg13g2_decap_8
XFILLER_50_133 VPWR VGND sg13g2_decap_8
XFILLER_23_336 VPWR VGND sg13g2_decap_8
XFILLER_35_196 VPWR VGND sg13g2_decap_8
XFILLER_2_207 VPWR VGND sg13g2_decap_8
XFILLER_105_658 VPWR VGND sg13g2_decap_8
XFILLER_104_168 VPWR VGND sg13g2_decap_8
XFILLER_59_712 VPWR VGND sg13g2_decap_8
XFILLER_101_875 VPWR VGND sg13g2_decap_8
XFILLER_86_564 VPWR VGND sg13g2_decap_8
XFILLER_74_715 VPWR VGND sg13g2_decap_8
XFILLER_59_789 VPWR VGND sg13g2_decap_8
XFILLER_58_266 VPWR VGND sg13g2_decap_8
XFILLER_19_609 VPWR VGND sg13g2_decap_8
XFILLER_100_385 VPWR VGND sg13g2_decap_8
XFILLER_73_214 VPWR VGND sg13g2_decap_8
XFILLER_46_417 VPWR VGND sg13g2_decap_8
XFILLER_18_119 VPWR VGND sg13g2_decap_8
XFILLER_27_620 VPWR VGND sg13g2_decap_8
XFILLER_39_480 VPWR VGND sg13g2_decap_8
XFILLER_82_770 VPWR VGND sg13g2_decap_8
XFILLER_70_910 VPWR VGND sg13g2_decap_8
XFILLER_55_973 VPWR VGND sg13g2_decap_8
XFILLER_15_837 VPWR VGND sg13g2_decap_8
XFILLER_27_697 VPWR VGND sg13g2_decap_8
XFILLER_81_291 VPWR VGND sg13g2_decap_8
XFILLER_54_494 VPWR VGND sg13g2_decap_8
XFILLER_42_634 VPWR VGND sg13g2_decap_8
XFILLER_14_336 VPWR VGND sg13g2_decap_8
XFILLER_25_42 VPWR VGND sg13g2_decap_8
XFILLER_26_196 VPWR VGND sg13g2_decap_8
XFILLER_70_987 VPWR VGND sg13g2_decap_8
XFILLER_41_133 VPWR VGND sg13g2_decap_8
XFILLER_10_564 VPWR VGND sg13g2_decap_8
XFILLER_41_63 VPWR VGND sg13g2_decap_8
XFILLER_6_546 VPWR VGND sg13g2_decap_8
XFILLER_29_1005 VPWR VGND sg13g2_decap_8
XFILLER_2_774 VPWR VGND sg13g2_decap_8
XFILLER_49_200 VPWR VGND sg13g2_decap_8
XFILLER_1_273 VPWR VGND sg13g2_decap_8
XFILLER_77_553 VPWR VGND sg13g2_decap_8
X_51_ net6 net14 _18_ VPWR VGND sg13g2_nor2_1
XFILLER_2_46 VPWR VGND sg13g2_decap_8
XFILLER_64_214 VPWR VGND sg13g2_decap_8
XFILLER_49_277 VPWR VGND sg13g2_decap_8
XFILLER_37_417 VPWR VGND sg13g2_decap_8
XFILLER_92_567 VPWR VGND sg13g2_decap_8
XFILLER_80_707 VPWR VGND sg13g2_decap_8
XFILLER_17_130 VPWR VGND sg13g2_decap_8
XFILLER_73_781 VPWR VGND sg13g2_decap_8
XFILLER_61_921 VPWR VGND sg13g2_decap_8
XFILLER_46_984 VPWR VGND sg13g2_decap_8
XFILLER_18_686 VPWR VGND sg13g2_decap_8
XFILLER_72_280 VPWR VGND sg13g2_decap_8
XFILLER_60_431 VPWR VGND sg13g2_decap_8
XFILLER_45_483 VPWR VGND sg13g2_decap_8
XFILLER_33_623 VPWR VGND sg13g2_decap_8
XFILLER_82_70 VPWR VGND sg13g2_decap_8
XFILLER_61_998 VPWR VGND sg13g2_decap_8
XFILLER_32_144 VPWR VGND sg13g2_decap_8
XFILLER_99_133 VPWR VGND sg13g2_decap_8
XFILLER_101_105 VPWR VGND sg13g2_decap_8
XFILLER_96_840 VPWR VGND sg13g2_decap_8
XFILLER_56_704 VPWR VGND sg13g2_decap_8
XFILLER_28_406 VPWR VGND sg13g2_decap_8
XFILLER_29_907 VPWR VGND sg13g2_decap_8
XFILLER_95_361 VPWR VGND sg13g2_decap_8
XFILLER_83_501 VPWR VGND sg13g2_decap_8
XFILLER_68_586 VPWR VGND sg13g2_decap_8
XFILLER_55_203 VPWR VGND sg13g2_decap_8
XFILLER_102_14 VPWR VGND sg13g2_decap_8
XFILLER_83_578 VPWR VGND sg13g2_decap_8
XFILLER_71_718 VPWR VGND sg13g2_decap_8
XFILLER_70_217 VPWR VGND sg13g2_decap_8
XFILLER_64_781 VPWR VGND sg13g2_decap_8
XFILLER_52_910 VPWR VGND sg13g2_decap_8
XFILLER_37_984 VPWR VGND sg13g2_decap_8
XFILLER_63_280 VPWR VGND sg13g2_decap_8
XFILLER_51_431 VPWR VGND sg13g2_decap_8
XFILLER_24_634 VPWR VGND sg13g2_decap_8
XFILLER_36_483 VPWR VGND sg13g2_decap_8
XFILLER_52_987 VPWR VGND sg13g2_decap_8
XFILLER_23_133 VPWR VGND sg13g2_decap_8
XFILLER_20_851 VPWR VGND sg13g2_decap_8
XFILLER_106_945 VPWR VGND sg13g2_decap_8
XFILLER_11_77 VPWR VGND sg13g2_decap_8
XFILLER_105_455 VPWR VGND sg13g2_decap_8
XFILLER_87_840 VPWR VGND sg13g2_decap_8
XFILLER_78_328 VPWR VGND sg13g2_decap_8
XFILLER_101_672 VPWR VGND sg13g2_decap_8
XFILLER_86_361 VPWR VGND sg13g2_decap_8
XFILLER_74_512 VPWR VGND sg13g2_decap_8
XFILLER_59_586 VPWR VGND sg13g2_decap_8
XFILLER_46_214 VPWR VGND sg13g2_decap_8
XFILLER_19_406 VPWR VGND sg13g2_decap_8
XFILLER_100_182 VPWR VGND sg13g2_decap_8
XFILLER_62_707 VPWR VGND sg13g2_decap_8
XFILLER_74_589 VPWR VGND sg13g2_decap_8
XFILLER_55_770 VPWR VGND sg13g2_decap_8
XFILLER_43_910 VPWR VGND sg13g2_decap_8
XFILLER_28_973 VPWR VGND sg13g2_decap_8
XFILLER_36_63 VPWR VGND sg13g2_decap_8
XFILLER_61_228 VPWR VGND sg13g2_decap_8
XFILLER_42_431 VPWR VGND sg13g2_decap_8
XFILLER_15_634 VPWR VGND sg13g2_decap_8
XFILLER_27_494 VPWR VGND sg13g2_decap_8
XFILLER_54_291 VPWR VGND sg13g2_decap_8
XFILLER_43_987 VPWR VGND sg13g2_decap_8
XFILLER_14_133 VPWR VGND sg13g2_decap_8
XFILLER_70_784 VPWR VGND sg13g2_decap_8
XFILLER_30_637 VPWR VGND sg13g2_decap_8
XFILLER_52_84 VPWR VGND sg13g2_decap_8
XFILLER_11_840 VPWR VGND sg13g2_decap_8
Xinput16 uio_in[7] net16 VPWR VGND sg13g2_buf_1
XFILLER_10_361 VPWR VGND sg13g2_decap_8
XFILLER_7_844 VPWR VGND sg13g2_decap_8
XFILLER_6_343 VPWR VGND sg13g2_decap_8
XFILLER_97_637 VPWR VGND sg13g2_decap_8
XFILLER_2_571 VPWR VGND sg13g2_decap_8
XFILLER_96_147 VPWR VGND sg13g2_decap_8
XFILLER_77_350 VPWR VGND sg13g2_decap_8
XFILLER_77_70 VPWR VGND sg13g2_decap_8
XFILLER_93_810 VPWR VGND sg13g2_decap_8
XFILLER_78_895 VPWR VGND sg13g2_decap_8
XFILLER_37_214 VPWR VGND sg13g2_decap_8
X_34_ net3 net11 _04_ VPWR VGND sg13g2_and2_1
XFILLER_53_707 VPWR VGND sg13g2_decap_8
XFILLER_93_887 VPWR VGND sg13g2_decap_8
XFILLER_92_364 VPWR VGND sg13g2_decap_8
XFILLER_80_504 VPWR VGND sg13g2_decap_8
XFILLER_65_567 VPWR VGND sg13g2_decap_8
XFILLER_52_217 VPWR VGND sg13g2_decap_8
XFILLER_19_973 VPWR VGND sg13g2_decap_8
XFILLER_46_781 VPWR VGND sg13g2_decap_8
XFILLER_45_280 VPWR VGND sg13g2_decap_8
XFILLER_18_483 VPWR VGND sg13g2_decap_8
Xheichips25_example_large_34 VPWR VGND uio_out[1] sg13g2_tielo
XFILLER_33_420 VPWR VGND sg13g2_decap_8
XFILLER_34_921 VPWR VGND sg13g2_decap_8
XFILLER_61_795 VPWR VGND sg13g2_decap_8
XFILLER_21_637 VPWR VGND sg13g2_decap_8
XFILLER_33_497 VPWR VGND sg13g2_decap_8
XFILLER_34_998 VPWR VGND sg13g2_decap_8
XFILLER_20_158 VPWR VGND sg13g2_decap_8
XFILLER_103_959 VPWR VGND sg13g2_decap_8
XFILLER_88_648 VPWR VGND sg13g2_decap_8
XFILLER_102_469 VPWR VGND sg13g2_decap_8
XFILLER_87_147 VPWR VGND sg13g2_decap_8
XFILLER_69_862 VPWR VGND sg13g2_decap_8
XFILLER_29_704 VPWR VGND sg13g2_decap_8
XFILLER_68_383 VPWR VGND sg13g2_decap_8
XFILLER_56_501 VPWR VGND sg13g2_decap_8
XFILLER_28_203 VPWR VGND sg13g2_decap_8
XFILLER_84_854 VPWR VGND sg13g2_decap_8
XFILLER_83_375 VPWR VGND sg13g2_decap_8
XFILLER_71_515 VPWR VGND sg13g2_decap_8
XFILLER_56_578 VPWR VGND sg13g2_decap_8
XFILLER_44_718 VPWR VGND sg13g2_decap_8
XFILLER_25_910 VPWR VGND sg13g2_decap_8
XFILLER_73_39 VPWR VGND sg13g2_decap_8
XFILLER_43_217 VPWR VGND sg13g2_decap_8
XFILLER_36_280 VPWR VGND sg13g2_decap_8
XFILLER_37_781 VPWR VGND sg13g2_decap_8
XFILLER_19_1015 VPWR VGND sg13g2_decap_8
XFILLER_24_431 VPWR VGND sg13g2_decap_8
XFILLER_25_987 VPWR VGND sg13g2_decap_8
XFILLER_52_784 VPWR VGND sg13g2_decap_8
XFILLER_40_924 VPWR VGND sg13g2_decap_8
XFILLER_11_147 VPWR VGND sg13g2_decap_8
XFILLER_12_648 VPWR VGND sg13g2_decap_8
XFILLER_22_32 VPWR VGND sg13g2_decap_8
XFILLER_98_25 VPWR VGND sg13g2_decap_8
XFILLER_106_742 VPWR VGND sg13g2_decap_8
XFILLER_4_847 VPWR VGND sg13g2_decap_8
XFILLER_105_252 VPWR VGND sg13g2_decap_8
XFILLER_3_357 VPWR VGND sg13g2_decap_8
XFILLER_79_648 VPWR VGND sg13g2_decap_8
XFILLER_78_125 VPWR VGND sg13g2_decap_8
XFILLER_26_1008 VPWR VGND sg13g2_decap_8
XFILLER_93_117 VPWR VGND sg13g2_decap_8
XFILLER_59_383 VPWR VGND sg13g2_decap_8
XFILLER_19_203 VPWR VGND sg13g2_decap_8
XFILLER_75_854 VPWR VGND sg13g2_decap_8
XFILLER_90_802 VPWR VGND sg13g2_decap_8
XFILLER_62_504 VPWR VGND sg13g2_decap_8
XFILLER_47_567 VPWR VGND sg13g2_decap_8
XFILLER_47_84 VPWR VGND sg13g2_decap_8
XFILLER_16_910 VPWR VGND sg13g2_decap_8
XFILLER_28_770 VPWR VGND sg13g2_decap_8
XFILLER_35_707 VPWR VGND sg13g2_decap_8
XFILLER_74_386 VPWR VGND sg13g2_decap_8
XFILLER_34_228 VPWR VGND sg13g2_decap_8
XFILLER_90_879 VPWR VGND sg13g2_decap_8
XFILLER_15_431 VPWR VGND sg13g2_decap_8
XFILLER_16_987 VPWR VGND sg13g2_decap_8
XFILLER_27_291 VPWR VGND sg13g2_decap_8
XFILLER_70_581 VPWR VGND sg13g2_decap_8
XFILLER_43_784 VPWR VGND sg13g2_decap_8
XFILLER_31_924 VPWR VGND sg13g2_decap_8
XFILLER_30_434 VPWR VGND sg13g2_decap_8
XFILLER_8_56 VPWR VGND sg13g2_decap_8
XFILLER_7_641 VPWR VGND sg13g2_decap_8
XFILLER_6_140 VPWR VGND sg13g2_decap_8
XFILLER_98_935 VPWR VGND sg13g2_decap_8
XFILLER_97_434 VPWR VGND sg13g2_decap_8
XFILLER_69_169 VPWR VGND sg13g2_decap_8
XFILLER_78_692 VPWR VGND sg13g2_decap_8
XFILLER_66_832 VPWR VGND sg13g2_decap_8
XFILLER_93_684 VPWR VGND sg13g2_decap_8
XFILLER_81_802 VPWR VGND sg13g2_decap_8
XFILLER_80_301 VPWR VGND sg13g2_decap_8
XFILLER_65_364 VPWR VGND sg13g2_decap_8
XFILLER_53_504 VPWR VGND sg13g2_decap_8
XFILLER_19_770 VPWR VGND sg13g2_decap_8
XFILLER_26_707 VPWR VGND sg13g2_decap_8
XFILLER_38_567 VPWR VGND sg13g2_decap_8
XFILLER_92_161 VPWR VGND sg13g2_decap_8
XFILLER_25_217 VPWR VGND sg13g2_decap_8
XFILLER_81_879 VPWR VGND sg13g2_decap_8
XFILLER_18_280 VPWR VGND sg13g2_decap_8
XFILLER_80_378 VPWR VGND sg13g2_decap_8
XFILLER_22_935 VPWR VGND sg13g2_decap_8
XFILLER_34_795 VPWR VGND sg13g2_decap_8
XFILLER_61_592 VPWR VGND sg13g2_decap_8
XFILLER_21_434 VPWR VGND sg13g2_decap_8
XFILLER_33_294 VPWR VGND sg13g2_decap_8
XFILLER_49_1019 VPWR VGND sg13g2_decap_8
XFILLER_89_924 VPWR VGND sg13g2_decap_8
XFILLER_68_39 VPWR VGND sg13g2_decap_8
XFILLER_103_756 VPWR VGND sg13g2_decap_8
XFILLER_88_445 VPWR VGND sg13g2_decap_8
XFILLER_102_266 VPWR VGND sg13g2_decap_8
XFILLER_29_501 VPWR VGND sg13g2_decap_8
XFILLER_68_180 VPWR VGND sg13g2_decap_8
XFILLER_57_854 VPWR VGND sg13g2_decap_8
XFILLER_90_109 VPWR VGND sg13g2_decap_8
XFILLER_84_651 VPWR VGND sg13g2_decap_8
XFILLER_84_49 VPWR VGND sg13g2_decap_8
XFILLER_44_515 VPWR VGND sg13g2_decap_8
XFILLER_17_32 VPWR VGND sg13g2_decap_8
XFILLER_17_718 VPWR VGND sg13g2_decap_8
XFILLER_29_578 VPWR VGND sg13g2_decap_8
XFILLER_95_1028 VPWR VGND sg13g2_fill_1
XFILLER_83_172 VPWR VGND sg13g2_decap_8
XFILLER_71_312 VPWR VGND sg13g2_decap_8
XFILLER_56_375 VPWR VGND sg13g2_decap_8
XFILLER_16_217 VPWR VGND sg13g2_decap_8
XFILLER_72_868 VPWR VGND sg13g2_decap_8
XFILLER_71_389 VPWR VGND sg13g2_decap_8
XFILLER_52_581 VPWR VGND sg13g2_decap_8
XFILLER_13_924 VPWR VGND sg13g2_decap_8
XFILLER_25_784 VPWR VGND sg13g2_decap_8
XFILLER_40_721 VPWR VGND sg13g2_decap_8
XFILLER_9_917 VPWR VGND sg13g2_decap_8
XFILLER_12_445 VPWR VGND sg13g2_decap_8
XFILLER_33_42 VPWR VGND sg13g2_decap_8
XFILLER_8_427 VPWR VGND sg13g2_decap_8
XFILLER_32_1012 VPWR VGND sg13g2_decap_8
XFILLER_40_798 VPWR VGND sg13g2_decap_8
XFILLER_4_644 VPWR VGND sg13g2_decap_8
XFILLER_3_154 VPWR VGND sg13g2_decap_8
XFILLER_79_445 VPWR VGND sg13g2_decap_8
XFILLER_95_949 VPWR VGND sg13g2_decap_8
XFILLER_0_861 VPWR VGND sg13g2_decap_8
XFILLER_94_448 VPWR VGND sg13g2_decap_8
XFILLER_66_139 VPWR VGND sg13g2_decap_8
XFILLER_59_180 VPWR VGND sg13g2_decap_8
XFILLER_48_854 VPWR VGND sg13g2_decap_8
XFILLER_81_109 VPWR VGND sg13g2_decap_8
XFILLER_75_651 VPWR VGND sg13g2_decap_8
XFILLER_47_364 VPWR VGND sg13g2_decap_8
XFILLER_35_504 VPWR VGND sg13g2_decap_8
XFILLER_74_183 VPWR VGND sg13g2_decap_8
XFILLER_62_301 VPWR VGND sg13g2_decap_8
XFILLER_90_676 VPWR VGND sg13g2_decap_8
XFILLER_74_71 VPWR VGND sg13g2_decap_8
XFILLER_63_868 VPWR VGND sg13g2_decap_8
XFILLER_62_378 VPWR VGND sg13g2_decap_8
XFILLER_50_518 VPWR VGND sg13g2_decap_8
XFILLER_16_784 VPWR VGND sg13g2_decap_8
XFILLER_31_721 VPWR VGND sg13g2_decap_8
XFILLER_43_581 VPWR VGND sg13g2_decap_8
XFILLER_30_231 VPWR VGND sg13g2_decap_8
XFILLER_90_81 VPWR VGND sg13g2_decap_8
XFILLER_88_4 VPWR VGND sg13g2_decap_8
XFILLER_31_798 VPWR VGND sg13g2_decap_8
XFILLER_8_994 VPWR VGND sg13g2_decap_8
XFILLER_98_732 VPWR VGND sg13g2_decap_8
XFILLER_97_231 VPWR VGND sg13g2_decap_8
XFILLER_31_0 VPWR VGND sg13g2_decap_8
XFILLER_86_949 VPWR VGND sg13g2_decap_8
XFILLER_85_448 VPWR VGND sg13g2_decap_8
XFILLER_54_802 VPWR VGND sg13g2_decap_8
XFILLER_26_504 VPWR VGND sg13g2_decap_8
XFILLER_38_364 VPWR VGND sg13g2_decap_8
XFILLER_39_865 VPWR VGND sg13g2_decap_8
XFILLER_93_481 VPWR VGND sg13g2_decap_8
XFILLER_65_161 VPWR VGND sg13g2_decap_8
XFILLER_53_301 VPWR VGND sg13g2_decap_8
XFILLER_54_879 VPWR VGND sg13g2_decap_8
XFILLER_81_676 VPWR VGND sg13g2_decap_8
XFILLER_80_175 VPWR VGND sg13g2_decap_8
XFILLER_55_1001 VPWR VGND sg13g2_decap_8
XFILLER_53_378 VPWR VGND sg13g2_decap_8
XFILLER_41_518 VPWR VGND sg13g2_decap_8
XFILLER_22_732 VPWR VGND sg13g2_decap_8
XFILLER_34_592 VPWR VGND sg13g2_decap_8
XFILLER_21_231 VPWR VGND sg13g2_decap_8
XFILLER_10_949 VPWR VGND sg13g2_decap_8
XFILLER_79_49 VPWR VGND sg13g2_decap_8
XFILLER_89_721 VPWR VGND sg13g2_decap_8
XFILLER_103_553 VPWR VGND sg13g2_decap_8
XFILLER_88_242 VPWR VGND sg13g2_decap_8
XFILLER_1_658 VPWR VGND sg13g2_decap_8
XFILLER_89_798 VPWR VGND sg13g2_decap_8
XFILLER_77_938 VPWR VGND sg13g2_decap_8
XFILLER_0_168 VPWR VGND sg13g2_decap_8
XFILLER_76_459 VPWR VGND sg13g2_decap_8
XFILLER_57_651 VPWR VGND sg13g2_decap_8
XFILLER_28_42 VPWR VGND sg13g2_decap_8
XFILLER_56_172 VPWR VGND sg13g2_decap_8
XFILLER_44_312 VPWR VGND sg13g2_decap_8
XFILLER_17_515 VPWR VGND sg13g2_decap_8
XFILLER_29_375 VPWR VGND sg13g2_decap_8
XFILLER_72_665 VPWR VGND sg13g2_decap_8
XFILLER_45_868 VPWR VGND sg13g2_decap_8
XFILLER_60_816 VPWR VGND sg13g2_decap_8
XFILLER_44_389 VPWR VGND sg13g2_decap_8
XFILLER_32_529 VPWR VGND sg13g2_decap_8
XFILLER_71_186 VPWR VGND sg13g2_decap_8
XFILLER_44_74 VPWR VGND sg13g2_decap_8
XFILLER_13_721 VPWR VGND sg13g2_decap_8
XFILLER_25_581 VPWR VGND sg13g2_decap_8
XFILLER_9_714 VPWR VGND sg13g2_decap_8
XFILLER_12_242 VPWR VGND sg13g2_decap_8
XFILLER_100_91 VPWR VGND sg13g2_decap_8
XFILLER_8_224 VPWR VGND sg13g2_decap_8
XFILLER_13_798 VPWR VGND sg13g2_decap_8
XFILLER_40_595 VPWR VGND sg13g2_decap_8
XFILLER_60_95 VPWR VGND sg13g2_decap_8
XFILLER_5_942 VPWR VGND sg13g2_decap_8
XFILLER_99_518 VPWR VGND sg13g2_decap_8
XFILLER_5_46 VPWR VGND sg13g2_decap_8
XFILLER_4_441 VPWR VGND sg13g2_decap_8
XFILLER_79_242 VPWR VGND sg13g2_decap_8
XFILLER_69_71 VPWR VGND sg13g2_decap_8
XFILLER_95_746 VPWR VGND sg13g2_decap_8
XFILLER_67_448 VPWR VGND sg13g2_decap_8
XFILLER_94_245 VPWR VGND sg13g2_decap_8
XFILLER_85_70 VPWR VGND sg13g2_decap_8
XFILLER_54_109 VPWR VGND sg13g2_decap_8
XFILLER_48_651 VPWR VGND sg13g2_decap_8
XFILLER_47_161 VPWR VGND sg13g2_decap_8
XFILLER_35_301 VPWR VGND sg13g2_decap_8
XFILLER_91_952 VPWR VGND sg13g2_decap_8
XFILLER_63_665 VPWR VGND sg13g2_decap_8
XFILLER_36_868 VPWR VGND sg13g2_decap_8
XFILLER_90_473 VPWR VGND sg13g2_decap_8
XFILLER_62_175 VPWR VGND sg13g2_decap_8
XFILLER_51_816 VPWR VGND sg13g2_decap_8
XFILLER_50_315 VPWR VGND sg13g2_decap_8
XFILLER_23_518 VPWR VGND sg13g2_decap_8
XFILLER_35_378 VPWR VGND sg13g2_decap_8
XFILLER_16_581 VPWR VGND sg13g2_decap_8
XFILLER_31_595 VPWR VGND sg13g2_decap_8
XFILLER_79_0 VPWR VGND sg13g2_decap_8
XFILLER_8_791 VPWR VGND sg13g2_decap_8
XFILLER_105_14 VPWR VGND sg13g2_decap_8
XFILLER_86_746 VPWR VGND sg13g2_decap_8
XFILLER_58_448 VPWR VGND sg13g2_decap_8
XFILLER_100_567 VPWR VGND sg13g2_decap_8
XFILLER_85_245 VPWR VGND sg13g2_decap_8
XFILLER_27_802 VPWR VGND sg13g2_decap_8
XFILLER_39_662 VPWR VGND sg13g2_decap_8
XFILLER_26_301 VPWR VGND sg13g2_decap_8
XFILLER_38_161 VPWR VGND sg13g2_decap_8
XFILLER_82_952 VPWR VGND sg13g2_decap_8
XFILLER_27_879 VPWR VGND sg13g2_decap_8
XFILLER_81_473 VPWR VGND sg13g2_decap_8
XFILLER_54_676 VPWR VGND sg13g2_decap_8
XFILLER_53_175 VPWR VGND sg13g2_decap_8
XFILLER_42_816 VPWR VGND sg13g2_decap_8
XFILLER_14_518 VPWR VGND sg13g2_decap_8
XFILLER_26_378 VPWR VGND sg13g2_decap_8
XFILLER_41_315 VPWR VGND sg13g2_decap_8
XFILLER_81_39 VPWR VGND sg13g2_decap_8
XFILLER_50_882 VPWR VGND sg13g2_decap_8
XFILLER_14_77 VPWR VGND sg13g2_decap_8
XFILLER_10_746 VPWR VGND sg13g2_decap_8
XFILLER_6_728 VPWR VGND sg13g2_decap_8
XFILLER_30_21 VPWR VGND sg13g2_decap_8
XFILLER_5_249 VPWR VGND sg13g2_decap_8
XFILLER_30_98 VPWR VGND sg13g2_decap_8
XFILLER_104_840 VPWR VGND sg13g2_decap_8
XFILLER_2_956 VPWR VGND sg13g2_decap_8
XFILLER_103_350 VPWR VGND sg13g2_decap_8
XFILLER_7_1005 VPWR VGND sg13g2_decap_8
XFILLER_1_455 VPWR VGND sg13g2_decap_8
XFILLER_89_595 VPWR VGND sg13g2_decap_8
XFILLER_77_735 VPWR VGND sg13g2_decap_8
XFILLER_39_74 VPWR VGND sg13g2_decap_8
XFILLER_76_256 VPWR VGND sg13g2_decap_8
XFILLER_49_459 VPWR VGND sg13g2_decap_8
XFILLER_92_749 VPWR VGND sg13g2_decap_8
XFILLER_17_312 VPWR VGND sg13g2_decap_8
XFILLER_29_172 VPWR VGND sg13g2_decap_8
XFILLER_91_259 VPWR VGND sg13g2_decap_8
XFILLER_73_963 VPWR VGND sg13g2_decap_8
XFILLER_18_868 VPWR VGND sg13g2_decap_8
XFILLER_72_462 VPWR VGND sg13g2_decap_8
XFILLER_60_613 VPWR VGND sg13g2_decap_8
XFILLER_55_84 VPWR VGND sg13g2_decap_8
XFILLER_45_665 VPWR VGND sg13g2_decap_8
XFILLER_17_389 VPWR VGND sg13g2_decap_8
XFILLER_33_805 VPWR VGND sg13g2_decap_8
XFILLER_44_186 VPWR VGND sg13g2_decap_8
XFILLER_32_326 VPWR VGND sg13g2_decap_8
XFILLER_41_882 VPWR VGND sg13g2_decap_8
XFILLER_9_511 VPWR VGND sg13g2_decap_8
XFILLER_13_595 VPWR VGND sg13g2_decap_8
XFILLER_72_7 VPWR VGND sg13g2_decap_8
XFILLER_40_392 VPWR VGND sg13g2_decap_8
XFILLER_9_588 VPWR VGND sg13g2_decap_8
XFILLER_99_315 VPWR VGND sg13g2_decap_8
XFILLER_45_1022 VPWR VGND sg13g2_decap_8
XFILLER_95_543 VPWR VGND sg13g2_decap_8
XFILLER_96_91 VPWR VGND sg13g2_decap_8
XFILLER_68_768 VPWR VGND sg13g2_decap_8
XFILLER_67_245 VPWR VGND sg13g2_decap_8
XFILLER_27_109 VPWR VGND sg13g2_decap_8
XFILLER_82_259 VPWR VGND sg13g2_decap_8
XFILLER_64_963 VPWR VGND sg13g2_decap_8
XFILLER_63_462 VPWR VGND sg13g2_decap_8
XFILLER_51_613 VPWR VGND sg13g2_decap_8
XFILLER_24_816 VPWR VGND sg13g2_decap_8
XFILLER_36_665 VPWR VGND sg13g2_decap_8
XFILLER_90_270 VPWR VGND sg13g2_decap_8
XFILLER_50_112 VPWR VGND sg13g2_decap_8
XFILLER_23_315 VPWR VGND sg13g2_decap_8
XFILLER_35_175 VPWR VGND sg13g2_decap_8
XFILLER_52_1015 VPWR VGND sg13g2_decap_8
XFILLER_50_189 VPWR VGND sg13g2_decap_8
XFILLER_32_893 VPWR VGND sg13g2_decap_8
XFILLER_31_392 VPWR VGND sg13g2_decap_8
XFILLER_105_637 VPWR VGND sg13g2_decap_8
XFILLER_104_147 VPWR VGND sg13g2_decap_8
XFILLER_99_882 VPWR VGND sg13g2_decap_8
XFILLER_76_39 VPWR VGND sg13g2_decap_8
XFILLER_101_854 VPWR VGND sg13g2_decap_8
XFILLER_86_543 VPWR VGND sg13g2_decap_8
XFILLER_59_768 VPWR VGND sg13g2_decap_8
XFILLER_58_245 VPWR VGND sg13g2_decap_8
XFILLER_100_364 VPWR VGND sg13g2_decap_8
XFILLER_55_952 VPWR VGND sg13g2_decap_8
XFILLER_92_49 VPWR VGND sg13g2_decap_8
XFILLER_54_473 VPWR VGND sg13g2_decap_8
XFILLER_42_613 VPWR VGND sg13g2_decap_8
XFILLER_15_816 VPWR VGND sg13g2_decap_8
XFILLER_25_21 VPWR VGND sg13g2_decap_8
XFILLER_27_676 VPWR VGND sg13g2_decap_8
XFILLER_81_270 VPWR VGND sg13g2_decap_8
XFILLER_14_315 VPWR VGND sg13g2_decap_8
XFILLER_26_175 VPWR VGND sg13g2_decap_8
XFILLER_41_112 VPWR VGND sg13g2_decap_8
XFILLER_70_966 VPWR VGND sg13g2_decap_8
XFILLER_30_819 VPWR VGND sg13g2_decap_8
XFILLER_23_882 VPWR VGND sg13g2_decap_8
XFILLER_25_98 VPWR VGND sg13g2_decap_8
XFILLER_41_189 VPWR VGND sg13g2_decap_8
XFILLER_10_543 VPWR VGND sg13g2_decap_8
XFILLER_6_525 VPWR VGND sg13g2_decap_8
XFILLER_41_42 VPWR VGND sg13g2_decap_8
XFILLER_9_0 VPWR VGND sg13g2_decap_8
XFILLER_29_1028 VPWR VGND sg13g2_fill_1
XFILLER_97_819 VPWR VGND sg13g2_decap_8
XFILLER_2_753 VPWR VGND sg13g2_decap_8
XFILLER_1_252 VPWR VGND sg13g2_decap_8
XFILLER_96_329 VPWR VGND sg13g2_decap_8
XFILLER_89_392 VPWR VGND sg13g2_decap_8
XFILLER_77_532 VPWR VGND sg13g2_decap_8
XFILLER_2_25 VPWR VGND sg13g2_decap_8
X_50_ net21 _13_ _16_ VPWR VGND sg13g2_xnor2_1
XFILLER_49_256 VPWR VGND sg13g2_decap_8
XFILLER_65_749 VPWR VGND sg13g2_decap_8
XFILLER_92_546 VPWR VGND sg13g2_decap_8
XFILLER_66_83 VPWR VGND sg13g2_decap_8
XFILLER_46_963 VPWR VGND sg13g2_decap_8
XFILLER_75_1015 VPWR VGND sg13g2_decap_8
XFILLER_73_760 VPWR VGND sg13g2_decap_8
XFILLER_61_900 VPWR VGND sg13g2_decap_8
XFILLER_45_462 VPWR VGND sg13g2_decap_8
XFILLER_18_665 VPWR VGND sg13g2_decap_8
XFILLER_33_602 VPWR VGND sg13g2_decap_8
XFILLER_60_410 VPWR VGND sg13g2_decap_8
XFILLER_17_186 VPWR VGND sg13g2_decap_8
XFILLER_32_123 VPWR VGND sg13g2_decap_8
XFILLER_61_977 VPWR VGND sg13g2_decap_8
XFILLER_21_819 VPWR VGND sg13g2_decap_8
XFILLER_33_679 VPWR VGND sg13g2_decap_8
XFILLER_60_487 VPWR VGND sg13g2_decap_8
XFILLER_14_882 VPWR VGND sg13g2_decap_8
XFILLER_13_392 VPWR VGND sg13g2_decap_8
XFILLER_9_385 VPWR VGND sg13g2_decap_8
XFILLER_99_112 VPWR VGND sg13g2_decap_8
XFILLER_82_1008 VPWR VGND sg13g2_decap_8
XFILLER_99_189 VPWR VGND sg13g2_decap_8
XFILLER_87_329 VPWR VGND sg13g2_decap_8
XFILLER_95_340 VPWR VGND sg13g2_decap_8
XFILLER_68_565 VPWR VGND sg13g2_decap_8
XFILLER_96_896 VPWR VGND sg13g2_decap_8
XFILLER_83_557 VPWR VGND sg13g2_decap_8
XFILLER_64_760 VPWR VGND sg13g2_decap_8
XFILLER_55_259 VPWR VGND sg13g2_decap_8
XFILLER_36_462 VPWR VGND sg13g2_decap_8
XFILLER_37_963 VPWR VGND sg13g2_decap_8
XFILLER_51_410 VPWR VGND sg13g2_decap_8
XFILLER_23_112 VPWR VGND sg13g2_decap_8
XFILLER_24_613 VPWR VGND sg13g2_decap_8
XFILLER_52_966 VPWR VGND sg13g2_decap_8
XFILLER_51_487 VPWR VGND sg13g2_decap_8
XFILLER_11_329 VPWR VGND sg13g2_decap_8
XFILLER_23_189 VPWR VGND sg13g2_decap_8
XFILLER_20_830 VPWR VGND sg13g2_decap_8
XFILLER_32_690 VPWR VGND sg13g2_decap_8
XFILLER_106_924 VPWR VGND sg13g2_decap_8
XFILLER_11_56 VPWR VGND sg13g2_decap_8
XFILLER_105_434 VPWR VGND sg13g2_decap_8
XFILLER_3_539 VPWR VGND sg13g2_decap_8
XFILLER_87_49 VPWR VGND sg13g2_decap_8
XFILLER_78_307 VPWR VGND sg13g2_decap_8
XFILLER_101_651 VPWR VGND sg13g2_decap_8
XFILLER_86_340 VPWR VGND sg13g2_decap_8
XFILLER_59_565 VPWR VGND sg13g2_decap_8
XFILLER_100_161 VPWR VGND sg13g2_decap_8
XFILLER_98_1026 VPWR VGND sg13g2_fill_2
XFILLER_87_896 VPWR VGND sg13g2_decap_8
XFILLER_4_1008 VPWR VGND sg13g2_decap_8
XFILLER_47_749 VPWR VGND sg13g2_decap_8
XFILLER_28_952 VPWR VGND sg13g2_decap_8
XFILLER_74_568 VPWR VGND sg13g2_decap_8
XFILLER_61_207 VPWR VGND sg13g2_decap_8
XFILLER_36_42 VPWR VGND sg13g2_decap_8
XFILLER_54_270 VPWR VGND sg13g2_decap_8
XFILLER_42_410 VPWR VGND sg13g2_decap_8
XFILLER_14_112 VPWR VGND sg13g2_decap_8
XFILLER_15_613 VPWR VGND sg13g2_decap_8
XFILLER_27_473 VPWR VGND sg13g2_decap_8
XFILLER_70_763 VPWR VGND sg13g2_decap_8
XFILLER_43_966 VPWR VGND sg13g2_decap_8
XFILLER_42_487 VPWR VGND sg13g2_decap_8
XFILLER_14_189 VPWR VGND sg13g2_decap_8
XFILLER_30_616 VPWR VGND sg13g2_decap_8
XFILLER_52_63 VPWR VGND sg13g2_decap_8
XFILLER_10_340 VPWR VGND sg13g2_decap_8
XFILLER_7_823 VPWR VGND sg13g2_decap_8
XFILLER_6_322 VPWR VGND sg13g2_decap_8
XFILLER_11_896 VPWR VGND sg13g2_decap_8
XFILLER_6_399 VPWR VGND sg13g2_decap_8
XFILLER_97_616 VPWR VGND sg13g2_decap_8
XFILLER_2_550 VPWR VGND sg13g2_decap_8
XFILLER_96_126 VPWR VGND sg13g2_decap_8
XFILLER_35_7 VPWR VGND sg13g2_decap_8
XFILLER_78_874 VPWR VGND sg13g2_decap_8
X_33_ VGND VPWR _01_ _03_ _02_ _00_ sg13g2_a21oi_2
XFILLER_93_866 VPWR VGND sg13g2_decap_8
XFILLER_92_343 VPWR VGND sg13g2_decap_8
XFILLER_65_546 VPWR VGND sg13g2_decap_8
XFILLER_19_952 VPWR VGND sg13g2_decap_8
XFILLER_38_749 VPWR VGND sg13g2_decap_8
XFILLER_46_760 VPWR VGND sg13g2_decap_8
XFILLER_18_462 VPWR VGND sg13g2_decap_8
XFILLER_34_900 VPWR VGND sg13g2_decap_8
Xheichips25_example_large_35 VPWR VGND uio_out[2] sg13g2_tielo
XFILLER_34_977 VPWR VGND sg13g2_decap_8
XFILLER_61_774 VPWR VGND sg13g2_decap_8
XFILLER_21_616 VPWR VGND sg13g2_decap_8
XFILLER_33_476 VPWR VGND sg13g2_decap_8
XFILLER_60_284 VPWR VGND sg13g2_decap_8
XFILLER_20_137 VPWR VGND sg13g2_decap_8
XFILLER_9_182 VPWR VGND sg13g2_decap_8
XFILLER_103_938 VPWR VGND sg13g2_decap_8
XFILLER_88_627 VPWR VGND sg13g2_decap_8
XFILLER_87_126 VPWR VGND sg13g2_decap_8
XFILLER_102_448 VPWR VGND sg13g2_decap_8
XFILLER_69_841 VPWR VGND sg13g2_decap_8
XFILLER_68_362 VPWR VGND sg13g2_decap_8
XFILLER_96_693 VPWR VGND sg13g2_decap_8
XFILLER_84_833 VPWR VGND sg13g2_decap_8
XFILLER_56_557 VPWR VGND sg13g2_decap_8
XFILLER_83_354 VPWR VGND sg13g2_decap_8
XFILLER_73_18 VPWR VGND sg13g2_decap_8
XFILLER_28_259 VPWR VGND sg13g2_decap_8
XFILLER_37_760 VPWR VGND sg13g2_decap_8
XFILLER_24_410 VPWR VGND sg13g2_decap_8
XFILLER_52_763 VPWR VGND sg13g2_decap_8
XFILLER_25_966 VPWR VGND sg13g2_decap_8
XFILLER_40_903 VPWR VGND sg13g2_decap_8
XFILLER_106_1008 VPWR VGND sg13g2_decap_8
XFILLER_12_627 VPWR VGND sg13g2_decap_8
XFILLER_24_487 VPWR VGND sg13g2_decap_8
XFILLER_51_284 VPWR VGND sg13g2_decap_8
XFILLER_8_609 VPWR VGND sg13g2_decap_8
XFILLER_11_126 VPWR VGND sg13g2_decap_8
XFILLER_22_11 VPWR VGND sg13g2_decap_8
XFILLER_4_826 VPWR VGND sg13g2_decap_8
XFILLER_22_88 VPWR VGND sg13g2_decap_8
XFILLER_106_721 VPWR VGND sg13g2_decap_8
XFILLER_3_336 VPWR VGND sg13g2_decap_8
XFILLER_105_231 VPWR VGND sg13g2_decap_8
XFILLER_106_798 VPWR VGND sg13g2_decap_8
XFILLER_79_627 VPWR VGND sg13g2_decap_8
XFILLER_78_104 VPWR VGND sg13g2_decap_8
XFILLER_59_362 VPWR VGND sg13g2_decap_8
XFILLER_87_693 VPWR VGND sg13g2_decap_8
XFILLER_75_833 VPWR VGND sg13g2_decap_8
XFILLER_47_546 VPWR VGND sg13g2_decap_8
XFILLER_47_63 VPWR VGND sg13g2_decap_8
XFILLER_74_365 VPWR VGND sg13g2_decap_8
XFILLER_19_259 VPWR VGND sg13g2_decap_8
XFILLER_34_207 VPWR VGND sg13g2_decap_8
XFILLER_90_858 VPWR VGND sg13g2_decap_8
XFILLER_15_410 VPWR VGND sg13g2_decap_8
XFILLER_27_270 VPWR VGND sg13g2_decap_8
XFILLER_103_91 VPWR VGND sg13g2_decap_8
XFILLER_43_763 VPWR VGND sg13g2_decap_8
XFILLER_16_966 VPWR VGND sg13g2_decap_8
XFILLER_31_903 VPWR VGND sg13g2_decap_8
XFILLER_70_560 VPWR VGND sg13g2_decap_8
XFILLER_63_84 VPWR VGND sg13g2_decap_8
XFILLER_15_487 VPWR VGND sg13g2_decap_8
XFILLER_30_413 VPWR VGND sg13g2_decap_8
XFILLER_42_284 VPWR VGND sg13g2_decap_8
XFILLER_8_35 VPWR VGND sg13g2_decap_8
XFILLER_7_620 VPWR VGND sg13g2_decap_8
XFILLER_11_693 VPWR VGND sg13g2_decap_8
XFILLER_7_697 VPWR VGND sg13g2_decap_8
XFILLER_98_914 VPWR VGND sg13g2_decap_8
XFILLER_6_196 VPWR VGND sg13g2_decap_8
XFILLER_97_413 VPWR VGND sg13g2_decap_8
XFILLER_88_81 VPWR VGND sg13g2_decap_8
XFILLER_69_148 VPWR VGND sg13g2_decap_8
XFILLER_78_671 VPWR VGND sg13g2_decap_8
XFILLER_66_811 VPWR VGND sg13g2_decap_8
XFILLER_38_546 VPWR VGND sg13g2_decap_8
XFILLER_93_663 VPWR VGND sg13g2_decap_8
XFILLER_92_140 VPWR VGND sg13g2_decap_8
XFILLER_66_888 VPWR VGND sg13g2_decap_8
XFILLER_65_343 VPWR VGND sg13g2_decap_8
XFILLER_81_858 VPWR VGND sg13g2_decap_8
XFILLER_80_357 VPWR VGND sg13g2_decap_8
XFILLER_61_571 VPWR VGND sg13g2_decap_8
XFILLER_21_413 VPWR VGND sg13g2_decap_8
XFILLER_22_914 VPWR VGND sg13g2_decap_8
XFILLER_34_774 VPWR VGND sg13g2_decap_8
XFILLER_33_273 VPWR VGND sg13g2_decap_8
XFILLER_30_980 VPWR VGND sg13g2_decap_8
XFILLER_89_903 VPWR VGND sg13g2_decap_8
XFILLER_103_735 VPWR VGND sg13g2_decap_8
XFILLER_88_424 VPWR VGND sg13g2_decap_8
XFILLER_68_18 VPWR VGND sg13g2_decap_8
XFILLER_102_245 VPWR VGND sg13g2_decap_8
XFILLER_97_980 VPWR VGND sg13g2_decap_8
XFILLER_96_490 VPWR VGND sg13g2_decap_8
XFILLER_84_630 VPWR VGND sg13g2_decap_8
XFILLER_84_28 VPWR VGND sg13g2_decap_8
XFILLER_57_833 VPWR VGND sg13g2_decap_8
XFILLER_83_151 VPWR VGND sg13g2_decap_8
XFILLER_56_354 VPWR VGND sg13g2_decap_8
XFILLER_17_11 VPWR VGND sg13g2_decap_8
XFILLER_29_557 VPWR VGND sg13g2_decap_8
XFILLER_72_847 VPWR VGND sg13g2_decap_8
XFILLER_17_88 VPWR VGND sg13g2_decap_8
XFILLER_71_368 VPWR VGND sg13g2_decap_8
XFILLER_52_560 VPWR VGND sg13g2_decap_8
XFILLER_13_903 VPWR VGND sg13g2_decap_8
XFILLER_25_763 VPWR VGND sg13g2_decap_8
XFILLER_40_700 VPWR VGND sg13g2_decap_8
XFILLER_12_424 VPWR VGND sg13g2_decap_8
XFILLER_24_284 VPWR VGND sg13g2_decap_8
XFILLER_33_21 VPWR VGND sg13g2_decap_8
XFILLER_8_406 VPWR VGND sg13g2_decap_8
XFILLER_40_777 VPWR VGND sg13g2_decap_8
XFILLER_21_980 VPWR VGND sg13g2_decap_8
XFILLER_33_98 VPWR VGND sg13g2_decap_8
XFILLER_4_623 VPWR VGND sg13g2_decap_8
XFILLER_3_133 VPWR VGND sg13g2_decap_8
XFILLER_79_424 VPWR VGND sg13g2_decap_8
XFILLER_106_595 VPWR VGND sg13g2_decap_8
XFILLER_0_840 VPWR VGND sg13g2_decap_8
XFILLER_95_928 VPWR VGND sg13g2_decap_8
XFILLER_94_427 VPWR VGND sg13g2_decap_8
XFILLER_66_118 VPWR VGND sg13g2_decap_8
XFILLER_88_991 VPWR VGND sg13g2_decap_8
XFILLER_87_490 VPWR VGND sg13g2_decap_8
XFILLER_75_630 VPWR VGND sg13g2_decap_8
XFILLER_58_84 VPWR VGND sg13g2_decap_8
XFILLER_48_833 VPWR VGND sg13g2_decap_8
XFILLER_47_343 VPWR VGND sg13g2_decap_8
XFILLER_74_162 VPWR VGND sg13g2_decap_8
XFILLER_63_847 VPWR VGND sg13g2_decap_8
XFILLER_90_655 VPWR VGND sg13g2_decap_8
XFILLER_62_357 VPWR VGND sg13g2_decap_8
XFILLER_43_560 VPWR VGND sg13g2_decap_8
XFILLER_16_763 VPWR VGND sg13g2_decap_8
XFILLER_31_700 VPWR VGND sg13g2_decap_8
XFILLER_15_284 VPWR VGND sg13g2_decap_8
XFILLER_30_210 VPWR VGND sg13g2_decap_8
XFILLER_90_60 VPWR VGND sg13g2_decap_8
XFILLER_31_777 VPWR VGND sg13g2_decap_8
XFILLER_12_991 VPWR VGND sg13g2_decap_8
XFILLER_30_287 VPWR VGND sg13g2_decap_8
XFILLER_8_973 VPWR VGND sg13g2_decap_8
XFILLER_11_490 VPWR VGND sg13g2_decap_8
XFILLER_7_494 VPWR VGND sg13g2_decap_8
XFILLER_99_91 VPWR VGND sg13g2_decap_8
XFILLER_98_711 VPWR VGND sg13g2_decap_8
XFILLER_97_210 VPWR VGND sg13g2_decap_8
XFILLER_98_788 VPWR VGND sg13g2_decap_8
XFILLER_86_928 VPWR VGND sg13g2_decap_8
XFILLER_100_749 VPWR VGND sg13g2_decap_8
XFILLER_97_287 VPWR VGND sg13g2_decap_8
XFILLER_85_427 VPWR VGND sg13g2_decap_8
XFILLER_79_991 VPWR VGND sg13g2_decap_8
XFILLER_39_844 VPWR VGND sg13g2_decap_8
XFILLER_65_140 VPWR VGND sg13g2_decap_8
XFILLER_38_343 VPWR VGND sg13g2_decap_8
XFILLER_94_994 VPWR VGND sg13g2_decap_8
XFILLER_93_460 VPWR VGND sg13g2_decap_8
XFILLER_66_685 VPWR VGND sg13g2_decap_8
XFILLER_81_655 VPWR VGND sg13g2_decap_8
XFILLER_54_858 VPWR VGND sg13g2_decap_8
XFILLER_53_357 VPWR VGND sg13g2_decap_8
XFILLER_0_1022 VPWR VGND sg13g2_decap_8
XFILLER_80_154 VPWR VGND sg13g2_decap_8
XFILLER_0_91 VPWR VGND sg13g2_decap_8
XFILLER_22_711 VPWR VGND sg13g2_decap_8
XFILLER_34_571 VPWR VGND sg13g2_decap_8
XFILLER_16_1008 VPWR VGND sg13g2_decap_8
XFILLER_21_210 VPWR VGND sg13g2_decap_8
XFILLER_10_928 VPWR VGND sg13g2_decap_8
XFILLER_21_287 VPWR VGND sg13g2_decap_8
XFILLER_22_788 VPWR VGND sg13g2_decap_8
XFILLER_102_7 VPWR VGND sg13g2_decap_8
XFILLER_79_28 VPWR VGND sg13g2_decap_8
XFILLER_89_700 VPWR VGND sg13g2_decap_8
XFILLER_103_532 VPWR VGND sg13g2_decap_8
XFILLER_88_221 VPWR VGND sg13g2_decap_8
XFILLER_1_637 VPWR VGND sg13g2_decap_8
XFILLER_89_777 VPWR VGND sg13g2_decap_8
XFILLER_77_917 VPWR VGND sg13g2_decap_8
XFILLER_0_147 VPWR VGND sg13g2_decap_8
XFILLER_88_298 VPWR VGND sg13g2_decap_8
XFILLER_76_438 VPWR VGND sg13g2_decap_8
XFILLER_57_630 VPWR VGND sg13g2_decap_8
XFILLER_28_21 VPWR VGND sg13g2_decap_8
XFILLER_29_354 VPWR VGND sg13g2_decap_8
XFILLER_85_994 VPWR VGND sg13g2_decap_8
XFILLER_56_151 VPWR VGND sg13g2_decap_8
XFILLER_45_847 VPWR VGND sg13g2_decap_8
XFILLER_28_98 VPWR VGND sg13g2_decap_8
XFILLER_72_644 VPWR VGND sg13g2_decap_8
XFILLER_71_165 VPWR VGND sg13g2_decap_8
XFILLER_44_368 VPWR VGND sg13g2_decap_8
XFILLER_44_53 VPWR VGND sg13g2_decap_8
XFILLER_13_700 VPWR VGND sg13g2_decap_8
XFILLER_25_560 VPWR VGND sg13g2_decap_8
XFILLER_32_508 VPWR VGND sg13g2_decap_8
XFILLER_12_221 VPWR VGND sg13g2_decap_8
XFILLER_8_203 VPWR VGND sg13g2_decap_8
XFILLER_13_777 VPWR VGND sg13g2_decap_8
XFILLER_100_70 VPWR VGND sg13g2_decap_8
XFILLER_40_574 VPWR VGND sg13g2_decap_8
XFILLER_60_74 VPWR VGND sg13g2_decap_8
XFILLER_12_298 VPWR VGND sg13g2_decap_8
XFILLER_5_921 VPWR VGND sg13g2_decap_8
XFILLER_5_25 VPWR VGND sg13g2_decap_8
XFILLER_4_420 VPWR VGND sg13g2_decap_8
XFILLER_5_998 VPWR VGND sg13g2_decap_8
XFILLER_106_392 VPWR VGND sg13g2_decap_8
XFILLER_79_221 VPWR VGND sg13g2_decap_8
XFILLER_4_497 VPWR VGND sg13g2_decap_8
XFILLER_95_725 VPWR VGND sg13g2_decap_8
XFILLER_94_224 VPWR VGND sg13g2_decap_8
XFILLER_79_298 VPWR VGND sg13g2_decap_8
XFILLER_67_427 VPWR VGND sg13g2_decap_8
XFILLER_48_630 VPWR VGND sg13g2_decap_8
XFILLER_47_140 VPWR VGND sg13g2_decap_8
XFILLER_91_931 VPWR VGND sg13g2_decap_8
XFILLER_63_644 VPWR VGND sg13g2_decap_8
XFILLER_36_847 VPWR VGND sg13g2_decap_8
XFILLER_39_1019 VPWR VGND sg13g2_decap_8
XFILLER_90_452 VPWR VGND sg13g2_decap_8
XFILLER_62_154 VPWR VGND sg13g2_decap_8
XFILLER_16_560 VPWR VGND sg13g2_decap_8
XFILLER_35_357 VPWR VGND sg13g2_decap_8
XFILLER_31_574 VPWR VGND sg13g2_decap_8
XFILLER_102_1022 VPWR VGND sg13g2_decap_8
XFILLER_8_770 VPWR VGND sg13g2_decap_8
XFILLER_105_819 VPWR VGND sg13g2_decap_8
XFILLER_7_291 VPWR VGND sg13g2_decap_8
XFILLER_104_329 VPWR VGND sg13g2_decap_8
XFILLER_86_725 VPWR VGND sg13g2_decap_8
XFILLER_98_585 VPWR VGND sg13g2_decap_8
XFILLER_85_224 VPWR VGND sg13g2_decap_8
XFILLER_58_427 VPWR VGND sg13g2_decap_8
XFILLER_100_546 VPWR VGND sg13g2_decap_8
XFILLER_22_1012 VPWR VGND sg13g2_decap_8
XFILLER_39_641 VPWR VGND sg13g2_decap_8
XFILLER_94_791 VPWR VGND sg13g2_decap_8
XFILLER_82_931 VPWR VGND sg13g2_decap_8
XFILLER_67_994 VPWR VGND sg13g2_decap_8
XFILLER_66_482 VPWR VGND sg13g2_decap_8
XFILLER_38_140 VPWR VGND sg13g2_decap_8
XFILLER_54_655 VPWR VGND sg13g2_decap_8
XFILLER_27_858 VPWR VGND sg13g2_decap_8
XFILLER_81_452 VPWR VGND sg13g2_decap_8
XFILLER_81_18 VPWR VGND sg13g2_decap_8
XFILLER_53_154 VPWR VGND sg13g2_decap_8
XFILLER_26_357 VPWR VGND sg13g2_decap_8
XFILLER_50_861 VPWR VGND sg13g2_decap_8
XFILLER_10_725 VPWR VGND sg13g2_decap_8
XFILLER_14_56 VPWR VGND sg13g2_decap_8
XFILLER_22_585 VPWR VGND sg13g2_decap_8
XFILLER_6_707 VPWR VGND sg13g2_decap_8
XFILLER_5_228 VPWR VGND sg13g2_decap_8
XFILLER_30_77 VPWR VGND sg13g2_decap_8
XFILLER_2_935 VPWR VGND sg13g2_decap_8
XFILLER_1_434 VPWR VGND sg13g2_decap_8
XFILLER_89_574 VPWR VGND sg13g2_decap_8
XFILLER_77_714 VPWR VGND sg13g2_decap_8
XFILLER_104_896 VPWR VGND sg13g2_decap_8
XFILLER_49_438 VPWR VGND sg13g2_decap_8
XFILLER_7_1028 VPWR VGND sg13g2_fill_1
XFILLER_39_53 VPWR VGND sg13g2_decap_8
XFILLER_76_235 VPWR VGND sg13g2_decap_8
XFILLER_92_728 VPWR VGND sg13g2_decap_8
XFILLER_58_994 VPWR VGND sg13g2_decap_8
XFILLER_29_151 VPWR VGND sg13g2_decap_8
XFILLER_91_238 VPWR VGND sg13g2_decap_8
XFILLER_85_791 VPWR VGND sg13g2_decap_8
XFILLER_73_942 VPWR VGND sg13g2_decap_8
XFILLER_45_644 VPWR VGND sg13g2_decap_8
XFILLER_18_847 VPWR VGND sg13g2_decap_8
XFILLER_72_441 VPWR VGND sg13g2_decap_8
XFILLER_55_63 VPWR VGND sg13g2_decap_8
XFILLER_44_165 VPWR VGND sg13g2_decap_8
XFILLER_17_368 VPWR VGND sg13g2_decap_8
XFILLER_32_305 VPWR VGND sg13g2_decap_8
XFILLER_60_669 VPWR VGND sg13g2_decap_8
XFILLER_41_861 VPWR VGND sg13g2_decap_8
XFILLER_13_574 VPWR VGND sg13g2_decap_8
XFILLER_40_371 VPWR VGND sg13g2_decap_8
XFILLER_71_95 VPWR VGND sg13g2_decap_8
XFILLER_9_567 VPWR VGND sg13g2_decap_8
XFILLER_65_7 VPWR VGND sg13g2_decap_8
XFILLER_45_1001 VPWR VGND sg13g2_decap_8
XFILLER_5_795 VPWR VGND sg13g2_decap_8
XFILLER_4_294 VPWR VGND sg13g2_decap_8
XFILLER_96_70 VPWR VGND sg13g2_decap_8
XFILLER_95_522 VPWR VGND sg13g2_decap_8
XFILLER_68_747 VPWR VGND sg13g2_decap_8
XFILLER_67_224 VPWR VGND sg13g2_decap_8
XFILLER_95_599 VPWR VGND sg13g2_decap_8
XFILLER_83_739 VPWR VGND sg13g2_decap_8
XFILLER_82_238 VPWR VGND sg13g2_decap_8
XFILLER_64_942 VPWR VGND sg13g2_decap_8
XFILLER_36_644 VPWR VGND sg13g2_decap_8
XFILLER_63_441 VPWR VGND sg13g2_decap_8
XFILLER_35_154 VPWR VGND sg13g2_decap_8
XFILLER_91_0 VPWR VGND sg13g2_decap_8
XFILLER_51_669 VPWR VGND sg13g2_decap_8
XFILLER_50_168 VPWR VGND sg13g2_decap_8
XFILLER_31_371 VPWR VGND sg13g2_decap_8
XFILLER_32_872 VPWR VGND sg13g2_decap_8
XFILLER_105_616 VPWR VGND sg13g2_decap_8
XFILLER_104_126 VPWR VGND sg13g2_decap_8
XFILLER_99_861 VPWR VGND sg13g2_decap_8
XFILLER_101_833 VPWR VGND sg13g2_decap_8
XFILLER_98_382 VPWR VGND sg13g2_decap_8
XFILLER_86_522 VPWR VGND sg13g2_decap_8
XFILLER_76_18 VPWR VGND sg13g2_decap_8
XFILLER_59_747 VPWR VGND sg13g2_decap_8
XFILLER_58_224 VPWR VGND sg13g2_decap_8
XFILLER_100_343 VPWR VGND sg13g2_decap_8
XFILLER_86_599 VPWR VGND sg13g2_decap_8
XFILLER_73_249 VPWR VGND sg13g2_decap_8
XFILLER_67_791 VPWR VGND sg13g2_decap_8
XFILLER_55_931 VPWR VGND sg13g2_decap_8
XFILLER_92_28 VPWR VGND sg13g2_decap_8
XFILLER_54_452 VPWR VGND sg13g2_decap_8
XFILLER_26_154 VPWR VGND sg13g2_decap_8
XFILLER_27_655 VPWR VGND sg13g2_decap_8
XFILLER_70_945 VPWR VGND sg13g2_decap_8
XFILLER_42_669 VPWR VGND sg13g2_decap_8
XFILLER_23_861 VPWR VGND sg13g2_decap_8
XFILLER_25_77 VPWR VGND sg13g2_decap_8
XFILLER_41_168 VPWR VGND sg13g2_decap_8
XFILLER_10_522 VPWR VGND sg13g2_decap_8
XFILLER_22_382 VPWR VGND sg13g2_decap_8
XFILLER_41_21 VPWR VGND sg13g2_decap_8
XFILLER_6_504 VPWR VGND sg13g2_decap_8
XFILLER_10_599 VPWR VGND sg13g2_decap_8
XFILLER_41_98 VPWR VGND sg13g2_decap_8
XFILLER_2_732 VPWR VGND sg13g2_decap_8
XFILLER_96_308 VPWR VGND sg13g2_decap_8
XFILLER_1_231 VPWR VGND sg13g2_decap_8
XFILLER_104_693 VPWR VGND sg13g2_decap_8
XFILLER_89_371 VPWR VGND sg13g2_decap_8
XFILLER_77_511 VPWR VGND sg13g2_decap_8
XFILLER_49_235 VPWR VGND sg13g2_decap_8
XFILLER_106_91 VPWR VGND sg13g2_decap_8
XFILLER_92_525 VPWR VGND sg13g2_decap_8
XFILLER_77_588 VPWR VGND sg13g2_decap_8
XFILLER_66_62 VPWR VGND sg13g2_decap_8
XFILLER_65_728 VPWR VGND sg13g2_decap_8
XFILLER_64_249 VPWR VGND sg13g2_decap_8
XFILLER_58_791 VPWR VGND sg13g2_decap_8
XFILLER_46_942 VPWR VGND sg13g2_decap_8
XFILLER_18_644 VPWR VGND sg13g2_decap_8
XFILLER_45_441 VPWR VGND sg13g2_decap_8
XFILLER_17_165 VPWR VGND sg13g2_decap_8
XFILLER_32_102 VPWR VGND sg13g2_decap_8
XFILLER_61_956 VPWR VGND sg13g2_decap_8
XFILLER_33_658 VPWR VGND sg13g2_decap_8
XFILLER_60_466 VPWR VGND sg13g2_decap_8
XFILLER_14_861 VPWR VGND sg13g2_decap_8
XFILLER_20_319 VPWR VGND sg13g2_decap_8
XFILLER_32_179 VPWR VGND sg13g2_decap_8
XFILLER_13_371 VPWR VGND sg13g2_decap_8
XFILLER_9_364 VPWR VGND sg13g2_decap_8
XFILLER_5_592 VPWR VGND sg13g2_decap_8
XFILLER_99_168 VPWR VGND sg13g2_decap_8
XFILLER_88_809 VPWR VGND sg13g2_decap_8
XFILLER_87_308 VPWR VGND sg13g2_decap_8
XFILLER_96_875 VPWR VGND sg13g2_decap_8
XFILLER_68_544 VPWR VGND sg13g2_decap_8
XFILLER_56_739 VPWR VGND sg13g2_decap_8
XFILLER_95_396 VPWR VGND sg13g2_decap_8
XFILLER_83_536 VPWR VGND sg13g2_decap_8
XFILLER_55_238 VPWR VGND sg13g2_decap_8
XFILLER_37_942 VPWR VGND sg13g2_decap_8
XFILLER_36_441 VPWR VGND sg13g2_decap_8
XFILLER_102_49 VPWR VGND sg13g2_decap_8
XFILLER_52_945 VPWR VGND sg13g2_decap_8
XFILLER_12_809 VPWR VGND sg13g2_decap_8
XFILLER_24_669 VPWR VGND sg13g2_decap_8
XFILLER_51_466 VPWR VGND sg13g2_decap_8
XFILLER_11_308 VPWR VGND sg13g2_decap_8
XFILLER_23_168 VPWR VGND sg13g2_decap_8
XFILLER_20_886 VPWR VGND sg13g2_decap_8
XFILLER_106_903 VPWR VGND sg13g2_decap_8
XFILLER_3_518 VPWR VGND sg13g2_decap_8
XFILLER_11_35 VPWR VGND sg13g2_decap_8
XFILLER_105_413 VPWR VGND sg13g2_decap_8
XFILLER_87_28 VPWR VGND sg13g2_decap_8
XFILLER_79_809 VPWR VGND sg13g2_decap_8
XFILLER_101_630 VPWR VGND sg13g2_decap_8
XFILLER_59_544 VPWR VGND sg13g2_decap_8
XFILLER_100_140 VPWR VGND sg13g2_decap_8
XFILLER_98_1005 VPWR VGND sg13g2_decap_8
XFILLER_87_875 VPWR VGND sg13g2_decap_8
XFILLER_47_728 VPWR VGND sg13g2_decap_8
XFILLER_86_396 VPWR VGND sg13g2_decap_8
XFILLER_74_547 VPWR VGND sg13g2_decap_8
XFILLER_46_249 VPWR VGND sg13g2_decap_8
XFILLER_28_931 VPWR VGND sg13g2_decap_8
XFILLER_36_21 VPWR VGND sg13g2_decap_8
XFILLER_27_452 VPWR VGND sg13g2_decap_8
XFILLER_43_945 VPWR VGND sg13g2_decap_8
XFILLER_70_742 VPWR VGND sg13g2_decap_8
XFILLER_15_669 VPWR VGND sg13g2_decap_8
XFILLER_36_98 VPWR VGND sg13g2_decap_8
XFILLER_52_42 VPWR VGND sg13g2_decap_8
XFILLER_42_466 VPWR VGND sg13g2_decap_8
XFILLER_14_168 VPWR VGND sg13g2_decap_8
XFILLER_35_1022 VPWR VGND sg13g2_decap_8
XFILLER_7_802 VPWR VGND sg13g2_decap_8
XFILLER_6_301 VPWR VGND sg13g2_decap_8
XFILLER_11_875 VPWR VGND sg13g2_decap_8
XFILLER_10_396 VPWR VGND sg13g2_decap_8
XFILLER_7_879 VPWR VGND sg13g2_decap_8
XFILLER_6_378 VPWR VGND sg13g2_decap_8
XFILLER_105_980 VPWR VGND sg13g2_decap_8
XFILLER_96_105 VPWR VGND sg13g2_decap_8
XFILLER_104_490 VPWR VGND sg13g2_decap_8
XFILLER_78_853 VPWR VGND sg13g2_decap_8
XFILLER_42_1026 VPWR VGND sg13g2_fill_2
XFILLER_28_7 VPWR VGND sg13g2_decap_8
X_32_ _02_ _00_ net18 VPWR VGND sg13g2_xor2_1
XFILLER_38_728 VPWR VGND sg13g2_decap_8
XFILLER_93_845 VPWR VGND sg13g2_decap_8
XFILLER_92_322 VPWR VGND sg13g2_decap_8
XFILLER_77_385 VPWR VGND sg13g2_decap_8
XFILLER_65_525 VPWR VGND sg13g2_decap_8
XFILLER_19_931 VPWR VGND sg13g2_decap_8
XFILLER_18_441 VPWR VGND sg13g2_decap_8
XFILLER_37_249 VPWR VGND sg13g2_decap_8
XFILLER_93_82 VPWR VGND sg13g2_decap_8
XFILLER_92_399 VPWR VGND sg13g2_decap_8
XFILLER_80_539 VPWR VGND sg13g2_decap_8
Xheichips25_example_large_25 VPWR VGND uio_oe[0] sg13g2_tielo
XFILLER_61_753 VPWR VGND sg13g2_decap_8
Xheichips25_example_large_36 VPWR VGND uio_out[3] sg13g2_tielo
XFILLER_33_455 VPWR VGND sg13g2_decap_8
XFILLER_34_956 VPWR VGND sg13g2_decap_8
XFILLER_60_263 VPWR VGND sg13g2_decap_8
XFILLER_20_116 VPWR VGND sg13g2_decap_8
XFILLER_9_161 VPWR VGND sg13g2_decap_8
XFILLER_103_917 VPWR VGND sg13g2_decap_8
XFILLER_88_606 VPWR VGND sg13g2_decap_8
XFILLER_102_427 VPWR VGND sg13g2_decap_8
XFILLER_87_105 VPWR VGND sg13g2_decap_8
XFILLER_69_820 VPWR VGND sg13g2_decap_8
XFILLER_96_672 VPWR VGND sg13g2_decap_8
XFILLER_84_812 VPWR VGND sg13g2_decap_8
XFILLER_69_897 VPWR VGND sg13g2_decap_8
XFILLER_68_341 VPWR VGND sg13g2_decap_8
XFILLER_3_91 VPWR VGND sg13g2_decap_8
XFILLER_95_193 VPWR VGND sg13g2_decap_8
XFILLER_83_333 VPWR VGND sg13g2_decap_8
XFILLER_56_536 VPWR VGND sg13g2_decap_8
XFILLER_28_238 VPWR VGND sg13g2_decap_8
XFILLER_29_739 VPWR VGND sg13g2_decap_8
XFILLER_84_889 VPWR VGND sg13g2_decap_8
XFILLER_58_1022 VPWR VGND sg13g2_decap_8
XFILLER_52_742 VPWR VGND sg13g2_decap_8
XFILLER_25_945 VPWR VGND sg13g2_decap_8
XFILLER_51_263 VPWR VGND sg13g2_decap_8
XFILLER_11_105 VPWR VGND sg13g2_decap_8
XFILLER_12_606 VPWR VGND sg13g2_decap_8
XFILLER_24_466 VPWR VGND sg13g2_decap_8
XFILLER_40_959 VPWR VGND sg13g2_decap_8
XFILLER_7_109 VPWR VGND sg13g2_decap_8
XFILLER_20_683 VPWR VGND sg13g2_decap_8
XFILLER_22_67 VPWR VGND sg13g2_decap_8
XFILLER_106_700 VPWR VGND sg13g2_decap_8
XFILLER_4_805 VPWR VGND sg13g2_decap_8
XFILLER_105_210 VPWR VGND sg13g2_decap_8
XFILLER_3_315 VPWR VGND sg13g2_decap_8
XFILLER_106_777 VPWR VGND sg13g2_decap_8
XFILLER_79_606 VPWR VGND sg13g2_decap_8
XFILLER_65_1015 VPWR VGND sg13g2_decap_8
XFILLER_105_287 VPWR VGND sg13g2_decap_8
XFILLER_94_609 VPWR VGND sg13g2_decap_8
XFILLER_87_672 VPWR VGND sg13g2_decap_8
XFILLER_75_812 VPWR VGND sg13g2_decap_8
XFILLER_59_341 VPWR VGND sg13g2_decap_8
XFILLER_102_994 VPWR VGND sg13g2_decap_8
XFILLER_47_525 VPWR VGND sg13g2_decap_8
XFILLER_47_42 VPWR VGND sg13g2_decap_8
XFILLER_19_238 VPWR VGND sg13g2_decap_8
XFILLER_86_193 VPWR VGND sg13g2_decap_8
XFILLER_75_889 VPWR VGND sg13g2_decap_8
XFILLER_74_344 VPWR VGND sg13g2_decap_8
XFILLER_90_837 VPWR VGND sg13g2_decap_8
XFILLER_62_539 VPWR VGND sg13g2_decap_8
XFILLER_103_70 VPWR VGND sg13g2_decap_8
XFILLER_43_742 VPWR VGND sg13g2_decap_8
XFILLER_16_945 VPWR VGND sg13g2_decap_8
XFILLER_72_1008 VPWR VGND sg13g2_decap_8
XFILLER_63_63 VPWR VGND sg13g2_decap_8
XFILLER_42_263 VPWR VGND sg13g2_decap_8
XFILLER_15_466 VPWR VGND sg13g2_decap_8
XFILLER_8_14 VPWR VGND sg13g2_decap_8
XFILLER_31_959 VPWR VGND sg13g2_decap_8
XFILLER_30_469 VPWR VGND sg13g2_decap_8
XFILLER_11_672 VPWR VGND sg13g2_decap_8
XFILLER_10_193 VPWR VGND sg13g2_decap_8
XFILLER_7_676 VPWR VGND sg13g2_decap_8
XFILLER_6_175 VPWR VGND sg13g2_decap_8
XFILLER_88_60 VPWR VGND sg13g2_decap_8
XFILLER_3_882 VPWR VGND sg13g2_decap_8
XFILLER_85_609 VPWR VGND sg13g2_decap_8
XFILLER_69_127 VPWR VGND sg13g2_decap_8
XFILLER_97_469 VPWR VGND sg13g2_decap_8
XFILLER_84_119 VPWR VGND sg13g2_decap_8
XFILLER_78_650 VPWR VGND sg13g2_decap_8
XFILLER_77_182 VPWR VGND sg13g2_decap_8
XFILLER_65_322 VPWR VGND sg13g2_decap_8
XFILLER_38_525 VPWR VGND sg13g2_decap_8
XFILLER_93_642 VPWR VGND sg13g2_decap_8
XFILLER_66_867 VPWR VGND sg13g2_decap_8
XFILLER_81_837 VPWR VGND sg13g2_decap_8
XFILLER_65_399 VPWR VGND sg13g2_decap_8
XFILLER_53_539 VPWR VGND sg13g2_decap_8
XFILLER_92_196 VPWR VGND sg13g2_decap_8
XFILLER_80_336 VPWR VGND sg13g2_decap_8
XFILLER_34_753 VPWR VGND sg13g2_decap_8
XFILLER_61_550 VPWR VGND sg13g2_decap_8
XFILLER_33_252 VPWR VGND sg13g2_decap_8
XFILLER_21_469 VPWR VGND sg13g2_decap_8
XFILLER_88_1026 VPWR VGND sg13g2_fill_2
XFILLER_103_714 VPWR VGND sg13g2_decap_8
XFILLER_88_403 VPWR VGND sg13g2_decap_8
XFILLER_1_819 VPWR VGND sg13g2_decap_8
XFILLER_102_224 VPWR VGND sg13g2_decap_8
XFILLER_89_959 VPWR VGND sg13g2_decap_8
XFILLER_0_329 VPWR VGND sg13g2_decap_8
XFILLER_57_812 VPWR VGND sg13g2_decap_8
XFILLER_75_119 VPWR VGND sg13g2_decap_8
XFILLER_69_694 VPWR VGND sg13g2_decap_8
XFILLER_29_536 VPWR VGND sg13g2_decap_8
XFILLER_83_130 VPWR VGND sg13g2_decap_8
XFILLER_57_889 VPWR VGND sg13g2_decap_8
XFILLER_56_333 VPWR VGND sg13g2_decap_8
XFILLER_95_1019 VPWR VGND sg13g2_decap_8
XFILLER_84_686 VPWR VGND sg13g2_decap_8
XFILLER_72_826 VPWR VGND sg13g2_decap_8
XFILLER_71_347 VPWR VGND sg13g2_decap_8
XFILLER_17_67 VPWR VGND sg13g2_decap_8
XFILLER_25_742 VPWR VGND sg13g2_decap_8
XFILLER_12_403 VPWR VGND sg13g2_decap_8
XFILLER_24_263 VPWR VGND sg13g2_decap_8
XFILLER_13_959 VPWR VGND sg13g2_decap_8
XFILLER_33_77 VPWR VGND sg13g2_decap_8
XFILLER_40_756 VPWR VGND sg13g2_decap_8
XFILLER_20_480 VPWR VGND sg13g2_decap_8
XFILLER_4_602 VPWR VGND sg13g2_decap_8
XFILLER_3_112 VPWR VGND sg13g2_decap_8
XFILLER_106_574 VPWR VGND sg13g2_decap_8
XFILLER_79_403 VPWR VGND sg13g2_decap_8
XFILLER_4_679 VPWR VGND sg13g2_decap_8
XFILLER_95_907 VPWR VGND sg13g2_decap_8
XFILLER_3_189 VPWR VGND sg13g2_decap_8
XFILLER_94_406 VPWR VGND sg13g2_decap_8
XFILLER_88_970 VPWR VGND sg13g2_decap_8
XFILLER_67_609 VPWR VGND sg13g2_decap_8
XFILLER_58_63 VPWR VGND sg13g2_decap_8
XFILLER_48_812 VPWR VGND sg13g2_decap_8
XFILLER_102_791 VPWR VGND sg13g2_decap_8
XFILLER_47_322 VPWR VGND sg13g2_decap_8
XFILLER_0_896 VPWR VGND sg13g2_decap_8
XFILLER_74_141 VPWR VGND sg13g2_decap_8
XFILLER_75_686 VPWR VGND sg13g2_decap_8
XFILLER_63_826 VPWR VGND sg13g2_decap_8
XFILLER_48_889 VPWR VGND sg13g2_decap_8
XFILLER_35_539 VPWR VGND sg13g2_decap_8
XFILLER_90_634 VPWR VGND sg13g2_decap_8
XFILLER_62_336 VPWR VGND sg13g2_decap_8
XFILLER_47_399 VPWR VGND sg13g2_decap_8
XFILLER_16_742 VPWR VGND sg13g2_decap_8
XFILLER_15_263 VPWR VGND sg13g2_decap_8
XFILLER_31_756 VPWR VGND sg13g2_decap_8
XFILLER_12_970 VPWR VGND sg13g2_decap_8
XFILLER_30_266 VPWR VGND sg13g2_decap_8
XFILLER_8_952 VPWR VGND sg13g2_decap_8
XFILLER_7_473 VPWR VGND sg13g2_decap_8
XFILLER_99_70 VPWR VGND sg13g2_decap_8
XFILLER_98_767 VPWR VGND sg13g2_decap_8
XFILLER_86_907 VPWR VGND sg13g2_decap_8
XFILLER_97_266 VPWR VGND sg13g2_decap_8
XFILLER_85_406 VPWR VGND sg13g2_decap_8
XFILLER_79_970 VPWR VGND sg13g2_decap_8
XFILLER_58_609 VPWR VGND sg13g2_decap_8
XFILLER_100_728 VPWR VGND sg13g2_decap_8
XFILLER_57_119 VPWR VGND sg13g2_decap_8
XFILLER_38_322 VPWR VGND sg13g2_decap_8
XFILLER_39_823 VPWR VGND sg13g2_decap_8
XFILLER_94_973 VPWR VGND sg13g2_decap_8
XFILLER_66_664 VPWR VGND sg13g2_decap_8
XFILLER_54_837 VPWR VGND sg13g2_decap_8
XFILLER_0_1001 VPWR VGND sg13g2_decap_8
XFILLER_81_634 VPWR VGND sg13g2_decap_8
XFILLER_80_133 VPWR VGND sg13g2_decap_8
XFILLER_65_196 VPWR VGND sg13g2_decap_8
XFILLER_53_336 VPWR VGND sg13g2_decap_8
XFILLER_0_70 VPWR VGND sg13g2_decap_8
XFILLER_26_539 VPWR VGND sg13g2_decap_8
XFILLER_38_399 VPWR VGND sg13g2_decap_8
XFILLER_34_550 VPWR VGND sg13g2_decap_8
XFILLER_10_907 VPWR VGND sg13g2_decap_8
XFILLER_22_767 VPWR VGND sg13g2_decap_8
XFILLER_21_266 VPWR VGND sg13g2_decap_8
XFILLER_88_200 VPWR VGND sg13g2_decap_8
XFILLER_1_616 VPWR VGND sg13g2_decap_8
XFILLER_103_511 VPWR VGND sg13g2_decap_8
XFILLER_89_756 VPWR VGND sg13g2_decap_8
XFILLER_0_126 VPWR VGND sg13g2_decap_8
XFILLER_95_39 VPWR VGND sg13g2_decap_8
XFILLER_76_417 VPWR VGND sg13g2_decap_8
XFILLER_103_588 VPWR VGND sg13g2_decap_8
XFILLER_88_277 VPWR VGND sg13g2_decap_8
XFILLER_48_119 VPWR VGND sg13g2_decap_8
XFILLER_85_973 VPWR VGND sg13g2_decap_8
XFILLER_69_491 VPWR VGND sg13g2_decap_8
XFILLER_56_130 VPWR VGND sg13g2_decap_8
XFILLER_29_333 VPWR VGND sg13g2_decap_8
XFILLER_84_483 VPWR VGND sg13g2_decap_8
XFILLER_72_623 VPWR VGND sg13g2_decap_8
XFILLER_57_686 VPWR VGND sg13g2_decap_8
XFILLER_45_826 VPWR VGND sg13g2_decap_8
XFILLER_28_77 VPWR VGND sg13g2_decap_8
XFILLER_44_347 VPWR VGND sg13g2_decap_8
XFILLER_71_144 VPWR VGND sg13g2_decap_8
XFILLER_44_32 VPWR VGND sg13g2_decap_8
XFILLER_12_200 VPWR VGND sg13g2_decap_8
XFILLER_13_756 VPWR VGND sg13g2_decap_8
XFILLER_40_553 VPWR VGND sg13g2_decap_8
XFILLER_9_749 VPWR VGND sg13g2_decap_8
XFILLER_12_277 VPWR VGND sg13g2_decap_8
XFILLER_60_53 VPWR VGND sg13g2_decap_8
XFILLER_8_259 VPWR VGND sg13g2_decap_8
XFILLER_5_900 VPWR VGND sg13g2_decap_8
XFILLER_79_200 VPWR VGND sg13g2_decap_8
XFILLER_5_977 VPWR VGND sg13g2_decap_8
XFILLER_4_476 VPWR VGND sg13g2_decap_8
XFILLER_106_371 VPWR VGND sg13g2_decap_8
XFILLER_95_704 VPWR VGND sg13g2_decap_8
XFILLER_68_929 VPWR VGND sg13g2_decap_8
XFILLER_67_406 VPWR VGND sg13g2_decap_8
XFILLER_94_203 VPWR VGND sg13g2_decap_8
XFILLER_79_277 VPWR VGND sg13g2_decap_8
XFILLER_0_693 VPWR VGND sg13g2_decap_8
XFILLER_91_910 VPWR VGND sg13g2_decap_8
XFILLER_78_1014 VPWR VGND sg13g2_decap_8
XFILLER_76_984 VPWR VGND sg13g2_decap_8
XFILLER_63_623 VPWR VGND sg13g2_decap_8
XFILLER_48_686 VPWR VGND sg13g2_decap_8
XFILLER_36_826 VPWR VGND sg13g2_decap_8
XFILLER_90_431 VPWR VGND sg13g2_decap_8
XFILLER_75_483 VPWR VGND sg13g2_decap_8
XFILLER_62_133 VPWR VGND sg13g2_decap_8
XFILLER_47_196 VPWR VGND sg13g2_decap_8
XFILLER_35_336 VPWR VGND sg13g2_decap_8
XFILLER_91_987 VPWR VGND sg13g2_decap_8
XFILLER_31_553 VPWR VGND sg13g2_decap_8
XFILLER_102_1001 VPWR VGND sg13g2_decap_8
XFILLER_7_270 VPWR VGND sg13g2_decap_8
XFILLER_104_308 VPWR VGND sg13g2_decap_8
XFILLER_98_564 VPWR VGND sg13g2_decap_8
XFILLER_86_704 VPWR VGND sg13g2_decap_8
XFILLER_59_929 VPWR VGND sg13g2_decap_8
XFILLER_58_406 VPWR VGND sg13g2_decap_8
XFILLER_100_525 VPWR VGND sg13g2_decap_8
XFILLER_85_203 VPWR VGND sg13g2_decap_8
XFILLER_39_620 VPWR VGND sg13g2_decap_8
XFILLER_105_49 VPWR VGND sg13g2_decap_8
XFILLER_94_770 VPWR VGND sg13g2_decap_8
XFILLER_82_910 VPWR VGND sg13g2_decap_8
XFILLER_67_973 VPWR VGND sg13g2_decap_8
XFILLER_66_461 VPWR VGND sg13g2_decap_8
XFILLER_27_837 VPWR VGND sg13g2_decap_8
XFILLER_81_431 VPWR VGND sg13g2_decap_8
XFILLER_54_634 VPWR VGND sg13g2_decap_8
XFILLER_26_336 VPWR VGND sg13g2_decap_8
XFILLER_38_196 VPWR VGND sg13g2_decap_8
XFILLER_39_697 VPWR VGND sg13g2_decap_8
XFILLER_82_987 VPWR VGND sg13g2_decap_8
XFILLER_53_133 VPWR VGND sg13g2_decap_8
XFILLER_50_840 VPWR VGND sg13g2_decap_8
XFILLER_14_35 VPWR VGND sg13g2_decap_8
XFILLER_10_704 VPWR VGND sg13g2_decap_8
XFILLER_22_564 VPWR VGND sg13g2_decap_8
XFILLER_5_207 VPWR VGND sg13g2_decap_8
XFILLER_30_56 VPWR VGND sg13g2_decap_8
XFILLER_2_914 VPWR VGND sg13g2_decap_8
XFILLER_1_413 VPWR VGND sg13g2_decap_8
XFILLER_104_875 VPWR VGND sg13g2_decap_8
XFILLER_89_553 VPWR VGND sg13g2_decap_8
XFILLER_39_32 VPWR VGND sg13g2_decap_8
XFILLER_103_385 VPWR VGND sg13g2_decap_8
XFILLER_76_214 VPWR VGND sg13g2_decap_8
XFILLER_49_417 VPWR VGND sg13g2_decap_8
XFILLER_92_707 VPWR VGND sg13g2_decap_8
XFILLER_29_130 VPWR VGND sg13g2_decap_8
XFILLER_91_217 VPWR VGND sg13g2_decap_8
XFILLER_85_770 VPWR VGND sg13g2_decap_8
XFILLER_73_921 VPWR VGND sg13g2_decap_8
XFILLER_58_973 VPWR VGND sg13g2_decap_8
XFILLER_18_826 VPWR VGND sg13g2_decap_8
XFILLER_84_280 VPWR VGND sg13g2_decap_8
XFILLER_72_420 VPWR VGND sg13g2_decap_8
XFILLER_57_483 VPWR VGND sg13g2_decap_8
XFILLER_55_42 VPWR VGND sg13g2_decap_8
XFILLER_45_623 VPWR VGND sg13g2_decap_8
XFILLER_73_998 VPWR VGND sg13g2_decap_8
XFILLER_44_144 VPWR VGND sg13g2_decap_8
XFILLER_17_347 VPWR VGND sg13g2_decap_8
XFILLER_72_497 VPWR VGND sg13g2_decap_8
XFILLER_60_648 VPWR VGND sg13g2_decap_8
XFILLER_41_840 VPWR VGND sg13g2_decap_8
XFILLER_13_553 VPWR VGND sg13g2_decap_8
XFILLER_71_74 VPWR VGND sg13g2_decap_8
XFILLER_40_350 VPWR VGND sg13g2_decap_8
XFILLER_9_546 VPWR VGND sg13g2_decap_8
XFILLER_58_7 VPWR VGND sg13g2_decap_8
XFILLER_5_774 VPWR VGND sg13g2_decap_8
XFILLER_4_273 VPWR VGND sg13g2_decap_8
XFILLER_95_501 VPWR VGND sg13g2_decap_8
XFILLER_68_726 VPWR VGND sg13g2_decap_8
XFILLER_67_203 VPWR VGND sg13g2_decap_8
XFILLER_1_980 VPWR VGND sg13g2_decap_8
XFILLER_0_490 VPWR VGND sg13g2_decap_8
XFILLER_95_578 VPWR VGND sg13g2_decap_8
XFILLER_83_718 VPWR VGND sg13g2_decap_8
XFILLER_82_217 VPWR VGND sg13g2_decap_8
XFILLER_76_781 VPWR VGND sg13g2_decap_8
XFILLER_64_921 VPWR VGND sg13g2_decap_8
XFILLER_49_984 VPWR VGND sg13g2_decap_8
XFILLER_75_280 VPWR VGND sg13g2_decap_8
XFILLER_63_420 VPWR VGND sg13g2_decap_8
XFILLER_48_483 VPWR VGND sg13g2_decap_8
XFILLER_36_623 VPWR VGND sg13g2_decap_8
XFILLER_35_133 VPWR VGND sg13g2_decap_8
XFILLER_91_784 VPWR VGND sg13g2_decap_8
XFILLER_64_998 VPWR VGND sg13g2_decap_8
XFILLER_63_497 VPWR VGND sg13g2_decap_8
XFILLER_91_1022 VPWR VGND sg13g2_decap_8
XFILLER_51_648 VPWR VGND sg13g2_decap_8
XFILLER_50_147 VPWR VGND sg13g2_decap_8
XFILLER_32_851 VPWR VGND sg13g2_decap_8
XFILLER_31_350 VPWR VGND sg13g2_decap_8
XFILLER_84_0 VPWR VGND sg13g2_decap_8
XFILLER_104_105 VPWR VGND sg13g2_decap_8
XFILLER_99_840 VPWR VGND sg13g2_decap_8
XFILLER_6_91 VPWR VGND sg13g2_decap_8
XFILLER_101_812 VPWR VGND sg13g2_decap_8
XFILLER_98_361 VPWR VGND sg13g2_decap_8
XFILLER_86_501 VPWR VGND sg13g2_decap_8
XFILLER_59_726 VPWR VGND sg13g2_decap_8
XFILLER_58_203 VPWR VGND sg13g2_decap_8
XFILLER_100_322 VPWR VGND sg13g2_decap_8
XFILLER_101_889 VPWR VGND sg13g2_decap_8
XFILLER_86_578 VPWR VGND sg13g2_decap_8
XFILLER_74_729 VPWR VGND sg13g2_decap_8
XFILLER_67_770 VPWR VGND sg13g2_decap_8
XFILLER_55_910 VPWR VGND sg13g2_decap_8
XFILLER_100_399 VPWR VGND sg13g2_decap_8
XFILLER_73_228 VPWR VGND sg13g2_decap_8
XFILLER_27_634 VPWR VGND sg13g2_decap_8
XFILLER_39_494 VPWR VGND sg13g2_decap_8
XFILLER_55_987 VPWR VGND sg13g2_decap_8
XFILLER_54_431 VPWR VGND sg13g2_decap_8
XFILLER_26_133 VPWR VGND sg13g2_decap_8
XFILLER_82_784 VPWR VGND sg13g2_decap_8
XFILLER_70_924 VPWR VGND sg13g2_decap_8
XFILLER_42_648 VPWR VGND sg13g2_decap_8
XFILLER_23_840 VPWR VGND sg13g2_decap_8
XFILLER_25_56 VPWR VGND sg13g2_decap_8
XFILLER_41_147 VPWR VGND sg13g2_decap_8
XFILLER_10_501 VPWR VGND sg13g2_decap_8
XFILLER_22_361 VPWR VGND sg13g2_decap_8
XFILLER_10_578 VPWR VGND sg13g2_decap_8
XFILLER_41_77 VPWR VGND sg13g2_decap_8
XFILLER_68_1013 VPWR VGND sg13g2_decap_8
XFILLER_2_711 VPWR VGND sg13g2_decap_8
XFILLER_1_210 VPWR VGND sg13g2_decap_8
XFILLER_29_1019 VPWR VGND sg13g2_decap_8
XFILLER_89_350 VPWR VGND sg13g2_decap_8
XFILLER_104_672 VPWR VGND sg13g2_decap_8
XFILLER_49_214 VPWR VGND sg13g2_decap_8
XFILLER_2_788 VPWR VGND sg13g2_decap_8
XFILLER_106_70 VPWR VGND sg13g2_decap_8
XFILLER_103_182 VPWR VGND sg13g2_decap_8
XFILLER_1_287 VPWR VGND sg13g2_decap_8
XFILLER_92_504 VPWR VGND sg13g2_decap_8
XFILLER_77_567 VPWR VGND sg13g2_decap_8
XFILLER_66_41 VPWR VGND sg13g2_decap_8
XFILLER_65_707 VPWR VGND sg13g2_decap_8
XFILLER_58_770 VPWR VGND sg13g2_decap_8
XFILLER_64_228 VPWR VGND sg13g2_decap_8
XFILLER_57_280 VPWR VGND sg13g2_decap_8
XFILLER_46_921 VPWR VGND sg13g2_decap_8
XFILLER_45_420 VPWR VGND sg13g2_decap_8
XFILLER_18_623 VPWR VGND sg13g2_decap_8
XFILLER_17_144 VPWR VGND sg13g2_decap_8
XFILLER_73_795 VPWR VGND sg13g2_decap_8
XFILLER_61_935 VPWR VGND sg13g2_decap_8
XFILLER_46_998 VPWR VGND sg13g2_decap_8
XFILLER_45_497 VPWR VGND sg13g2_decap_8
XFILLER_33_637 VPWR VGND sg13g2_decap_8
XFILLER_82_84 VPWR VGND sg13g2_decap_8
XFILLER_72_294 VPWR VGND sg13g2_decap_8
XFILLER_60_445 VPWR VGND sg13g2_decap_8
XFILLER_14_840 VPWR VGND sg13g2_decap_8
XFILLER_13_350 VPWR VGND sg13g2_decap_8
XFILLER_32_158 VPWR VGND sg13g2_decap_8
XFILLER_9_343 VPWR VGND sg13g2_decap_8
XFILLER_12_1012 VPWR VGND sg13g2_decap_8
XFILLER_56_4 VPWR VGND sg13g2_decap_8
XFILLER_5_571 VPWR VGND sg13g2_decap_8
XFILLER_102_609 VPWR VGND sg13g2_decap_8
XFILLER_99_147 VPWR VGND sg13g2_decap_8
XFILLER_101_119 VPWR VGND sg13g2_decap_8
XFILLER_68_523 VPWR VGND sg13g2_decap_8
XFILLER_96_854 VPWR VGND sg13g2_decap_8
XFILLER_95_375 VPWR VGND sg13g2_decap_8
XFILLER_83_515 VPWR VGND sg13g2_decap_8
XFILLER_56_718 VPWR VGND sg13g2_decap_8
XFILLER_55_217 VPWR VGND sg13g2_decap_8
XFILLER_49_781 VPWR VGND sg13g2_decap_8
XFILLER_48_280 VPWR VGND sg13g2_decap_8
XFILLER_36_420 VPWR VGND sg13g2_decap_8
XFILLER_37_921 VPWR VGND sg13g2_decap_8
XFILLER_102_28 VPWR VGND sg13g2_decap_8
XFILLER_91_581 VPWR VGND sg13g2_decap_8
XFILLER_64_795 VPWR VGND sg13g2_decap_8
XFILLER_52_924 VPWR VGND sg13g2_decap_8
XFILLER_36_497 VPWR VGND sg13g2_decap_8
XFILLER_37_998 VPWR VGND sg13g2_decap_8
XFILLER_63_294 VPWR VGND sg13g2_decap_8
XFILLER_51_445 VPWR VGND sg13g2_decap_8
XFILLER_23_147 VPWR VGND sg13g2_decap_8
XFILLER_24_648 VPWR VGND sg13g2_decap_8
XFILLER_20_865 VPWR VGND sg13g2_decap_8
XFILLER_11_14 VPWR VGND sg13g2_decap_8
XFILLER_106_959 VPWR VGND sg13g2_decap_8
XFILLER_105_469 VPWR VGND sg13g2_decap_8
XFILLER_87_854 VPWR VGND sg13g2_decap_8
XFILLER_59_523 VPWR VGND sg13g2_decap_8
XFILLER_86_375 VPWR VGND sg13g2_decap_8
XFILLER_47_707 VPWR VGND sg13g2_decap_8
XFILLER_28_910 VPWR VGND sg13g2_decap_8
XFILLER_101_686 VPWR VGND sg13g2_decap_8
XFILLER_98_1028 VPWR VGND sg13g2_fill_1
XFILLER_74_526 VPWR VGND sg13g2_decap_8
XFILLER_46_228 VPWR VGND sg13g2_decap_8
XFILLER_100_196 VPWR VGND sg13g2_decap_8
XFILLER_27_431 VPWR VGND sg13g2_decap_8
XFILLER_39_291 VPWR VGND sg13g2_decap_8
XFILLER_82_581 VPWR VGND sg13g2_decap_8
XFILLER_70_721 VPWR VGND sg13g2_decap_8
XFILLER_55_784 VPWR VGND sg13g2_decap_8
XFILLER_43_924 VPWR VGND sg13g2_decap_8
XFILLER_28_987 VPWR VGND sg13g2_decap_8
XFILLER_36_77 VPWR VGND sg13g2_decap_8
XFILLER_42_445 VPWR VGND sg13g2_decap_8
XFILLER_15_648 VPWR VGND sg13g2_decap_8
XFILLER_70_798 VPWR VGND sg13g2_decap_8
XFILLER_52_21 VPWR VGND sg13g2_decap_8
XFILLER_14_147 VPWR VGND sg13g2_decap_8
XFILLER_35_1001 VPWR VGND sg13g2_decap_8
XFILLER_52_98 VPWR VGND sg13g2_decap_8
XFILLER_11_854 VPWR VGND sg13g2_decap_8
XFILLER_10_375 VPWR VGND sg13g2_decap_8
XFILLER_7_858 VPWR VGND sg13g2_decap_8
XFILLER_6_357 VPWR VGND sg13g2_decap_8
XFILLER_69_309 VPWR VGND sg13g2_decap_8
XFILLER_78_832 VPWR VGND sg13g2_decap_8
XFILLER_42_1005 VPWR VGND sg13g2_decap_8
XFILLER_2_585 VPWR VGND sg13g2_decap_8
XFILLER_93_824 VPWR VGND sg13g2_decap_8
XFILLER_77_364 VPWR VGND sg13g2_decap_8
XFILLER_77_84 VPWR VGND sg13g2_decap_8
XFILLER_65_504 VPWR VGND sg13g2_decap_8
X_31_ net10 net2 _02_ VPWR VGND sg13g2_xor2_1
XFILLER_38_707 VPWR VGND sg13g2_decap_8
XFILLER_92_301 VPWR VGND sg13g2_decap_8
XFILLER_19_910 VPWR VGND sg13g2_decap_8
XFILLER_37_228 VPWR VGND sg13g2_decap_8
XFILLER_18_420 VPWR VGND sg13g2_decap_8
XFILLER_93_61 VPWR VGND sg13g2_decap_8
XFILLER_92_378 VPWR VGND sg13g2_decap_8
XFILLER_80_518 VPWR VGND sg13g2_decap_8
XFILLER_46_795 VPWR VGND sg13g2_decap_8
XFILLER_19_987 VPWR VGND sg13g2_decap_8
XFILLER_34_935 VPWR VGND sg13g2_decap_8
XFILLER_73_592 VPWR VGND sg13g2_decap_8
XFILLER_61_732 VPWR VGND sg13g2_decap_8
XFILLER_45_294 VPWR VGND sg13g2_decap_8
Xheichips25_example_large_26 VPWR VGND uio_oe[1] sg13g2_tielo
XFILLER_18_497 VPWR VGND sg13g2_decap_8
Xheichips25_example_large_37 VPWR VGND uio_out[4] sg13g2_tielo
XFILLER_33_434 VPWR VGND sg13g2_decap_8
XFILLER_60_242 VPWR VGND sg13g2_decap_8
XFILLER_9_140 VPWR VGND sg13g2_decap_8
XFILLER_47_0 VPWR VGND sg13g2_decap_8
XFILLER_102_406 VPWR VGND sg13g2_decap_8
XFILLER_68_320 VPWR VGND sg13g2_decap_8
XFILLER_96_651 VPWR VGND sg13g2_decap_8
XFILLER_69_876 VPWR VGND sg13g2_decap_8
XFILLER_3_70 VPWR VGND sg13g2_decap_8
XFILLER_29_718 VPWR VGND sg13g2_decap_8
XFILLER_95_172 VPWR VGND sg13g2_decap_8
XFILLER_83_312 VPWR VGND sg13g2_decap_8
XFILLER_68_397 VPWR VGND sg13g2_decap_8
XFILLER_56_515 VPWR VGND sg13g2_decap_8
XFILLER_28_217 VPWR VGND sg13g2_decap_8
XFILLER_84_868 VPWR VGND sg13g2_decap_8
XFILLER_83_389 VPWR VGND sg13g2_decap_8
XFILLER_71_529 VPWR VGND sg13g2_decap_8
XFILLER_58_1001 VPWR VGND sg13g2_decap_8
XFILLER_52_721 VPWR VGND sg13g2_decap_8
XFILLER_25_924 VPWR VGND sg13g2_decap_8
XFILLER_37_795 VPWR VGND sg13g2_decap_8
XFILLER_64_592 VPWR VGND sg13g2_decap_8
XFILLER_24_445 VPWR VGND sg13g2_decap_8
XFILLER_36_294 VPWR VGND sg13g2_decap_8
XFILLER_51_242 VPWR VGND sg13g2_decap_8
XFILLER_52_798 VPWR VGND sg13g2_decap_8
XFILLER_40_938 VPWR VGND sg13g2_decap_8
XFILLER_20_662 VPWR VGND sg13g2_decap_8
XFILLER_22_46 VPWR VGND sg13g2_decap_8
XFILLER_98_39 VPWR VGND sg13g2_decap_8
XFILLER_106_756 VPWR VGND sg13g2_decap_8
XFILLER_105_266 VPWR VGND sg13g2_decap_8
XFILLER_78_139 VPWR VGND sg13g2_decap_8
XFILLER_59_320 VPWR VGND sg13g2_decap_8
XFILLER_102_973 VPWR VGND sg13g2_decap_8
XFILLER_87_651 VPWR VGND sg13g2_decap_8
XFILLER_47_504 VPWR VGND sg13g2_decap_8
XFILLER_47_21 VPWR VGND sg13g2_decap_8
XFILLER_101_483 VPWR VGND sg13g2_decap_8
XFILLER_86_172 VPWR VGND sg13g2_decap_8
XFILLER_74_323 VPWR VGND sg13g2_decap_8
XFILLER_59_397 VPWR VGND sg13g2_decap_8
XFILLER_19_217 VPWR VGND sg13g2_decap_8
XFILLER_90_816 VPWR VGND sg13g2_decap_8
XFILLER_75_868 VPWR VGND sg13g2_decap_8
XFILLER_47_98 VPWR VGND sg13g2_decap_8
XFILLER_62_518 VPWR VGND sg13g2_decap_8
XFILLER_16_924 VPWR VGND sg13g2_decap_8
XFILLER_28_784 VPWR VGND sg13g2_decap_8
XFILLER_63_42 VPWR VGND sg13g2_decap_8
XFILLER_55_581 VPWR VGND sg13g2_decap_8
XFILLER_43_721 VPWR VGND sg13g2_decap_8
XFILLER_15_445 VPWR VGND sg13g2_decap_8
XFILLER_42_242 VPWR VGND sg13g2_decap_8
XFILLER_70_595 VPWR VGND sg13g2_decap_8
XFILLER_43_798 VPWR VGND sg13g2_decap_8
XFILLER_31_938 VPWR VGND sg13g2_decap_8
XFILLER_11_651 VPWR VGND sg13g2_decap_8
XFILLER_30_448 VPWR VGND sg13g2_decap_8
XFILLER_10_172 VPWR VGND sg13g2_decap_8
XFILLER_7_655 VPWR VGND sg13g2_decap_8
XFILLER_6_154 VPWR VGND sg13g2_decap_8
XFILLER_98_949 VPWR VGND sg13g2_decap_8
XFILLER_69_106 VPWR VGND sg13g2_decap_8
XFILLER_3_861 VPWR VGND sg13g2_decap_8
XFILLER_40_7 VPWR VGND sg13g2_decap_8
XFILLER_97_448 VPWR VGND sg13g2_decap_8
XFILLER_2_382 VPWR VGND sg13g2_decap_8
XFILLER_38_504 VPWR VGND sg13g2_decap_8
XFILLER_93_621 VPWR VGND sg13g2_decap_8
XFILLER_77_161 VPWR VGND sg13g2_decap_8
XFILLER_66_846 VPWR VGND sg13g2_decap_8
XFILLER_65_301 VPWR VGND sg13g2_decap_8
XFILLER_93_698 VPWR VGND sg13g2_decap_8
XFILLER_92_175 VPWR VGND sg13g2_decap_8
XFILLER_81_816 VPWR VGND sg13g2_decap_8
XFILLER_80_315 VPWR VGND sg13g2_decap_8
XFILLER_65_378 VPWR VGND sg13g2_decap_8
XFILLER_53_518 VPWR VGND sg13g2_decap_8
XFILLER_19_784 VPWR VGND sg13g2_decap_8
XFILLER_74_890 VPWR VGND sg13g2_decap_8
XFILLER_46_592 VPWR VGND sg13g2_decap_8
XFILLER_18_294 VPWR VGND sg13g2_decap_8
XFILLER_34_732 VPWR VGND sg13g2_decap_8
XFILLER_33_231 VPWR VGND sg13g2_decap_8
XFILLER_22_949 VPWR VGND sg13g2_decap_8
XFILLER_21_448 VPWR VGND sg13g2_decap_8
XFILLER_88_1005 VPWR VGND sg13g2_decap_8
XFILLER_102_203 VPWR VGND sg13g2_decap_8
XFILLER_89_938 VPWR VGND sg13g2_decap_8
XFILLER_0_308 VPWR VGND sg13g2_decap_8
XFILLER_88_459 VPWR VGND sg13g2_decap_8
XFILLER_25_1022 VPWR VGND sg13g2_decap_8
XFILLER_69_673 VPWR VGND sg13g2_decap_8
XFILLER_56_312 VPWR VGND sg13g2_decap_8
XFILLER_29_515 VPWR VGND sg13g2_decap_8
XFILLER_84_665 VPWR VGND sg13g2_decap_8
XFILLER_72_805 VPWR VGND sg13g2_decap_8
XFILLER_68_194 VPWR VGND sg13g2_decap_8
XFILLER_57_868 VPWR VGND sg13g2_decap_8
XFILLER_56_389 VPWR VGND sg13g2_decap_8
XFILLER_44_529 VPWR VGND sg13g2_decap_8
XFILLER_17_46 VPWR VGND sg13g2_decap_8
XFILLER_83_186 VPWR VGND sg13g2_decap_8
XFILLER_71_326 VPWR VGND sg13g2_decap_8
XFILLER_25_721 VPWR VGND sg13g2_decap_8
XFILLER_37_592 VPWR VGND sg13g2_decap_8
XFILLER_24_242 VPWR VGND sg13g2_decap_8
XFILLER_80_882 VPWR VGND sg13g2_decap_8
XFILLER_52_595 VPWR VGND sg13g2_decap_8
XFILLER_13_938 VPWR VGND sg13g2_decap_8
XFILLER_25_798 VPWR VGND sg13g2_decap_8
XFILLER_40_735 VPWR VGND sg13g2_decap_8
XFILLER_12_459 VPWR VGND sg13g2_decap_8
XFILLER_33_56 VPWR VGND sg13g2_decap_8
XFILLER_32_1026 VPWR VGND sg13g2_fill_2
XFILLER_4_658 VPWR VGND sg13g2_decap_8
XFILLER_106_553 VPWR VGND sg13g2_decap_8
XFILLER_3_168 VPWR VGND sg13g2_decap_8
XFILLER_79_459 VPWR VGND sg13g2_decap_8
XFILLER_58_42 VPWR VGND sg13g2_decap_8
XFILLER_0_875 VPWR VGND sg13g2_decap_8
XFILLER_102_770 VPWR VGND sg13g2_decap_8
XFILLER_47_301 VPWR VGND sg13g2_decap_8
XFILLER_101_280 VPWR VGND sg13g2_decap_8
XFILLER_75_665 VPWR VGND sg13g2_decap_8
XFILLER_74_120 VPWR VGND sg13g2_decap_8
XFILLER_63_805 VPWR VGND sg13g2_decap_8
XFILLER_59_194 VPWR VGND sg13g2_decap_8
XFILLER_48_868 VPWR VGND sg13g2_decap_8
XFILLER_90_613 VPWR VGND sg13g2_decap_8
XFILLER_62_315 VPWR VGND sg13g2_decap_8
XFILLER_47_378 VPWR VGND sg13g2_decap_8
XFILLER_35_518 VPWR VGND sg13g2_decap_8
XFILLER_74_197 VPWR VGND sg13g2_decap_8
XFILLER_74_85 VPWR VGND sg13g2_decap_8
XFILLER_16_721 VPWR VGND sg13g2_decap_8
XFILLER_28_581 VPWR VGND sg13g2_decap_8
XFILLER_15_242 VPWR VGND sg13g2_decap_8
XFILLER_71_893 VPWR VGND sg13g2_decap_8
XFILLER_43_595 VPWR VGND sg13g2_decap_8
XFILLER_16_798 VPWR VGND sg13g2_decap_8
XFILLER_31_735 VPWR VGND sg13g2_decap_8
XFILLER_70_392 VPWR VGND sg13g2_decap_8
XFILLER_30_245 VPWR VGND sg13g2_decap_8
XFILLER_90_95 VPWR VGND sg13g2_decap_8
XFILLER_8_931 VPWR VGND sg13g2_decap_8
XFILLER_7_452 VPWR VGND sg13g2_decap_8
XFILLER_48_1022 VPWR VGND sg13g2_decap_8
XFILLER_98_746 VPWR VGND sg13g2_decap_8
XFILLER_100_707 VPWR VGND sg13g2_decap_8
XFILLER_97_245 VPWR VGND sg13g2_decap_8
XFILLER_39_802 VPWR VGND sg13g2_decap_8
XFILLER_38_301 VPWR VGND sg13g2_decap_8
XFILLER_94_952 VPWR VGND sg13g2_decap_8
XFILLER_66_643 VPWR VGND sg13g2_decap_8
XFILLER_39_879 VPWR VGND sg13g2_decap_8
XFILLER_81_613 VPWR VGND sg13g2_decap_8
XFILLER_54_816 VPWR VGND sg13g2_decap_8
XFILLER_53_315 VPWR VGND sg13g2_decap_8
XFILLER_26_518 VPWR VGND sg13g2_decap_8
XFILLER_38_378 VPWR VGND sg13g2_decap_8
XFILLER_93_495 VPWR VGND sg13g2_decap_8
XFILLER_80_112 VPWR VGND sg13g2_decap_8
XFILLER_65_175 VPWR VGND sg13g2_decap_8
XFILLER_19_581 VPWR VGND sg13g2_decap_8
XFILLER_80_189 VPWR VGND sg13g2_decap_8
XFILLER_62_882 VPWR VGND sg13g2_decap_8
XFILLER_55_1015 VPWR VGND sg13g2_decap_8
XFILLER_21_245 VPWR VGND sg13g2_decap_8
XFILLER_22_746 VPWR VGND sg13g2_decap_8
XFILLER_9_91 VPWR VGND sg13g2_decap_8
XFILLER_89_735 VPWR VGND sg13g2_decap_8
XFILLER_62_1008 VPWR VGND sg13g2_decap_8
XFILLER_0_105 VPWR VGND sg13g2_decap_8
XFILLER_103_567 VPWR VGND sg13g2_decap_8
XFILLER_95_18 VPWR VGND sg13g2_decap_8
XFILLER_88_256 VPWR VGND sg13g2_decap_8
XFILLER_69_470 VPWR VGND sg13g2_decap_8
XFILLER_29_312 VPWR VGND sg13g2_decap_8
XFILLER_85_952 VPWR VGND sg13g2_decap_8
XFILLER_28_56 VPWR VGND sg13g2_decap_8
XFILLER_84_462 VPWR VGND sg13g2_decap_8
XFILLER_72_602 VPWR VGND sg13g2_decap_8
XFILLER_57_665 VPWR VGND sg13g2_decap_8
XFILLER_45_805 VPWR VGND sg13g2_decap_8
XFILLER_17_529 VPWR VGND sg13g2_decap_8
XFILLER_71_123 VPWR VGND sg13g2_decap_8
XFILLER_56_186 VPWR VGND sg13g2_decap_8
XFILLER_44_326 VPWR VGND sg13g2_decap_8
XFILLER_29_389 VPWR VGND sg13g2_decap_8
XFILLER_72_679 VPWR VGND sg13g2_decap_8
XFILLER_44_11 VPWR VGND sg13g2_decap_8
XFILLER_53_882 VPWR VGND sg13g2_decap_8
XFILLER_13_735 VPWR VGND sg13g2_decap_8
XFILLER_25_595 VPWR VGND sg13g2_decap_8
XFILLER_52_392 VPWR VGND sg13g2_decap_8
XFILLER_44_88 VPWR VGND sg13g2_decap_8
XFILLER_40_532 VPWR VGND sg13g2_decap_8
XFILLER_9_728 VPWR VGND sg13g2_decap_8
XFILLER_12_256 VPWR VGND sg13g2_decap_8
XFILLER_60_32 VPWR VGND sg13g2_decap_8
XFILLER_8_238 VPWR VGND sg13g2_decap_8
XFILLER_5_956 VPWR VGND sg13g2_decap_8
XFILLER_106_350 VPWR VGND sg13g2_decap_8
XFILLER_4_455 VPWR VGND sg13g2_decap_8
XFILLER_79_256 VPWR VGND sg13g2_decap_8
XFILLER_69_85 VPWR VGND sg13g2_decap_8
XFILLER_68_908 VPWR VGND sg13g2_decap_8
XFILLER_0_672 VPWR VGND sg13g2_decap_8
XFILLER_39_109 VPWR VGND sg13g2_decap_8
XFILLER_94_259 VPWR VGND sg13g2_decap_8
XFILLER_76_963 VPWR VGND sg13g2_decap_8
XFILLER_85_84 VPWR VGND sg13g2_decap_8
XFILLER_75_462 VPWR VGND sg13g2_decap_8
XFILLER_63_602 VPWR VGND sg13g2_decap_8
XFILLER_48_665 VPWR VGND sg13g2_decap_8
XFILLER_36_805 VPWR VGND sg13g2_decap_8
XFILLER_90_410 VPWR VGND sg13g2_decap_8
XFILLER_62_112 VPWR VGND sg13g2_decap_8
XFILLER_47_175 VPWR VGND sg13g2_decap_8
XFILLER_35_315 VPWR VGND sg13g2_decap_8
XFILLER_91_966 VPWR VGND sg13g2_decap_8
XFILLER_63_679 VPWR VGND sg13g2_decap_8
XFILLER_90_487 VPWR VGND sg13g2_decap_8
XFILLER_62_189 VPWR VGND sg13g2_decap_8
XFILLER_50_329 VPWR VGND sg13g2_decap_8
XFILLER_44_893 VPWR VGND sg13g2_decap_8
XFILLER_93_5 VPWR VGND sg13g2_decap_8
XFILLER_71_690 VPWR VGND sg13g2_decap_8
XFILLER_43_392 VPWR VGND sg13g2_decap_8
XFILLER_16_595 VPWR VGND sg13g2_decap_8
XFILLER_31_532 VPWR VGND sg13g2_decap_8
XFILLER_86_4 VPWR VGND sg13g2_decap_8
XFILLER_85_1008 VPWR VGND sg13g2_decap_8
XFILLER_98_543 VPWR VGND sg13g2_decap_8
XFILLER_59_908 VPWR VGND sg13g2_decap_8
XFILLER_105_28 VPWR VGND sg13g2_decap_8
XFILLER_100_504 VPWR VGND sg13g2_decap_8
XFILLER_85_259 VPWR VGND sg13g2_decap_8
XFILLER_67_952 VPWR VGND sg13g2_decap_8
XFILLER_66_440 VPWR VGND sg13g2_decap_8
XFILLER_54_613 VPWR VGND sg13g2_decap_8
XFILLER_27_816 VPWR VGND sg13g2_decap_8
XFILLER_39_676 VPWR VGND sg13g2_decap_8
XFILLER_93_292 VPWR VGND sg13g2_decap_8
XFILLER_81_410 VPWR VGND sg13g2_decap_8
XFILLER_53_112 VPWR VGND sg13g2_decap_8
XFILLER_26_315 VPWR VGND sg13g2_decap_8
XFILLER_38_175 VPWR VGND sg13g2_decap_8
XFILLER_82_966 VPWR VGND sg13g2_decap_8
XFILLER_81_487 VPWR VGND sg13g2_decap_8
XFILLER_53_189 VPWR VGND sg13g2_decap_8
XFILLER_35_882 VPWR VGND sg13g2_decap_8
XFILLER_41_329 VPWR VGND sg13g2_decap_8
XFILLER_14_14 VPWR VGND sg13g2_decap_8
XFILLER_22_543 VPWR VGND sg13g2_decap_8
XFILLER_50_896 VPWR VGND sg13g2_decap_8
XFILLER_30_35 VPWR VGND sg13g2_decap_8
XFILLER_89_532 VPWR VGND sg13g2_decap_8
XFILLER_104_854 VPWR VGND sg13g2_decap_8
XFILLER_39_11 VPWR VGND sg13g2_decap_8
XFILLER_103_364 VPWR VGND sg13g2_decap_8
XFILLER_77_749 VPWR VGND sg13g2_decap_8
XFILLER_7_1019 VPWR VGND sg13g2_decap_8
XFILLER_1_469 VPWR VGND sg13g2_decap_8
XFILLER_58_952 VPWR VGND sg13g2_decap_8
XFILLER_39_88 VPWR VGND sg13g2_decap_8
XFILLER_73_900 VPWR VGND sg13g2_decap_8
XFILLER_57_462 VPWR VGND sg13g2_decap_8
XFILLER_45_602 VPWR VGND sg13g2_decap_8
XFILLER_18_805 VPWR VGND sg13g2_decap_8
XFILLER_55_21 VPWR VGND sg13g2_decap_8
XFILLER_17_326 VPWR VGND sg13g2_decap_8
XFILLER_29_186 VPWR VGND sg13g2_decap_8
XFILLER_73_977 VPWR VGND sg13g2_decap_8
XFILLER_45_679 VPWR VGND sg13g2_decap_8
XFILLER_44_123 VPWR VGND sg13g2_decap_8
XFILLER_33_819 VPWR VGND sg13g2_decap_8
XFILLER_72_476 VPWR VGND sg13g2_decap_8
XFILLER_60_627 VPWR VGND sg13g2_decap_8
XFILLER_55_98 VPWR VGND sg13g2_decap_8
XFILLER_26_882 VPWR VGND sg13g2_decap_8
XFILLER_13_532 VPWR VGND sg13g2_decap_8
XFILLER_25_392 VPWR VGND sg13g2_decap_8
XFILLER_71_53 VPWR VGND sg13g2_decap_8
XFILLER_9_525 VPWR VGND sg13g2_decap_8
XFILLER_41_896 VPWR VGND sg13g2_decap_8
XFILLER_5_753 VPWR VGND sg13g2_decap_8
XFILLER_99_329 VPWR VGND sg13g2_decap_8
XFILLER_4_252 VPWR VGND sg13g2_decap_8
XFILLER_68_705 VPWR VGND sg13g2_decap_8
XFILLER_95_557 VPWR VGND sg13g2_decap_8
XFILLER_76_760 VPWR VGND sg13g2_decap_8
XFILLER_67_259 VPWR VGND sg13g2_decap_8
XFILLER_64_900 VPWR VGND sg13g2_decap_8
XFILLER_49_963 VPWR VGND sg13g2_decap_8
XFILLER_48_462 VPWR VGND sg13g2_decap_8
XFILLER_36_602 VPWR VGND sg13g2_decap_8
XFILLER_35_112 VPWR VGND sg13g2_decap_8
XFILLER_91_763 VPWR VGND sg13g2_decap_8
XFILLER_64_977 VPWR VGND sg13g2_decap_8
XFILLER_36_679 VPWR VGND sg13g2_decap_8
XFILLER_91_1001 VPWR VGND sg13g2_decap_8
XFILLER_63_476 VPWR VGND sg13g2_decap_8
XFILLER_51_627 VPWR VGND sg13g2_decap_8
XFILLER_17_893 VPWR VGND sg13g2_decap_8
XFILLER_23_329 VPWR VGND sg13g2_decap_8
XFILLER_35_189 VPWR VGND sg13g2_decap_8
XFILLER_90_284 VPWR VGND sg13g2_decap_8
XFILLER_50_126 VPWR VGND sg13g2_decap_8
XFILLER_44_690 VPWR VGND sg13g2_decap_8
XFILLER_16_392 VPWR VGND sg13g2_decap_8
XFILLER_32_830 VPWR VGND sg13g2_decap_8
XFILLER_77_0 VPWR VGND sg13g2_decap_8
XFILLER_6_70 VPWR VGND sg13g2_decap_8
XFILLER_98_340 VPWR VGND sg13g2_decap_8
XFILLER_59_705 VPWR VGND sg13g2_decap_8
XFILLER_100_301 VPWR VGND sg13g2_decap_8
XFILLER_99_896 VPWR VGND sg13g2_decap_8
XFILLER_101_868 VPWR VGND sg13g2_decap_8
XFILLER_86_557 VPWR VGND sg13g2_decap_8
XFILLER_100_378 VPWR VGND sg13g2_decap_8
XFILLER_74_708 VPWR VGND sg13g2_decap_8
XFILLER_73_207 VPWR VGND sg13g2_decap_8
XFILLER_58_259 VPWR VGND sg13g2_decap_8
XFILLER_54_410 VPWR VGND sg13g2_decap_8
XFILLER_26_112 VPWR VGND sg13g2_decap_8
XFILLER_27_613 VPWR VGND sg13g2_decap_8
XFILLER_39_473 VPWR VGND sg13g2_decap_8
XFILLER_82_763 VPWR VGND sg13g2_decap_8
XFILLER_70_903 VPWR VGND sg13g2_decap_8
XFILLER_55_966 VPWR VGND sg13g2_decap_8
XFILLER_54_487 VPWR VGND sg13g2_decap_8
XFILLER_42_627 VPWR VGND sg13g2_decap_8
XFILLER_14_329 VPWR VGND sg13g2_decap_8
XFILLER_25_35 VPWR VGND sg13g2_decap_8
XFILLER_26_189 VPWR VGND sg13g2_decap_8
XFILLER_81_284 VPWR VGND sg13g2_decap_8
XFILLER_41_126 VPWR VGND sg13g2_decap_8
XFILLER_22_340 VPWR VGND sg13g2_decap_8
XFILLER_50_693 VPWR VGND sg13g2_decap_8
XFILLER_23_896 VPWR VGND sg13g2_decap_8
XFILLER_10_557 VPWR VGND sg13g2_decap_8
XFILLER_41_56 VPWR VGND sg13g2_decap_8
XFILLER_6_539 VPWR VGND sg13g2_decap_8
XFILLER_104_651 VPWR VGND sg13g2_decap_8
XFILLER_2_767 VPWR VGND sg13g2_decap_8
XFILLER_1_266 VPWR VGND sg13g2_decap_8
XFILLER_103_161 VPWR VGND sg13g2_decap_8
XFILLER_77_546 VPWR VGND sg13g2_decap_8
XFILLER_2_39 VPWR VGND sg13g2_decap_8
XFILLER_64_207 VPWR VGND sg13g2_decap_8
XFILLER_46_900 VPWR VGND sg13g2_decap_8
XFILLER_18_602 VPWR VGND sg13g2_decap_8
XFILLER_66_97 VPWR VGND sg13g2_decap_8
XFILLER_46_977 VPWR VGND sg13g2_decap_8
XFILLER_17_123 VPWR VGND sg13g2_decap_8
XFILLER_73_774 VPWR VGND sg13g2_decap_8
XFILLER_72_273 VPWR VGND sg13g2_decap_8
XFILLER_61_914 VPWR VGND sg13g2_decap_8
XFILLER_45_476 VPWR VGND sg13g2_decap_8
XFILLER_18_679 VPWR VGND sg13g2_decap_8
XFILLER_33_616 VPWR VGND sg13g2_decap_8
XFILLER_82_63 VPWR VGND sg13g2_decap_8
XFILLER_60_424 VPWR VGND sg13g2_decap_8
XFILLER_32_137 VPWR VGND sg13g2_decap_8
XFILLER_41_693 VPWR VGND sg13g2_decap_8
XFILLER_9_322 VPWR VGND sg13g2_decap_8
XFILLER_14_896 VPWR VGND sg13g2_decap_8
XFILLER_70_7 VPWR VGND sg13g2_decap_8
XFILLER_9_399 VPWR VGND sg13g2_decap_8
XFILLER_5_550 VPWR VGND sg13g2_decap_8
XFILLER_99_126 VPWR VGND sg13g2_decap_8
XFILLER_49_4 VPWR VGND sg13g2_decap_8
XFILLER_68_502 VPWR VGND sg13g2_decap_8
XFILLER_96_833 VPWR VGND sg13g2_decap_8
XFILLER_95_354 VPWR VGND sg13g2_decap_8
XFILLER_68_579 VPWR VGND sg13g2_decap_8
XFILLER_49_760 VPWR VGND sg13g2_decap_8
XFILLER_37_900 VPWR VGND sg13g2_decap_8
XFILLER_52_903 VPWR VGND sg13g2_decap_8
XFILLER_37_977 VPWR VGND sg13g2_decap_8
XFILLER_91_560 VPWR VGND sg13g2_decap_8
XFILLER_64_774 VPWR VGND sg13g2_decap_8
XFILLER_63_273 VPWR VGND sg13g2_decap_8
XFILLER_24_627 VPWR VGND sg13g2_decap_8
XFILLER_36_476 VPWR VGND sg13g2_decap_8
XFILLER_51_424 VPWR VGND sg13g2_decap_8
XFILLER_17_690 VPWR VGND sg13g2_decap_8
XFILLER_23_126 VPWR VGND sg13g2_decap_8
XFILLER_60_991 VPWR VGND sg13g2_decap_8
XFILLER_20_844 VPWR VGND sg13g2_decap_8
XFILLER_106_938 VPWR VGND sg13g2_decap_8
XFILLER_105_448 VPWR VGND sg13g2_decap_8
XFILLER_59_502 VPWR VGND sg13g2_decap_8
XFILLER_99_693 VPWR VGND sg13g2_decap_8
XFILLER_87_833 VPWR VGND sg13g2_decap_8
XFILLER_101_665 VPWR VGND sg13g2_decap_8
XFILLER_86_354 VPWR VGND sg13g2_decap_8
XFILLER_74_505 VPWR VGND sg13g2_decap_8
XFILLER_59_579 VPWR VGND sg13g2_decap_8
XFILLER_100_175 VPWR VGND sg13g2_decap_8
XFILLER_46_207 VPWR VGND sg13g2_decap_8
XFILLER_27_410 VPWR VGND sg13g2_decap_8
XFILLER_39_270 VPWR VGND sg13g2_decap_8
XFILLER_55_763 VPWR VGND sg13g2_decap_8
XFILLER_43_903 VPWR VGND sg13g2_decap_8
XFILLER_28_966 VPWR VGND sg13g2_decap_8
XFILLER_82_560 VPWR VGND sg13g2_decap_8
XFILLER_70_700 VPWR VGND sg13g2_decap_8
XFILLER_15_627 VPWR VGND sg13g2_decap_8
XFILLER_27_487 VPWR VGND sg13g2_decap_8
XFILLER_36_56 VPWR VGND sg13g2_decap_8
XFILLER_54_284 VPWR VGND sg13g2_decap_8
XFILLER_42_424 VPWR VGND sg13g2_decap_8
XFILLER_14_126 VPWR VGND sg13g2_decap_8
XFILLER_70_777 VPWR VGND sg13g2_decap_8
XFILLER_51_991 VPWR VGND sg13g2_decap_8
XFILLER_11_833 VPWR VGND sg13g2_decap_8
XFILLER_23_693 VPWR VGND sg13g2_decap_8
XFILLER_52_77 VPWR VGND sg13g2_decap_8
XFILLER_50_490 VPWR VGND sg13g2_decap_8
XFILLER_10_354 VPWR VGND sg13g2_decap_8
XFILLER_7_837 VPWR VGND sg13g2_decap_8
XFILLER_6_336 VPWR VGND sg13g2_decap_8
XFILLER_78_811 VPWR VGND sg13g2_decap_8
XFILLER_2_564 VPWR VGND sg13g2_decap_8
XFILLER_77_63 VPWR VGND sg13g2_decap_8
XFILLER_93_803 VPWR VGND sg13g2_decap_8
XFILLER_78_888 VPWR VGND sg13g2_decap_8
XFILLER_77_343 VPWR VGND sg13g2_decap_8
X_30_ net2 net10 _01_ VPWR VGND sg13g2_and2_1
XFILLER_42_1028 VPWR VGND sg13g2_fill_1
XFILLER_37_207 VPWR VGND sg13g2_decap_8
XFILLER_93_40 VPWR VGND sg13g2_decap_8
XFILLER_92_357 VPWR VGND sg13g2_decap_8
XFILLER_19_966 VPWR VGND sg13g2_decap_8
XFILLER_73_571 VPWR VGND sg13g2_decap_8
XFILLER_61_711 VPWR VGND sg13g2_decap_8
XFILLER_46_774 VPWR VGND sg13g2_decap_8
XFILLER_18_476 VPWR VGND sg13g2_decap_8
XFILLER_34_914 VPWR VGND sg13g2_decap_8
XFILLER_60_221 VPWR VGND sg13g2_decap_8
Xheichips25_example_large_27 VPWR VGND uio_oe[2] sg13g2_tielo
XFILLER_45_273 VPWR VGND sg13g2_decap_8
XFILLER_33_413 VPWR VGND sg13g2_decap_8
Xheichips25_example_large_38 VPWR VGND uio_out[5] sg13g2_tielo
XFILLER_61_788 VPWR VGND sg13g2_decap_8
XFILLER_60_298 VPWR VGND sg13g2_decap_8
XFILLER_42_991 VPWR VGND sg13g2_decap_8
XFILLER_14_693 VPWR VGND sg13g2_decap_8
XFILLER_41_490 VPWR VGND sg13g2_decap_8
XFILLER_9_196 VPWR VGND sg13g2_decap_8
XFILLER_96_630 VPWR VGND sg13g2_decap_8
XFILLER_69_855 VPWR VGND sg13g2_decap_8
XFILLER_95_151 VPWR VGND sg13g2_decap_8
XFILLER_84_847 VPWR VGND sg13g2_decap_8
XFILLER_68_376 VPWR VGND sg13g2_decap_8
XFILLER_3_1022 VPWR VGND sg13g2_decap_8
XFILLER_83_368 VPWR VGND sg13g2_decap_8
XFILLER_71_508 VPWR VGND sg13g2_decap_8
XFILLER_64_571 VPWR VGND sg13g2_decap_8
XFILLER_52_700 VPWR VGND sg13g2_decap_8
XFILLER_25_903 VPWR VGND sg13g2_decap_8
XFILLER_37_774 VPWR VGND sg13g2_decap_8
XFILLER_51_221 VPWR VGND sg13g2_decap_8
XFILLER_19_1008 VPWR VGND sg13g2_decap_8
XFILLER_24_424 VPWR VGND sg13g2_decap_8
XFILLER_36_273 VPWR VGND sg13g2_decap_8
XFILLER_52_777 VPWR VGND sg13g2_decap_8
XFILLER_40_917 VPWR VGND sg13g2_decap_8
XFILLER_51_298 VPWR VGND sg13g2_decap_8
XFILLER_33_980 VPWR VGND sg13g2_decap_8
XFILLER_20_641 VPWR VGND sg13g2_decap_8
XFILLER_22_25 VPWR VGND sg13g2_decap_8
XFILLER_98_18 VPWR VGND sg13g2_decap_8
XFILLER_106_735 VPWR VGND sg13g2_decap_8
XFILLER_105_245 VPWR VGND sg13g2_decap_8
XFILLER_0_7 VPWR VGND sg13g2_decap_8
XFILLER_99_490 VPWR VGND sg13g2_decap_8
XFILLER_87_630 VPWR VGND sg13g2_decap_8
XFILLER_78_118 VPWR VGND sg13g2_decap_8
XFILLER_102_952 VPWR VGND sg13g2_decap_8
XFILLER_101_462 VPWR VGND sg13g2_decap_8
XFILLER_86_151 VPWR VGND sg13g2_decap_8
XFILLER_75_847 VPWR VGND sg13g2_decap_8
XFILLER_74_302 VPWR VGND sg13g2_decap_8
XFILLER_59_376 VPWR VGND sg13g2_decap_8
XFILLER_47_77 VPWR VGND sg13g2_decap_8
XFILLER_74_379 VPWR VGND sg13g2_decap_8
XFILLER_55_560 VPWR VGND sg13g2_decap_8
XFILLER_43_700 VPWR VGND sg13g2_decap_8
XFILLER_16_903 VPWR VGND sg13g2_decap_8
XFILLER_28_763 VPWR VGND sg13g2_decap_8
XFILLER_63_21 VPWR VGND sg13g2_decap_8
XFILLER_42_221 VPWR VGND sg13g2_decap_8
XFILLER_15_424 VPWR VGND sg13g2_decap_8
XFILLER_27_284 VPWR VGND sg13g2_decap_8
XFILLER_43_777 VPWR VGND sg13g2_decap_8
XFILLER_31_917 VPWR VGND sg13g2_decap_8
XFILLER_70_574 VPWR VGND sg13g2_decap_8
XFILLER_63_98 VPWR VGND sg13g2_decap_8
XFILLER_24_991 VPWR VGND sg13g2_decap_8
XFILLER_30_427 VPWR VGND sg13g2_decap_8
XFILLER_42_298 VPWR VGND sg13g2_decap_8
XFILLER_8_49 VPWR VGND sg13g2_decap_8
XFILLER_11_630 VPWR VGND sg13g2_decap_8
XFILLER_23_490 VPWR VGND sg13g2_decap_8
XFILLER_10_151 VPWR VGND sg13g2_decap_8
XFILLER_7_634 VPWR VGND sg13g2_decap_8
XFILLER_6_133 VPWR VGND sg13g2_decap_8
XFILLER_3_840 VPWR VGND sg13g2_decap_8
XFILLER_98_928 VPWR VGND sg13g2_decap_8
XFILLER_97_427 VPWR VGND sg13g2_decap_8
XFILLER_88_95 VPWR VGND sg13g2_decap_8
XFILLER_2_361 VPWR VGND sg13g2_decap_8
XFILLER_33_7 VPWR VGND sg13g2_decap_8
XFILLER_77_140 VPWR VGND sg13g2_decap_8
XFILLER_93_600 VPWR VGND sg13g2_decap_8
XFILLER_78_685 VPWR VGND sg13g2_decap_8
XFILLER_66_825 VPWR VGND sg13g2_decap_8
XFILLER_65_357 VPWR VGND sg13g2_decap_8
XFILLER_93_677 VPWR VGND sg13g2_decap_8
XFILLER_92_154 VPWR VGND sg13g2_decap_8
XFILLER_19_763 VPWR VGND sg13g2_decap_8
XFILLER_34_711 VPWR VGND sg13g2_decap_8
XFILLER_46_571 VPWR VGND sg13g2_decap_8
XFILLER_18_273 VPWR VGND sg13g2_decap_8
XFILLER_33_210 VPWR VGND sg13g2_decap_8
XFILLER_61_585 VPWR VGND sg13g2_decap_8
XFILLER_15_991 VPWR VGND sg13g2_decap_8
XFILLER_21_427 VPWR VGND sg13g2_decap_8
XFILLER_22_928 VPWR VGND sg13g2_decap_8
XFILLER_33_287 VPWR VGND sg13g2_decap_8
XFILLER_34_788 VPWR VGND sg13g2_decap_8
XFILLER_105_1022 VPWR VGND sg13g2_decap_8
XFILLER_14_490 VPWR VGND sg13g2_decap_8
XFILLER_88_1028 VPWR VGND sg13g2_fill_1
XFILLER_30_994 VPWR VGND sg13g2_decap_8
XFILLER_89_917 VPWR VGND sg13g2_decap_8
XFILLER_103_749 VPWR VGND sg13g2_decap_8
XFILLER_88_438 VPWR VGND sg13g2_decap_8
XFILLER_25_1001 VPWR VGND sg13g2_decap_8
XFILLER_102_259 VPWR VGND sg13g2_decap_8
XFILLER_69_652 VPWR VGND sg13g2_decap_8
XFILLER_97_994 VPWR VGND sg13g2_decap_8
XFILLER_68_173 VPWR VGND sg13g2_decap_8
XFILLER_84_644 VPWR VGND sg13g2_decap_8
XFILLER_57_847 VPWR VGND sg13g2_decap_8
XFILLER_83_165 VPWR VGND sg13g2_decap_8
XFILLER_71_305 VPWR VGND sg13g2_decap_8
XFILLER_56_368 VPWR VGND sg13g2_decap_8
XFILLER_44_508 VPWR VGND sg13g2_decap_8
XFILLER_17_25 VPWR VGND sg13g2_decap_8
XFILLER_25_700 VPWR VGND sg13g2_decap_8
XFILLER_37_571 VPWR VGND sg13g2_decap_8
XFILLER_80_861 VPWR VGND sg13g2_decap_8
XFILLER_13_917 VPWR VGND sg13g2_decap_8
XFILLER_24_221 VPWR VGND sg13g2_decap_8
XFILLER_25_777 VPWR VGND sg13g2_decap_8
XFILLER_52_574 VPWR VGND sg13g2_decap_8
XFILLER_40_714 VPWR VGND sg13g2_decap_8
XFILLER_12_438 VPWR VGND sg13g2_decap_8
XFILLER_24_298 VPWR VGND sg13g2_decap_8
XFILLER_33_35 VPWR VGND sg13g2_decap_8
XFILLER_32_1005 VPWR VGND sg13g2_decap_8
XFILLER_21_994 VPWR VGND sg13g2_decap_8
XFILLER_106_532 VPWR VGND sg13g2_decap_8
XFILLER_4_637 VPWR VGND sg13g2_decap_8
XFILLER_3_147 VPWR VGND sg13g2_decap_8
XFILLER_79_438 VPWR VGND sg13g2_decap_8
XFILLER_58_21 VPWR VGND sg13g2_decap_8
XFILLER_0_854 VPWR VGND sg13g2_decap_8
XFILLER_59_173 VPWR VGND sg13g2_decap_8
XFILLER_58_98 VPWR VGND sg13g2_decap_8
XFILLER_75_644 VPWR VGND sg13g2_decap_8
XFILLER_48_847 VPWR VGND sg13g2_decap_8
XFILLER_74_42 VPWR VGND sg13g2_decap_8
XFILLER_47_357 VPWR VGND sg13g2_decap_8
XFILLER_16_700 VPWR VGND sg13g2_decap_8
XFILLER_28_560 VPWR VGND sg13g2_decap_8
XFILLER_74_176 VPWR VGND sg13g2_decap_8
XFILLER_74_53 VPWR VGND sg13g2_fill_1
XFILLER_90_669 VPWR VGND sg13g2_decap_8
XFILLER_15_221 VPWR VGND sg13g2_decap_8
XFILLER_16_777 VPWR VGND sg13g2_decap_8
XFILLER_71_872 VPWR VGND sg13g2_decap_8
XFILLER_70_371 VPWR VGND sg13g2_decap_8
XFILLER_43_574 VPWR VGND sg13g2_decap_8
XFILLER_31_714 VPWR VGND sg13g2_decap_8
XFILLER_15_298 VPWR VGND sg13g2_decap_8
XFILLER_30_224 VPWR VGND sg13g2_decap_8
XFILLER_90_74 VPWR VGND sg13g2_decap_8
XFILLER_8_910 VPWR VGND sg13g2_decap_8
XFILLER_7_431 VPWR VGND sg13g2_decap_8
XFILLER_8_987 VPWR VGND sg13g2_decap_8
XFILLER_48_1001 VPWR VGND sg13g2_decap_8
XFILLER_98_725 VPWR VGND sg13g2_decap_8
XFILLER_97_224 VPWR VGND sg13g2_decap_8
XFILLER_94_931 VPWR VGND sg13g2_decap_8
XFILLER_66_622 VPWR VGND sg13g2_decap_8
XFILLER_78_482 VPWR VGND sg13g2_decap_8
XFILLER_39_858 VPWR VGND sg13g2_decap_8
XFILLER_93_474 VPWR VGND sg13g2_decap_8
XFILLER_65_154 VPWR VGND sg13g2_decap_8
XFILLER_19_560 VPWR VGND sg13g2_decap_8
XFILLER_38_357 VPWR VGND sg13g2_decap_8
XFILLER_66_699 VPWR VGND sg13g2_decap_8
XFILLER_81_669 VPWR VGND sg13g2_decap_8
XFILLER_62_861 VPWR VGND sg13g2_decap_8
XFILLER_80_168 VPWR VGND sg13g2_decap_8
XFILLER_22_725 VPWR VGND sg13g2_decap_8
XFILLER_34_585 VPWR VGND sg13g2_decap_8
XFILLER_61_382 VPWR VGND sg13g2_decap_8
XFILLER_21_224 VPWR VGND sg13g2_decap_8
XFILLER_9_70 VPWR VGND sg13g2_decap_8
XFILLER_30_791 VPWR VGND sg13g2_decap_8
XFILLER_89_714 VPWR VGND sg13g2_decap_8
XFILLER_103_546 VPWR VGND sg13g2_decap_8
XFILLER_88_235 VPWR VGND sg13g2_decap_8
XFILLER_97_791 VPWR VGND sg13g2_decap_8
XFILLER_85_931 VPWR VGND sg13g2_decap_8
XFILLER_57_644 VPWR VGND sg13g2_decap_8
XFILLER_28_35 VPWR VGND sg13g2_decap_8
XFILLER_84_441 VPWR VGND sg13g2_decap_8
XFILLER_56_165 VPWR VGND sg13g2_decap_8
XFILLER_44_305 VPWR VGND sg13g2_decap_8
XFILLER_17_508 VPWR VGND sg13g2_decap_8
XFILLER_29_368 VPWR VGND sg13g2_decap_8
XFILLER_71_102 VPWR VGND sg13g2_decap_8
XFILLER_72_658 VPWR VGND sg13g2_decap_8
XFILLER_60_809 VPWR VGND sg13g2_decap_8
XFILLER_53_861 VPWR VGND sg13g2_decap_8
XFILLER_71_179 VPWR VGND sg13g2_decap_8
XFILLER_52_371 VPWR VGND sg13g2_decap_8
XFILLER_44_67 VPWR VGND sg13g2_decap_8
XFILLER_13_714 VPWR VGND sg13g2_decap_8
XFILLER_25_574 VPWR VGND sg13g2_decap_8
XFILLER_40_511 VPWR VGND sg13g2_decap_8
XFILLER_9_707 VPWR VGND sg13g2_decap_8
XFILLER_12_235 VPWR VGND sg13g2_decap_8
XFILLER_8_217 VPWR VGND sg13g2_decap_8
XFILLER_40_588 VPWR VGND sg13g2_decap_8
XFILLER_100_84 VPWR VGND sg13g2_decap_8
XFILLER_21_791 VPWR VGND sg13g2_decap_8
XFILLER_60_88 VPWR VGND sg13g2_decap_8
XFILLER_5_935 VPWR VGND sg13g2_decap_8
XFILLER_4_434 VPWR VGND sg13g2_decap_8
XFILLER_5_39 VPWR VGND sg13g2_decap_8
XFILLER_69_64 VPWR VGND sg13g2_decap_8
XFILLER_69_42 VPWR VGND sg13g2_decap_8
XFILLER_79_235 VPWR VGND sg13g2_decap_8
XFILLER_95_739 VPWR VGND sg13g2_decap_8
XFILLER_0_651 VPWR VGND sg13g2_decap_8
XFILLER_94_238 VPWR VGND sg13g2_decap_8
XFILLER_76_942 VPWR VGND sg13g2_decap_8
XFILLER_48_644 VPWR VGND sg13g2_decap_8
XFILLER_85_63 VPWR VGND sg13g2_decap_8
XFILLER_75_441 VPWR VGND sg13g2_decap_8
XFILLER_47_154 VPWR VGND sg13g2_decap_8
XFILLER_91_945 VPWR VGND sg13g2_decap_8
XFILLER_90_466 VPWR VGND sg13g2_decap_8
XFILLER_63_658 VPWR VGND sg13g2_decap_8
XFILLER_51_809 VPWR VGND sg13g2_decap_8
XFILLER_62_168 VPWR VGND sg13g2_decap_8
XFILLER_50_308 VPWR VGND sg13g2_decap_8
XFILLER_44_872 VPWR VGND sg13g2_decap_8
XFILLER_43_371 VPWR VGND sg13g2_decap_8
XFILLER_16_574 VPWR VGND sg13g2_decap_8
XFILLER_31_511 VPWR VGND sg13g2_decap_8
XFILLER_31_588 VPWR VGND sg13g2_decap_8
XFILLER_8_784 VPWR VGND sg13g2_decap_8
XFILLER_98_522 VPWR VGND sg13g2_decap_8
XFILLER_98_599 VPWR VGND sg13g2_decap_8
XFILLER_86_739 VPWR VGND sg13g2_decap_8
XFILLER_85_238 VPWR VGND sg13g2_decap_8
XFILLER_67_931 VPWR VGND sg13g2_decap_8
XFILLER_22_1026 VPWR VGND sg13g2_fill_2
XFILLER_38_154 VPWR VGND sg13g2_decap_8
XFILLER_39_655 VPWR VGND sg13g2_decap_8
XFILLER_93_271 VPWR VGND sg13g2_decap_8
XFILLER_82_945 VPWR VGND sg13g2_decap_8
XFILLER_66_496 VPWR VGND sg13g2_decap_8
XFILLER_81_466 VPWR VGND sg13g2_decap_8
XFILLER_54_669 VPWR VGND sg13g2_decap_8
XFILLER_42_809 VPWR VGND sg13g2_decap_8
XFILLER_53_168 VPWR VGND sg13g2_decap_8
XFILLER_35_861 VPWR VGND sg13g2_decap_8
XFILLER_41_308 VPWR VGND sg13g2_decap_8
XFILLER_22_522 VPWR VGND sg13g2_decap_8
XFILLER_34_382 VPWR VGND sg13g2_decap_8
XFILLER_50_875 VPWR VGND sg13g2_decap_8
XFILLER_10_739 VPWR VGND sg13g2_decap_8
XFILLER_22_599 VPWR VGND sg13g2_decap_8
XFILLER_30_14 VPWR VGND sg13g2_decap_8
XFILLER_100_7 VPWR VGND sg13g2_decap_8
XFILLER_104_833 VPWR VGND sg13g2_decap_8
XFILLER_89_511 VPWR VGND sg13g2_decap_8
XFILLER_2_949 VPWR VGND sg13g2_decap_8
XFILLER_103_343 VPWR VGND sg13g2_decap_8
XFILLER_1_448 VPWR VGND sg13g2_decap_8
XFILLER_89_588 VPWR VGND sg13g2_decap_8
XFILLER_77_728 VPWR VGND sg13g2_decap_8
XFILLER_76_249 VPWR VGND sg13g2_decap_8
XFILLER_58_931 VPWR VGND sg13g2_decap_8
XFILLER_39_67 VPWR VGND sg13g2_decap_8
XFILLER_57_441 VPWR VGND sg13g2_decap_8
XFILLER_44_102 VPWR VGND sg13g2_decap_8
XFILLER_17_305 VPWR VGND sg13g2_decap_8
XFILLER_29_165 VPWR VGND sg13g2_decap_8
XFILLER_73_956 VPWR VGND sg13g2_decap_8
XFILLER_72_455 VPWR VGND sg13g2_decap_8
XFILLER_55_77 VPWR VGND sg13g2_decap_8
XFILLER_45_658 VPWR VGND sg13g2_decap_8
XFILLER_60_606 VPWR VGND sg13g2_decap_8
XFILLER_44_179 VPWR VGND sg13g2_decap_8
XFILLER_26_861 VPWR VGND sg13g2_decap_8
XFILLER_32_319 VPWR VGND sg13g2_decap_8
XFILLER_38_1022 VPWR VGND sg13g2_decap_8
XFILLER_13_511 VPWR VGND sg13g2_decap_8
XFILLER_25_371 VPWR VGND sg13g2_decap_8
XFILLER_71_32 VPWR VGND sg13g2_decap_8
XFILLER_41_875 VPWR VGND sg13g2_decap_8
XFILLER_9_504 VPWR VGND sg13g2_decap_8
XFILLER_13_588 VPWR VGND sg13g2_decap_8
XFILLER_40_385 VPWR VGND sg13g2_decap_8
XFILLER_5_732 VPWR VGND sg13g2_decap_8
XFILLER_99_308 VPWR VGND sg13g2_decap_8
XFILLER_4_231 VPWR VGND sg13g2_decap_8
XFILLER_45_1015 VPWR VGND sg13g2_decap_8
XFILLER_96_84 VPWR VGND sg13g2_decap_8
XFILLER_95_536 VPWR VGND sg13g2_decap_8
XFILLER_67_238 VPWR VGND sg13g2_decap_8
XFILLER_49_942 VPWR VGND sg13g2_decap_8
XFILLER_48_441 VPWR VGND sg13g2_decap_8
XFILLER_91_742 VPWR VGND sg13g2_decap_8
XFILLER_64_956 VPWR VGND sg13g2_decap_8
XFILLER_63_455 VPWR VGND sg13g2_decap_8
XFILLER_24_809 VPWR VGND sg13g2_decap_8
XFILLER_36_658 VPWR VGND sg13g2_decap_8
XFILLER_90_263 VPWR VGND sg13g2_decap_8
XFILLER_51_606 VPWR VGND sg13g2_decap_8
XFILLER_50_105 VPWR VGND sg13g2_decap_8
XFILLER_17_872 VPWR VGND sg13g2_decap_8
XFILLER_23_308 VPWR VGND sg13g2_decap_8
XFILLER_35_168 VPWR VGND sg13g2_decap_8
XFILLER_16_371 VPWR VGND sg13g2_decap_8
XFILLER_52_1008 VPWR VGND sg13g2_decap_8
XFILLER_32_886 VPWR VGND sg13g2_decap_8
XFILLER_31_385 VPWR VGND sg13g2_decap_8
XFILLER_8_581 VPWR VGND sg13g2_decap_8
XFILLER_99_875 VPWR VGND sg13g2_decap_8
XFILLER_101_847 VPWR VGND sg13g2_decap_8
XFILLER_98_396 VPWR VGND sg13g2_decap_8
XFILLER_86_536 VPWR VGND sg13g2_decap_8
XFILLER_58_238 VPWR VGND sg13g2_decap_8
XFILLER_100_357 VPWR VGND sg13g2_decap_8
XFILLER_39_452 VPWR VGND sg13g2_decap_8
XFILLER_55_945 VPWR VGND sg13g2_decap_8
XFILLER_82_742 VPWR VGND sg13g2_decap_8
XFILLER_66_293 VPWR VGND sg13g2_decap_8
XFILLER_15_809 VPWR VGND sg13g2_decap_8
XFILLER_27_669 VPWR VGND sg13g2_decap_8
XFILLER_81_263 VPWR VGND sg13g2_decap_8
XFILLER_54_466 VPWR VGND sg13g2_decap_8
XFILLER_42_606 VPWR VGND sg13g2_decap_8
XFILLER_14_308 VPWR VGND sg13g2_decap_8
XFILLER_25_14 VPWR VGND sg13g2_decap_8
XFILLER_26_168 VPWR VGND sg13g2_decap_8
XFILLER_41_105 VPWR VGND sg13g2_decap_8
XFILLER_70_959 VPWR VGND sg13g2_decap_8
XFILLER_23_875 VPWR VGND sg13g2_decap_8
XFILLER_50_672 VPWR VGND sg13g2_decap_8
XFILLER_10_536 VPWR VGND sg13g2_decap_8
XFILLER_6_518 VPWR VGND sg13g2_decap_8
XFILLER_22_396 VPWR VGND sg13g2_decap_8
XFILLER_41_35 VPWR VGND sg13g2_decap_8
XFILLER_104_630 VPWR VGND sg13g2_decap_8
XFILLER_2_746 VPWR VGND sg13g2_decap_8
XFILLER_103_140 VPWR VGND sg13g2_decap_8
XFILLER_1_245 VPWR VGND sg13g2_decap_8
XFILLER_89_385 VPWR VGND sg13g2_decap_8
XFILLER_77_525 VPWR VGND sg13g2_decap_8
XFILLER_2_18 VPWR VGND sg13g2_decap_8
XFILLER_49_249 VPWR VGND sg13g2_decap_8
XFILLER_92_539 VPWR VGND sg13g2_decap_8
XFILLER_66_76 VPWR VGND sg13g2_decap_8
XFILLER_17_102 VPWR VGND sg13g2_decap_8
XFILLER_73_753 VPWR VGND sg13g2_decap_8
XFILLER_46_956 VPWR VGND sg13g2_decap_8
XFILLER_45_455 VPWR VGND sg13g2_decap_8
XFILLER_18_658 VPWR VGND sg13g2_decap_8
XFILLER_75_1008 VPWR VGND sg13g2_decap_8
XFILLER_72_252 VPWR VGND sg13g2_decap_8
XFILLER_60_403 VPWR VGND sg13g2_decap_8
XFILLER_17_179 VPWR VGND sg13g2_decap_8
XFILLER_82_42 VPWR VGND sg13g2_decap_8
XFILLER_32_116 VPWR VGND sg13g2_decap_8
XFILLER_9_301 VPWR VGND sg13g2_decap_8
XFILLER_14_875 VPWR VGND sg13g2_decap_8
XFILLER_41_672 VPWR VGND sg13g2_decap_8
XFILLER_13_385 VPWR VGND sg13g2_decap_8
XFILLER_40_182 VPWR VGND sg13g2_decap_8
XFILLER_9_378 VPWR VGND sg13g2_decap_8
XFILLER_63_7 VPWR VGND sg13g2_decap_8
XFILLER_99_105 VPWR VGND sg13g2_decap_8
XFILLER_96_812 VPWR VGND sg13g2_decap_8
XFILLER_95_333 VPWR VGND sg13g2_decap_8
XFILLER_96_889 VPWR VGND sg13g2_decap_8
XFILLER_68_558 VPWR VGND sg13g2_decap_8
XFILLER_64_753 VPWR VGND sg13g2_decap_8
XFILLER_37_956 VPWR VGND sg13g2_decap_8
XFILLER_63_252 VPWR VGND sg13g2_decap_8
XFILLER_51_403 VPWR VGND sg13g2_decap_8
XFILLER_24_606 VPWR VGND sg13g2_decap_8
XFILLER_36_455 VPWR VGND sg13g2_decap_8
XFILLER_52_959 VPWR VGND sg13g2_decap_8
XFILLER_23_105 VPWR VGND sg13g2_decap_8
XFILLER_60_970 VPWR VGND sg13g2_decap_8
XFILLER_20_823 VPWR VGND sg13g2_decap_8
XFILLER_32_683 VPWR VGND sg13g2_decap_8
XFILLER_31_182 VPWR VGND sg13g2_decap_8
XFILLER_106_917 VPWR VGND sg13g2_decap_8
XFILLER_11_49 VPWR VGND sg13g2_decap_8
XFILLER_105_427 VPWR VGND sg13g2_decap_8
XFILLER_99_672 VPWR VGND sg13g2_decap_8
XFILLER_87_812 VPWR VGND sg13g2_decap_8
XFILLER_101_644 VPWR VGND sg13g2_decap_8
XFILLER_98_193 VPWR VGND sg13g2_decap_8
XFILLER_87_889 VPWR VGND sg13g2_decap_8
XFILLER_86_333 VPWR VGND sg13g2_decap_8
XFILLER_59_558 VPWR VGND sg13g2_decap_8
XFILLER_100_154 VPWR VGND sg13g2_decap_8
XFILLER_98_1019 VPWR VGND sg13g2_decap_8
XFILLER_55_742 VPWR VGND sg13g2_decap_8
XFILLER_28_945 VPWR VGND sg13g2_decap_8
XFILLER_36_35 VPWR VGND sg13g2_decap_8
XFILLER_54_263 VPWR VGND sg13g2_decap_8
XFILLER_42_403 VPWR VGND sg13g2_decap_8
XFILLER_15_606 VPWR VGND sg13g2_decap_8
XFILLER_27_466 VPWR VGND sg13g2_decap_8
XFILLER_43_959 VPWR VGND sg13g2_decap_8
XFILLER_14_105 VPWR VGND sg13g2_decap_8
XFILLER_70_756 VPWR VGND sg13g2_decap_8
XFILLER_30_609 VPWR VGND sg13g2_decap_8
XFILLER_52_56 VPWR VGND sg13g2_decap_8
XFILLER_51_970 VPWR VGND sg13g2_decap_8
XFILLER_11_812 VPWR VGND sg13g2_decap_8
XFILLER_23_672 VPWR VGND sg13g2_decap_8
XFILLER_10_333 VPWR VGND sg13g2_decap_8
XFILLER_7_816 VPWR VGND sg13g2_decap_8
XFILLER_22_193 VPWR VGND sg13g2_decap_8
XFILLER_6_315 VPWR VGND sg13g2_decap_8
XFILLER_11_889 VPWR VGND sg13g2_decap_8
XFILLER_97_609 VPWR VGND sg13g2_decap_8
XFILLER_81_1012 VPWR VGND sg13g2_decap_8
XFILLER_2_543 VPWR VGND sg13g2_decap_8
XFILLER_105_994 VPWR VGND sg13g2_decap_8
XFILLER_96_119 VPWR VGND sg13g2_decap_8
XFILLER_89_182 VPWR VGND sg13g2_decap_8
XFILLER_77_322 VPWR VGND sg13g2_decap_8
XFILLER_77_42 VPWR VGND sg13g2_decap_8
XFILLER_78_867 VPWR VGND sg13g2_decap_8
XFILLER_77_399 VPWR VGND sg13g2_decap_8
XFILLER_65_539 VPWR VGND sg13g2_decap_8
XFILLER_93_859 VPWR VGND sg13g2_decap_8
XFILLER_92_336 VPWR VGND sg13g2_decap_8
XFILLER_46_753 VPWR VGND sg13g2_decap_8
XFILLER_19_945 VPWR VGND sg13g2_decap_8
XFILLER_73_550 VPWR VGND sg13g2_decap_8
XFILLER_45_252 VPWR VGND sg13g2_decap_8
XFILLER_18_455 VPWR VGND sg13g2_decap_8
XFILLER_93_96 VPWR VGND sg13g2_decap_8
XFILLER_60_200 VPWR VGND sg13g2_decap_8
Xheichips25_example_large_28 VPWR VGND uio_oe[3] sg13g2_tielo
Xheichips25_example_large_39 VPWR VGND uio_out[6] sg13g2_tielo
XFILLER_61_767 VPWR VGND sg13g2_decap_8
XFILLER_21_609 VPWR VGND sg13g2_decap_8
XFILLER_33_469 VPWR VGND sg13g2_decap_8
XFILLER_60_277 VPWR VGND sg13g2_decap_8
XFILLER_42_970 VPWR VGND sg13g2_decap_8
XFILLER_14_672 VPWR VGND sg13g2_decap_8
XFILLER_13_182 VPWR VGND sg13g2_decap_8
XFILLER_9_175 VPWR VGND sg13g2_decap_8
XFILLER_61_4 VPWR VGND sg13g2_decap_8
XFILLER_6_882 VPWR VGND sg13g2_decap_8
XFILLER_87_119 VPWR VGND sg13g2_decap_8
XFILLER_69_834 VPWR VGND sg13g2_decap_8
XFILLER_95_130 VPWR VGND sg13g2_decap_8
XFILLER_68_355 VPWR VGND sg13g2_decap_8
XFILLER_96_686 VPWR VGND sg13g2_decap_8
XFILLER_84_826 VPWR VGND sg13g2_decap_8
XFILLER_3_1001 VPWR VGND sg13g2_decap_8
XFILLER_83_347 VPWR VGND sg13g2_decap_8
XFILLER_64_550 VPWR VGND sg13g2_decap_8
XFILLER_24_403 VPWR VGND sg13g2_decap_8
XFILLER_36_252 VPWR VGND sg13g2_decap_8
XFILLER_37_753 VPWR VGND sg13g2_decap_8
XFILLER_51_200 VPWR VGND sg13g2_decap_8
XFILLER_25_959 VPWR VGND sg13g2_decap_8
XFILLER_52_756 VPWR VGND sg13g2_decap_8
XFILLER_51_277 VPWR VGND sg13g2_decap_8
XFILLER_11_119 VPWR VGND sg13g2_decap_8
XFILLER_20_620 VPWR VGND sg13g2_decap_8
XFILLER_32_480 VPWR VGND sg13g2_decap_8
XFILLER_20_697 VPWR VGND sg13g2_decap_8
XFILLER_106_714 VPWR VGND sg13g2_decap_8
XFILLER_4_819 VPWR VGND sg13g2_decap_8
XFILLER_105_224 VPWR VGND sg13g2_decap_8
XFILLER_3_329 VPWR VGND sg13g2_decap_8
XFILLER_102_931 VPWR VGND sg13g2_decap_8
XFILLER_101_441 VPWR VGND sg13g2_decap_8
XFILLER_86_130 VPWR VGND sg13g2_decap_8
XFILLER_59_355 VPWR VGND sg13g2_decap_8
XFILLER_87_686 VPWR VGND sg13g2_decap_8
XFILLER_75_826 VPWR VGND sg13g2_decap_8
XFILLER_47_539 VPWR VGND sg13g2_decap_8
XFILLER_47_56 VPWR VGND sg13g2_decap_8
XFILLER_28_742 VPWR VGND sg13g2_decap_8
XFILLER_74_358 VPWR VGND sg13g2_decap_8
XFILLER_103_84 VPWR VGND sg13g2_decap_8
XFILLER_42_200 VPWR VGND sg13g2_decap_8
XFILLER_15_403 VPWR VGND sg13g2_decap_8
XFILLER_16_959 VPWR VGND sg13g2_decap_8
XFILLER_27_263 VPWR VGND sg13g2_decap_8
XFILLER_70_553 VPWR VGND sg13g2_decap_8
XFILLER_43_756 VPWR VGND sg13g2_decap_8
XFILLER_63_77 VPWR VGND sg13g2_decap_8
XFILLER_42_277 VPWR VGND sg13g2_decap_8
XFILLER_24_970 VPWR VGND sg13g2_decap_8
XFILLER_30_406 VPWR VGND sg13g2_decap_8
XFILLER_8_28 VPWR VGND sg13g2_decap_8
XFILLER_10_130 VPWR VGND sg13g2_decap_8
XFILLER_7_613 VPWR VGND sg13g2_decap_8
XFILLER_6_112 VPWR VGND sg13g2_decap_8
XFILLER_11_686 VPWR VGND sg13g2_decap_8
XFILLER_12_81 VPWR VGND sg13g2_decap_8
XFILLER_98_907 VPWR VGND sg13g2_decap_8
XFILLER_6_189 VPWR VGND sg13g2_decap_8
XFILLER_97_406 VPWR VGND sg13g2_decap_8
XFILLER_2_340 VPWR VGND sg13g2_decap_8
XFILLER_105_791 VPWR VGND sg13g2_decap_8
XFILLER_88_74 VPWR VGND sg13g2_decap_8
XFILLER_3_896 VPWR VGND sg13g2_decap_8
XFILLER_78_664 VPWR VGND sg13g2_decap_8
XFILLER_66_804 VPWR VGND sg13g2_decap_8
XFILLER_26_7 VPWR VGND sg13g2_decap_8
XFILLER_93_656 VPWR VGND sg13g2_decap_8
XFILLER_92_133 VPWR VGND sg13g2_decap_8
XFILLER_77_196 VPWR VGND sg13g2_decap_8
XFILLER_65_336 VPWR VGND sg13g2_decap_8
XFILLER_19_742 VPWR VGND sg13g2_decap_8
XFILLER_38_539 VPWR VGND sg13g2_decap_8
XFILLER_46_550 VPWR VGND sg13g2_decap_8
XFILLER_18_252 VPWR VGND sg13g2_decap_8
XFILLER_22_907 VPWR VGND sg13g2_decap_8
XFILLER_34_767 VPWR VGND sg13g2_decap_8
XFILLER_61_564 VPWR VGND sg13g2_decap_8
XFILLER_15_970 VPWR VGND sg13g2_decap_8
XFILLER_21_406 VPWR VGND sg13g2_decap_8
XFILLER_33_266 VPWR VGND sg13g2_decap_8
XFILLER_105_1001 VPWR VGND sg13g2_decap_8
XFILLER_30_973 VPWR VGND sg13g2_decap_8
XFILLER_52_0 VPWR VGND sg13g2_decap_8
XFILLER_103_728 VPWR VGND sg13g2_decap_8
XFILLER_88_417 VPWR VGND sg13g2_decap_8
XFILLER_102_238 VPWR VGND sg13g2_decap_8
XFILLER_69_631 VPWR VGND sg13g2_decap_8
XFILLER_97_973 VPWR VGND sg13g2_decap_8
XFILLER_84_623 VPWR VGND sg13g2_decap_8
XFILLER_68_152 VPWR VGND sg13g2_decap_8
XFILLER_57_826 VPWR VGND sg13g2_decap_8
XFILLER_96_483 VPWR VGND sg13g2_decap_8
XFILLER_56_347 VPWR VGND sg13g2_decap_8
XFILLER_83_144 VPWR VGND sg13g2_decap_8
XFILLER_37_550 VPWR VGND sg13g2_decap_8
XFILLER_24_200 VPWR VGND sg13g2_decap_8
XFILLER_80_840 VPWR VGND sg13g2_decap_8
XFILLER_52_553 VPWR VGND sg13g2_decap_8
XFILLER_25_756 VPWR VGND sg13g2_decap_8
XFILLER_12_417 VPWR VGND sg13g2_decap_8
XFILLER_24_277 VPWR VGND sg13g2_decap_8
XFILLER_33_14 VPWR VGND sg13g2_decap_8
XFILLER_21_973 VPWR VGND sg13g2_decap_8
XFILLER_32_1028 VPWR VGND sg13g2_fill_1
XFILLER_20_494 VPWR VGND sg13g2_decap_8
XFILLER_4_616 VPWR VGND sg13g2_decap_8
XFILLER_106_511 VPWR VGND sg13g2_decap_8
XFILLER_3_126 VPWR VGND sg13g2_decap_8
XFILLER_106_588 VPWR VGND sg13g2_decap_8
XFILLER_79_417 VPWR VGND sg13g2_decap_8
XFILLER_0_833 VPWR VGND sg13g2_decap_8
XFILLER_88_984 VPWR VGND sg13g2_decap_8
XFILLER_59_152 VPWR VGND sg13g2_decap_8
XFILLER_58_77 VPWR VGND sg13g2_decap_8
XFILLER_48_826 VPWR VGND sg13g2_decap_8
XFILLER_87_483 VPWR VGND sg13g2_decap_8
XFILLER_75_623 VPWR VGND sg13g2_decap_8
XFILLER_47_336 VPWR VGND sg13g2_decap_8
XFILLER_74_155 VPWR VGND sg13g2_decap_8
XFILLER_74_21 VPWR VGND sg13g2_decap_8
XFILLER_90_648 VPWR VGND sg13g2_decap_8
XFILLER_15_200 VPWR VGND sg13g2_decap_8
XFILLER_71_851 VPWR VGND sg13g2_decap_8
XFILLER_43_553 VPWR VGND sg13g2_decap_8
XFILLER_16_756 VPWR VGND sg13g2_decap_8
XFILLER_70_350 VPWR VGND sg13g2_decap_8
XFILLER_15_277 VPWR VGND sg13g2_decap_8
XFILLER_30_203 VPWR VGND sg13g2_decap_8
XFILLER_90_53 VPWR VGND sg13g2_decap_8
XFILLER_8_966 VPWR VGND sg13g2_decap_8
XFILLER_7_410 VPWR VGND sg13g2_decap_8
XFILLER_11_483 VPWR VGND sg13g2_decap_8
XFILLER_12_984 VPWR VGND sg13g2_decap_8
XFILLER_23_91 VPWR VGND sg13g2_decap_8
XFILLER_7_487 VPWR VGND sg13g2_decap_8
XFILLER_99_84 VPWR VGND sg13g2_decap_8
XFILLER_98_704 VPWR VGND sg13g2_decap_8
XFILLER_97_203 VPWR VGND sg13g2_decap_8
XFILLER_3_693 VPWR VGND sg13g2_decap_8
XFILLER_94_910 VPWR VGND sg13g2_decap_8
XFILLER_79_984 VPWR VGND sg13g2_decap_8
XFILLER_78_461 VPWR VGND sg13g2_decap_8
XFILLER_66_601 VPWR VGND sg13g2_decap_8
XFILLER_24_4 VPWR VGND sg13g2_decap_8
XFILLER_38_336 VPWR VGND sg13g2_decap_8
XFILLER_39_837 VPWR VGND sg13g2_decap_8
XFILLER_94_987 VPWR VGND sg13g2_decap_8
XFILLER_93_453 VPWR VGND sg13g2_decap_8
XFILLER_66_678 VPWR VGND sg13g2_decap_8
XFILLER_65_133 VPWR VGND sg13g2_decap_8
XFILLER_81_648 VPWR VGND sg13g2_decap_8
XFILLER_0_1015 VPWR VGND sg13g2_decap_8
XFILLER_94_1022 VPWR VGND sg13g2_decap_8
XFILLER_80_147 VPWR VGND sg13g2_decap_8
XFILLER_62_840 VPWR VGND sg13g2_decap_8
XFILLER_0_84 VPWR VGND sg13g2_decap_8
XFILLER_61_361 VPWR VGND sg13g2_decap_8
XFILLER_21_203 VPWR VGND sg13g2_decap_8
XFILLER_22_704 VPWR VGND sg13g2_decap_8
XFILLER_34_564 VPWR VGND sg13g2_decap_8
XFILLER_30_770 VPWR VGND sg13g2_decap_8
XFILLER_103_525 VPWR VGND sg13g2_decap_8
XFILLER_88_214 VPWR VGND sg13g2_decap_8
XFILLER_97_770 VPWR VGND sg13g2_decap_8
XFILLER_85_910 VPWR VGND sg13g2_decap_8
XFILLER_28_14 VPWR VGND sg13g2_decap_8
XFILLER_96_280 VPWR VGND sg13g2_decap_8
XFILLER_84_420 VPWR VGND sg13g2_decap_8
XFILLER_57_623 VPWR VGND sg13g2_decap_8
XFILLER_85_987 VPWR VGND sg13g2_decap_8
XFILLER_56_144 VPWR VGND sg13g2_decap_8
XFILLER_29_347 VPWR VGND sg13g2_decap_8
XFILLER_84_497 VPWR VGND sg13g2_decap_8
XFILLER_72_637 VPWR VGND sg13g2_decap_8
XFILLER_71_158 VPWR VGND sg13g2_decap_8
XFILLER_53_840 VPWR VGND sg13g2_decap_8
XFILLER_52_350 VPWR VGND sg13g2_decap_8
XFILLER_44_46 VPWR VGND sg13g2_decap_8
XFILLER_25_553 VPWR VGND sg13g2_decap_8
XFILLER_12_214 VPWR VGND sg13g2_decap_8
XFILLER_100_63 VPWR VGND sg13g2_decap_8
XFILLER_40_567 VPWR VGND sg13g2_decap_8
XFILLER_21_770 VPWR VGND sg13g2_decap_8
XFILLER_60_67 VPWR VGND sg13g2_decap_8
XFILLER_5_914 VPWR VGND sg13g2_decap_8
XFILLER_20_291 VPWR VGND sg13g2_decap_8
XFILLER_5_18 VPWR VGND sg13g2_decap_8
XFILLER_4_413 VPWR VGND sg13g2_decap_8
XFILLER_69_21 VPWR VGND sg13g2_decap_8
XFILLER_106_385 VPWR VGND sg13g2_decap_8
XFILLER_79_214 VPWR VGND sg13g2_decap_8
XFILLER_0_630 VPWR VGND sg13g2_decap_8
XFILLER_95_718 VPWR VGND sg13g2_decap_8
XFILLER_94_217 VPWR VGND sg13g2_decap_8
XFILLER_76_921 VPWR VGND sg13g2_decap_8
XFILLER_88_781 VPWR VGND sg13g2_decap_8
XFILLER_87_280 VPWR VGND sg13g2_decap_8
XFILLER_85_42 VPWR VGND sg13g2_decap_8
XFILLER_75_420 VPWR VGND sg13g2_decap_8
XFILLER_48_623 VPWR VGND sg13g2_decap_8
XFILLER_47_133 VPWR VGND sg13g2_decap_8
XFILLER_91_924 VPWR VGND sg13g2_decap_8
XFILLER_78_1028 VPWR VGND sg13g2_fill_1
XFILLER_76_998 VPWR VGND sg13g2_decap_8
XFILLER_75_497 VPWR VGND sg13g2_decap_8
XFILLER_63_637 VPWR VGND sg13g2_decap_8
XFILLER_90_445 VPWR VGND sg13g2_decap_8
XFILLER_62_147 VPWR VGND sg13g2_decap_8
XFILLER_44_851 VPWR VGND sg13g2_decap_8
XFILLER_18_91 VPWR VGND sg13g2_decap_8
XFILLER_43_350 VPWR VGND sg13g2_decap_8
XFILLER_16_553 VPWR VGND sg13g2_decap_8
XFILLER_15_1012 VPWR VGND sg13g2_decap_8
XFILLER_31_567 VPWR VGND sg13g2_decap_8
XFILLER_12_781 VPWR VGND sg13g2_decap_8
XFILLER_102_1015 VPWR VGND sg13g2_decap_8
XFILLER_8_763 VPWR VGND sg13g2_decap_8
XFILLER_11_280 VPWR VGND sg13g2_decap_8
XFILLER_7_284 VPWR VGND sg13g2_decap_8
XFILLER_98_501 VPWR VGND sg13g2_decap_8
XFILLER_4_980 VPWR VGND sg13g2_decap_8
XFILLER_3_490 VPWR VGND sg13g2_decap_8
XFILLER_98_578 VPWR VGND sg13g2_decap_8
XFILLER_86_718 VPWR VGND sg13g2_decap_8
XFILLER_85_217 VPWR VGND sg13g2_decap_8
XFILLER_67_910 VPWR VGND sg13g2_decap_8
XFILLER_100_539 VPWR VGND sg13g2_decap_8
XFILLER_79_781 VPWR VGND sg13g2_decap_8
XFILLER_22_1005 VPWR VGND sg13g2_decap_8
XFILLER_39_634 VPWR VGND sg13g2_decap_8
XFILLER_67_987 VPWR VGND sg13g2_decap_8
XFILLER_38_133 VPWR VGND sg13g2_decap_8
XFILLER_94_784 VPWR VGND sg13g2_decap_8
XFILLER_93_250 VPWR VGND sg13g2_decap_8
XFILLER_82_924 VPWR VGND sg13g2_decap_8
XFILLER_66_475 VPWR VGND sg13g2_decap_8
XFILLER_81_445 VPWR VGND sg13g2_decap_8
XFILLER_54_648 VPWR VGND sg13g2_decap_8
XFILLER_53_147 VPWR VGND sg13g2_decap_8
XFILLER_35_840 VPWR VGND sg13g2_decap_8
XFILLER_22_501 VPWR VGND sg13g2_decap_8
XFILLER_34_361 VPWR VGND sg13g2_decap_8
XFILLER_50_854 VPWR VGND sg13g2_decap_8
XFILLER_10_718 VPWR VGND sg13g2_decap_8
XFILLER_14_49 VPWR VGND sg13g2_decap_8
XFILLER_22_578 VPWR VGND sg13g2_decap_8
XFILLER_104_812 VPWR VGND sg13g2_decap_8
XFILLER_2_928 VPWR VGND sg13g2_decap_8
XFILLER_103_322 VPWR VGND sg13g2_decap_8
XFILLER_1_427 VPWR VGND sg13g2_decap_8
XFILLER_104_889 VPWR VGND sg13g2_decap_8
XFILLER_89_567 VPWR VGND sg13g2_decap_8
XFILLER_77_707 VPWR VGND sg13g2_decap_8
XFILLER_58_910 VPWR VGND sg13g2_decap_8
XFILLER_39_46 VPWR VGND sg13g2_decap_8
XFILLER_103_399 VPWR VGND sg13g2_decap_8
XFILLER_76_228 VPWR VGND sg13g2_decap_8
XFILLER_57_420 VPWR VGND sg13g2_decap_8
XFILLER_58_987 VPWR VGND sg13g2_decap_8
XFILLER_29_144 VPWR VGND sg13g2_decap_8
XFILLER_85_784 VPWR VGND sg13g2_decap_8
XFILLER_73_935 VPWR VGND sg13g2_decap_8
XFILLER_57_497 VPWR VGND sg13g2_decap_8
XFILLER_45_637 VPWR VGND sg13g2_decap_8
XFILLER_84_294 VPWR VGND sg13g2_decap_8
XFILLER_72_434 VPWR VGND sg13g2_decap_8
XFILLER_55_56 VPWR VGND sg13g2_decap_8
XFILLER_26_840 VPWR VGND sg13g2_decap_8
XFILLER_44_158 VPWR VGND sg13g2_decap_8
XFILLER_25_350 VPWR VGND sg13g2_decap_8
XFILLER_38_1001 VPWR VGND sg13g2_decap_8
XFILLER_71_11 VPWR VGND sg13g2_decap_8
XFILLER_41_854 VPWR VGND sg13g2_decap_8
XFILLER_13_567 VPWR VGND sg13g2_decap_8
XFILLER_71_88 VPWR VGND sg13g2_decap_8
XFILLER_40_364 VPWR VGND sg13g2_decap_8
XFILLER_5_711 VPWR VGND sg13g2_decap_8
XFILLER_4_210 VPWR VGND sg13g2_decap_8
XFILLER_5_788 VPWR VGND sg13g2_decap_8
XFILLER_106_182 VPWR VGND sg13g2_decap_8
XFILLER_4_287 VPWR VGND sg13g2_decap_8
XFILLER_20_81 VPWR VGND sg13g2_decap_8
XFILLER_95_515 VPWR VGND sg13g2_decap_8
XFILLER_96_63 VPWR VGND sg13g2_decap_8
XFILLER_67_217 VPWR VGND sg13g2_decap_8
XFILLER_49_921 VPWR VGND sg13g2_decap_8
XFILLER_48_420 VPWR VGND sg13g2_decap_8
XFILLER_1_994 VPWR VGND sg13g2_decap_8
XFILLER_91_721 VPWR VGND sg13g2_decap_8
XFILLER_76_795 VPWR VGND sg13g2_decap_8
XFILLER_64_935 VPWR VGND sg13g2_decap_8
XFILLER_49_998 VPWR VGND sg13g2_decap_8
XFILLER_36_637 VPWR VGND sg13g2_decap_8
XFILLER_75_294 VPWR VGND sg13g2_decap_8
XFILLER_63_434 VPWR VGND sg13g2_decap_8
XFILLER_48_497 VPWR VGND sg13g2_decap_8
XFILLER_35_147 VPWR VGND sg13g2_decap_8
XFILLER_91_798 VPWR VGND sg13g2_decap_8
XFILLER_90_242 VPWR VGND sg13g2_decap_8
XFILLER_16_350 VPWR VGND sg13g2_decap_8
XFILLER_17_851 VPWR VGND sg13g2_decap_8
XFILLER_32_865 VPWR VGND sg13g2_decap_8
XFILLER_31_364 VPWR VGND sg13g2_decap_8
XFILLER_8_560 VPWR VGND sg13g2_decap_8
XFILLER_105_609 VPWR VGND sg13g2_decap_8
XFILLER_104_119 VPWR VGND sg13g2_decap_8
XFILLER_99_854 VPWR VGND sg13g2_decap_8
XFILLER_98_375 VPWR VGND sg13g2_decap_8
XFILLER_86_515 VPWR VGND sg13g2_decap_8
XFILLER_101_826 VPWR VGND sg13g2_decap_8
XFILLER_58_217 VPWR VGND sg13g2_decap_8
XFILLER_100_336 VPWR VGND sg13g2_decap_8
XFILLER_39_431 VPWR VGND sg13g2_decap_8
XFILLER_94_581 VPWR VGND sg13g2_decap_8
XFILLER_82_721 VPWR VGND sg13g2_decap_8
XFILLER_67_784 VPWR VGND sg13g2_decap_8
XFILLER_66_272 VPWR VGND sg13g2_decap_8
XFILLER_55_924 VPWR VGND sg13g2_decap_8
XFILLER_54_445 VPWR VGND sg13g2_decap_8
XFILLER_27_648 VPWR VGND sg13g2_decap_8
XFILLER_82_798 VPWR VGND sg13g2_decap_8
XFILLER_81_242 VPWR VGND sg13g2_decap_8
XFILLER_70_938 VPWR VGND sg13g2_decap_8
XFILLER_26_147 VPWR VGND sg13g2_decap_8
XFILLER_50_651 VPWR VGND sg13g2_decap_8
XFILLER_23_854 VPWR VGND sg13g2_decap_8
XFILLER_10_515 VPWR VGND sg13g2_decap_8
XFILLER_22_375 VPWR VGND sg13g2_decap_8
XFILLER_41_14 VPWR VGND sg13g2_decap_8
XFILLER_68_1027 VPWR VGND sg13g2_fill_2
XFILLER_2_725 VPWR VGND sg13g2_decap_8
XFILLER_1_224 VPWR VGND sg13g2_decap_8
XFILLER_89_364 VPWR VGND sg13g2_decap_8
XFILLER_77_504 VPWR VGND sg13g2_decap_8
XFILLER_104_686 VPWR VGND sg13g2_decap_8
XFILLER_66_11 VPWR VGND sg13g2_decap_8
XFILLER_49_228 VPWR VGND sg13g2_decap_8
XFILLER_106_84 VPWR VGND sg13g2_decap_8
XFILLER_103_196 VPWR VGND sg13g2_decap_8
XFILLER_92_518 VPWR VGND sg13g2_decap_8
XFILLER_85_581 VPWR VGND sg13g2_decap_8
XFILLER_66_55 VPWR VGND sg13g2_decap_8
XFILLER_58_784 VPWR VGND sg13g2_decap_8
XFILLER_46_935 VPWR VGND sg13g2_decap_8
XFILLER_73_732 VPWR VGND sg13g2_decap_8
XFILLER_72_231 VPWR VGND sg13g2_decap_8
XFILLER_57_294 VPWR VGND sg13g2_decap_8
XFILLER_45_434 VPWR VGND sg13g2_decap_8
XFILLER_18_637 VPWR VGND sg13g2_decap_8
XFILLER_82_21 VPWR VGND sg13g2_decap_8
XFILLER_17_158 VPWR VGND sg13g2_decap_8
XFILLER_61_949 VPWR VGND sg13g2_decap_8
XFILLER_82_98 VPWR VGND sg13g2_decap_8
XFILLER_60_459 VPWR VGND sg13g2_decap_8
XFILLER_41_651 VPWR VGND sg13g2_decap_8
XFILLER_14_854 VPWR VGND sg13g2_decap_8
XFILLER_13_364 VPWR VGND sg13g2_decap_8
XFILLER_15_81 VPWR VGND sg13g2_decap_8
XFILLER_40_161 VPWR VGND sg13g2_decap_8
XFILLER_9_357 VPWR VGND sg13g2_decap_8
XFILLER_12_1026 VPWR VGND sg13g2_fill_2
XFILLER_31_91 VPWR VGND sg13g2_decap_8
XFILLER_5_585 VPWR VGND sg13g2_decap_8
XFILLER_95_312 VPWR VGND sg13g2_decap_8
XFILLER_68_537 VPWR VGND sg13g2_decap_8
XFILLER_96_868 VPWR VGND sg13g2_decap_8
XFILLER_1_791 VPWR VGND sg13g2_decap_8
XFILLER_95_389 VPWR VGND sg13g2_decap_8
XFILLER_83_529 VPWR VGND sg13g2_decap_8
XFILLER_49_795 VPWR VGND sg13g2_decap_8
XFILLER_37_935 VPWR VGND sg13g2_decap_8
XFILLER_76_592 VPWR VGND sg13g2_decap_8
XFILLER_64_732 VPWR VGND sg13g2_decap_8
XFILLER_48_294 VPWR VGND sg13g2_decap_8
XFILLER_36_434 VPWR VGND sg13g2_decap_8
XFILLER_63_231 VPWR VGND sg13g2_decap_8
XFILLER_91_595 VPWR VGND sg13g2_decap_8
XFILLER_52_938 VPWR VGND sg13g2_decap_8
XFILLER_51_459 VPWR VGND sg13g2_decap_8
XFILLER_20_802 VPWR VGND sg13g2_decap_8
XFILLER_31_161 VPWR VGND sg13g2_decap_8
XFILLER_32_662 VPWR VGND sg13g2_decap_8
XFILLER_82_0 VPWR VGND sg13g2_decap_8
XFILLER_20_879 VPWR VGND sg13g2_decap_8
XFILLER_11_28 VPWR VGND sg13g2_decap_8
XFILLER_105_406 VPWR VGND sg13g2_decap_8
XFILLER_99_651 VPWR VGND sg13g2_decap_8
XFILLER_28_1022 VPWR VGND sg13g2_decap_8
XFILLER_101_623 VPWR VGND sg13g2_decap_8
XFILLER_98_172 VPWR VGND sg13g2_decap_8
XFILLER_86_312 VPWR VGND sg13g2_decap_8
XFILLER_59_537 VPWR VGND sg13g2_decap_8
XFILLER_100_133 VPWR VGND sg13g2_decap_8
XFILLER_87_868 VPWR VGND sg13g2_decap_8
XFILLER_86_389 VPWR VGND sg13g2_decap_8
XFILLER_28_924 VPWR VGND sg13g2_decap_8
XFILLER_67_581 VPWR VGND sg13g2_decap_8
XFILLER_55_721 VPWR VGND sg13g2_decap_8
XFILLER_36_14 VPWR VGND sg13g2_decap_8
XFILLER_54_242 VPWR VGND sg13g2_decap_8
XFILLER_27_445 VPWR VGND sg13g2_decap_8
XFILLER_82_595 VPWR VGND sg13g2_decap_8
XFILLER_70_735 VPWR VGND sg13g2_decap_8
XFILLER_55_798 VPWR VGND sg13g2_decap_8
XFILLER_43_938 VPWR VGND sg13g2_decap_8
XFILLER_42_459 VPWR VGND sg13g2_decap_8
XFILLER_23_651 VPWR VGND sg13g2_decap_8
XFILLER_52_35 VPWR VGND sg13g2_decap_8
XFILLER_35_1015 VPWR VGND sg13g2_decap_8
XFILLER_10_312 VPWR VGND sg13g2_decap_8
XFILLER_22_172 VPWR VGND sg13g2_decap_8
XFILLER_11_868 VPWR VGND sg13g2_decap_8
XFILLER_10_389 VPWR VGND sg13g2_decap_8
XFILLER_2_522 VPWR VGND sg13g2_decap_8
XFILLER_105_973 VPWR VGND sg13g2_decap_8
XFILLER_77_21 VPWR VGND sg13g2_decap_8
XFILLER_104_483 VPWR VGND sg13g2_decap_8
XFILLER_89_161 VPWR VGND sg13g2_decap_8
XFILLER_78_846 VPWR VGND sg13g2_decap_8
XFILLER_77_301 VPWR VGND sg13g2_decap_8
XFILLER_2_599 VPWR VGND sg13g2_decap_8
XFILLER_42_1019 VPWR VGND sg13g2_decap_8
XFILLER_93_838 VPWR VGND sg13g2_decap_8
XFILLER_92_315 VPWR VGND sg13g2_decap_8
XFILLER_77_378 VPWR VGND sg13g2_decap_8
XFILLER_77_98 VPWR VGND sg13g2_decap_8
XFILLER_65_518 VPWR VGND sg13g2_decap_8
XFILLER_19_924 VPWR VGND sg13g2_decap_8
XFILLER_58_581 VPWR VGND sg13g2_decap_8
XFILLER_46_732 VPWR VGND sg13g2_decap_8
XFILLER_18_434 VPWR VGND sg13g2_decap_8
XFILLER_93_75 VPWR VGND sg13g2_decap_8
XFILLER_45_231 VPWR VGND sg13g2_decap_8
XFILLER_61_746 VPWR VGND sg13g2_decap_8
Xheichips25_example_large_29 VPWR VGND uio_oe[4] sg13g2_tielo
XFILLER_34_949 VPWR VGND sg13g2_decap_8
XFILLER_60_256 VPWR VGND sg13g2_decap_8
XFILLER_26_91 VPWR VGND sg13g2_decap_8
XFILLER_33_448 VPWR VGND sg13g2_decap_8
XFILLER_14_651 VPWR VGND sg13g2_decap_8
XFILLER_20_109 VPWR VGND sg13g2_decap_8
XFILLER_13_161 VPWR VGND sg13g2_decap_8
XFILLER_9_154 VPWR VGND sg13g2_decap_8
XFILLER_6_861 VPWR VGND sg13g2_decap_8
XFILLER_54_4 VPWR VGND sg13g2_decap_8
XFILLER_5_382 VPWR VGND sg13g2_decap_8
XFILLER_69_813 VPWR VGND sg13g2_decap_8
XFILLER_96_665 VPWR VGND sg13g2_decap_8
XFILLER_84_805 VPWR VGND sg13g2_decap_8
XFILLER_68_334 VPWR VGND sg13g2_decap_8
XFILLER_56_529 VPWR VGND sg13g2_decap_8
XFILLER_3_84 VPWR VGND sg13g2_decap_8
XFILLER_95_186 VPWR VGND sg13g2_decap_8
XFILLER_83_326 VPWR VGND sg13g2_decap_8
XFILLER_49_592 VPWR VGND sg13g2_decap_8
XFILLER_37_732 VPWR VGND sg13g2_decap_8
XFILLER_58_1015 VPWR VGND sg13g2_decap_8
XFILLER_36_231 VPWR VGND sg13g2_decap_8
XFILLER_92_882 VPWR VGND sg13g2_decap_8
XFILLER_52_735 VPWR VGND sg13g2_decap_8
XFILLER_25_938 VPWR VGND sg13g2_decap_8
XFILLER_91_392 VPWR VGND sg13g2_decap_8
XFILLER_24_459 VPWR VGND sg13g2_decap_8
XFILLER_51_256 VPWR VGND sg13g2_decap_8
XFILLER_20_676 VPWR VGND sg13g2_decap_8
XFILLER_3_308 VPWR VGND sg13g2_decap_8
XFILLER_105_203 VPWR VGND sg13g2_decap_8
XFILLER_65_1008 VPWR VGND sg13g2_decap_8
XFILLER_102_910 VPWR VGND sg13g2_decap_8
XFILLER_101_420 VPWR VGND sg13g2_decap_8
XFILLER_75_805 VPWR VGND sg13g2_decap_8
XFILLER_59_334 VPWR VGND sg13g2_decap_8
XFILLER_102_987 VPWR VGND sg13g2_decap_8
XFILLER_87_665 VPWR VGND sg13g2_decap_8
XFILLER_47_518 VPWR VGND sg13g2_decap_8
XFILLER_47_35 VPWR VGND sg13g2_decap_8
XFILLER_101_497 VPWR VGND sg13g2_decap_8
XFILLER_86_186 VPWR VGND sg13g2_decap_8
XFILLER_74_337 VPWR VGND sg13g2_decap_8
XFILLER_28_721 VPWR VGND sg13g2_decap_8
XFILLER_27_242 VPWR VGND sg13g2_decap_8
XFILLER_103_63 VPWR VGND sg13g2_decap_8
XFILLER_83_893 VPWR VGND sg13g2_decap_8
XFILLER_55_595 VPWR VGND sg13g2_decap_8
XFILLER_43_735 VPWR VGND sg13g2_decap_8
XFILLER_16_938 VPWR VGND sg13g2_decap_8
XFILLER_28_798 VPWR VGND sg13g2_decap_8
XFILLER_82_392 VPWR VGND sg13g2_decap_8
XFILLER_70_532 VPWR VGND sg13g2_decap_8
XFILLER_63_56 VPWR VGND sg13g2_decap_8
XFILLER_15_459 VPWR VGND sg13g2_decap_8
XFILLER_42_256 VPWR VGND sg13g2_decap_8
XFILLER_11_665 VPWR VGND sg13g2_decap_8
XFILLER_10_186 VPWR VGND sg13g2_decap_8
XFILLER_7_669 VPWR VGND sg13g2_decap_8
XFILLER_6_168 VPWR VGND sg13g2_decap_8
XFILLER_12_60 VPWR VGND sg13g2_decap_8
XFILLER_88_53 VPWR VGND sg13g2_decap_8
XFILLER_105_770 VPWR VGND sg13g2_decap_8
XFILLER_3_875 VPWR VGND sg13g2_decap_8
XFILLER_104_280 VPWR VGND sg13g2_decap_8
XFILLER_78_643 VPWR VGND sg13g2_decap_8
XFILLER_2_396 VPWR VGND sg13g2_decap_8
XFILLER_38_518 VPWR VGND sg13g2_decap_8
XFILLER_93_635 VPWR VGND sg13g2_decap_8
XFILLER_92_112 VPWR VGND sg13g2_decap_8
XFILLER_77_175 VPWR VGND sg13g2_decap_8
XFILLER_65_315 VPWR VGND sg13g2_decap_8
XFILLER_19_7 VPWR VGND sg13g2_decap_8
XFILLER_19_721 VPWR VGND sg13g2_decap_8
XFILLER_18_231 VPWR VGND sg13g2_decap_8
XFILLER_92_189 VPWR VGND sg13g2_decap_8
XFILLER_80_329 VPWR VGND sg13g2_decap_8
XFILLER_19_798 VPWR VGND sg13g2_decap_8
XFILLER_61_543 VPWR VGND sg13g2_decap_8
XFILLER_33_245 VPWR VGND sg13g2_decap_8
XFILLER_34_746 VPWR VGND sg13g2_decap_8
XFILLER_30_952 VPWR VGND sg13g2_decap_8
XFILLER_88_1019 VPWR VGND sg13g2_decap_8
XFILLER_103_707 VPWR VGND sg13g2_decap_8
XFILLER_45_0 VPWR VGND sg13g2_decap_8
XFILLER_102_217 VPWR VGND sg13g2_decap_8
XFILLER_69_610 VPWR VGND sg13g2_decap_8
XFILLER_97_952 VPWR VGND sg13g2_decap_8
XFILLER_68_131 VPWR VGND sg13g2_decap_8
XFILLER_96_462 VPWR VGND sg13g2_decap_8
XFILLER_84_602 VPWR VGND sg13g2_decap_8
XFILLER_69_687 VPWR VGND sg13g2_decap_8
XFILLER_57_805 VPWR VGND sg13g2_decap_8
XFILLER_83_123 VPWR VGND sg13g2_decap_8
XFILLER_56_326 VPWR VGND sg13g2_decap_8
XFILLER_29_529 VPWR VGND sg13g2_decap_8
XFILLER_84_679 VPWR VGND sg13g2_decap_8
XFILLER_72_819 VPWR VGND sg13g2_decap_8
XFILLER_65_882 VPWR VGND sg13g2_decap_8
XFILLER_25_735 VPWR VGND sg13g2_decap_8
XFILLER_52_532 VPWR VGND sg13g2_decap_8
XFILLER_80_896 VPWR VGND sg13g2_decap_8
XFILLER_24_256 VPWR VGND sg13g2_decap_8
XFILLER_71_1012 VPWR VGND sg13g2_decap_8
XFILLER_40_749 VPWR VGND sg13g2_decap_8
XFILLER_21_952 VPWR VGND sg13g2_decap_8
XFILLER_20_473 VPWR VGND sg13g2_decap_8
XFILLER_3_105 VPWR VGND sg13g2_decap_8
XFILLER_106_567 VPWR VGND sg13g2_decap_8
XFILLER_0_812 VPWR VGND sg13g2_decap_8
XFILLER_88_963 VPWR VGND sg13g2_decap_8
XFILLER_59_120 VPWR VGND sg13g2_decap_8
XFILLER_58_56 VPWR VGND sg13g2_decap_8
XFILLER_87_462 VPWR VGND sg13g2_decap_8
XFILLER_75_602 VPWR VGND sg13g2_decap_8
XFILLER_48_805 VPWR VGND sg13g2_decap_8
XFILLER_0_889 VPWR VGND sg13g2_decap_8
XFILLER_102_784 VPWR VGND sg13g2_decap_8
XFILLER_47_315 VPWR VGND sg13g2_decap_8
XFILLER_101_294 VPWR VGND sg13g2_decap_8
XFILLER_75_679 VPWR VGND sg13g2_decap_8
XFILLER_74_134 VPWR VGND sg13g2_decap_8
XFILLER_63_819 VPWR VGND sg13g2_decap_8
XFILLER_90_627 VPWR VGND sg13g2_decap_8
XFILLER_62_329 VPWR VGND sg13g2_decap_8
XFILLER_56_893 VPWR VGND sg13g2_decap_8
XFILLER_83_690 VPWR VGND sg13g2_decap_8
XFILLER_74_99 VPWR VGND sg13g2_decap_8
XFILLER_71_830 VPWR VGND sg13g2_decap_8
XFILLER_55_392 VPWR VGND sg13g2_decap_8
XFILLER_43_532 VPWR VGND sg13g2_decap_8
XFILLER_16_735 VPWR VGND sg13g2_decap_8
XFILLER_28_595 VPWR VGND sg13g2_decap_8
XFILLER_15_256 VPWR VGND sg13g2_decap_8
XFILLER_90_32 VPWR VGND sg13g2_decap_8
XFILLER_31_749 VPWR VGND sg13g2_decap_8
XFILLER_12_963 VPWR VGND sg13g2_decap_8
XFILLER_30_259 VPWR VGND sg13g2_decap_8
XFILLER_8_945 VPWR VGND sg13g2_decap_8
XFILLER_11_462 VPWR VGND sg13g2_decap_8
XFILLER_23_70 VPWR VGND sg13g2_decap_8
XFILLER_7_466 VPWR VGND sg13g2_decap_8
XFILLER_99_63 VPWR VGND sg13g2_decap_8
XFILLER_3_672 VPWR VGND sg13g2_decap_8
XFILLER_97_259 VPWR VGND sg13g2_decap_8
XFILLER_79_963 VPWR VGND sg13g2_decap_8
XFILLER_78_440 VPWR VGND sg13g2_decap_8
XFILLER_2_193 VPWR VGND sg13g2_decap_8
XFILLER_39_816 VPWR VGND sg13g2_decap_8
XFILLER_93_432 VPWR VGND sg13g2_decap_8
XFILLER_65_112 VPWR VGND sg13g2_decap_8
XFILLER_17_4 VPWR VGND sg13g2_decap_8
XFILLER_38_315 VPWR VGND sg13g2_decap_8
XFILLER_94_966 VPWR VGND sg13g2_decap_8
XFILLER_66_657 VPWR VGND sg13g2_decap_8
XFILLER_94_1001 VPWR VGND sg13g2_decap_8
XFILLER_81_627 VPWR VGND sg13g2_decap_8
XFILLER_65_189 VPWR VGND sg13g2_decap_8
XFILLER_53_329 VPWR VGND sg13g2_decap_8
XFILLER_47_882 VPWR VGND sg13g2_decap_8
XFILLER_80_126 VPWR VGND sg13g2_decap_8
XFILLER_0_63 VPWR VGND sg13g2_decap_8
XFILLER_19_595 VPWR VGND sg13g2_decap_8
XFILLER_34_543 VPWR VGND sg13g2_decap_8
XFILLER_61_340 VPWR VGND sg13g2_decap_8
XFILLER_62_896 VPWR VGND sg13g2_decap_8
XFILLER_21_259 VPWR VGND sg13g2_decap_8
XFILLER_103_504 VPWR VGND sg13g2_decap_8
XFILLER_1_609 VPWR VGND sg13g2_decap_8
XFILLER_89_749 VPWR VGND sg13g2_decap_8
XFILLER_0_119 VPWR VGND sg13g2_decap_8
XFILLER_57_602 VPWR VGND sg13g2_decap_8
XFILLER_69_484 VPWR VGND sg13g2_decap_8
XFILLER_29_326 VPWR VGND sg13g2_decap_8
XFILLER_85_966 VPWR VGND sg13g2_decap_8
XFILLER_57_679 VPWR VGND sg13g2_decap_8
XFILLER_56_123 VPWR VGND sg13g2_decap_8
XFILLER_45_819 VPWR VGND sg13g2_decap_8
XFILLER_84_476 VPWR VGND sg13g2_decap_8
XFILLER_72_616 VPWR VGND sg13g2_decap_8
XFILLER_38_882 VPWR VGND sg13g2_decap_8
XFILLER_71_137 VPWR VGND sg13g2_decap_8
XFILLER_44_25 VPWR VGND sg13g2_decap_8
XFILLER_25_532 VPWR VGND sg13g2_decap_8
XFILLER_80_693 VPWR VGND sg13g2_decap_8
XFILLER_53_896 VPWR VGND sg13g2_decap_8
XFILLER_13_749 VPWR VGND sg13g2_decap_8
XFILLER_100_42 VPWR VGND sg13g2_decap_8
XFILLER_40_546 VPWR VGND sg13g2_decap_8
XFILLER_60_46 VPWR VGND sg13g2_decap_8
XFILLER_20_270 VPWR VGND sg13g2_decap_8
XFILLER_106_364 VPWR VGND sg13g2_decap_8
XFILLER_4_469 VPWR VGND sg13g2_decap_8
XFILLER_69_99 VPWR VGND sg13g2_decap_8
XFILLER_88_760 VPWR VGND sg13g2_decap_8
XFILLER_76_900 VPWR VGND sg13g2_decap_8
XFILLER_48_602 VPWR VGND sg13g2_decap_8
XFILLER_102_581 VPWR VGND sg13g2_decap_8
XFILLER_85_21 VPWR VGND sg13g2_decap_8
XFILLER_47_112 VPWR VGND sg13g2_decap_8
XFILLER_0_686 VPWR VGND sg13g2_decap_8
XFILLER_91_903 VPWR VGND sg13g2_decap_8
XFILLER_78_1007 VPWR VGND sg13g2_decap_8
XFILLER_76_977 VPWR VGND sg13g2_decap_8
XFILLER_48_679 VPWR VGND sg13g2_decap_8
XFILLER_36_819 VPWR VGND sg13g2_decap_8
XFILLER_85_98 VPWR VGND sg13g2_decap_8
XFILLER_75_476 VPWR VGND sg13g2_decap_8
XFILLER_63_616 VPWR VGND sg13g2_decap_8
XFILLER_47_189 VPWR VGND sg13g2_decap_8
XFILLER_18_70 VPWR VGND sg13g2_decap_8
XFILLER_35_329 VPWR VGND sg13g2_decap_8
XFILLER_90_424 VPWR VGND sg13g2_decap_8
XFILLER_62_126 VPWR VGND sg13g2_decap_8
XFILLER_56_690 VPWR VGND sg13g2_decap_8
XFILLER_44_830 VPWR VGND sg13g2_decap_8
XFILLER_16_532 VPWR VGND sg13g2_decap_8
XFILLER_28_392 VPWR VGND sg13g2_decap_8
XFILLER_29_893 VPWR VGND sg13g2_decap_8
XFILLER_31_546 VPWR VGND sg13g2_decap_8
XFILLER_12_760 VPWR VGND sg13g2_decap_8
XFILLER_8_742 VPWR VGND sg13g2_decap_8
XFILLER_7_263 VPWR VGND sg13g2_decap_8
XFILLER_98_557 VPWR VGND sg13g2_decap_8
XFILLER_79_760 VPWR VGND sg13g2_decap_8
XFILLER_100_518 VPWR VGND sg13g2_decap_8
XFILLER_38_112 VPWR VGND sg13g2_decap_8
XFILLER_39_613 VPWR VGND sg13g2_decap_8
XFILLER_94_763 VPWR VGND sg13g2_decap_8
XFILLER_82_903 VPWR VGND sg13g2_decap_8
XFILLER_67_966 VPWR VGND sg13g2_decap_8
XFILLER_66_454 VPWR VGND sg13g2_decap_8
XFILLER_22_1028 VPWR VGND sg13g2_fill_1
XFILLER_54_627 VPWR VGND sg13g2_decap_8
XFILLER_26_329 VPWR VGND sg13g2_decap_8
XFILLER_81_424 VPWR VGND sg13g2_decap_8
XFILLER_53_126 VPWR VGND sg13g2_decap_8
XFILLER_19_392 VPWR VGND sg13g2_decap_8
XFILLER_38_189 VPWR VGND sg13g2_decap_8
XFILLER_34_340 VPWR VGND sg13g2_decap_8
XFILLER_90_991 VPWR VGND sg13g2_decap_8
XFILLER_62_693 VPWR VGND sg13g2_decap_8
XFILLER_50_833 VPWR VGND sg13g2_decap_8
XFILLER_35_896 VPWR VGND sg13g2_decap_8
XFILLER_14_28 VPWR VGND sg13g2_decap_8
XFILLER_22_557 VPWR VGND sg13g2_decap_8
XFILLER_2_907 VPWR VGND sg13g2_decap_8
XFILLER_30_49 VPWR VGND sg13g2_decap_8
XFILLER_1_406 VPWR VGND sg13g2_decap_8
XFILLER_103_301 VPWR VGND sg13g2_decap_8
XFILLER_89_546 VPWR VGND sg13g2_decap_8
XFILLER_104_868 VPWR VGND sg13g2_decap_8
XFILLER_76_207 VPWR VGND sg13g2_decap_8
XFILLER_39_25 VPWR VGND sg13g2_decap_8
XFILLER_103_378 VPWR VGND sg13g2_decap_8
XFILLER_85_763 VPWR VGND sg13g2_decap_8
XFILLER_69_281 VPWR VGND sg13g2_decap_8
XFILLER_58_966 VPWR VGND sg13g2_decap_8
XFILLER_29_123 VPWR VGND sg13g2_decap_8
XFILLER_84_273 VPWR VGND sg13g2_decap_8
XFILLER_73_914 VPWR VGND sg13g2_decap_8
XFILLER_72_413 VPWR VGND sg13g2_decap_8
XFILLER_57_476 VPWR VGND sg13g2_decap_8
XFILLER_55_35 VPWR VGND sg13g2_decap_8
XFILLER_45_616 VPWR VGND sg13g2_decap_8
XFILLER_18_819 VPWR VGND sg13g2_decap_8
XFILLER_44_137 VPWR VGND sg13g2_decap_8
XFILLER_81_991 VPWR VGND sg13g2_decap_8
XFILLER_53_693 VPWR VGND sg13g2_decap_8
XFILLER_41_833 VPWR VGND sg13g2_decap_8
XFILLER_26_896 VPWR VGND sg13g2_decap_8
XFILLER_80_490 VPWR VGND sg13g2_decap_8
XFILLER_13_546 VPWR VGND sg13g2_decap_8
XFILLER_40_343 VPWR VGND sg13g2_decap_8
XFILLER_71_67 VPWR VGND sg13g2_decap_8
XFILLER_9_539 VPWR VGND sg13g2_decap_8
XFILLER_84_1022 VPWR VGND sg13g2_decap_8
XFILLER_5_767 VPWR VGND sg13g2_decap_8
XFILLER_4_266 VPWR VGND sg13g2_decap_8
XFILLER_20_60 VPWR VGND sg13g2_decap_8
XFILLER_106_161 VPWR VGND sg13g2_decap_8
XFILLER_96_42 VPWR VGND sg13g2_decap_8
XFILLER_68_719 VPWR VGND sg13g2_decap_8
XFILLER_49_900 VPWR VGND sg13g2_decap_8
XFILLER_1_973 VPWR VGND sg13g2_decap_8
XFILLER_49_977 VPWR VGND sg13g2_decap_8
XFILLER_0_483 VPWR VGND sg13g2_decap_8
XFILLER_91_700 VPWR VGND sg13g2_decap_8
XFILLER_76_774 VPWR VGND sg13g2_decap_8
XFILLER_75_273 VPWR VGND sg13g2_decap_8
XFILLER_64_914 VPWR VGND sg13g2_decap_8
XFILLER_63_413 VPWR VGND sg13g2_decap_8
XFILLER_48_476 VPWR VGND sg13g2_decap_8
XFILLER_36_616 VPWR VGND sg13g2_decap_8
XFILLER_90_221 VPWR VGND sg13g2_decap_8
XFILLER_17_830 VPWR VGND sg13g2_decap_8
XFILLER_29_690 VPWR VGND sg13g2_decap_8
XFILLER_35_126 VPWR VGND sg13g2_decap_8
XFILLER_91_777 VPWR VGND sg13g2_decap_8
XFILLER_91_1015 VPWR VGND sg13g2_decap_8
XFILLER_90_298 VPWR VGND sg13g2_decap_8
XFILLER_72_980 VPWR VGND sg13g2_decap_8
XFILLER_31_343 VPWR VGND sg13g2_decap_8
XFILLER_32_844 VPWR VGND sg13g2_decap_8
XFILLER_6_84 VPWR VGND sg13g2_decap_8
XFILLER_99_833 VPWR VGND sg13g2_decap_8
XFILLER_101_805 VPWR VGND sg13g2_decap_8
XFILLER_98_354 VPWR VGND sg13g2_decap_8
XFILLER_59_719 VPWR VGND sg13g2_decap_8
XFILLER_100_315 VPWR VGND sg13g2_decap_8
XFILLER_39_410 VPWR VGND sg13g2_decap_8
XFILLER_6_1022 VPWR VGND sg13g2_decap_8
XFILLER_94_560 VPWR VGND sg13g2_decap_8
XFILLER_82_700 VPWR VGND sg13g2_decap_8
XFILLER_67_763 VPWR VGND sg13g2_decap_8
XFILLER_66_251 VPWR VGND sg13g2_decap_8
XFILLER_55_903 VPWR VGND sg13g2_decap_8
XFILLER_27_627 VPWR VGND sg13g2_decap_8
XFILLER_39_487 VPWR VGND sg13g2_decap_8
XFILLER_81_221 VPWR VGND sg13g2_decap_8
XFILLER_54_424 VPWR VGND sg13g2_decap_8
XFILLER_26_126 VPWR VGND sg13g2_decap_8
XFILLER_82_777 VPWR VGND sg13g2_decap_8
XFILLER_70_917 VPWR VGND sg13g2_decap_8
XFILLER_81_298 VPWR VGND sg13g2_decap_8
XFILLER_63_980 VPWR VGND sg13g2_decap_8
XFILLER_23_833 VPWR VGND sg13g2_decap_8
XFILLER_25_49 VPWR VGND sg13g2_decap_8
XFILLER_35_693 VPWR VGND sg13g2_decap_8
XFILLER_62_490 VPWR VGND sg13g2_decap_8
XFILLER_50_630 VPWR VGND sg13g2_decap_8
XFILLER_22_354 VPWR VGND sg13g2_decap_8
XFILLER_68_1006 VPWR VGND sg13g2_decap_8
XFILLER_2_704 VPWR VGND sg13g2_decap_8
XFILLER_1_203 VPWR VGND sg13g2_decap_8
XFILLER_104_665 VPWR VGND sg13g2_decap_8
XFILLER_89_343 VPWR VGND sg13g2_decap_8
XFILLER_106_63 VPWR VGND sg13g2_decap_8
XFILLER_103_175 VPWR VGND sg13g2_decap_8
XFILLER_49_207 VPWR VGND sg13g2_decap_8
XFILLER_66_34 VPWR VGND sg13g2_decap_8
XFILLER_100_882 VPWR VGND sg13g2_decap_8
XFILLER_85_560 VPWR VGND sg13g2_decap_8
XFILLER_73_711 VPWR VGND sg13g2_decap_8
XFILLER_58_763 VPWR VGND sg13g2_decap_8
XFILLER_46_914 VPWR VGND sg13g2_decap_8
XFILLER_18_616 VPWR VGND sg13g2_decap_8
XFILLER_72_210 VPWR VGND sg13g2_decap_8
XFILLER_57_273 VPWR VGND sg13g2_decap_8
XFILLER_45_413 VPWR VGND sg13g2_decap_8
XFILLER_17_137 VPWR VGND sg13g2_decap_8
XFILLER_73_788 VPWR VGND sg13g2_decap_8
XFILLER_61_928 VPWR VGND sg13g2_decap_8
XFILLER_72_287 VPWR VGND sg13g2_decap_8
XFILLER_60_438 VPWR VGND sg13g2_decap_8
XFILLER_54_991 VPWR VGND sg13g2_decap_8
XFILLER_14_833 VPWR VGND sg13g2_decap_8
XFILLER_26_693 VPWR VGND sg13g2_decap_8
XFILLER_82_77 VPWR VGND sg13g2_decap_8
XFILLER_53_490 VPWR VGND sg13g2_decap_8
XFILLER_41_630 VPWR VGND sg13g2_decap_8
XFILLER_13_343 VPWR VGND sg13g2_decap_8
XFILLER_15_60 VPWR VGND sg13g2_decap_8
XFILLER_40_140 VPWR VGND sg13g2_decap_8
XFILLER_9_336 VPWR VGND sg13g2_decap_8
XFILLER_12_1005 VPWR VGND sg13g2_decap_8
XFILLER_31_70 VPWR VGND sg13g2_decap_8
XFILLER_5_564 VPWR VGND sg13g2_decap_8
XFILLER_96_847 VPWR VGND sg13g2_decap_8
XFILLER_68_516 VPWR VGND sg13g2_decap_8
XFILLER_1_770 VPWR VGND sg13g2_decap_8
XFILLER_0_280 VPWR VGND sg13g2_decap_8
XFILLER_95_368 VPWR VGND sg13g2_decap_8
XFILLER_83_508 VPWR VGND sg13g2_decap_8
XFILLER_76_571 VPWR VGND sg13g2_decap_8
XFILLER_64_711 VPWR VGND sg13g2_decap_8
XFILLER_49_774 VPWR VGND sg13g2_decap_8
XFILLER_37_914 VPWR VGND sg13g2_decap_8
XFILLER_63_210 VPWR VGND sg13g2_decap_8
XFILLER_48_273 VPWR VGND sg13g2_decap_8
XFILLER_36_413 VPWR VGND sg13g2_decap_8
XFILLER_64_788 VPWR VGND sg13g2_decap_8
XFILLER_52_917 VPWR VGND sg13g2_decap_8
XFILLER_91_574 VPWR VGND sg13g2_decap_8
XFILLER_63_287 VPWR VGND sg13g2_decap_8
XFILLER_51_438 VPWR VGND sg13g2_decap_8
XFILLER_45_980 VPWR VGND sg13g2_decap_8
XFILLER_32_641 VPWR VGND sg13g2_decap_8
XFILLER_31_140 VPWR VGND sg13g2_decap_8
XFILLER_20_858 VPWR VGND sg13g2_decap_8
XFILLER_75_0 VPWR VGND sg13g2_decap_8
XFILLER_99_630 VPWR VGND sg13g2_decap_8
XFILLER_28_1001 VPWR VGND sg13g2_decap_8
XFILLER_101_602 VPWR VGND sg13g2_decap_8
XFILLER_98_151 VPWR VGND sg13g2_decap_8
XFILLER_87_847 VPWR VGND sg13g2_decap_8
XFILLER_59_516 VPWR VGND sg13g2_decap_8
XFILLER_100_112 VPWR VGND sg13g2_decap_8
XFILLER_101_679 VPWR VGND sg13g2_decap_8
XFILLER_86_368 VPWR VGND sg13g2_decap_8
XFILLER_74_519 VPWR VGND sg13g2_decap_8
XFILLER_67_560 VPWR VGND sg13g2_decap_8
XFILLER_55_700 VPWR VGND sg13g2_decap_8
XFILLER_28_903 VPWR VGND sg13g2_decap_8
XFILLER_100_189 VPWR VGND sg13g2_decap_8
XFILLER_54_221 VPWR VGND sg13g2_decap_8
XFILLER_27_424 VPWR VGND sg13g2_decap_8
XFILLER_39_284 VPWR VGND sg13g2_decap_8
XFILLER_55_777 VPWR VGND sg13g2_decap_8
XFILLER_43_917 VPWR VGND sg13g2_decap_8
XFILLER_82_574 VPWR VGND sg13g2_decap_8
XFILLER_70_714 VPWR VGND sg13g2_decap_8
XFILLER_36_980 VPWR VGND sg13g2_decap_8
XFILLER_54_298 VPWR VGND sg13g2_decap_8
XFILLER_52_14 VPWR VGND sg13g2_decap_8
XFILLER_42_438 VPWR VGND sg13g2_decap_8
XFILLER_23_630 VPWR VGND sg13g2_decap_8
XFILLER_35_490 VPWR VGND sg13g2_decap_8
XFILLER_22_151 VPWR VGND sg13g2_decap_8
XFILLER_11_847 VPWR VGND sg13g2_decap_8
XFILLER_10_368 VPWR VGND sg13g2_decap_8
XFILLER_2_501 VPWR VGND sg13g2_decap_8
XFILLER_105_952 VPWR VGND sg13g2_decap_8
XFILLER_89_140 VPWR VGND sg13g2_decap_8
XFILLER_104_462 VPWR VGND sg13g2_decap_8
XFILLER_78_825 VPWR VGND sg13g2_decap_8
XFILLER_2_578 VPWR VGND sg13g2_decap_8
XFILLER_77_77 VPWR VGND sg13g2_decap_8
XFILLER_93_817 VPWR VGND sg13g2_decap_8
XFILLER_77_357 VPWR VGND sg13g2_decap_8
XFILLER_58_560 VPWR VGND sg13g2_decap_8
XFILLER_19_903 VPWR VGND sg13g2_decap_8
XFILLER_46_711 VPWR VGND sg13g2_decap_8
XFILLER_45_210 VPWR VGND sg13g2_decap_8
XFILLER_18_413 VPWR VGND sg13g2_decap_8
XFILLER_93_54 VPWR VGND sg13g2_decap_8
XFILLER_73_585 VPWR VGND sg13g2_decap_8
XFILLER_61_725 VPWR VGND sg13g2_decap_8
XFILLER_46_788 VPWR VGND sg13g2_decap_8
XFILLER_45_287 VPWR VGND sg13g2_decap_8
XFILLER_27_991 VPWR VGND sg13g2_decap_8
XFILLER_33_427 VPWR VGND sg13g2_decap_8
XFILLER_34_928 VPWR VGND sg13g2_decap_8
XFILLER_60_235 VPWR VGND sg13g2_decap_8
XFILLER_14_630 VPWR VGND sg13g2_decap_8
XFILLER_26_70 VPWR VGND sg13g2_decap_8
XFILLER_26_490 VPWR VGND sg13g2_decap_8
XFILLER_13_140 VPWR VGND sg13g2_decap_8
XFILLER_9_133 VPWR VGND sg13g2_decap_8
XFILLER_6_840 VPWR VGND sg13g2_decap_8
XFILLER_5_361 VPWR VGND sg13g2_decap_8
XFILLER_68_313 VPWR VGND sg13g2_decap_8
XFILLER_96_644 VPWR VGND sg13g2_decap_8
XFILLER_69_869 VPWR VGND sg13g2_decap_8
XFILLER_3_63 VPWR VGND sg13g2_decap_8
XFILLER_95_165 VPWR VGND sg13g2_decap_8
XFILLER_83_305 VPWR VGND sg13g2_decap_8
XFILLER_56_508 VPWR VGND sg13g2_decap_8
XFILLER_49_571 VPWR VGND sg13g2_decap_8
XFILLER_36_210 VPWR VGND sg13g2_decap_8
XFILLER_37_711 VPWR VGND sg13g2_decap_8
XFILLER_92_861 VPWR VGND sg13g2_decap_8
XFILLER_25_917 VPWR VGND sg13g2_decap_8
XFILLER_91_371 VPWR VGND sg13g2_decap_8
XFILLER_64_585 VPWR VGND sg13g2_decap_8
XFILLER_52_714 VPWR VGND sg13g2_decap_8
XFILLER_18_980 VPWR VGND sg13g2_decap_8
XFILLER_36_287 VPWR VGND sg13g2_decap_8
XFILLER_37_788 VPWR VGND sg13g2_decap_8
XFILLER_51_235 VPWR VGND sg13g2_decap_8
XFILLER_24_438 VPWR VGND sg13g2_decap_8
XFILLER_33_994 VPWR VGND sg13g2_decap_8
XFILLER_20_655 VPWR VGND sg13g2_decap_8
XFILLER_22_39 VPWR VGND sg13g2_decap_8
XFILLER_106_749 VPWR VGND sg13g2_decap_8
XFILLER_105_259 VPWR VGND sg13g2_decap_8
XFILLER_59_313 VPWR VGND sg13g2_decap_8
XFILLER_87_644 VPWR VGND sg13g2_decap_8
XFILLER_102_966 VPWR VGND sg13g2_decap_8
XFILLER_86_165 VPWR VGND sg13g2_decap_8
XFILLER_47_14 VPWR VGND sg13g2_decap_8
XFILLER_28_700 VPWR VGND sg13g2_decap_8
XFILLER_101_476 VPWR VGND sg13g2_decap_8
XFILLER_74_316 VPWR VGND sg13g2_decap_8
XFILLER_68_880 VPWR VGND sg13g2_decap_8
XFILLER_103_42 VPWR VGND sg13g2_decap_8
XFILLER_90_809 VPWR VGND sg13g2_decap_8
XFILLER_16_917 VPWR VGND sg13g2_decap_8
XFILLER_27_221 VPWR VGND sg13g2_decap_8
XFILLER_28_777 VPWR VGND sg13g2_decap_8
XFILLER_83_872 VPWR VGND sg13g2_decap_8
XFILLER_82_371 VPWR VGND sg13g2_decap_8
XFILLER_70_511 VPWR VGND sg13g2_decap_8
XFILLER_55_574 VPWR VGND sg13g2_decap_8
XFILLER_43_714 VPWR VGND sg13g2_decap_8
XFILLER_63_35 VPWR VGND sg13g2_decap_8
XFILLER_42_235 VPWR VGND sg13g2_decap_8
XFILLER_15_438 VPWR VGND sg13g2_decap_8
XFILLER_27_298 VPWR VGND sg13g2_decap_8
XFILLER_70_588 VPWR VGND sg13g2_decap_8
XFILLER_11_644 VPWR VGND sg13g2_decap_8
XFILLER_10_165 VPWR VGND sg13g2_decap_8
XFILLER_7_648 VPWR VGND sg13g2_decap_8
XFILLER_6_147 VPWR VGND sg13g2_decap_8
XFILLER_88_32 VPWR VGND sg13g2_decap_8
XFILLER_3_854 VPWR VGND sg13g2_decap_8
XFILLER_2_375 VPWR VGND sg13g2_decap_8
XFILLER_78_622 VPWR VGND sg13g2_decap_8
XFILLER_93_614 VPWR VGND sg13g2_decap_8
XFILLER_77_154 VPWR VGND sg13g2_decap_8
XFILLER_19_700 VPWR VGND sg13g2_decap_8
XFILLER_78_699 VPWR VGND sg13g2_decap_8
XFILLER_66_839 VPWR VGND sg13g2_decap_8
XFILLER_59_880 VPWR VGND sg13g2_decap_8
XFILLER_18_210 VPWR VGND sg13g2_decap_8
XFILLER_81_809 VPWR VGND sg13g2_decap_8
XFILLER_92_168 VPWR VGND sg13g2_decap_8
XFILLER_80_308 VPWR VGND sg13g2_decap_8
XFILLER_74_883 VPWR VGND sg13g2_decap_8
XFILLER_46_585 VPWR VGND sg13g2_decap_8
XFILLER_19_777 VPWR VGND sg13g2_decap_8
XFILLER_34_725 VPWR VGND sg13g2_decap_8
XFILLER_73_382 VPWR VGND sg13g2_decap_8
XFILLER_61_522 VPWR VGND sg13g2_decap_8
XFILLER_18_287 VPWR VGND sg13g2_decap_8
XFILLER_33_224 VPWR VGND sg13g2_decap_8
XFILLER_18_1022 VPWR VGND sg13g2_decap_8
XFILLER_61_599 VPWR VGND sg13g2_decap_8
XFILLER_30_931 VPWR VGND sg13g2_decap_8
XFILLER_97_931 VPWR VGND sg13g2_decap_8
XFILLER_68_110 VPWR VGND sg13g2_decap_8
XFILLER_25_1015 VPWR VGND sg13g2_decap_8
XFILLER_38_0 VPWR VGND sg13g2_decap_8
XFILLER_96_441 VPWR VGND sg13g2_decap_8
XFILLER_69_666 VPWR VGND sg13g2_decap_8
XFILLER_56_305 VPWR VGND sg13g2_decap_8
XFILLER_29_508 VPWR VGND sg13g2_decap_8
XFILLER_83_102 VPWR VGND sg13g2_decap_8
XFILLER_68_187 VPWR VGND sg13g2_decap_8
XFILLER_84_658 VPWR VGND sg13g2_decap_8
XFILLER_65_861 VPWR VGND sg13g2_decap_8
XFILLER_83_179 VPWR VGND sg13g2_decap_8
XFILLER_71_319 VPWR VGND sg13g2_decap_8
XFILLER_52_511 VPWR VGND sg13g2_decap_8
XFILLER_17_39 VPWR VGND sg13g2_decap_8
XFILLER_25_714 VPWR VGND sg13g2_decap_8
XFILLER_37_585 VPWR VGND sg13g2_decap_8
XFILLER_64_382 VPWR VGND sg13g2_decap_8
XFILLER_24_235 VPWR VGND sg13g2_decap_8
XFILLER_80_875 VPWR VGND sg13g2_decap_8
XFILLER_40_728 VPWR VGND sg13g2_decap_8
XFILLER_52_588 VPWR VGND sg13g2_decap_8
XFILLER_21_931 VPWR VGND sg13g2_decap_8
XFILLER_33_49 VPWR VGND sg13g2_decap_8
XFILLER_33_791 VPWR VGND sg13g2_decap_8
XFILLER_32_1019 VPWR VGND sg13g2_decap_8
XFILLER_20_452 VPWR VGND sg13g2_decap_8
XFILLER_106_546 VPWR VGND sg13g2_decap_8
XFILLER_88_942 VPWR VGND sg13g2_decap_8
XFILLER_58_35 VPWR VGND sg13g2_decap_8
XFILLER_102_763 VPWR VGND sg13g2_decap_8
XFILLER_87_441 VPWR VGND sg13g2_decap_8
XFILLER_0_868 VPWR VGND sg13g2_decap_8
XFILLER_101_273 VPWR VGND sg13g2_decap_8
XFILLER_74_113 VPWR VGND sg13g2_decap_8
XFILLER_59_187 VPWR VGND sg13g2_decap_8
XFILLER_90_606 VPWR VGND sg13g2_decap_8
XFILLER_75_658 VPWR VGND sg13g2_decap_8
XFILLER_62_308 VPWR VGND sg13g2_decap_8
XFILLER_56_872 VPWR VGND sg13g2_decap_8
XFILLER_43_511 VPWR VGND sg13g2_decap_8
XFILLER_16_714 VPWR VGND sg13g2_decap_8
XFILLER_28_574 VPWR VGND sg13g2_decap_8
XFILLER_74_78 VPWR VGND sg13g2_decap_8
XFILLER_55_371 VPWR VGND sg13g2_decap_8
XFILLER_15_235 VPWR VGND sg13g2_decap_8
XFILLER_90_11 VPWR VGND sg13g2_decap_8
XFILLER_71_886 VPWR VGND sg13g2_decap_8
XFILLER_70_385 VPWR VGND sg13g2_decap_8
XFILLER_43_588 VPWR VGND sg13g2_decap_8
XFILLER_31_728 VPWR VGND sg13g2_decap_8
XFILLER_90_88 VPWR VGND sg13g2_decap_8
XFILLER_11_441 VPWR VGND sg13g2_decap_8
XFILLER_12_942 VPWR VGND sg13g2_decap_8
XFILLER_30_238 VPWR VGND sg13g2_decap_8
XFILLER_8_924 VPWR VGND sg13g2_decap_8
XFILLER_7_445 VPWR VGND sg13g2_decap_8
XFILLER_99_42 VPWR VGND sg13g2_decap_8
XFILLER_48_1015 VPWR VGND sg13g2_decap_8
XFILLER_98_739 VPWR VGND sg13g2_decap_8
XFILLER_3_651 VPWR VGND sg13g2_decap_8
XFILLER_97_238 VPWR VGND sg13g2_decap_8
XFILLER_79_942 VPWR VGND sg13g2_decap_8
XFILLER_2_172 VPWR VGND sg13g2_decap_8
XFILLER_31_7 VPWR VGND sg13g2_decap_8
XFILLER_94_945 VPWR VGND sg13g2_decap_8
XFILLER_93_411 VPWR VGND sg13g2_decap_8
XFILLER_78_496 VPWR VGND sg13g2_decap_8
XFILLER_66_636 VPWR VGND sg13g2_decap_8
XFILLER_81_606 VPWR VGND sg13g2_decap_8
XFILLER_54_809 VPWR VGND sg13g2_decap_8
XFILLER_93_488 VPWR VGND sg13g2_decap_8
XFILLER_80_105 VPWR VGND sg13g2_decap_8
XFILLER_65_168 VPWR VGND sg13g2_decap_8
XFILLER_53_308 VPWR VGND sg13g2_decap_8
XFILLER_47_861 VPWR VGND sg13g2_decap_8
XFILLER_0_42 VPWR VGND sg13g2_decap_8
XFILLER_19_574 VPWR VGND sg13g2_decap_8
XFILLER_74_680 VPWR VGND sg13g2_decap_8
XFILLER_46_382 VPWR VGND sg13g2_decap_8
XFILLER_34_522 VPWR VGND sg13g2_decap_8
XFILLER_62_875 VPWR VGND sg13g2_decap_8
XFILLER_55_1008 VPWR VGND sg13g2_decap_8
XFILLER_61_396 VPWR VGND sg13g2_decap_8
XFILLER_22_739 VPWR VGND sg13g2_decap_8
XFILLER_34_599 VPWR VGND sg13g2_decap_8
XFILLER_21_238 VPWR VGND sg13g2_decap_8
XFILLER_9_84 VPWR VGND sg13g2_decap_8
XFILLER_89_728 VPWR VGND sg13g2_decap_8
XFILLER_88_249 VPWR VGND sg13g2_decap_8
XFILLER_69_463 VPWR VGND sg13g2_decap_8
XFILLER_85_945 VPWR VGND sg13g2_decap_8
XFILLER_56_102 VPWR VGND sg13g2_decap_8
XFILLER_29_305 VPWR VGND sg13g2_decap_8
XFILLER_84_455 VPWR VGND sg13g2_decap_8
XFILLER_57_658 VPWR VGND sg13g2_decap_8
XFILLER_28_49 VPWR VGND sg13g2_decap_8
XFILLER_56_179 VPWR VGND sg13g2_decap_8
XFILLER_44_319 VPWR VGND sg13g2_decap_8
XFILLER_38_861 VPWR VGND sg13g2_decap_8
XFILLER_71_116 VPWR VGND sg13g2_decap_8
XFILLER_25_511 VPWR VGND sg13g2_decap_8
XFILLER_37_382 VPWR VGND sg13g2_decap_8
XFILLER_53_875 VPWR VGND sg13g2_decap_8
XFILLER_100_21 VPWR VGND sg13g2_decap_8
XFILLER_80_672 VPWR VGND sg13g2_decap_8
XFILLER_52_385 VPWR VGND sg13g2_decap_8
XFILLER_13_728 VPWR VGND sg13g2_decap_8
XFILLER_25_588 VPWR VGND sg13g2_decap_8
XFILLER_40_525 VPWR VGND sg13g2_decap_8
XFILLER_12_249 VPWR VGND sg13g2_decap_8
XFILLER_100_98 VPWR VGND sg13g2_decap_8
XFILLER_60_25 VPWR VGND sg13g2_decap_8
XFILLER_60_14 VPWR VGND sg13g2_decap_4
XFILLER_5_949 VPWR VGND sg13g2_decap_8
XFILLER_4_448 VPWR VGND sg13g2_decap_8
XFILLER_106_343 VPWR VGND sg13g2_decap_8
XFILLER_69_56 VPWR VGND sg13g2_decap_4
XFILLER_79_249 VPWR VGND sg13g2_decap_8
XFILLER_69_78 VPWR VGND sg13g2_decap_8
XFILLER_0_665 VPWR VGND sg13g2_decap_8
XFILLER_102_560 VPWR VGND sg13g2_decap_8
XFILLER_85_77 VPWR VGND sg13g2_decap_8
XFILLER_76_956 VPWR VGND sg13g2_decap_8
XFILLER_75_455 VPWR VGND sg13g2_decap_8
XFILLER_48_658 VPWR VGND sg13g2_decap_8
XFILLER_90_403 VPWR VGND sg13g2_decap_8
XFILLER_62_105 VPWR VGND sg13g2_decap_8
XFILLER_47_168 VPWR VGND sg13g2_decap_8
XFILLER_29_872 VPWR VGND sg13g2_decap_8
XFILLER_35_308 VPWR VGND sg13g2_decap_8
XFILLER_91_959 VPWR VGND sg13g2_decap_8
XFILLER_16_511 VPWR VGND sg13g2_decap_8
XFILLER_28_371 VPWR VGND sg13g2_decap_8
XFILLER_71_683 VPWR VGND sg13g2_decap_8
XFILLER_44_886 VPWR VGND sg13g2_decap_8
XFILLER_43_385 VPWR VGND sg13g2_decap_8
XFILLER_16_588 VPWR VGND sg13g2_decap_8
XFILLER_31_525 VPWR VGND sg13g2_decap_8
XFILLER_70_182 VPWR VGND sg13g2_decap_8
XFILLER_34_81 VPWR VGND sg13g2_decap_8
XFILLER_8_721 VPWR VGND sg13g2_decap_8
XFILLER_79_7 VPWR VGND sg13g2_decap_8
XFILLER_8_798 VPWR VGND sg13g2_decap_8
XFILLER_7_242 VPWR VGND sg13g2_decap_8
XFILLER_50_91 VPWR VGND sg13g2_decap_8
XFILLER_98_536 VPWR VGND sg13g2_decap_8
XFILLER_61_1012 VPWR VGND sg13g2_decap_8
XFILLER_67_945 VPWR VGND sg13g2_decap_8
XFILLER_94_742 VPWR VGND sg13g2_decap_8
XFILLER_78_293 VPWR VGND sg13g2_decap_8
XFILLER_66_433 VPWR VGND sg13g2_decap_8
XFILLER_27_809 VPWR VGND sg13g2_decap_8
XFILLER_39_669 VPWR VGND sg13g2_decap_8
XFILLER_81_403 VPWR VGND sg13g2_decap_8
XFILLER_54_606 VPWR VGND sg13g2_decap_8
XFILLER_53_105 VPWR VGND sg13g2_decap_8
XFILLER_26_308 VPWR VGND sg13g2_decap_8
XFILLER_38_168 VPWR VGND sg13g2_decap_8
XFILLER_93_285 VPWR VGND sg13g2_decap_8
XFILLER_82_959 VPWR VGND sg13g2_decap_8
XFILLER_19_371 VPWR VGND sg13g2_decap_8
XFILLER_90_970 VPWR VGND sg13g2_decap_8
XFILLER_35_875 VPWR VGND sg13g2_decap_8
XFILLER_62_672 VPWR VGND sg13g2_decap_8
XFILLER_50_812 VPWR VGND sg13g2_decap_8
XFILLER_61_193 VPWR VGND sg13g2_decap_8
XFILLER_22_536 VPWR VGND sg13g2_decap_8
XFILLER_34_396 VPWR VGND sg13g2_decap_8
XFILLER_50_889 VPWR VGND sg13g2_decap_8
XFILLER_30_28 VPWR VGND sg13g2_decap_8
XFILLER_104_847 VPWR VGND sg13g2_decap_8
XFILLER_89_525 VPWR VGND sg13g2_decap_8
XFILLER_103_357 VPWR VGND sg13g2_decap_8
XFILLER_69_260 VPWR VGND sg13g2_decap_8
XFILLER_29_102 VPWR VGND sg13g2_decap_8
XFILLER_85_742 VPWR VGND sg13g2_decap_8
XFILLER_58_945 VPWR VGND sg13g2_decap_8
XFILLER_84_252 VPWR VGND sg13g2_decap_8
XFILLER_57_455 VPWR VGND sg13g2_decap_8
XFILLER_55_14 VPWR VGND sg13g2_decap_8
XFILLER_17_319 VPWR VGND sg13g2_decap_8
XFILLER_29_179 VPWR VGND sg13g2_decap_8
XFILLER_44_116 VPWR VGND sg13g2_decap_8
XFILLER_81_970 VPWR VGND sg13g2_decap_8
XFILLER_72_469 VPWR VGND sg13g2_decap_8
XFILLER_26_875 VPWR VGND sg13g2_decap_8
XFILLER_53_672 VPWR VGND sg13g2_decap_8
XFILLER_41_812 VPWR VGND sg13g2_decap_8
XFILLER_13_525 VPWR VGND sg13g2_decap_8
XFILLER_25_385 VPWR VGND sg13g2_decap_8
XFILLER_71_46 VPWR VGND sg13g2_decap_8
XFILLER_52_182 VPWR VGND sg13g2_decap_8
XFILLER_40_322 VPWR VGND sg13g2_decap_8
XFILLER_41_889 VPWR VGND sg13g2_decap_8
XFILLER_9_518 VPWR VGND sg13g2_decap_8
XFILLER_40_399 VPWR VGND sg13g2_decap_8
XFILLER_5_746 VPWR VGND sg13g2_decap_8
XFILLER_106_140 VPWR VGND sg13g2_decap_8
XFILLER_105_0 VPWR VGND sg13g2_decap_8
XFILLER_84_1001 VPWR VGND sg13g2_decap_8
XFILLER_4_245 VPWR VGND sg13g2_decap_8
XFILLER_96_21 VPWR VGND sg13g2_decap_8
XFILLER_1_952 VPWR VGND sg13g2_decap_8
XFILLER_0_462 VPWR VGND sg13g2_decap_8
XFILLER_96_98 VPWR VGND sg13g2_decap_8
XFILLER_76_753 VPWR VGND sg13g2_decap_8
XFILLER_49_956 VPWR VGND sg13g2_decap_8
XFILLER_75_252 VPWR VGND sg13g2_decap_8
XFILLER_48_455 VPWR VGND sg13g2_decap_8
XFILLER_29_81 VPWR VGND sg13g2_decap_8
XFILLER_91_756 VPWR VGND sg13g2_decap_8
XFILLER_90_200 VPWR VGND sg13g2_decap_8
XFILLER_35_105 VPWR VGND sg13g2_decap_8
XFILLER_63_469 VPWR VGND sg13g2_decap_8
XFILLER_90_277 VPWR VGND sg13g2_decap_8
XFILLER_50_119 VPWR VGND sg13g2_decap_8
XFILLER_45_91 VPWR VGND sg13g2_decap_8
XFILLER_44_683 VPWR VGND sg13g2_decap_8
XFILLER_16_385 VPWR VGND sg13g2_decap_8
XFILLER_17_886 VPWR VGND sg13g2_decap_8
XFILLER_32_823 VPWR VGND sg13g2_decap_8
XFILLER_71_480 VPWR VGND sg13g2_decap_8
XFILLER_43_182 VPWR VGND sg13g2_decap_8
XFILLER_31_322 VPWR VGND sg13g2_decap_8
XFILLER_31_399 VPWR VGND sg13g2_decap_8
XFILLER_8_595 VPWR VGND sg13g2_decap_8
XFILLER_99_812 VPWR VGND sg13g2_decap_8
XFILLER_6_63 VPWR VGND sg13g2_decap_8
XFILLER_99_889 VPWR VGND sg13g2_decap_8
XFILLER_98_333 VPWR VGND sg13g2_decap_8
XFILLER_6_1001 VPWR VGND sg13g2_decap_8
XFILLER_67_742 VPWR VGND sg13g2_decap_8
XFILLER_66_230 VPWR VGND sg13g2_decap_8
XFILLER_54_403 VPWR VGND sg13g2_decap_8
XFILLER_27_606 VPWR VGND sg13g2_decap_8
XFILLER_39_466 VPWR VGND sg13g2_decap_8
XFILLER_81_200 VPWR VGND sg13g2_decap_8
XFILLER_55_959 VPWR VGND sg13g2_decap_8
XFILLER_26_105 VPWR VGND sg13g2_decap_8
XFILLER_82_756 VPWR VGND sg13g2_decap_8
XFILLER_81_277 VPWR VGND sg13g2_decap_8
XFILLER_23_812 VPWR VGND sg13g2_decap_8
XFILLER_25_28 VPWR VGND sg13g2_decap_8
XFILLER_35_672 VPWR VGND sg13g2_decap_8
XFILLER_41_119 VPWR VGND sg13g2_decap_8
XFILLER_22_333 VPWR VGND sg13g2_decap_8
XFILLER_34_193 VPWR VGND sg13g2_decap_8
XFILLER_50_686 VPWR VGND sg13g2_decap_8
XFILLER_23_889 VPWR VGND sg13g2_decap_8
XFILLER_41_49 VPWR VGND sg13g2_decap_8
XFILLER_89_322 VPWR VGND sg13g2_decap_8
XFILLER_9_7 VPWR VGND sg13g2_decap_8
XFILLER_104_644 VPWR VGND sg13g2_decap_8
XFILLER_1_259 VPWR VGND sg13g2_decap_8
XFILLER_106_42 VPWR VGND sg13g2_decap_8
XFILLER_103_154 VPWR VGND sg13g2_decap_8
XFILLER_89_399 VPWR VGND sg13g2_decap_8
XFILLER_77_539 VPWR VGND sg13g2_decap_8
XFILLER_58_742 VPWR VGND sg13g2_decap_8
XFILLER_100_861 VPWR VGND sg13g2_decap_8
XFILLER_57_252 VPWR VGND sg13g2_decap_8
XFILLER_17_116 VPWR VGND sg13g2_decap_8
XFILLER_73_767 VPWR VGND sg13g2_decap_8
XFILLER_61_907 VPWR VGND sg13g2_decap_8
XFILLER_45_469 VPWR VGND sg13g2_decap_8
XFILLER_33_609 VPWR VGND sg13g2_decap_8
XFILLER_82_56 VPWR VGND sg13g2_decap_8
XFILLER_72_266 VPWR VGND sg13g2_decap_8
XFILLER_60_417 VPWR VGND sg13g2_decap_8
XFILLER_54_970 VPWR VGND sg13g2_decap_8
XFILLER_14_812 VPWR VGND sg13g2_decap_8
XFILLER_26_672 VPWR VGND sg13g2_decap_8
XFILLER_13_322 VPWR VGND sg13g2_decap_8
XFILLER_25_182 VPWR VGND sg13g2_decap_8
XFILLER_41_686 VPWR VGND sg13g2_decap_8
XFILLER_9_315 VPWR VGND sg13g2_decap_8
XFILLER_14_889 VPWR VGND sg13g2_decap_8
XFILLER_13_399 VPWR VGND sg13g2_decap_8
XFILLER_40_196 VPWR VGND sg13g2_decap_8
XFILLER_12_1028 VPWR VGND sg13g2_fill_1
XFILLER_5_543 VPWR VGND sg13g2_decap_8
XFILLER_99_119 VPWR VGND sg13g2_decap_8
XFILLER_96_826 VPWR VGND sg13g2_decap_8
XFILLER_95_347 VPWR VGND sg13g2_decap_8
XFILLER_76_550 VPWR VGND sg13g2_decap_8
XFILLER_49_753 VPWR VGND sg13g2_decap_8
XFILLER_48_252 VPWR VGND sg13g2_decap_8
XFILLER_91_553 VPWR VGND sg13g2_decap_8
XFILLER_64_767 VPWR VGND sg13g2_decap_8
XFILLER_36_469 VPWR VGND sg13g2_decap_8
XFILLER_63_266 VPWR VGND sg13g2_decap_8
XFILLER_51_417 VPWR VGND sg13g2_decap_8
XFILLER_17_683 VPWR VGND sg13g2_decap_8
XFILLER_23_119 VPWR VGND sg13g2_decap_8
XFILLER_44_480 VPWR VGND sg13g2_decap_8
XFILLER_16_182 VPWR VGND sg13g2_decap_8
XFILLER_32_620 VPWR VGND sg13g2_decap_8
XFILLER_60_984 VPWR VGND sg13g2_decap_8
XFILLER_20_837 VPWR VGND sg13g2_decap_8
XFILLER_32_697 VPWR VGND sg13g2_decap_8
XFILLER_31_196 VPWR VGND sg13g2_decap_8
XFILLER_9_882 VPWR VGND sg13g2_decap_8
XFILLER_8_392 VPWR VGND sg13g2_decap_8
XFILLER_98_130 VPWR VGND sg13g2_decap_8
XFILLER_99_686 VPWR VGND sg13g2_decap_8
XFILLER_87_826 VPWR VGND sg13g2_decap_8
XFILLER_101_658 VPWR VGND sg13g2_decap_8
XFILLER_86_347 VPWR VGND sg13g2_decap_8
XFILLER_100_168 VPWR VGND sg13g2_decap_8
XFILLER_54_200 VPWR VGND sg13g2_decap_8
XFILLER_27_403 VPWR VGND sg13g2_decap_8
XFILLER_28_959 VPWR VGND sg13g2_decap_8
XFILLER_39_263 VPWR VGND sg13g2_decap_8
XFILLER_82_553 VPWR VGND sg13g2_decap_8
XFILLER_55_756 VPWR VGND sg13g2_decap_8
XFILLER_36_49 VPWR VGND sg13g2_decap_8
XFILLER_54_277 VPWR VGND sg13g2_decap_8
XFILLER_42_417 VPWR VGND sg13g2_decap_8
XFILLER_14_119 VPWR VGND sg13g2_decap_8
XFILLER_51_984 VPWR VGND sg13g2_decap_8
XFILLER_22_130 VPWR VGND sg13g2_decap_8
XFILLER_50_483 VPWR VGND sg13g2_decap_8
XFILLER_11_826 VPWR VGND sg13g2_decap_8
XFILLER_23_686 VPWR VGND sg13g2_decap_8
XFILLER_10_347 VPWR VGND sg13g2_decap_8
XFILLER_6_329 VPWR VGND sg13g2_decap_8
XFILLER_105_931 VPWR VGND sg13g2_decap_8
XFILLER_104_441 VPWR VGND sg13g2_decap_8
XFILLER_78_804 VPWR VGND sg13g2_decap_8
XFILLER_7_4 VPWR VGND sg13g2_decap_8
XFILLER_2_557 VPWR VGND sg13g2_decap_8
XFILLER_81_1026 VPWR VGND sg13g2_fill_2
XFILLER_89_196 VPWR VGND sg13g2_decap_8
XFILLER_77_336 VPWR VGND sg13g2_decap_8
XFILLER_77_56 VPWR VGND sg13g2_decap_8
XFILLER_93_33 VPWR VGND sg13g2_decap_8
XFILLER_19_959 VPWR VGND sg13g2_decap_8
XFILLER_46_767 VPWR VGND sg13g2_decap_8
XFILLER_18_469 VPWR VGND sg13g2_decap_8
XFILLER_34_907 VPWR VGND sg13g2_decap_8
XFILLER_73_564 VPWR VGND sg13g2_decap_8
XFILLER_61_704 VPWR VGND sg13g2_decap_8
XFILLER_45_266 VPWR VGND sg13g2_decap_8
XFILLER_27_970 VPWR VGND sg13g2_decap_8
XFILLER_33_406 VPWR VGND sg13g2_decap_8
XFILLER_60_214 VPWR VGND sg13g2_decap_8
XFILLER_42_984 VPWR VGND sg13g2_decap_8
XFILLER_9_112 VPWR VGND sg13g2_decap_8
XFILLER_14_686 VPWR VGND sg13g2_decap_8
XFILLER_41_483 VPWR VGND sg13g2_decap_8
XFILLER_13_196 VPWR VGND sg13g2_decap_8
XFILLER_42_81 VPWR VGND sg13g2_decap_8
XFILLER_9_189 VPWR VGND sg13g2_decap_8
XFILLER_5_340 VPWR VGND sg13g2_decap_8
XFILLER_6_896 VPWR VGND sg13g2_decap_8
XFILLER_96_623 VPWR VGND sg13g2_decap_8
XFILLER_69_848 VPWR VGND sg13g2_decap_8
XFILLER_3_42 VPWR VGND sg13g2_decap_8
XFILLER_95_144 VPWR VGND sg13g2_decap_8
XFILLER_68_369 VPWR VGND sg13g2_decap_8
XFILLER_49_550 VPWR VGND sg13g2_decap_8
XFILLER_3_1015 VPWR VGND sg13g2_decap_8
XFILLER_97_1022 VPWR VGND sg13g2_decap_8
XFILLER_92_840 VPWR VGND sg13g2_decap_8
XFILLER_37_767 VPWR VGND sg13g2_decap_8
XFILLER_91_350 VPWR VGND sg13g2_decap_8
XFILLER_64_564 VPWR VGND sg13g2_decap_8
XFILLER_24_417 VPWR VGND sg13g2_decap_8
XFILLER_36_266 VPWR VGND sg13g2_decap_8
XFILLER_51_214 VPWR VGND sg13g2_decap_8
XFILLER_17_480 VPWR VGND sg13g2_decap_8
XFILLER_33_973 VPWR VGND sg13g2_decap_8
XFILLER_60_781 VPWR VGND sg13g2_decap_8
XFILLER_20_634 VPWR VGND sg13g2_decap_8
XFILLER_22_18 VPWR VGND sg13g2_decap_8
XFILLER_32_494 VPWR VGND sg13g2_decap_8
XFILLER_106_728 VPWR VGND sg13g2_decap_8
XFILLER_105_238 VPWR VGND sg13g2_decap_8
XFILLER_102_945 VPWR VGND sg13g2_decap_8
XFILLER_99_483 VPWR VGND sg13g2_decap_8
XFILLER_87_623 VPWR VGND sg13g2_decap_8
XFILLER_101_455 VPWR VGND sg13g2_decap_8
XFILLER_86_144 VPWR VGND sg13g2_decap_8
XFILLER_59_369 VPWR VGND sg13g2_decap_8
XFILLER_27_200 VPWR VGND sg13g2_decap_8
XFILLER_103_21 VPWR VGND sg13g2_decap_8
XFILLER_83_851 VPWR VGND sg13g2_decap_8
XFILLER_55_553 VPWR VGND sg13g2_decap_8
XFILLER_28_756 VPWR VGND sg13g2_decap_8
XFILLER_82_350 VPWR VGND sg13g2_decap_8
XFILLER_63_14 VPWR VGND sg13g2_decap_8
XFILLER_15_417 VPWR VGND sg13g2_decap_8
XFILLER_27_277 VPWR VGND sg13g2_decap_8
XFILLER_103_98 VPWR VGND sg13g2_decap_8
XFILLER_42_214 VPWR VGND sg13g2_decap_8
XFILLER_70_567 VPWR VGND sg13g2_decap_8
XFILLER_51_781 VPWR VGND sg13g2_decap_8
XFILLER_11_623 VPWR VGND sg13g2_decap_8
XFILLER_23_483 VPWR VGND sg13g2_decap_8
XFILLER_24_984 VPWR VGND sg13g2_decap_8
XFILLER_50_280 VPWR VGND sg13g2_decap_8
XFILLER_10_144 VPWR VGND sg13g2_decap_8
XFILLER_7_627 VPWR VGND sg13g2_decap_8
XFILLER_6_126 VPWR VGND sg13g2_decap_8
XFILLER_88_11 VPWR VGND sg13g2_decap_8
XFILLER_12_95 VPWR VGND sg13g2_decap_8
XFILLER_3_833 VPWR VGND sg13g2_decap_8
XFILLER_88_88 VPWR VGND sg13g2_decap_8
XFILLER_78_601 VPWR VGND sg13g2_decap_8
XFILLER_2_354 VPWR VGND sg13g2_decap_8
XFILLER_78_678 VPWR VGND sg13g2_decap_8
XFILLER_77_133 VPWR VGND sg13g2_decap_8
XFILLER_66_818 VPWR VGND sg13g2_decap_8
XFILLER_92_147 VPWR VGND sg13g2_decap_8
XFILLER_19_756 VPWR VGND sg13g2_decap_8
XFILLER_74_862 VPWR VGND sg13g2_decap_8
XFILLER_73_361 VPWR VGND sg13g2_decap_8
XFILLER_61_501 VPWR VGND sg13g2_decap_8
XFILLER_46_564 VPWR VGND sg13g2_decap_8
XFILLER_18_266 VPWR VGND sg13g2_decap_8
XFILLER_33_203 VPWR VGND sg13g2_decap_8
XFILLER_34_704 VPWR VGND sg13g2_decap_8
XFILLER_37_81 VPWR VGND sg13g2_decap_8
XFILLER_61_578 VPWR VGND sg13g2_decap_8
XFILLER_18_1001 VPWR VGND sg13g2_decap_8
XFILLER_42_781 VPWR VGND sg13g2_decap_8
XFILLER_14_483 VPWR VGND sg13g2_decap_8
XFILLER_15_984 VPWR VGND sg13g2_decap_8
XFILLER_30_910 VPWR VGND sg13g2_decap_8
XFILLER_105_1015 VPWR VGND sg13g2_decap_8
XFILLER_53_91 VPWR VGND sg13g2_decap_8
XFILLER_41_280 VPWR VGND sg13g2_decap_8
XFILLER_30_987 VPWR VGND sg13g2_decap_8
XFILLER_6_693 VPWR VGND sg13g2_decap_8
XFILLER_97_910 VPWR VGND sg13g2_decap_8
XFILLER_96_420 VPWR VGND sg13g2_decap_8
XFILLER_69_645 VPWR VGND sg13g2_decap_8
XFILLER_97_987 VPWR VGND sg13g2_decap_8
XFILLER_96_497 VPWR VGND sg13g2_decap_8
XFILLER_84_637 VPWR VGND sg13g2_decap_8
XFILLER_68_166 VPWR VGND sg13g2_decap_8
XFILLER_65_840 VPWR VGND sg13g2_decap_8
XFILLER_17_18 VPWR VGND sg13g2_decap_8
XFILLER_83_158 VPWR VGND sg13g2_decap_8
XFILLER_64_361 VPWR VGND sg13g2_decap_8
XFILLER_37_564 VPWR VGND sg13g2_decap_8
XFILLER_80_854 VPWR VGND sg13g2_decap_8
XFILLER_24_214 VPWR VGND sg13g2_decap_8
XFILLER_52_567 VPWR VGND sg13g2_decap_8
XFILLER_40_707 VPWR VGND sg13g2_decap_8
XFILLER_21_910 VPWR VGND sg13g2_decap_8
XFILLER_33_28 VPWR VGND sg13g2_decap_8
XFILLER_33_770 VPWR VGND sg13g2_decap_8
XFILLER_20_431 VPWR VGND sg13g2_decap_8
XFILLER_32_291 VPWR VGND sg13g2_decap_8
XFILLER_21_987 VPWR VGND sg13g2_decap_8
XFILLER_106_525 VPWR VGND sg13g2_decap_8
XFILLER_99_280 VPWR VGND sg13g2_decap_8
XFILLER_88_921 VPWR VGND sg13g2_decap_8
XFILLER_87_420 VPWR VGND sg13g2_decap_8
XFILLER_58_14 VPWR VGND sg13g2_decap_8
XFILLER_0_847 VPWR VGND sg13g2_decap_8
XFILLER_102_742 VPWR VGND sg13g2_decap_8
XFILLER_101_252 VPWR VGND sg13g2_decap_8
XFILLER_88_998 VPWR VGND sg13g2_decap_8
XFILLER_87_497 VPWR VGND sg13g2_decap_8
XFILLER_75_637 VPWR VGND sg13g2_decap_8
XFILLER_59_166 VPWR VGND sg13g2_decap_8
XFILLER_56_851 VPWR VGND sg13g2_decap_8
XFILLER_74_169 VPWR VGND sg13g2_decap_8
XFILLER_74_35 VPWR VGND sg13g2_decap_8
XFILLER_55_350 VPWR VGND sg13g2_decap_8
XFILLER_28_553 VPWR VGND sg13g2_decap_8
XFILLER_15_214 VPWR VGND sg13g2_decap_8
XFILLER_71_865 VPWR VGND sg13g2_decap_8
XFILLER_43_567 VPWR VGND sg13g2_decap_8
XFILLER_31_707 VPWR VGND sg13g2_decap_8
XFILLER_70_364 VPWR VGND sg13g2_decap_8
XFILLER_12_921 VPWR VGND sg13g2_decap_8
XFILLER_24_781 VPWR VGND sg13g2_decap_8
XFILLER_30_217 VPWR VGND sg13g2_decap_8
XFILLER_90_67 VPWR VGND sg13g2_decap_8
XFILLER_8_903 VPWR VGND sg13g2_decap_8
XFILLER_11_420 VPWR VGND sg13g2_decap_8
XFILLER_23_280 VPWR VGND sg13g2_decap_8
XFILLER_7_424 VPWR VGND sg13g2_decap_8
XFILLER_12_998 VPWR VGND sg13g2_decap_8
XFILLER_99_21 VPWR VGND sg13g2_decap_8
XFILLER_11_497 VPWR VGND sg13g2_decap_8
XFILLER_99_98 VPWR VGND sg13g2_decap_8
XFILLER_3_630 VPWR VGND sg13g2_decap_8
XFILLER_98_718 VPWR VGND sg13g2_decap_8
XFILLER_97_217 VPWR VGND sg13g2_decap_8
XFILLER_79_921 VPWR VGND sg13g2_decap_8
XFILLER_2_151 VPWR VGND sg13g2_decap_8
XFILLER_94_924 VPWR VGND sg13g2_decap_8
XFILLER_79_998 VPWR VGND sg13g2_decap_8
XFILLER_78_475 VPWR VGND sg13g2_decap_8
XFILLER_66_615 VPWR VGND sg13g2_decap_8
XFILLER_65_147 VPWR VGND sg13g2_decap_8
XFILLER_47_840 VPWR VGND sg13g2_decap_8
XFILLER_48_91 VPWR VGND sg13g2_decap_8
XFILLER_93_467 VPWR VGND sg13g2_decap_8
XFILLER_46_361 VPWR VGND sg13g2_decap_8
XFILLER_0_21 VPWR VGND sg13g2_decap_8
XFILLER_19_553 VPWR VGND sg13g2_decap_8
XFILLER_34_501 VPWR VGND sg13g2_decap_8
XFILLER_62_854 VPWR VGND sg13g2_decap_8
XFILLER_0_98 VPWR VGND sg13g2_decap_8
XFILLER_22_718 VPWR VGND sg13g2_decap_8
XFILLER_61_375 VPWR VGND sg13g2_decap_8
XFILLER_15_781 VPWR VGND sg13g2_decap_8
XFILLER_21_217 VPWR VGND sg13g2_decap_8
XFILLER_34_578 VPWR VGND sg13g2_decap_8
XFILLER_9_63 VPWR VGND sg13g2_decap_8
XFILLER_14_280 VPWR VGND sg13g2_decap_8
XFILLER_30_784 VPWR VGND sg13g2_decap_8
XFILLER_50_0 VPWR VGND sg13g2_decap_8
XFILLER_7_991 VPWR VGND sg13g2_decap_8
XFILLER_6_490 VPWR VGND sg13g2_decap_8
XFILLER_89_707 VPWR VGND sg13g2_decap_8
XFILLER_103_539 VPWR VGND sg13g2_decap_8
XFILLER_88_228 VPWR VGND sg13g2_decap_8
XFILLER_69_442 VPWR VGND sg13g2_decap_8
XFILLER_97_784 VPWR VGND sg13g2_decap_8
XFILLER_85_924 VPWR VGND sg13g2_decap_8
XFILLER_57_637 VPWR VGND sg13g2_decap_8
XFILLER_28_28 VPWR VGND sg13g2_decap_8
XFILLER_96_294 VPWR VGND sg13g2_decap_8
XFILLER_84_434 VPWR VGND sg13g2_decap_8
XFILLER_38_840 VPWR VGND sg13g2_decap_8
XFILLER_56_158 VPWR VGND sg13g2_decap_8
XFILLER_37_361 VPWR VGND sg13g2_decap_8
XFILLER_80_651 VPWR VGND sg13g2_decap_8
XFILLER_53_854 VPWR VGND sg13g2_decap_8
XFILLER_13_707 VPWR VGND sg13g2_decap_8
XFILLER_25_567 VPWR VGND sg13g2_decap_8
XFILLER_52_364 VPWR VGND sg13g2_decap_8
XFILLER_40_504 VPWR VGND sg13g2_decap_8
XFILLER_12_228 VPWR VGND sg13g2_decap_8
XFILLER_100_77 VPWR VGND sg13g2_decap_8
XFILLER_21_784 VPWR VGND sg13g2_decap_8
XFILLER_5_928 VPWR VGND sg13g2_decap_8
XFILLER_106_322 VPWR VGND sg13g2_decap_8
XFILLER_4_427 VPWR VGND sg13g2_decap_8
XFILLER_69_35 VPWR VGND sg13g2_decap_8
XFILLER_106_399 VPWR VGND sg13g2_decap_8
XFILLER_79_228 VPWR VGND sg13g2_decap_8
XFILLER_0_644 VPWR VGND sg13g2_decap_8
XFILLER_88_795 VPWR VGND sg13g2_decap_8
XFILLER_76_935 VPWR VGND sg13g2_decap_8
XFILLER_87_294 VPWR VGND sg13g2_decap_8
XFILLER_85_56 VPWR VGND sg13g2_decap_8
XFILLER_75_434 VPWR VGND sg13g2_decap_8
XFILLER_48_637 VPWR VGND sg13g2_decap_8
XFILLER_91_938 VPWR VGND sg13g2_decap_8
XFILLER_47_147 VPWR VGND sg13g2_decap_8
XFILLER_28_350 VPWR VGND sg13g2_decap_8
XFILLER_29_851 VPWR VGND sg13g2_decap_8
XFILLER_90_459 VPWR VGND sg13g2_decap_8
XFILLER_71_662 VPWR VGND sg13g2_decap_8
XFILLER_44_865 VPWR VGND sg13g2_decap_8
XFILLER_16_567 VPWR VGND sg13g2_decap_8
XFILLER_70_161 VPWR VGND sg13g2_decap_8
XFILLER_43_364 VPWR VGND sg13g2_decap_8
XFILLER_31_504 VPWR VGND sg13g2_decap_8
XFILLER_34_60 VPWR VGND sg13g2_decap_8
XFILLER_8_700 VPWR VGND sg13g2_decap_8
XFILLER_15_1026 VPWR VGND sg13g2_fill_2
XFILLER_7_221 VPWR VGND sg13g2_decap_8
XFILLER_12_795 VPWR VGND sg13g2_decap_8
XFILLER_8_777 VPWR VGND sg13g2_decap_8
XFILLER_11_294 VPWR VGND sg13g2_decap_8
XFILLER_50_70 VPWR VGND sg13g2_decap_8
XFILLER_7_298 VPWR VGND sg13g2_decap_8
XFILLER_98_515 VPWR VGND sg13g2_decap_8
XFILLER_4_994 VPWR VGND sg13g2_decap_8
XFILLER_94_721 VPWR VGND sg13g2_decap_8
XFILLER_79_795 VPWR VGND sg13g2_decap_8
XFILLER_78_272 VPWR VGND sg13g2_decap_8
XFILLER_67_924 VPWR VGND sg13g2_decap_8
XFILLER_66_412 VPWR VGND sg13g2_decap_8
XFILLER_22_4 VPWR VGND sg13g2_decap_8
XFILLER_22_1019 VPWR VGND sg13g2_decap_8
XFILLER_39_648 VPWR VGND sg13g2_decap_8
XFILLER_93_264 VPWR VGND sg13g2_decap_8
XFILLER_82_938 VPWR VGND sg13g2_decap_8
XFILLER_19_350 VPWR VGND sg13g2_decap_8
XFILLER_38_147 VPWR VGND sg13g2_decap_8
XFILLER_94_798 VPWR VGND sg13g2_decap_8
XFILLER_66_489 VPWR VGND sg13g2_decap_8
XFILLER_81_459 VPWR VGND sg13g2_decap_8
XFILLER_62_651 VPWR VGND sg13g2_decap_8
XFILLER_35_854 VPWR VGND sg13g2_decap_8
XFILLER_22_515 VPWR VGND sg13g2_decap_8
XFILLER_34_375 VPWR VGND sg13g2_decap_8
XFILLER_61_172 VPWR VGND sg13g2_decap_8
XFILLER_50_868 VPWR VGND sg13g2_decap_8
XFILLER_30_581 VPWR VGND sg13g2_decap_8
XFILLER_89_504 VPWR VGND sg13g2_decap_8
XFILLER_104_826 VPWR VGND sg13g2_decap_8
XFILLER_103_336 VPWR VGND sg13g2_decap_8
XFILLER_85_721 VPWR VGND sg13g2_decap_8
XFILLER_58_924 VPWR VGND sg13g2_decap_8
XFILLER_97_581 VPWR VGND sg13g2_decap_8
XFILLER_57_434 VPWR VGND sg13g2_decap_8
XFILLER_84_231 VPWR VGND sg13g2_decap_8
XFILLER_29_158 VPWR VGND sg13g2_decap_8
XFILLER_85_798 VPWR VGND sg13g2_decap_8
XFILLER_73_949 VPWR VGND sg13g2_decap_8
XFILLER_72_448 VPWR VGND sg13g2_decap_8
XFILLER_53_651 VPWR VGND sg13g2_decap_8
XFILLER_26_854 VPWR VGND sg13g2_decap_8
XFILLER_52_161 VPWR VGND sg13g2_decap_8
XFILLER_13_504 VPWR VGND sg13g2_decap_8
XFILLER_25_364 VPWR VGND sg13g2_decap_8
XFILLER_38_1015 VPWR VGND sg13g2_decap_8
XFILLER_40_301 VPWR VGND sg13g2_decap_8
XFILLER_71_25 VPWR VGND sg13g2_decap_8
XFILLER_41_868 VPWR VGND sg13g2_decap_8
XFILLER_40_378 VPWR VGND sg13g2_decap_8
XFILLER_21_581 VPWR VGND sg13g2_decap_8
XFILLER_5_725 VPWR VGND sg13g2_decap_8
XFILLER_4_224 VPWR VGND sg13g2_decap_8
XFILLER_45_1008 VPWR VGND sg13g2_decap_8
XFILLER_20_95 VPWR VGND sg13g2_decap_8
XFILLER_106_196 VPWR VGND sg13g2_decap_8
XFILLER_1_931 VPWR VGND sg13g2_decap_8
XFILLER_96_77 VPWR VGND sg13g2_decap_8
XFILLER_95_529 VPWR VGND sg13g2_decap_8
XFILLER_49_935 VPWR VGND sg13g2_decap_8
XFILLER_0_441 VPWR VGND sg13g2_decap_8
XFILLER_88_592 VPWR VGND sg13g2_decap_8
XFILLER_76_732 VPWR VGND sg13g2_decap_8
XFILLER_48_434 VPWR VGND sg13g2_decap_8
XFILLER_29_60 VPWR VGND sg13g2_decap_8
XFILLER_75_231 VPWR VGND sg13g2_decap_8
XFILLER_91_735 VPWR VGND sg13g2_decap_8
XFILLER_64_949 VPWR VGND sg13g2_decap_8
XFILLER_90_256 VPWR VGND sg13g2_decap_8
XFILLER_63_448 VPWR VGND sg13g2_decap_8
XFILLER_17_865 VPWR VGND sg13g2_decap_8
XFILLER_45_70 VPWR VGND sg13g2_decap_8
XFILLER_44_662 VPWR VGND sg13g2_decap_8
XFILLER_43_161 VPWR VGND sg13g2_decap_8
XFILLER_16_364 VPWR VGND sg13g2_decap_8
XFILLER_31_301 VPWR VGND sg13g2_decap_8
XFILLER_32_802 VPWR VGND sg13g2_decap_8
XFILLER_91_7 VPWR VGND sg13g2_decap_8
XFILLER_31_378 VPWR VGND sg13g2_decap_8
XFILLER_32_879 VPWR VGND sg13g2_decap_8
XFILLER_8_574 VPWR VGND sg13g2_decap_8
XFILLER_12_592 VPWR VGND sg13g2_decap_8
XFILLER_6_42 VPWR VGND sg13g2_decap_8
XFILLER_98_312 VPWR VGND sg13g2_decap_8
XFILLER_99_868 VPWR VGND sg13g2_decap_8
XFILLER_4_791 VPWR VGND sg13g2_decap_8
XFILLER_98_389 VPWR VGND sg13g2_decap_8
XFILLER_86_529 VPWR VGND sg13g2_decap_8
XFILLER_79_592 VPWR VGND sg13g2_decap_8
XFILLER_67_721 VPWR VGND sg13g2_decap_8
XFILLER_13_0 VPWR VGND sg13g2_decap_8
XFILLER_39_445 VPWR VGND sg13g2_decap_8
XFILLER_94_595 VPWR VGND sg13g2_decap_8
XFILLER_82_735 VPWR VGND sg13g2_decap_8
XFILLER_67_798 VPWR VGND sg13g2_decap_8
XFILLER_66_286 VPWR VGND sg13g2_decap_8
XFILLER_55_938 VPWR VGND sg13g2_decap_8
XFILLER_81_256 VPWR VGND sg13g2_decap_8
XFILLER_54_459 VPWR VGND sg13g2_decap_8
XFILLER_35_651 VPWR VGND sg13g2_decap_8
XFILLER_22_312 VPWR VGND sg13g2_decap_8
XFILLER_34_172 VPWR VGND sg13g2_decap_8
XFILLER_50_665 VPWR VGND sg13g2_decap_8
XFILLER_23_868 VPWR VGND sg13g2_decap_8
XFILLER_10_529 VPWR VGND sg13g2_decap_8
XFILLER_22_389 VPWR VGND sg13g2_decap_8
XFILLER_41_28 VPWR VGND sg13g2_decap_8
XFILLER_104_623 VPWR VGND sg13g2_decap_8
XFILLER_89_301 VPWR VGND sg13g2_decap_8
XFILLER_2_739 VPWR VGND sg13g2_decap_8
XFILLER_103_133 VPWR VGND sg13g2_decap_8
XFILLER_1_238 VPWR VGND sg13g2_decap_8
XFILLER_106_21 VPWR VGND sg13g2_decap_8
XFILLER_89_378 VPWR VGND sg13g2_decap_8
XFILLER_77_518 VPWR VGND sg13g2_decap_8
XFILLER_58_721 VPWR VGND sg13g2_decap_8
XFILLER_106_98 VPWR VGND sg13g2_decap_8
XFILLER_100_840 VPWR VGND sg13g2_decap_8
XFILLER_66_69 VPWR VGND sg13g2_decap_8
XFILLER_57_231 VPWR VGND sg13g2_decap_8
XFILLER_85_595 VPWR VGND sg13g2_decap_8
XFILLER_58_798 VPWR VGND sg13g2_decap_8
XFILLER_46_949 VPWR VGND sg13g2_decap_8
XFILLER_73_746 VPWR VGND sg13g2_decap_8
XFILLER_72_245 VPWR VGND sg13g2_decap_8
XFILLER_45_448 VPWR VGND sg13g2_decap_8
XFILLER_82_35 VPWR VGND sg13g2_decap_8
XFILLER_26_651 VPWR VGND sg13g2_decap_8
XFILLER_32_109 VPWR VGND sg13g2_decap_8
XFILLER_13_301 VPWR VGND sg13g2_decap_8
XFILLER_25_161 VPWR VGND sg13g2_decap_8
XFILLER_41_665 VPWR VGND sg13g2_decap_8
XFILLER_14_868 VPWR VGND sg13g2_decap_8
XFILLER_51_1012 VPWR VGND sg13g2_decap_8
XFILLER_13_378 VPWR VGND sg13g2_decap_8
XFILLER_15_95 VPWR VGND sg13g2_decap_8
XFILLER_40_175 VPWR VGND sg13g2_decap_8
XFILLER_5_522 VPWR VGND sg13g2_decap_8
XFILLER_5_599 VPWR VGND sg13g2_decap_8
XFILLER_96_805 VPWR VGND sg13g2_decap_8
XFILLER_95_326 VPWR VGND sg13g2_decap_8
XFILLER_49_732 VPWR VGND sg13g2_decap_8
XFILLER_48_231 VPWR VGND sg13g2_decap_8
XFILLER_37_949 VPWR VGND sg13g2_decap_8
XFILLER_91_532 VPWR VGND sg13g2_decap_8
XFILLER_64_746 VPWR VGND sg13g2_decap_8
XFILLER_63_245 VPWR VGND sg13g2_decap_8
XFILLER_36_448 VPWR VGND sg13g2_decap_8
XFILLER_17_662 VPWR VGND sg13g2_decap_8
XFILLER_16_161 VPWR VGND sg13g2_decap_8
XFILLER_60_963 VPWR VGND sg13g2_decap_8
XFILLER_20_816 VPWR VGND sg13g2_decap_8
XFILLER_32_676 VPWR VGND sg13g2_decap_8
XFILLER_31_175 VPWR VGND sg13g2_decap_8
XFILLER_9_861 VPWR VGND sg13g2_decap_8
XFILLER_8_371 VPWR VGND sg13g2_decap_8
XFILLER_99_665 VPWR VGND sg13g2_decap_8
XFILLER_87_805 VPWR VGND sg13g2_decap_8
XFILLER_101_637 VPWR VGND sg13g2_decap_8
XFILLER_98_186 VPWR VGND sg13g2_decap_8
XFILLER_86_326 VPWR VGND sg13g2_decap_8
XFILLER_100_147 VPWR VGND sg13g2_decap_8
XFILLER_39_242 VPWR VGND sg13g2_decap_8
XFILLER_95_893 VPWR VGND sg13g2_decap_8
XFILLER_67_595 VPWR VGND sg13g2_decap_8
XFILLER_55_735 VPWR VGND sg13g2_decap_8
XFILLER_28_938 VPWR VGND sg13g2_decap_8
XFILLER_36_28 VPWR VGND sg13g2_decap_8
XFILLER_94_392 VPWR VGND sg13g2_decap_8
XFILLER_82_532 VPWR VGND sg13g2_decap_8
XFILLER_27_459 VPWR VGND sg13g2_decap_8
XFILLER_54_256 VPWR VGND sg13g2_decap_8
XFILLER_74_1023 VPWR VGND sg13g2_decap_4
XFILLER_70_749 VPWR VGND sg13g2_decap_8
XFILLER_51_963 VPWR VGND sg13g2_decap_8
XFILLER_11_805 VPWR VGND sg13g2_decap_8
XFILLER_23_665 VPWR VGND sg13g2_decap_8
XFILLER_52_49 VPWR VGND sg13g2_decap_8
XFILLER_50_462 VPWR VGND sg13g2_decap_8
XFILLER_10_326 VPWR VGND sg13g2_decap_8
XFILLER_7_809 VPWR VGND sg13g2_decap_8
XFILLER_6_308 VPWR VGND sg13g2_decap_8
XFILLER_22_186 VPWR VGND sg13g2_decap_8
XFILLER_105_910 VPWR VGND sg13g2_decap_8
XFILLER_104_420 VPWR VGND sg13g2_decap_8
XFILLER_81_1005 VPWR VGND sg13g2_decap_8
XFILLER_2_536 VPWR VGND sg13g2_decap_8
XFILLER_105_987 VPWR VGND sg13g2_decap_8
XFILLER_77_35 VPWR VGND sg13g2_decap_8
XFILLER_104_497 VPWR VGND sg13g2_decap_8
XFILLER_89_175 VPWR VGND sg13g2_decap_8
XFILLER_77_315 VPWR VGND sg13g2_decap_8
XFILLER_93_12 VPWR VGND sg13g2_decap_8
XFILLER_92_329 VPWR VGND sg13g2_decap_8
XFILLER_86_893 VPWR VGND sg13g2_decap_8
XFILLER_58_595 VPWR VGND sg13g2_decap_8
XFILLER_19_938 VPWR VGND sg13g2_decap_8
XFILLER_85_392 VPWR VGND sg13g2_decap_8
XFILLER_73_543 VPWR VGND sg13g2_decap_8
XFILLER_46_746 VPWR VGND sg13g2_decap_8
XFILLER_45_245 VPWR VGND sg13g2_decap_8
XFILLER_18_448 VPWR VGND sg13g2_decap_8
XFILLER_93_89 VPWR VGND sg13g2_decap_8
XFILLER_42_963 VPWR VGND sg13g2_decap_8
XFILLER_14_665 VPWR VGND sg13g2_decap_8
XFILLER_13_175 VPWR VGND sg13g2_decap_8
XFILLER_41_462 VPWR VGND sg13g2_decap_8
XFILLER_42_60 VPWR VGND sg13g2_decap_8
XFILLER_9_168 VPWR VGND sg13g2_decap_8
XFILLER_10_893 VPWR VGND sg13g2_decap_8
XFILLER_6_875 VPWR VGND sg13g2_decap_8
XFILLER_5_396 VPWR VGND sg13g2_decap_8
XFILLER_96_602 VPWR VGND sg13g2_decap_8
XFILLER_69_827 VPWR VGND sg13g2_decap_8
XFILLER_3_21 VPWR VGND sg13g2_decap_8
XFILLER_95_123 VPWR VGND sg13g2_decap_8
XFILLER_96_679 VPWR VGND sg13g2_decap_8
XFILLER_84_819 VPWR VGND sg13g2_decap_8
XFILLER_68_348 VPWR VGND sg13g2_decap_8
XFILLER_3_98 VPWR VGND sg13g2_decap_8
XFILLER_97_1001 VPWR VGND sg13g2_decap_8
XFILLER_77_882 VPWR VGND sg13g2_decap_8
XFILLER_64_543 VPWR VGND sg13g2_decap_8
XFILLER_37_746 VPWR VGND sg13g2_decap_8
XFILLER_92_896 VPWR VGND sg13g2_decap_8
XFILLER_36_245 VPWR VGND sg13g2_decap_8
XFILLER_52_749 VPWR VGND sg13g2_decap_8
XFILLER_60_760 VPWR VGND sg13g2_decap_8
XFILLER_33_952 VPWR VGND sg13g2_decap_8
XFILLER_20_613 VPWR VGND sg13g2_decap_8
XFILLER_32_473 VPWR VGND sg13g2_decap_8
XFILLER_80_0 VPWR VGND sg13g2_decap_8
XFILLER_106_707 VPWR VGND sg13g2_decap_8
XFILLER_105_217 VPWR VGND sg13g2_decap_8
XFILLER_99_462 VPWR VGND sg13g2_decap_8
XFILLER_87_602 VPWR VGND sg13g2_decap_8
XFILLER_102_924 VPWR VGND sg13g2_decap_8
XFILLER_86_123 VPWR VGND sg13g2_decap_8
XFILLER_101_434 VPWR VGND sg13g2_decap_8
XFILLER_87_679 VPWR VGND sg13g2_decap_8
XFILLER_75_819 VPWR VGND sg13g2_decap_8
XFILLER_59_348 VPWR VGND sg13g2_decap_8
XFILLER_47_49 VPWR VGND sg13g2_decap_8
XFILLER_41_1022 VPWR VGND sg13g2_decap_8
XFILLER_95_690 VPWR VGND sg13g2_decap_8
XFILLER_83_830 VPWR VGND sg13g2_decap_8
XFILLER_67_392 VPWR VGND sg13g2_decap_8
XFILLER_55_532 VPWR VGND sg13g2_decap_8
XFILLER_28_735 VPWR VGND sg13g2_decap_8
XFILLER_27_256 VPWR VGND sg13g2_decap_8
XFILLER_103_77 VPWR VGND sg13g2_decap_8
XFILLER_70_546 VPWR VGND sg13g2_decap_8
XFILLER_43_749 VPWR VGND sg13g2_decap_8
XFILLER_24_963 VPWR VGND sg13g2_decap_8
XFILLER_51_760 VPWR VGND sg13g2_decap_8
XFILLER_11_602 VPWR VGND sg13g2_decap_8
XFILLER_23_462 VPWR VGND sg13g2_decap_8
XFILLER_10_123 VPWR VGND sg13g2_decap_8
XFILLER_7_606 VPWR VGND sg13g2_decap_8
XFILLER_6_105 VPWR VGND sg13g2_decap_8
XFILLER_11_679 VPWR VGND sg13g2_decap_8
XFILLER_3_812 VPWR VGND sg13g2_decap_8
XFILLER_12_74 VPWR VGND sg13g2_decap_8
XFILLER_88_67 VPWR VGND sg13g2_decap_8
XFILLER_3_889 VPWR VGND sg13g2_decap_8
XFILLER_2_333 VPWR VGND sg13g2_decap_8
XFILLER_105_784 VPWR VGND sg13g2_decap_8
XFILLER_77_112 VPWR VGND sg13g2_decap_8
XFILLER_104_294 VPWR VGND sg13g2_decap_8
XFILLER_78_657 VPWR VGND sg13g2_decap_8
XFILLER_77_189 VPWR VGND sg13g2_decap_8
XFILLER_65_329 VPWR VGND sg13g2_decap_8
XFILLER_93_649 VPWR VGND sg13g2_decap_8
XFILLER_92_126 VPWR VGND sg13g2_decap_8
XFILLER_86_690 VPWR VGND sg13g2_decap_8
XFILLER_74_841 VPWR VGND sg13g2_decap_8
XFILLER_58_392 VPWR VGND sg13g2_decap_8
XFILLER_46_543 VPWR VGND sg13g2_decap_8
XFILLER_19_735 VPWR VGND sg13g2_decap_8
XFILLER_37_60 VPWR VGND sg13g2_decap_8
XFILLER_73_340 VPWR VGND sg13g2_decap_8
XFILLER_18_245 VPWR VGND sg13g2_decap_8
XFILLER_61_557 VPWR VGND sg13g2_decap_8
XFILLER_15_963 VPWR VGND sg13g2_decap_8
XFILLER_33_259 VPWR VGND sg13g2_decap_8
XFILLER_53_70 VPWR VGND sg13g2_decap_8
XFILLER_42_760 VPWR VGND sg13g2_decap_8
XFILLER_14_462 VPWR VGND sg13g2_decap_8
XFILLER_30_966 VPWR VGND sg13g2_decap_8
XFILLER_10_690 VPWR VGND sg13g2_decap_8
XFILLER_6_672 VPWR VGND sg13g2_decap_8
XFILLER_5_193 VPWR VGND sg13g2_decap_8
XFILLER_69_624 VPWR VGND sg13g2_decap_8
XFILLER_97_966 VPWR VGND sg13g2_decap_8
XFILLER_68_145 VPWR VGND sg13g2_decap_8
XFILLER_57_819 VPWR VGND sg13g2_decap_8
XFILLER_96_476 VPWR VGND sg13g2_decap_8
XFILLER_84_616 VPWR VGND sg13g2_decap_8
XFILLER_83_137 VPWR VGND sg13g2_decap_8
XFILLER_37_543 VPWR VGND sg13g2_decap_8
XFILLER_64_340 VPWR VGND sg13g2_decap_8
XFILLER_92_693 VPWR VGND sg13g2_decap_8
XFILLER_80_833 VPWR VGND sg13g2_decap_8
XFILLER_65_896 VPWR VGND sg13g2_decap_8
XFILLER_25_749 VPWR VGND sg13g2_decap_8
XFILLER_52_546 VPWR VGND sg13g2_decap_8
XFILLER_71_1026 VPWR VGND sg13g2_fill_2
XFILLER_20_410 VPWR VGND sg13g2_decap_8
XFILLER_21_966 VPWR VGND sg13g2_decap_8
XFILLER_32_270 VPWR VGND sg13g2_decap_8
XFILLER_20_487 VPWR VGND sg13g2_decap_8
XFILLER_106_504 VPWR VGND sg13g2_decap_8
XFILLER_4_609 VPWR VGND sg13g2_decap_8
XFILLER_3_119 VPWR VGND sg13g2_decap_8
XFILLER_88_900 VPWR VGND sg13g2_decap_8
XFILLER_102_721 VPWR VGND sg13g2_decap_8
XFILLER_0_826 VPWR VGND sg13g2_decap_8
XFILLER_101_231 VPWR VGND sg13g2_decap_8
XFILLER_88_977 VPWR VGND sg13g2_decap_8
XFILLER_59_145 VPWR VGND sg13g2_decap_8
XFILLER_59_134 VPWR VGND sg13g2_decap_4
XFILLER_48_819 VPWR VGND sg13g2_decap_8
XFILLER_102_798 VPWR VGND sg13g2_decap_8
XFILLER_87_476 VPWR VGND sg13g2_decap_8
XFILLER_75_616 VPWR VGND sg13g2_decap_8
XFILLER_47_329 VPWR VGND sg13g2_decap_8
XFILLER_74_148 VPWR VGND sg13g2_decap_8
XFILLER_74_14 VPWR VGND sg13g2_decap_8
XFILLER_56_830 VPWR VGND sg13g2_decap_8
XFILLER_28_532 VPWR VGND sg13g2_decap_8
XFILLER_71_844 VPWR VGND sg13g2_decap_8
XFILLER_16_749 VPWR VGND sg13g2_decap_8
XFILLER_70_343 VPWR VGND sg13g2_decap_8
XFILLER_43_546 VPWR VGND sg13g2_decap_8
XFILLER_90_46 VPWR VGND sg13g2_decap_8
XFILLER_12_900 VPWR VGND sg13g2_decap_8
XFILLER_24_760 VPWR VGND sg13g2_decap_8
XFILLER_7_403 VPWR VGND sg13g2_decap_8
XFILLER_12_977 VPWR VGND sg13g2_decap_8
XFILLER_8_959 VPWR VGND sg13g2_decap_8
XFILLER_11_476 VPWR VGND sg13g2_decap_8
XFILLER_23_84 VPWR VGND sg13g2_decap_8
XFILLER_87_1022 VPWR VGND sg13g2_decap_8
XFILLER_99_77 VPWR VGND sg13g2_decap_8
XFILLER_79_900 VPWR VGND sg13g2_decap_8
XFILLER_2_130 VPWR VGND sg13g2_decap_8
XFILLER_105_581 VPWR VGND sg13g2_decap_8
XFILLER_3_686 VPWR VGND sg13g2_decap_8
XFILLER_94_903 VPWR VGND sg13g2_decap_8
XFILLER_79_977 VPWR VGND sg13g2_decap_8
XFILLER_78_454 VPWR VGND sg13g2_decap_8
XFILLER_48_70 VPWR VGND sg13g2_decap_8
XFILLER_93_446 VPWR VGND sg13g2_decap_8
XFILLER_65_126 VPWR VGND sg13g2_decap_8
XFILLER_19_532 VPWR VGND sg13g2_decap_8
XFILLER_38_329 VPWR VGND sg13g2_decap_8
XFILLER_46_340 VPWR VGND sg13g2_decap_8
XFILLER_0_1008 VPWR VGND sg13g2_decap_8
XFILLER_94_1015 VPWR VGND sg13g2_decap_8
XFILLER_62_833 VPWR VGND sg13g2_decap_8
XFILLER_47_896 VPWR VGND sg13g2_decap_8
XFILLER_0_77 VPWR VGND sg13g2_decap_8
XFILLER_61_354 VPWR VGND sg13g2_decap_8
XFILLER_34_557 VPWR VGND sg13g2_decap_8
XFILLER_15_760 VPWR VGND sg13g2_decap_8
XFILLER_9_42 VPWR VGND sg13g2_decap_8
XFILLER_30_763 VPWR VGND sg13g2_decap_8
XFILLER_7_970 VPWR VGND sg13g2_decap_8
XFILLER_88_207 VPWR VGND sg13g2_decap_8
XFILLER_43_0 VPWR VGND sg13g2_decap_8
XFILLER_103_518 VPWR VGND sg13g2_decap_8
XFILLER_9_1022 VPWR VGND sg13g2_decap_8
XFILLER_97_763 VPWR VGND sg13g2_decap_8
XFILLER_85_903 VPWR VGND sg13g2_decap_8
XFILLER_69_421 VPWR VGND sg13g2_decap_8
XFILLER_96_273 VPWR VGND sg13g2_decap_8
XFILLER_84_413 VPWR VGND sg13g2_decap_8
XFILLER_57_616 VPWR VGND sg13g2_decap_8
XFILLER_69_498 VPWR VGND sg13g2_decap_8
XFILLER_56_137 VPWR VGND sg13g2_decap_8
XFILLER_37_340 VPWR VGND sg13g2_decap_8
XFILLER_65_693 VPWR VGND sg13g2_decap_8
XFILLER_53_833 VPWR VGND sg13g2_decap_8
XFILLER_38_896 VPWR VGND sg13g2_decap_8
XFILLER_92_490 VPWR VGND sg13g2_decap_8
XFILLER_80_630 VPWR VGND sg13g2_decap_8
XFILLER_52_343 VPWR VGND sg13g2_decap_8
XFILLER_44_39 VPWR VGND sg13g2_decap_8
XFILLER_25_546 VPWR VGND sg13g2_decap_8
XFILLER_12_207 VPWR VGND sg13g2_decap_8
XFILLER_100_56 VPWR VGND sg13g2_decap_8
XFILLER_21_763 VPWR VGND sg13g2_decap_8
XFILLER_20_284 VPWR VGND sg13g2_decap_8
XFILLER_5_907 VPWR VGND sg13g2_decap_8
XFILLER_4_406 VPWR VGND sg13g2_decap_8
XFILLER_106_301 VPWR VGND sg13g2_decap_8
XFILLER_69_14 VPWR VGND sg13g2_decap_8
XFILLER_106_378 VPWR VGND sg13g2_decap_8
XFILLER_79_207 VPWR VGND sg13g2_decap_8
XFILLER_0_623 VPWR VGND sg13g2_decap_8
XFILLER_88_774 VPWR VGND sg13g2_decap_8
XFILLER_85_35 VPWR VGND sg13g2_decap_8
XFILLER_76_914 VPWR VGND sg13g2_decap_8
XFILLER_75_413 VPWR VGND sg13g2_decap_8
XFILLER_48_616 VPWR VGND sg13g2_decap_8
XFILLER_102_595 VPWR VGND sg13g2_decap_8
XFILLER_87_273 VPWR VGND sg13g2_decap_8
XFILLER_47_126 VPWR VGND sg13g2_decap_8
XFILLER_29_830 VPWR VGND sg13g2_decap_8
XFILLER_91_917 VPWR VGND sg13g2_decap_8
XFILLER_90_438 VPWR VGND sg13g2_decap_8
XFILLER_84_980 VPWR VGND sg13g2_decap_8
XFILLER_18_84 VPWR VGND sg13g2_decap_8
XFILLER_71_641 VPWR VGND sg13g2_decap_8
XFILLER_44_844 VPWR VGND sg13g2_decap_8
XFILLER_43_343 VPWR VGND sg13g2_decap_8
XFILLER_16_546 VPWR VGND sg13g2_decap_8
XFILLER_70_140 VPWR VGND sg13g2_decap_8
XFILLER_12_774 VPWR VGND sg13g2_decap_8
XFILLER_15_1005 VPWR VGND sg13g2_decap_8
XFILLER_102_1008 VPWR VGND sg13g2_decap_8
XFILLER_8_756 VPWR VGND sg13g2_decap_8
XFILLER_7_200 VPWR VGND sg13g2_decap_8
XFILLER_11_273 VPWR VGND sg13g2_decap_8
XFILLER_7_277 VPWR VGND sg13g2_decap_8
XFILLER_4_973 VPWR VGND sg13g2_decap_8
XFILLER_3_483 VPWR VGND sg13g2_decap_8
XFILLER_94_700 VPWR VGND sg13g2_decap_8
XFILLER_79_774 VPWR VGND sg13g2_decap_8
XFILLER_78_251 VPWR VGND sg13g2_decap_8
XFILLER_67_903 VPWR VGND sg13g2_decap_8
XFILLER_39_627 VPWR VGND sg13g2_decap_8
XFILLER_15_4 VPWR VGND sg13g2_decap_8
XFILLER_38_126 VPWR VGND sg13g2_decap_8
XFILLER_94_777 VPWR VGND sg13g2_decap_8
XFILLER_93_243 VPWR VGND sg13g2_decap_8
XFILLER_82_917 VPWR VGND sg13g2_decap_8
XFILLER_66_468 VPWR VGND sg13g2_decap_8
XFILLER_81_438 VPWR VGND sg13g2_decap_8
XFILLER_75_980 VPWR VGND sg13g2_decap_8
XFILLER_47_693 VPWR VGND sg13g2_decap_8
XFILLER_35_833 VPWR VGND sg13g2_decap_8
XFILLER_62_630 VPWR VGND sg13g2_decap_8
XFILLER_61_151 VPWR VGND sg13g2_decap_8
XFILLER_34_354 VPWR VGND sg13g2_decap_8
XFILLER_50_847 VPWR VGND sg13g2_decap_8
XFILLER_30_560 VPWR VGND sg13g2_decap_8
XFILLER_104_805 VPWR VGND sg13g2_decap_8
XFILLER_103_315 VPWR VGND sg13g2_decap_8
XFILLER_39_39 VPWR VGND sg13g2_decap_8
XFILLER_97_560 VPWR VGND sg13g2_decap_8
XFILLER_85_700 VPWR VGND sg13g2_decap_8
XFILLER_58_903 VPWR VGND sg13g2_decap_8
XFILLER_84_210 VPWR VGND sg13g2_decap_8
XFILLER_69_295 VPWR VGND sg13g2_decap_8
XFILLER_57_413 VPWR VGND sg13g2_decap_8
XFILLER_85_777 VPWR VGND sg13g2_decap_8
XFILLER_73_928 VPWR VGND sg13g2_decap_8
XFILLER_29_137 VPWR VGND sg13g2_decap_8
XFILLER_84_287 VPWR VGND sg13g2_decap_8
XFILLER_72_427 VPWR VGND sg13g2_decap_8
XFILLER_55_49 VPWR VGND sg13g2_decap_8
XFILLER_26_833 VPWR VGND sg13g2_decap_8
XFILLER_65_490 VPWR VGND sg13g2_decap_8
XFILLER_53_630 VPWR VGND sg13g2_decap_8
XFILLER_25_343 VPWR VGND sg13g2_decap_8
XFILLER_38_693 VPWR VGND sg13g2_decap_8
XFILLER_52_140 VPWR VGND sg13g2_decap_8
XFILLER_41_847 VPWR VGND sg13g2_decap_8
XFILLER_40_357 VPWR VGND sg13g2_decap_8
XFILLER_21_560 VPWR VGND sg13g2_decap_8
XFILLER_5_704 VPWR VGND sg13g2_decap_8
XFILLER_4_203 VPWR VGND sg13g2_decap_8
XFILLER_106_175 VPWR VGND sg13g2_decap_8
XFILLER_1_910 VPWR VGND sg13g2_decap_8
XFILLER_20_74 VPWR VGND sg13g2_decap_8
XFILLER_0_420 VPWR VGND sg13g2_decap_8
XFILLER_96_56 VPWR VGND sg13g2_decap_8
XFILLER_95_508 VPWR VGND sg13g2_decap_8
XFILLER_88_571 VPWR VGND sg13g2_decap_8
XFILLER_76_711 VPWR VGND sg13g2_decap_8
XFILLER_49_914 VPWR VGND sg13g2_decap_8
XFILLER_1_987 VPWR VGND sg13g2_decap_8
XFILLER_103_882 VPWR VGND sg13g2_decap_8
XFILLER_75_210 VPWR VGND sg13g2_decap_8
XFILLER_48_413 VPWR VGND sg13g2_decap_8
XFILLER_0_497 VPWR VGND sg13g2_decap_8
XFILLER_102_392 VPWR VGND sg13g2_decap_8
XFILLER_64_928 VPWR VGND sg13g2_decap_8
XFILLER_91_714 VPWR VGND sg13g2_decap_8
XFILLER_76_788 VPWR VGND sg13g2_decap_8
XFILLER_75_287 VPWR VGND sg13g2_decap_8
XFILLER_63_427 VPWR VGND sg13g2_decap_8
XFILLER_57_980 VPWR VGND sg13g2_decap_8
XFILLER_90_235 VPWR VGND sg13g2_decap_8
XFILLER_44_641 VPWR VGND sg13g2_decap_8
XFILLER_17_844 VPWR VGND sg13g2_decap_8
XFILLER_72_994 VPWR VGND sg13g2_decap_8
XFILLER_43_140 VPWR VGND sg13g2_decap_8
XFILLER_16_343 VPWR VGND sg13g2_decap_8
XFILLER_32_858 VPWR VGND sg13g2_decap_8
XFILLER_31_357 VPWR VGND sg13g2_decap_8
XFILLER_84_7 VPWR VGND sg13g2_decap_8
XFILLER_12_571 VPWR VGND sg13g2_decap_8
XFILLER_61_81 VPWR VGND sg13g2_decap_8
XFILLER_8_553 VPWR VGND sg13g2_decap_8
XFILLER_6_21 VPWR VGND sg13g2_decap_8
XFILLER_99_847 VPWR VGND sg13g2_decap_8
XFILLER_6_98 VPWR VGND sg13g2_decap_8
XFILLER_4_770 VPWR VGND sg13g2_decap_8
XFILLER_3_280 VPWR VGND sg13g2_decap_8
XFILLER_101_819 VPWR VGND sg13g2_decap_8
XFILLER_98_368 VPWR VGND sg13g2_decap_8
XFILLER_86_508 VPWR VGND sg13g2_decap_8
XFILLER_67_700 VPWR VGND sg13g2_decap_8
XFILLER_100_329 VPWR VGND sg13g2_decap_8
XFILLER_79_571 VPWR VGND sg13g2_decap_8
XFILLER_39_424 VPWR VGND sg13g2_decap_8
XFILLER_67_777 VPWR VGND sg13g2_decap_8
XFILLER_55_917 VPWR VGND sg13g2_decap_8
XFILLER_94_574 VPWR VGND sg13g2_decap_8
XFILLER_82_714 VPWR VGND sg13g2_decap_8
XFILLER_66_265 VPWR VGND sg13g2_decap_8
XFILLER_48_980 VPWR VGND sg13g2_decap_8
XFILLER_81_235 VPWR VGND sg13g2_decap_8
XFILLER_54_438 VPWR VGND sg13g2_decap_8
XFILLER_47_490 VPWR VGND sg13g2_decap_8
XFILLER_35_630 VPWR VGND sg13g2_decap_8
XFILLER_34_151 VPWR VGND sg13g2_decap_8
XFILLER_63_994 VPWR VGND sg13g2_decap_8
XFILLER_23_847 VPWR VGND sg13g2_decap_8
XFILLER_50_644 VPWR VGND sg13g2_decap_8
XFILLER_10_508 VPWR VGND sg13g2_decap_8
XFILLER_22_368 VPWR VGND sg13g2_decap_8
XFILLER_104_602 VPWR VGND sg13g2_decap_8
XFILLER_2_718 VPWR VGND sg13g2_decap_8
XFILLER_103_112 VPWR VGND sg13g2_decap_8
XFILLER_1_217 VPWR VGND sg13g2_decap_8
XFILLER_104_679 VPWR VGND sg13g2_decap_8
XFILLER_89_357 VPWR VGND sg13g2_decap_8
XFILLER_58_700 VPWR VGND sg13g2_decap_8
XFILLER_106_77 VPWR VGND sg13g2_decap_8
XFILLER_103_189 VPWR VGND sg13g2_decap_8
XFILLER_57_210 VPWR VGND sg13g2_decap_8
XFILLER_66_48 VPWR VGND sg13g2_decap_8
XFILLER_58_777 VPWR VGND sg13g2_decap_8
XFILLER_100_896 VPWR VGND sg13g2_decap_8
XFILLER_85_574 VPWR VGND sg13g2_decap_8
XFILLER_73_725 VPWR VGND sg13g2_decap_8
XFILLER_57_287 VPWR VGND sg13g2_decap_8
XFILLER_46_928 VPWR VGND sg13g2_decap_8
XFILLER_45_427 VPWR VGND sg13g2_decap_8
XFILLER_39_991 VPWR VGND sg13g2_decap_8
XFILLER_82_14 VPWR VGND sg13g2_decap_8
XFILLER_72_224 VPWR VGND sg13g2_decap_8
XFILLER_26_630 VPWR VGND sg13g2_decap_8
XFILLER_38_490 VPWR VGND sg13g2_decap_8
XFILLER_25_140 VPWR VGND sg13g2_decap_8
XFILLER_14_847 VPWR VGND sg13g2_decap_8
XFILLER_41_644 VPWR VGND sg13g2_decap_8
XFILLER_13_357 VPWR VGND sg13g2_decap_8
XFILLER_15_74 VPWR VGND sg13g2_decap_8
XFILLER_40_154 VPWR VGND sg13g2_decap_8
XFILLER_5_501 VPWR VGND sg13g2_decap_8
XFILLER_12_1019 VPWR VGND sg13g2_decap_8
XFILLER_31_84 VPWR VGND sg13g2_decap_8
XFILLER_5_578 VPWR VGND sg13g2_decap_8
XFILLER_95_305 VPWR VGND sg13g2_decap_8
XFILLER_49_711 VPWR VGND sg13g2_decap_8
XFILLER_48_210 VPWR VGND sg13g2_decap_8
XFILLER_1_784 VPWR VGND sg13g2_decap_8
XFILLER_0_294 VPWR VGND sg13g2_decap_8
XFILLER_91_511 VPWR VGND sg13g2_decap_8
XFILLER_76_585 VPWR VGND sg13g2_decap_8
XFILLER_64_725 VPWR VGND sg13g2_decap_8
XFILLER_49_788 VPWR VGND sg13g2_decap_8
XFILLER_48_287 VPWR VGND sg13g2_decap_8
XFILLER_36_427 VPWR VGND sg13g2_decap_8
XFILLER_37_928 VPWR VGND sg13g2_decap_8
XFILLER_63_224 VPWR VGND sg13g2_decap_8
XFILLER_56_81 VPWR VGND sg13g2_decap_8
XFILLER_17_641 VPWR VGND sg13g2_decap_8
XFILLER_91_588 VPWR VGND sg13g2_decap_8
XFILLER_16_140 VPWR VGND sg13g2_decap_8
XFILLER_72_791 VPWR VGND sg13g2_decap_8
XFILLER_60_942 VPWR VGND sg13g2_decap_8
XFILLER_45_994 VPWR VGND sg13g2_decap_8
XFILLER_32_655 VPWR VGND sg13g2_decap_8
XFILLER_72_91 VPWR VGND sg13g2_decap_8
XFILLER_31_154 VPWR VGND sg13g2_decap_8
XFILLER_9_840 VPWR VGND sg13g2_decap_8
XFILLER_8_350 VPWR VGND sg13g2_decap_8
XFILLER_99_644 VPWR VGND sg13g2_decap_8
XFILLER_28_1015 VPWR VGND sg13g2_decap_8
XFILLER_98_165 VPWR VGND sg13g2_decap_8
XFILLER_86_305 VPWR VGND sg13g2_decap_8
XFILLER_101_616 VPWR VGND sg13g2_decap_8
XFILLER_100_126 VPWR VGND sg13g2_decap_8
XFILLER_39_221 VPWR VGND sg13g2_decap_8
XFILLER_95_872 VPWR VGND sg13g2_decap_8
XFILLER_94_371 VPWR VGND sg13g2_decap_8
XFILLER_82_511 VPWR VGND sg13g2_decap_8
XFILLER_67_574 VPWR VGND sg13g2_decap_8
XFILLER_55_714 VPWR VGND sg13g2_decap_8
XFILLER_28_917 VPWR VGND sg13g2_decap_8
XFILLER_54_235 VPWR VGND sg13g2_decap_8
XFILLER_27_438 VPWR VGND sg13g2_decap_8
XFILLER_39_298 VPWR VGND sg13g2_decap_8
XFILLER_82_588 VPWR VGND sg13g2_decap_8
XFILLER_74_1002 VPWR VGND sg13g2_decap_8
XFILLER_70_728 VPWR VGND sg13g2_decap_8
XFILLER_63_791 VPWR VGND sg13g2_decap_8
XFILLER_51_942 VPWR VGND sg13g2_decap_8
XFILLER_36_994 VPWR VGND sg13g2_decap_8
XFILLER_52_28 VPWR VGND sg13g2_decap_8
XFILLER_50_441 VPWR VGND sg13g2_decap_8
XFILLER_23_644 VPWR VGND sg13g2_decap_8
XFILLER_35_1008 VPWR VGND sg13g2_decap_8
XFILLER_10_305 VPWR VGND sg13g2_decap_8
XFILLER_22_165 VPWR VGND sg13g2_decap_8
XFILLER_2_515 VPWR VGND sg13g2_decap_8
XFILLER_105_966 VPWR VGND sg13g2_decap_8
XFILLER_89_154 VPWR VGND sg13g2_decap_8
XFILLER_81_1028 VPWR VGND sg13g2_fill_1
XFILLER_77_14 VPWR VGND sg13g2_decap_8
XFILLER_104_476 VPWR VGND sg13g2_decap_8
XFILLER_78_839 VPWR VGND sg13g2_decap_8
XFILLER_92_308 VPWR VGND sg13g2_decap_8
XFILLER_86_872 VPWR VGND sg13g2_decap_8
XFILLER_85_371 VPWR VGND sg13g2_decap_8
XFILLER_58_574 VPWR VGND sg13g2_decap_8
XFILLER_46_725 VPWR VGND sg13g2_decap_8
XFILLER_19_917 VPWR VGND sg13g2_decap_8
XFILLER_100_693 VPWR VGND sg13g2_decap_8
XFILLER_73_522 VPWR VGND sg13g2_decap_8
XFILLER_45_224 VPWR VGND sg13g2_decap_8
XFILLER_18_427 VPWR VGND sg13g2_decap_8
XFILLER_93_68 VPWR VGND sg13g2_decap_8
XFILLER_73_599 VPWR VGND sg13g2_decap_8
XFILLER_61_739 VPWR VGND sg13g2_decap_8
XFILLER_26_84 VPWR VGND sg13g2_decap_8
XFILLER_60_249 VPWR VGND sg13g2_decap_8
XFILLER_42_942 VPWR VGND sg13g2_decap_8
XFILLER_14_644 VPWR VGND sg13g2_decap_8
XFILLER_41_441 VPWR VGND sg13g2_decap_8
XFILLER_13_154 VPWR VGND sg13g2_decap_8
XFILLER_9_147 VPWR VGND sg13g2_decap_8
XFILLER_10_872 VPWR VGND sg13g2_decap_8
XFILLER_6_854 VPWR VGND sg13g2_decap_8
XFILLER_47_7 VPWR VGND sg13g2_decap_8
XFILLER_5_375 VPWR VGND sg13g2_decap_8
XFILLER_69_806 VPWR VGND sg13g2_decap_8
XFILLER_95_102 VPWR VGND sg13g2_decap_8
XFILLER_68_327 VPWR VGND sg13g2_decap_8
XFILLER_96_658 VPWR VGND sg13g2_decap_8
XFILLER_3_77 VPWR VGND sg13g2_decap_8
XFILLER_1_581 VPWR VGND sg13g2_decap_8
XFILLER_95_179 VPWR VGND sg13g2_decap_8
XFILLER_83_319 VPWR VGND sg13g2_decap_8
XFILLER_77_861 VPWR VGND sg13g2_decap_8
XFILLER_67_91 VPWR VGND sg13g2_decap_8
XFILLER_49_585 VPWR VGND sg13g2_decap_8
XFILLER_37_725 VPWR VGND sg13g2_decap_8
XFILLER_76_382 VPWR VGND sg13g2_decap_8
XFILLER_64_522 VPWR VGND sg13g2_decap_8
XFILLER_36_224 VPWR VGND sg13g2_decap_8
XFILLER_92_875 VPWR VGND sg13g2_decap_8
XFILLER_58_1008 VPWR VGND sg13g2_decap_8
XFILLER_91_385 VPWR VGND sg13g2_decap_8
XFILLER_64_599 VPWR VGND sg13g2_decap_8
XFILLER_52_728 VPWR VGND sg13g2_decap_8
XFILLER_45_791 VPWR VGND sg13g2_decap_8
XFILLER_18_994 VPWR VGND sg13g2_decap_8
XFILLER_33_931 VPWR VGND sg13g2_decap_8
XFILLER_51_249 VPWR VGND sg13g2_decap_8
XFILLER_32_452 VPWR VGND sg13g2_decap_8
XFILLER_20_669 VPWR VGND sg13g2_decap_8
XFILLER_102_903 VPWR VGND sg13g2_decap_8
XFILLER_99_441 VPWR VGND sg13g2_decap_8
XFILLER_101_413 VPWR VGND sg13g2_decap_8
XFILLER_86_102 VPWR VGND sg13g2_decap_8
XFILLER_59_327 VPWR VGND sg13g2_decap_8
XFILLER_87_658 VPWR VGND sg13g2_decap_8
XFILLER_47_28 VPWR VGND sg13g2_decap_8
XFILLER_41_1001 VPWR VGND sg13g2_decap_8
XFILLER_86_179 VPWR VGND sg13g2_decap_8
XFILLER_68_894 VPWR VGND sg13g2_decap_8
XFILLER_28_714 VPWR VGND sg13g2_decap_8
XFILLER_67_371 VPWR VGND sg13g2_decap_8
XFILLER_55_511 VPWR VGND sg13g2_decap_8
XFILLER_27_235 VPWR VGND sg13g2_decap_8
XFILLER_103_56 VPWR VGND sg13g2_decap_8
XFILLER_83_886 VPWR VGND sg13g2_decap_8
XFILLER_82_385 VPWR VGND sg13g2_decap_8
XFILLER_70_525 VPWR VGND sg13g2_decap_8
XFILLER_63_49 VPWR VGND sg13g2_decap_8
XFILLER_55_588 VPWR VGND sg13g2_decap_8
XFILLER_43_728 VPWR VGND sg13g2_decap_8
XFILLER_36_791 VPWR VGND sg13g2_decap_8
XFILLER_42_249 VPWR VGND sg13g2_decap_8
XFILLER_23_441 VPWR VGND sg13g2_decap_8
XFILLER_24_942 VPWR VGND sg13g2_decap_8
XFILLER_10_102 VPWR VGND sg13g2_decap_8
XFILLER_11_658 VPWR VGND sg13g2_decap_8
XFILLER_10_179 VPWR VGND sg13g2_decap_8
XFILLER_12_53 VPWR VGND sg13g2_decap_8
XFILLER_88_46 VPWR VGND sg13g2_decap_8
XFILLER_2_312 VPWR VGND sg13g2_decap_8
XFILLER_105_763 VPWR VGND sg13g2_decap_8
XFILLER_3_868 VPWR VGND sg13g2_decap_8
XFILLER_104_273 VPWR VGND sg13g2_decap_8
XFILLER_78_636 VPWR VGND sg13g2_decap_8
XFILLER_2_389 VPWR VGND sg13g2_decap_8
XFILLER_93_628 VPWR VGND sg13g2_decap_8
XFILLER_92_105 VPWR VGND sg13g2_decap_8
XFILLER_77_168 VPWR VGND sg13g2_decap_8
XFILLER_65_308 VPWR VGND sg13g2_decap_8
XFILLER_19_714 VPWR VGND sg13g2_decap_8
XFILLER_101_980 VPWR VGND sg13g2_decap_8
XFILLER_74_820 VPWR VGND sg13g2_decap_8
XFILLER_59_894 VPWR VGND sg13g2_decap_8
XFILLER_58_371 VPWR VGND sg13g2_decap_8
XFILLER_46_522 VPWR VGND sg13g2_decap_8
XFILLER_18_224 VPWR VGND sg13g2_decap_8
XFILLER_100_490 VPWR VGND sg13g2_decap_8
XFILLER_74_897 VPWR VGND sg13g2_decap_8
XFILLER_73_396 VPWR VGND sg13g2_decap_8
XFILLER_61_536 VPWR VGND sg13g2_decap_8
XFILLER_46_599 VPWR VGND sg13g2_decap_8
XFILLER_34_739 VPWR VGND sg13g2_decap_8
XFILLER_14_441 VPWR VGND sg13g2_decap_8
XFILLER_15_942 VPWR VGND sg13g2_decap_8
XFILLER_33_238 VPWR VGND sg13g2_decap_8
XFILLER_30_945 VPWR VGND sg13g2_decap_8
XFILLER_6_651 VPWR VGND sg13g2_decap_8
XFILLER_5_172 VPWR VGND sg13g2_decap_8
XFILLER_69_603 VPWR VGND sg13g2_decap_8
XFILLER_64_1012 VPWR VGND sg13g2_decap_8
XFILLER_97_945 VPWR VGND sg13g2_decap_8
XFILLER_96_455 VPWR VGND sg13g2_decap_8
XFILLER_78_90 VPWR VGND sg13g2_decap_8
XFILLER_68_124 VPWR VGND sg13g2_decap_8
XFILLER_56_319 VPWR VGND sg13g2_decap_8
XFILLER_83_116 VPWR VGND sg13g2_decap_8
XFILLER_49_382 VPWR VGND sg13g2_decap_8
XFILLER_37_522 VPWR VGND sg13g2_decap_8
XFILLER_65_875 VPWR VGND sg13g2_decap_8
XFILLER_92_672 VPWR VGND sg13g2_decap_8
XFILLER_80_812 VPWR VGND sg13g2_decap_8
XFILLER_52_525 VPWR VGND sg13g2_decap_8
XFILLER_25_728 VPWR VGND sg13g2_decap_8
XFILLER_37_599 VPWR VGND sg13g2_decap_8
XFILLER_91_182 VPWR VGND sg13g2_decap_8
XFILLER_64_396 VPWR VGND sg13g2_decap_8
XFILLER_18_791 VPWR VGND sg13g2_decap_8
XFILLER_24_249 VPWR VGND sg13g2_decap_8
XFILLER_80_889 VPWR VGND sg13g2_decap_8
XFILLER_71_1005 VPWR VGND sg13g2_decap_8
XFILLER_21_945 VPWR VGND sg13g2_decap_8
XFILLER_20_466 VPWR VGND sg13g2_decap_8
XFILLER_0_805 VPWR VGND sg13g2_decap_8
XFILLER_102_700 VPWR VGND sg13g2_decap_8
XFILLER_101_210 VPWR VGND sg13g2_decap_8
XFILLER_88_956 VPWR VGND sg13g2_decap_8
XFILLER_87_455 VPWR VGND sg13g2_decap_8
XFILLER_59_113 VPWR VGND sg13g2_decap_8
XFILLER_58_49 VPWR VGND sg13g2_decap_8
XFILLER_102_777 VPWR VGND sg13g2_decap_8
XFILLER_47_308 VPWR VGND sg13g2_decap_8
XFILLER_101_287 VPWR VGND sg13g2_decap_8
XFILLER_74_127 VPWR VGND sg13g2_decap_8
XFILLER_68_691 VPWR VGND sg13g2_decap_8
XFILLER_28_511 VPWR VGND sg13g2_decap_8
XFILLER_83_683 VPWR VGND sg13g2_decap_8
XFILLER_71_823 VPWR VGND sg13g2_decap_8
XFILLER_56_886 VPWR VGND sg13g2_decap_8
XFILLER_55_385 VPWR VGND sg13g2_decap_8
XFILLER_43_525 VPWR VGND sg13g2_decap_8
XFILLER_16_728 VPWR VGND sg13g2_decap_8
XFILLER_28_588 VPWR VGND sg13g2_decap_8
XFILLER_82_182 VPWR VGND sg13g2_decap_8
XFILLER_70_322 VPWR VGND sg13g2_decap_8
XFILLER_15_249 VPWR VGND sg13g2_decap_8
XFILLER_90_25 VPWR VGND sg13g2_decap_8
XFILLER_70_399 VPWR VGND sg13g2_decap_8
XFILLER_12_956 VPWR VGND sg13g2_decap_8
XFILLER_8_938 VPWR VGND sg13g2_decap_8
XFILLER_11_455 VPWR VGND sg13g2_decap_8
XFILLER_23_63 VPWR VGND sg13g2_decap_8
XFILLER_99_56 VPWR VGND sg13g2_decap_8
XFILLER_87_1001 VPWR VGND sg13g2_decap_8
XFILLER_7_459 VPWR VGND sg13g2_decap_8
XFILLER_3_0 VPWR VGND sg13g2_decap_8
XFILLER_105_560 VPWR VGND sg13g2_decap_8
XFILLER_3_665 VPWR VGND sg13g2_decap_8
XFILLER_79_956 VPWR VGND sg13g2_decap_8
XFILLER_78_433 VPWR VGND sg13g2_decap_8
XFILLER_2_186 VPWR VGND sg13g2_decap_8
XFILLER_39_809 VPWR VGND sg13g2_decap_8
XFILLER_65_105 VPWR VGND sg13g2_decap_8
XFILLER_38_308 VPWR VGND sg13g2_decap_8
XFILLER_94_959 VPWR VGND sg13g2_decap_8
XFILLER_93_425 VPWR VGND sg13g2_decap_8
XFILLER_59_691 VPWR VGND sg13g2_decap_8
XFILLER_19_511 VPWR VGND sg13g2_decap_8
XFILLER_47_875 VPWR VGND sg13g2_decap_8
XFILLER_80_119 VPWR VGND sg13g2_decap_8
XFILLER_74_694 VPWR VGND sg13g2_decap_8
XFILLER_62_812 VPWR VGND sg13g2_decap_8
XFILLER_0_56 VPWR VGND sg13g2_decap_8
XFILLER_19_588 VPWR VGND sg13g2_decap_8
XFILLER_73_193 VPWR VGND sg13g2_decap_8
XFILLER_64_81 VPWR VGND sg13g2_decap_8
XFILLER_61_333 VPWR VGND sg13g2_decap_8
XFILLER_46_396 VPWR VGND sg13g2_decap_8
XFILLER_34_536 VPWR VGND sg13g2_decap_8
XFILLER_62_889 VPWR VGND sg13g2_decap_8
XFILLER_9_21 VPWR VGND sg13g2_decap_8
XFILLER_30_742 VPWR VGND sg13g2_decap_8
XFILLER_80_91 VPWR VGND sg13g2_decap_8
XFILLER_9_98 VPWR VGND sg13g2_decap_8
XFILLER_31_1022 VPWR VGND sg13g2_decap_8
XFILLER_69_400 VPWR VGND sg13g2_decap_8
XFILLER_9_1001 VPWR VGND sg13g2_decap_8
XFILLER_97_742 VPWR VGND sg13g2_decap_8
XFILLER_36_0 VPWR VGND sg13g2_decap_8
XFILLER_96_252 VPWR VGND sg13g2_decap_8
XFILLER_69_477 VPWR VGND sg13g2_decap_8
XFILLER_29_319 VPWR VGND sg13g2_decap_8
XFILLER_85_959 VPWR VGND sg13g2_decap_8
XFILLER_56_116 VPWR VGND sg13g2_decap_8
XFILLER_84_469 VPWR VGND sg13g2_decap_8
XFILLER_72_609 VPWR VGND sg13g2_decap_8
XFILLER_38_875 VPWR VGND sg13g2_decap_8
XFILLER_93_992 VPWR VGND sg13g2_decap_8
XFILLER_65_672 VPWR VGND sg13g2_decap_8
XFILLER_53_812 VPWR VGND sg13g2_decap_8
XFILLER_25_525 VPWR VGND sg13g2_decap_8
XFILLER_64_193 VPWR VGND sg13g2_decap_8
XFILLER_52_322 VPWR VGND sg13g2_decap_8
XFILLER_44_18 VPWR VGND sg13g2_decap_8
XFILLER_37_396 VPWR VGND sg13g2_decap_8
XFILLER_80_686 VPWR VGND sg13g2_decap_8
XFILLER_53_889 VPWR VGND sg13g2_decap_8
XFILLER_100_35 VPWR VGND sg13g2_decap_8
XFILLER_52_399 VPWR VGND sg13g2_decap_8
XFILLER_40_539 VPWR VGND sg13g2_decap_8
XFILLER_21_742 VPWR VGND sg13g2_decap_8
XFILLER_60_39 VPWR VGND sg13g2_decap_8
XFILLER_20_263 VPWR VGND sg13g2_decap_8
XFILLER_106_357 VPWR VGND sg13g2_decap_8
XFILLER_0_602 VPWR VGND sg13g2_decap_8
XFILLER_88_753 VPWR VGND sg13g2_decap_8
XFILLER_87_252 VPWR VGND sg13g2_decap_8
XFILLER_85_14 VPWR VGND sg13g2_decap_8
XFILLER_0_679 VPWR VGND sg13g2_decap_8
XFILLER_102_574 VPWR VGND sg13g2_decap_8
XFILLER_47_105 VPWR VGND sg13g2_decap_8
XFILLER_75_469 VPWR VGND sg13g2_decap_8
XFILLER_63_609 VPWR VGND sg13g2_decap_8
XFILLER_90_417 VPWR VGND sg13g2_decap_8
XFILLER_62_119 VPWR VGND sg13g2_decap_8
XFILLER_56_683 VPWR VGND sg13g2_decap_8
XFILLER_44_823 VPWR VGND sg13g2_decap_8
XFILLER_16_525 VPWR VGND sg13g2_decap_8
XFILLER_18_63 VPWR VGND sg13g2_decap_8
XFILLER_29_886 VPWR VGND sg13g2_decap_8
XFILLER_83_480 VPWR VGND sg13g2_decap_8
XFILLER_71_620 VPWR VGND sg13g2_decap_8
XFILLER_55_182 VPWR VGND sg13g2_decap_8
XFILLER_43_322 VPWR VGND sg13g2_decap_8
XFILLER_28_385 VPWR VGND sg13g2_decap_8
XFILLER_71_697 VPWR VGND sg13g2_decap_8
XFILLER_70_196 VPWR VGND sg13g2_decap_8
XFILLER_43_399 VPWR VGND sg13g2_decap_8
XFILLER_31_539 VPWR VGND sg13g2_decap_8
XFILLER_12_753 VPWR VGND sg13g2_decap_8
XFILLER_15_1028 VPWR VGND sg13g2_fill_1
XFILLER_34_95 VPWR VGND sg13g2_decap_8
XFILLER_8_735 VPWR VGND sg13g2_decap_8
XFILLER_11_252 VPWR VGND sg13g2_decap_8
XFILLER_7_256 VPWR VGND sg13g2_decap_8
XFILLER_4_952 VPWR VGND sg13g2_decap_8
XFILLER_3_462 VPWR VGND sg13g2_decap_8
XFILLER_79_753 VPWR VGND sg13g2_decap_8
XFILLER_78_230 VPWR VGND sg13g2_decap_8
XFILLER_61_1026 VPWR VGND sg13g2_fill_2
XFILLER_59_92 VPWR VGND sg13g2_decap_8
XFILLER_39_606 VPWR VGND sg13g2_decap_8
XFILLER_93_222 VPWR VGND sg13g2_decap_8
XFILLER_67_959 VPWR VGND sg13g2_decap_8
XFILLER_38_105 VPWR VGND sg13g2_decap_8
XFILLER_94_756 VPWR VGND sg13g2_decap_8
XFILLER_66_447 VPWR VGND sg13g2_decap_8
XFILLER_81_417 VPWR VGND sg13g2_decap_8
XFILLER_75_91 VPWR VGND sg13g2_decap_8
XFILLER_53_119 VPWR VGND sg13g2_decap_8
XFILLER_47_672 VPWR VGND sg13g2_decap_8
XFILLER_35_812 VPWR VGND sg13g2_decap_8
XFILLER_93_299 VPWR VGND sg13g2_decap_8
XFILLER_74_491 VPWR VGND sg13g2_decap_8
XFILLER_46_193 VPWR VGND sg13g2_decap_8
XFILLER_19_385 VPWR VGND sg13g2_decap_8
XFILLER_34_333 VPWR VGND sg13g2_decap_8
XFILLER_90_984 VPWR VGND sg13g2_decap_8
XFILLER_62_686 VPWR VGND sg13g2_decap_8
XFILLER_50_826 VPWR VGND sg13g2_decap_8
XFILLER_35_889 VPWR VGND sg13g2_decap_8
XFILLER_89_539 VPWR VGND sg13g2_decap_8
XFILLER_39_18 VPWR VGND sg13g2_decap_8
XFILLER_69_274 VPWR VGND sg13g2_decap_8
XFILLER_58_959 VPWR VGND sg13g2_decap_8
XFILLER_29_116 VPWR VGND sg13g2_decap_8
XFILLER_85_756 VPWR VGND sg13g2_decap_8
XFILLER_73_907 VPWR VGND sg13g2_decap_8
XFILLER_57_469 VPWR VGND sg13g2_decap_8
XFILLER_45_609 VPWR VGND sg13g2_decap_8
XFILLER_84_266 VPWR VGND sg13g2_decap_8
XFILLER_72_406 VPWR VGND sg13g2_decap_8
XFILLER_55_28 VPWR VGND sg13g2_decap_8
XFILLER_26_812 VPWR VGND sg13g2_decap_8
XFILLER_38_672 VPWR VGND sg13g2_decap_8
XFILLER_77_1022 VPWR VGND sg13g2_decap_8
XFILLER_25_322 VPWR VGND sg13g2_decap_8
XFILLER_37_193 VPWR VGND sg13g2_decap_8
XFILLER_81_984 VPWR VGND sg13g2_decap_8
XFILLER_26_889 VPWR VGND sg13g2_decap_8
XFILLER_80_483 VPWR VGND sg13g2_decap_8
XFILLER_53_686 VPWR VGND sg13g2_decap_8
XFILLER_41_826 VPWR VGND sg13g2_decap_8
XFILLER_13_539 VPWR VGND sg13g2_decap_8
XFILLER_25_399 VPWR VGND sg13g2_decap_8
XFILLER_52_196 VPWR VGND sg13g2_decap_8
XFILLER_40_336 VPWR VGND sg13g2_decap_8
XFILLER_84_1015 VPWR VGND sg13g2_decap_8
XFILLER_106_154 VPWR VGND sg13g2_decap_8
XFILLER_4_259 VPWR VGND sg13g2_decap_8
XFILLER_20_53 VPWR VGND sg13g2_decap_8
XFILLER_96_35 VPWR VGND sg13g2_decap_8
XFILLER_103_861 VPWR VGND sg13g2_decap_8
XFILLER_88_550 VPWR VGND sg13g2_decap_8
XFILLER_1_966 VPWR VGND sg13g2_decap_8
XFILLER_102_371 VPWR VGND sg13g2_decap_8
XFILLER_0_476 VPWR VGND sg13g2_decap_8
XFILLER_76_767 VPWR VGND sg13g2_decap_8
XFILLER_64_907 VPWR VGND sg13g2_decap_8
XFILLER_48_469 VPWR VGND sg13g2_decap_8
XFILLER_29_95 VPWR VGND sg13g2_decap_8
XFILLER_36_609 VPWR VGND sg13g2_decap_8
XFILLER_90_214 VPWR VGND sg13g2_decap_8
XFILLER_75_266 VPWR VGND sg13g2_decap_8
XFILLER_63_406 VPWR VGND sg13g2_decap_8
XFILLER_17_823 VPWR VGND sg13g2_decap_8
XFILLER_29_683 VPWR VGND sg13g2_decap_8
XFILLER_35_119 VPWR VGND sg13g2_decap_8
XFILLER_56_480 VPWR VGND sg13g2_decap_8
XFILLER_44_620 VPWR VGND sg13g2_decap_8
XFILLER_16_322 VPWR VGND sg13g2_decap_8
XFILLER_28_182 VPWR VGND sg13g2_decap_8
XFILLER_91_1008 VPWR VGND sg13g2_decap_8
XFILLER_72_973 VPWR VGND sg13g2_decap_8
XFILLER_71_494 VPWR VGND sg13g2_decap_8
XFILLER_44_697 VPWR VGND sg13g2_decap_8
XFILLER_16_399 VPWR VGND sg13g2_decap_8
XFILLER_32_837 VPWR VGND sg13g2_decap_8
XFILLER_43_196 VPWR VGND sg13g2_decap_8
XFILLER_31_336 VPWR VGND sg13g2_decap_8
XFILLER_12_550 VPWR VGND sg13g2_decap_8
XFILLER_77_7 VPWR VGND sg13g2_decap_8
XFILLER_8_532 VPWR VGND sg13g2_decap_8
XFILLER_99_826 VPWR VGND sg13g2_decap_8
XFILLER_6_77 VPWR VGND sg13g2_decap_8
XFILLER_98_347 VPWR VGND sg13g2_decap_8
XFILLER_100_308 VPWR VGND sg13g2_decap_8
XFILLER_79_550 VPWR VGND sg13g2_decap_8
XFILLER_6_1015 VPWR VGND sg13g2_decap_8
XFILLER_39_403 VPWR VGND sg13g2_decap_8
XFILLER_94_553 VPWR VGND sg13g2_decap_8
XFILLER_67_756 VPWR VGND sg13g2_decap_8
XFILLER_66_244 VPWR VGND sg13g2_decap_8
XFILLER_54_417 VPWR VGND sg13g2_decap_8
XFILLER_26_119 VPWR VGND sg13g2_decap_8
XFILLER_81_214 VPWR VGND sg13g2_decap_8
XFILLER_19_182 VPWR VGND sg13g2_decap_8
XFILLER_63_973 VPWR VGND sg13g2_decap_8
XFILLER_34_130 VPWR VGND sg13g2_decap_8
XFILLER_90_781 VPWR VGND sg13g2_decap_8
XFILLER_62_483 VPWR VGND sg13g2_decap_8
XFILLER_50_623 VPWR VGND sg13g2_decap_8
XFILLER_23_826 VPWR VGND sg13g2_decap_8
XFILLER_35_686 VPWR VGND sg13g2_decap_8
XFILLER_22_347 VPWR VGND sg13g2_decap_8
XFILLER_89_336 VPWR VGND sg13g2_decap_8
XFILLER_104_658 VPWR VGND sg13g2_decap_8
XFILLER_106_56 VPWR VGND sg13g2_decap_8
XFILLER_103_168 VPWR VGND sg13g2_decap_8
XFILLER_66_27 VPWR VGND sg13g2_decap_8
XFILLER_85_553 VPWR VGND sg13g2_decap_8
XFILLER_58_756 VPWR VGND sg13g2_decap_8
XFILLER_46_907 VPWR VGND sg13g2_decap_8
XFILLER_18_609 VPWR VGND sg13g2_decap_8
XFILLER_100_875 VPWR VGND sg13g2_decap_8
XFILLER_73_704 VPWR VGND sg13g2_decap_8
XFILLER_72_203 VPWR VGND sg13g2_decap_8
XFILLER_57_266 VPWR VGND sg13g2_decap_8
XFILLER_45_406 VPWR VGND sg13g2_decap_8
XFILLER_39_970 VPWR VGND sg13g2_decap_8
XFILLER_54_984 VPWR VGND sg13g2_decap_8
XFILLER_81_781 VPWR VGND sg13g2_decap_8
XFILLER_53_483 VPWR VGND sg13g2_decap_8
XFILLER_41_623 VPWR VGND sg13g2_decap_8
XFILLER_14_826 VPWR VGND sg13g2_decap_8
XFILLER_26_686 VPWR VGND sg13g2_decap_8
XFILLER_80_280 VPWR VGND sg13g2_decap_8
XFILLER_13_336 VPWR VGND sg13g2_decap_8
XFILLER_15_53 VPWR VGND sg13g2_decap_8
XFILLER_25_196 VPWR VGND sg13g2_decap_8
XFILLER_40_133 VPWR VGND sg13g2_decap_8
XFILLER_9_329 VPWR VGND sg13g2_decap_8
XFILLER_31_63 VPWR VGND sg13g2_decap_8
XFILLER_103_0 VPWR VGND sg13g2_decap_8
XFILLER_5_557 VPWR VGND sg13g2_decap_8
XFILLER_68_509 VPWR VGND sg13g2_decap_8
XFILLER_1_763 VPWR VGND sg13g2_decap_8
XFILLER_0_273 VPWR VGND sg13g2_decap_8
XFILLER_49_767 VPWR VGND sg13g2_decap_8
XFILLER_37_907 VPWR VGND sg13g2_decap_8
XFILLER_76_564 VPWR VGND sg13g2_decap_8
XFILLER_64_704 VPWR VGND sg13g2_decap_8
XFILLER_63_203 VPWR VGND sg13g2_decap_8
XFILLER_48_266 VPWR VGND sg13g2_decap_8
XFILLER_36_406 VPWR VGND sg13g2_decap_8
XFILLER_56_60 VPWR VGND sg13g2_decap_8
XFILLER_17_620 VPWR VGND sg13g2_decap_8
XFILLER_29_480 VPWR VGND sg13g2_decap_8
XFILLER_91_567 VPWR VGND sg13g2_decap_8
XFILLER_45_973 VPWR VGND sg13g2_decap_8
XFILLER_72_770 VPWR VGND sg13g2_decap_8
XFILLER_60_921 VPWR VGND sg13g2_decap_8
XFILLER_17_697 VPWR VGND sg13g2_decap_8
XFILLER_72_70 VPWR VGND sg13g2_decap_8
XFILLER_71_291 VPWR VGND sg13g2_decap_8
XFILLER_44_494 VPWR VGND sg13g2_decap_8
XFILLER_16_196 VPWR VGND sg13g2_decap_8
XFILLER_31_133 VPWR VGND sg13g2_decap_8
XFILLER_32_634 VPWR VGND sg13g2_decap_8
XFILLER_60_998 VPWR VGND sg13g2_decap_8
XFILLER_9_896 VPWR VGND sg13g2_decap_8
XFILLER_99_623 VPWR VGND sg13g2_decap_8
XFILLER_98_144 VPWR VGND sg13g2_decap_8
XFILLER_59_509 VPWR VGND sg13g2_decap_8
XFILLER_100_105 VPWR VGND sg13g2_decap_8
XFILLER_39_200 VPWR VGND sg13g2_decap_8
.ends

