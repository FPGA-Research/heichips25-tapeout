module heichips25_example_small (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net25;

 sg13g2_and2_1 _29_ (.A(net1),
    .B(net9),
    .X(_00_));
 sg13g2_and2_1 _30_ (.A(net2),
    .B(net10),
    .X(_01_));
 sg13g2_xor2_1 _31_ (.B(net10),
    .A(net2),
    .X(_02_));
 sg13g2_xor2_1 _32_ (.B(_02_),
    .A(_00_),
    .X(net18));
 sg13g2_a21oi_2 _33_ (.B1(_01_),
    .Y(_03_),
    .A2(_02_),
    .A1(_00_));
 sg13g2_and2_1 _34_ (.A(net3),
    .B(net11),
    .X(_04_));
 sg13g2_xnor2_1 _35_ (.Y(_05_),
    .A(net3),
    .B(net11));
 sg13g2_nor2_1 _36_ (.A(_03_),
    .B(_05_),
    .Y(_06_));
 sg13g2_xor2_1 _37_ (.B(_05_),
    .A(_03_),
    .X(net19));
 sg13g2_or2_1 _38_ (.X(_07_),
    .B(net12),
    .A(net4));
 sg13g2_and2_1 _39_ (.A(net4),
    .B(net12),
    .X(_08_));
 sg13g2_xor2_1 _40_ (.B(net12),
    .A(net4),
    .X(_09_));
 sg13g2_nor2_1 _41_ (.A(_04_),
    .B(_06_),
    .Y(_10_));
 sg13g2_xnor2_1 _42_ (.Y(net20),
    .A(_09_),
    .B(_10_));
 sg13g2_nand2b_1 _43_ (.Y(_11_),
    .B(_09_),
    .A_N(_05_));
 sg13g2_a21oi_1 _44_ (.A1(_04_),
    .A2(_07_),
    .Y(_12_),
    .B1(_08_));
 sg13g2_o21ai_1 _45_ (.B1(_12_),
    .Y(_13_),
    .A1(_03_),
    .A2(_11_));
 sg13g2_nand2_1 _46_ (.Y(_14_),
    .A(net5),
    .B(net13));
 sg13g2_xor2_1 _47_ (.B(net13),
    .A(net5),
    .X(_15_));
 sg13g2_inv_1 _48_ (.Y(_16_),
    .A(_15_));
 sg13g2_nand2_1 _49_ (.Y(_17_),
    .A(_13_),
    .B(_15_));
 sg13g2_xnor2_1 _50_ (.Y(net21),
    .A(_13_),
    .B(_16_));
 sg13g2_nor2_1 _51_ (.A(net6),
    .B(net14),
    .Y(_18_));
 sg13g2_xnor2_1 _52_ (.Y(_19_),
    .A(net6),
    .B(net14));
 sg13g2_nand2_1 _53_ (.Y(_20_),
    .A(_14_),
    .B(_17_));
 sg13g2_xnor2_1 _54_ (.Y(net22),
    .A(_19_),
    .B(_20_));
 sg13g2_nor2_1 _55_ (.A(_16_),
    .B(_19_),
    .Y(_21_));
 sg13g2_nor2_1 _56_ (.A(_14_),
    .B(_18_),
    .Y(_22_));
 sg13g2_a221oi_1 _57_ (.B2(_21_),
    .C1(_22_),
    .B1(_13_),
    .A1(net6),
    .Y(_23_),
    .A2(net14));
 sg13g2_nand2_1 _58_ (.Y(_24_),
    .A(net7),
    .B(net15));
 sg13g2_nor2_1 _59_ (.A(net7),
    .B(net15),
    .Y(_25_));
 sg13g2_xor2_1 _60_ (.B(net15),
    .A(net7),
    .X(_26_));
 sg13g2_xnor2_1 _61_ (.Y(net23),
    .A(_23_),
    .B(_26_));
 sg13g2_o21ai_1 _62_ (.B1(_24_),
    .Y(_27_),
    .A1(_23_),
    .A2(_25_));
 sg13g2_xnor2_1 _63_ (.Y(_28_),
    .A(net8),
    .B(net16));
 sg13g2_xnor2_1 _64_ (.Y(net24),
    .A(_27_),
    .B(_28_));
 sg13g2_xor2_1 _65_ (.B(net9),
    .A(net1),
    .X(net17));
 sg13g2_tielo heichips25_example_small_26 (.L_LO(net26));
 sg13g2_tielo heichips25_example_small_27 (.L_LO(net27));
 sg13g2_tielo heichips25_example_small_28 (.L_LO(net28));
 sg13g2_tielo heichips25_example_small_29 (.L_LO(net29));
 sg13g2_tielo heichips25_example_small_30 (.L_LO(net30));
 sg13g2_tielo heichips25_example_small_31 (.L_LO(net31));
 sg13g2_tielo heichips25_example_small_32 (.L_LO(net32));
 sg13g2_tielo heichips25_example_small_33 (.L_LO(net33));
 sg13g2_tielo heichips25_example_small_34 (.L_LO(net34));
 sg13g2_tielo heichips25_example_small_35 (.L_LO(net35));
 sg13g2_tielo heichips25_example_small_36 (.L_LO(net36));
 sg13g2_tielo heichips25_example_small_37 (.L_LO(net37));
 sg13g2_tielo heichips25_example_small_38 (.L_LO(net38));
 sg13g2_tielo heichips25_example_small_39 (.L_LO(net39));
 sg13g2_tielo heichips25_example_small_40 (.L_LO(net40));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[4]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[5]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(uio_in[6]),
    .X(net15));
 sg13g2_buf_1 input16 (.A(uio_in[7]),
    .X(net16));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[0]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[1]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[2]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[3]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[4]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[5]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[6]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[7]));
 sg13g2_tielo heichips25_example_small_25 (.L_LO(net25));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_decap_8 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_0_868 ();
 sg13g2_decap_8 FILLER_0_875 ();
 sg13g2_decap_8 FILLER_0_882 ();
 sg13g2_decap_8 FILLER_0_889 ();
 sg13g2_decap_8 FILLER_0_896 ();
 sg13g2_decap_8 FILLER_0_903 ();
 sg13g2_decap_8 FILLER_0_910 ();
 sg13g2_decap_8 FILLER_0_917 ();
 sg13g2_fill_1 FILLER_0_924 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_decap_8 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_1_868 ();
 sg13g2_decap_8 FILLER_1_875 ();
 sg13g2_decap_8 FILLER_1_882 ();
 sg13g2_decap_8 FILLER_1_889 ();
 sg13g2_decap_8 FILLER_1_896 ();
 sg13g2_decap_8 FILLER_1_903 ();
 sg13g2_decap_8 FILLER_1_910 ();
 sg13g2_decap_8 FILLER_1_917 ();
 sg13g2_fill_1 FILLER_1_924 ();
 sg13g2_decap_8 FILLER_2_4 ();
 sg13g2_decap_8 FILLER_2_11 ();
 sg13g2_decap_8 FILLER_2_18 ();
 sg13g2_decap_8 FILLER_2_25 ();
 sg13g2_decap_8 FILLER_2_32 ();
 sg13g2_decap_8 FILLER_2_39 ();
 sg13g2_decap_8 FILLER_2_46 ();
 sg13g2_decap_8 FILLER_2_53 ();
 sg13g2_decap_8 FILLER_2_60 ();
 sg13g2_decap_8 FILLER_2_67 ();
 sg13g2_decap_8 FILLER_2_74 ();
 sg13g2_decap_8 FILLER_2_81 ();
 sg13g2_decap_8 FILLER_2_88 ();
 sg13g2_decap_8 FILLER_2_95 ();
 sg13g2_decap_8 FILLER_2_102 ();
 sg13g2_decap_8 FILLER_2_109 ();
 sg13g2_decap_8 FILLER_2_116 ();
 sg13g2_decap_8 FILLER_2_123 ();
 sg13g2_decap_8 FILLER_2_130 ();
 sg13g2_decap_8 FILLER_2_137 ();
 sg13g2_decap_8 FILLER_2_144 ();
 sg13g2_decap_8 FILLER_2_151 ();
 sg13g2_decap_8 FILLER_2_158 ();
 sg13g2_decap_8 FILLER_2_165 ();
 sg13g2_decap_8 FILLER_2_172 ();
 sg13g2_decap_8 FILLER_2_179 ();
 sg13g2_decap_8 FILLER_2_186 ();
 sg13g2_decap_8 FILLER_2_193 ();
 sg13g2_decap_8 FILLER_2_200 ();
 sg13g2_decap_8 FILLER_2_207 ();
 sg13g2_decap_8 FILLER_2_214 ();
 sg13g2_decap_8 FILLER_2_221 ();
 sg13g2_decap_8 FILLER_2_228 ();
 sg13g2_decap_8 FILLER_2_235 ();
 sg13g2_decap_8 FILLER_2_242 ();
 sg13g2_decap_8 FILLER_2_249 ();
 sg13g2_decap_8 FILLER_2_256 ();
 sg13g2_decap_8 FILLER_2_263 ();
 sg13g2_decap_8 FILLER_2_270 ();
 sg13g2_decap_8 FILLER_2_277 ();
 sg13g2_decap_8 FILLER_2_284 ();
 sg13g2_decap_8 FILLER_2_291 ();
 sg13g2_decap_8 FILLER_2_298 ();
 sg13g2_decap_8 FILLER_2_305 ();
 sg13g2_decap_8 FILLER_2_312 ();
 sg13g2_decap_8 FILLER_2_319 ();
 sg13g2_decap_8 FILLER_2_326 ();
 sg13g2_decap_8 FILLER_2_333 ();
 sg13g2_decap_8 FILLER_2_340 ();
 sg13g2_decap_8 FILLER_2_347 ();
 sg13g2_decap_8 FILLER_2_354 ();
 sg13g2_decap_8 FILLER_2_361 ();
 sg13g2_decap_8 FILLER_2_368 ();
 sg13g2_decap_8 FILLER_2_375 ();
 sg13g2_decap_8 FILLER_2_382 ();
 sg13g2_decap_8 FILLER_2_389 ();
 sg13g2_decap_8 FILLER_2_396 ();
 sg13g2_decap_8 FILLER_2_403 ();
 sg13g2_decap_8 FILLER_2_410 ();
 sg13g2_decap_8 FILLER_2_417 ();
 sg13g2_decap_8 FILLER_2_424 ();
 sg13g2_decap_8 FILLER_2_431 ();
 sg13g2_decap_8 FILLER_2_438 ();
 sg13g2_decap_8 FILLER_2_445 ();
 sg13g2_decap_8 FILLER_2_452 ();
 sg13g2_decap_8 FILLER_2_459 ();
 sg13g2_decap_8 FILLER_2_466 ();
 sg13g2_decap_8 FILLER_2_473 ();
 sg13g2_decap_8 FILLER_2_480 ();
 sg13g2_decap_8 FILLER_2_487 ();
 sg13g2_decap_8 FILLER_2_494 ();
 sg13g2_decap_8 FILLER_2_501 ();
 sg13g2_decap_8 FILLER_2_508 ();
 sg13g2_decap_8 FILLER_2_515 ();
 sg13g2_decap_8 FILLER_2_522 ();
 sg13g2_decap_8 FILLER_2_529 ();
 sg13g2_decap_8 FILLER_2_536 ();
 sg13g2_decap_8 FILLER_2_543 ();
 sg13g2_decap_8 FILLER_2_550 ();
 sg13g2_decap_8 FILLER_2_557 ();
 sg13g2_decap_8 FILLER_2_564 ();
 sg13g2_decap_8 FILLER_2_571 ();
 sg13g2_decap_8 FILLER_2_578 ();
 sg13g2_decap_8 FILLER_2_585 ();
 sg13g2_decap_8 FILLER_2_592 ();
 sg13g2_decap_8 FILLER_2_599 ();
 sg13g2_decap_8 FILLER_2_606 ();
 sg13g2_decap_8 FILLER_2_613 ();
 sg13g2_decap_8 FILLER_2_620 ();
 sg13g2_decap_8 FILLER_2_627 ();
 sg13g2_decap_8 FILLER_2_634 ();
 sg13g2_decap_8 FILLER_2_641 ();
 sg13g2_decap_8 FILLER_2_648 ();
 sg13g2_decap_8 FILLER_2_655 ();
 sg13g2_decap_8 FILLER_2_662 ();
 sg13g2_decap_8 FILLER_2_669 ();
 sg13g2_decap_8 FILLER_2_676 ();
 sg13g2_decap_8 FILLER_2_683 ();
 sg13g2_decap_8 FILLER_2_690 ();
 sg13g2_decap_8 FILLER_2_697 ();
 sg13g2_decap_8 FILLER_2_704 ();
 sg13g2_decap_8 FILLER_2_711 ();
 sg13g2_decap_8 FILLER_2_718 ();
 sg13g2_decap_8 FILLER_2_725 ();
 sg13g2_decap_8 FILLER_2_732 ();
 sg13g2_decap_8 FILLER_2_739 ();
 sg13g2_decap_8 FILLER_2_746 ();
 sg13g2_decap_8 FILLER_2_753 ();
 sg13g2_decap_8 FILLER_2_760 ();
 sg13g2_decap_8 FILLER_2_767 ();
 sg13g2_decap_8 FILLER_2_774 ();
 sg13g2_decap_8 FILLER_2_781 ();
 sg13g2_decap_8 FILLER_2_788 ();
 sg13g2_decap_8 FILLER_2_795 ();
 sg13g2_decap_8 FILLER_2_802 ();
 sg13g2_decap_8 FILLER_2_809 ();
 sg13g2_decap_8 FILLER_2_816 ();
 sg13g2_decap_8 FILLER_2_823 ();
 sg13g2_decap_8 FILLER_2_830 ();
 sg13g2_decap_8 FILLER_2_837 ();
 sg13g2_decap_8 FILLER_2_844 ();
 sg13g2_decap_8 FILLER_2_851 ();
 sg13g2_decap_8 FILLER_2_858 ();
 sg13g2_decap_8 FILLER_2_865 ();
 sg13g2_decap_8 FILLER_2_872 ();
 sg13g2_decap_8 FILLER_2_879 ();
 sg13g2_decap_8 FILLER_2_886 ();
 sg13g2_decap_8 FILLER_2_893 ();
 sg13g2_decap_8 FILLER_2_900 ();
 sg13g2_decap_8 FILLER_2_907 ();
 sg13g2_decap_8 FILLER_2_914 ();
 sg13g2_decap_4 FILLER_2_921 ();
 sg13g2_decap_8 FILLER_3_4 ();
 sg13g2_decap_8 FILLER_3_11 ();
 sg13g2_decap_8 FILLER_3_18 ();
 sg13g2_decap_8 FILLER_3_25 ();
 sg13g2_decap_8 FILLER_3_32 ();
 sg13g2_decap_8 FILLER_3_39 ();
 sg13g2_decap_8 FILLER_3_46 ();
 sg13g2_decap_8 FILLER_3_53 ();
 sg13g2_decap_8 FILLER_3_60 ();
 sg13g2_decap_8 FILLER_3_67 ();
 sg13g2_decap_8 FILLER_3_74 ();
 sg13g2_decap_8 FILLER_3_81 ();
 sg13g2_decap_8 FILLER_3_88 ();
 sg13g2_decap_8 FILLER_3_95 ();
 sg13g2_decap_8 FILLER_3_102 ();
 sg13g2_decap_8 FILLER_3_109 ();
 sg13g2_decap_8 FILLER_3_116 ();
 sg13g2_decap_8 FILLER_3_123 ();
 sg13g2_decap_8 FILLER_3_130 ();
 sg13g2_decap_8 FILLER_3_137 ();
 sg13g2_decap_8 FILLER_3_144 ();
 sg13g2_decap_8 FILLER_3_151 ();
 sg13g2_decap_8 FILLER_3_158 ();
 sg13g2_decap_8 FILLER_3_165 ();
 sg13g2_decap_8 FILLER_3_172 ();
 sg13g2_decap_8 FILLER_3_179 ();
 sg13g2_decap_8 FILLER_3_186 ();
 sg13g2_decap_8 FILLER_3_193 ();
 sg13g2_decap_8 FILLER_3_200 ();
 sg13g2_decap_8 FILLER_3_207 ();
 sg13g2_decap_8 FILLER_3_214 ();
 sg13g2_decap_8 FILLER_3_221 ();
 sg13g2_decap_8 FILLER_3_228 ();
 sg13g2_decap_8 FILLER_3_235 ();
 sg13g2_decap_8 FILLER_3_242 ();
 sg13g2_decap_8 FILLER_3_249 ();
 sg13g2_decap_8 FILLER_3_256 ();
 sg13g2_decap_8 FILLER_3_263 ();
 sg13g2_decap_8 FILLER_3_270 ();
 sg13g2_decap_8 FILLER_3_277 ();
 sg13g2_decap_8 FILLER_3_284 ();
 sg13g2_decap_8 FILLER_3_291 ();
 sg13g2_decap_8 FILLER_3_298 ();
 sg13g2_decap_8 FILLER_3_305 ();
 sg13g2_decap_8 FILLER_3_312 ();
 sg13g2_decap_8 FILLER_3_319 ();
 sg13g2_decap_8 FILLER_3_326 ();
 sg13g2_decap_8 FILLER_3_333 ();
 sg13g2_decap_8 FILLER_3_340 ();
 sg13g2_decap_8 FILLER_3_347 ();
 sg13g2_decap_8 FILLER_3_354 ();
 sg13g2_decap_8 FILLER_3_361 ();
 sg13g2_decap_8 FILLER_3_368 ();
 sg13g2_decap_8 FILLER_3_375 ();
 sg13g2_decap_8 FILLER_3_382 ();
 sg13g2_decap_8 FILLER_3_389 ();
 sg13g2_decap_8 FILLER_3_396 ();
 sg13g2_decap_8 FILLER_3_403 ();
 sg13g2_decap_8 FILLER_3_410 ();
 sg13g2_decap_8 FILLER_3_417 ();
 sg13g2_decap_8 FILLER_3_424 ();
 sg13g2_decap_8 FILLER_3_431 ();
 sg13g2_decap_8 FILLER_3_438 ();
 sg13g2_decap_8 FILLER_3_445 ();
 sg13g2_decap_8 FILLER_3_452 ();
 sg13g2_decap_8 FILLER_3_459 ();
 sg13g2_decap_8 FILLER_3_466 ();
 sg13g2_decap_8 FILLER_3_473 ();
 sg13g2_decap_8 FILLER_3_480 ();
 sg13g2_decap_8 FILLER_3_487 ();
 sg13g2_decap_8 FILLER_3_494 ();
 sg13g2_decap_8 FILLER_3_501 ();
 sg13g2_decap_8 FILLER_3_508 ();
 sg13g2_decap_8 FILLER_3_515 ();
 sg13g2_decap_8 FILLER_3_522 ();
 sg13g2_decap_8 FILLER_3_529 ();
 sg13g2_decap_8 FILLER_3_536 ();
 sg13g2_decap_8 FILLER_3_543 ();
 sg13g2_decap_8 FILLER_3_550 ();
 sg13g2_decap_8 FILLER_3_557 ();
 sg13g2_decap_8 FILLER_3_564 ();
 sg13g2_decap_8 FILLER_3_571 ();
 sg13g2_decap_8 FILLER_3_578 ();
 sg13g2_decap_8 FILLER_3_585 ();
 sg13g2_decap_8 FILLER_3_592 ();
 sg13g2_decap_8 FILLER_3_599 ();
 sg13g2_decap_8 FILLER_3_606 ();
 sg13g2_decap_8 FILLER_3_613 ();
 sg13g2_decap_8 FILLER_3_620 ();
 sg13g2_decap_8 FILLER_3_627 ();
 sg13g2_decap_8 FILLER_3_634 ();
 sg13g2_decap_8 FILLER_3_641 ();
 sg13g2_decap_8 FILLER_3_648 ();
 sg13g2_decap_8 FILLER_3_655 ();
 sg13g2_decap_8 FILLER_3_662 ();
 sg13g2_decap_8 FILLER_3_669 ();
 sg13g2_decap_8 FILLER_3_676 ();
 sg13g2_decap_8 FILLER_3_683 ();
 sg13g2_decap_8 FILLER_3_690 ();
 sg13g2_decap_8 FILLER_3_697 ();
 sg13g2_decap_8 FILLER_3_704 ();
 sg13g2_decap_8 FILLER_3_711 ();
 sg13g2_decap_8 FILLER_3_718 ();
 sg13g2_decap_8 FILLER_3_725 ();
 sg13g2_decap_8 FILLER_3_732 ();
 sg13g2_decap_8 FILLER_3_739 ();
 sg13g2_decap_8 FILLER_3_746 ();
 sg13g2_decap_8 FILLER_3_753 ();
 sg13g2_decap_8 FILLER_3_760 ();
 sg13g2_decap_8 FILLER_3_767 ();
 sg13g2_decap_8 FILLER_3_774 ();
 sg13g2_decap_8 FILLER_3_781 ();
 sg13g2_decap_8 FILLER_3_788 ();
 sg13g2_decap_8 FILLER_3_795 ();
 sg13g2_decap_8 FILLER_3_802 ();
 sg13g2_decap_8 FILLER_3_809 ();
 sg13g2_decap_8 FILLER_3_816 ();
 sg13g2_decap_8 FILLER_3_823 ();
 sg13g2_decap_8 FILLER_3_830 ();
 sg13g2_decap_8 FILLER_3_837 ();
 sg13g2_decap_8 FILLER_3_844 ();
 sg13g2_decap_8 FILLER_3_851 ();
 sg13g2_decap_8 FILLER_3_858 ();
 sg13g2_decap_8 FILLER_3_865 ();
 sg13g2_decap_8 FILLER_3_872 ();
 sg13g2_decap_8 FILLER_3_879 ();
 sg13g2_decap_8 FILLER_3_886 ();
 sg13g2_decap_8 FILLER_3_893 ();
 sg13g2_decap_8 FILLER_3_900 ();
 sg13g2_decap_8 FILLER_3_907 ();
 sg13g2_decap_8 FILLER_3_914 ();
 sg13g2_decap_4 FILLER_3_921 ();
 sg13g2_decap_8 FILLER_4_4 ();
 sg13g2_decap_8 FILLER_4_11 ();
 sg13g2_decap_8 FILLER_4_18 ();
 sg13g2_decap_8 FILLER_4_25 ();
 sg13g2_decap_8 FILLER_4_32 ();
 sg13g2_decap_8 FILLER_4_39 ();
 sg13g2_decap_8 FILLER_4_46 ();
 sg13g2_decap_8 FILLER_4_53 ();
 sg13g2_decap_8 FILLER_4_60 ();
 sg13g2_decap_8 FILLER_4_67 ();
 sg13g2_decap_8 FILLER_4_74 ();
 sg13g2_decap_8 FILLER_4_81 ();
 sg13g2_decap_8 FILLER_4_88 ();
 sg13g2_decap_8 FILLER_4_95 ();
 sg13g2_decap_8 FILLER_4_102 ();
 sg13g2_decap_8 FILLER_4_109 ();
 sg13g2_decap_8 FILLER_4_116 ();
 sg13g2_decap_8 FILLER_4_123 ();
 sg13g2_decap_8 FILLER_4_130 ();
 sg13g2_decap_8 FILLER_4_137 ();
 sg13g2_decap_8 FILLER_4_144 ();
 sg13g2_decap_8 FILLER_4_151 ();
 sg13g2_decap_8 FILLER_4_158 ();
 sg13g2_decap_8 FILLER_4_165 ();
 sg13g2_decap_8 FILLER_4_172 ();
 sg13g2_decap_8 FILLER_4_179 ();
 sg13g2_decap_8 FILLER_4_186 ();
 sg13g2_decap_8 FILLER_4_193 ();
 sg13g2_decap_8 FILLER_4_200 ();
 sg13g2_decap_8 FILLER_4_207 ();
 sg13g2_decap_8 FILLER_4_214 ();
 sg13g2_decap_8 FILLER_4_221 ();
 sg13g2_decap_8 FILLER_4_228 ();
 sg13g2_decap_8 FILLER_4_235 ();
 sg13g2_decap_8 FILLER_4_242 ();
 sg13g2_decap_8 FILLER_4_249 ();
 sg13g2_decap_8 FILLER_4_256 ();
 sg13g2_decap_8 FILLER_4_263 ();
 sg13g2_decap_8 FILLER_4_270 ();
 sg13g2_decap_8 FILLER_4_277 ();
 sg13g2_decap_8 FILLER_4_284 ();
 sg13g2_decap_8 FILLER_4_291 ();
 sg13g2_decap_8 FILLER_4_298 ();
 sg13g2_decap_8 FILLER_4_305 ();
 sg13g2_decap_8 FILLER_4_312 ();
 sg13g2_decap_8 FILLER_4_319 ();
 sg13g2_decap_8 FILLER_4_326 ();
 sg13g2_decap_8 FILLER_4_333 ();
 sg13g2_decap_8 FILLER_4_340 ();
 sg13g2_decap_8 FILLER_4_347 ();
 sg13g2_decap_8 FILLER_4_354 ();
 sg13g2_decap_8 FILLER_4_361 ();
 sg13g2_decap_8 FILLER_4_368 ();
 sg13g2_decap_8 FILLER_4_375 ();
 sg13g2_decap_8 FILLER_4_382 ();
 sg13g2_decap_8 FILLER_4_389 ();
 sg13g2_decap_8 FILLER_4_396 ();
 sg13g2_decap_8 FILLER_4_403 ();
 sg13g2_decap_8 FILLER_4_410 ();
 sg13g2_decap_8 FILLER_4_417 ();
 sg13g2_decap_8 FILLER_4_424 ();
 sg13g2_decap_8 FILLER_4_431 ();
 sg13g2_decap_8 FILLER_4_438 ();
 sg13g2_decap_8 FILLER_4_445 ();
 sg13g2_decap_8 FILLER_4_452 ();
 sg13g2_decap_8 FILLER_4_459 ();
 sg13g2_decap_8 FILLER_4_466 ();
 sg13g2_decap_8 FILLER_4_473 ();
 sg13g2_decap_8 FILLER_4_480 ();
 sg13g2_decap_8 FILLER_4_487 ();
 sg13g2_decap_8 FILLER_4_494 ();
 sg13g2_decap_8 FILLER_4_501 ();
 sg13g2_decap_8 FILLER_4_508 ();
 sg13g2_decap_8 FILLER_4_515 ();
 sg13g2_decap_8 FILLER_4_522 ();
 sg13g2_decap_8 FILLER_4_529 ();
 sg13g2_decap_8 FILLER_4_536 ();
 sg13g2_decap_8 FILLER_4_543 ();
 sg13g2_decap_8 FILLER_4_550 ();
 sg13g2_decap_8 FILLER_4_557 ();
 sg13g2_decap_8 FILLER_4_564 ();
 sg13g2_decap_8 FILLER_4_571 ();
 sg13g2_decap_8 FILLER_4_578 ();
 sg13g2_decap_8 FILLER_4_585 ();
 sg13g2_decap_8 FILLER_4_592 ();
 sg13g2_decap_8 FILLER_4_599 ();
 sg13g2_decap_8 FILLER_4_606 ();
 sg13g2_decap_8 FILLER_4_613 ();
 sg13g2_decap_8 FILLER_4_620 ();
 sg13g2_decap_8 FILLER_4_627 ();
 sg13g2_decap_8 FILLER_4_634 ();
 sg13g2_decap_8 FILLER_4_641 ();
 sg13g2_decap_8 FILLER_4_648 ();
 sg13g2_decap_8 FILLER_4_655 ();
 sg13g2_decap_8 FILLER_4_662 ();
 sg13g2_decap_8 FILLER_4_669 ();
 sg13g2_decap_8 FILLER_4_676 ();
 sg13g2_decap_8 FILLER_4_683 ();
 sg13g2_decap_8 FILLER_4_690 ();
 sg13g2_decap_8 FILLER_4_697 ();
 sg13g2_decap_8 FILLER_4_704 ();
 sg13g2_decap_8 FILLER_4_711 ();
 sg13g2_decap_8 FILLER_4_718 ();
 sg13g2_decap_8 FILLER_4_725 ();
 sg13g2_decap_8 FILLER_4_732 ();
 sg13g2_decap_8 FILLER_4_739 ();
 sg13g2_decap_8 FILLER_4_746 ();
 sg13g2_decap_8 FILLER_4_753 ();
 sg13g2_decap_8 FILLER_4_760 ();
 sg13g2_decap_8 FILLER_4_767 ();
 sg13g2_decap_8 FILLER_4_774 ();
 sg13g2_decap_8 FILLER_4_781 ();
 sg13g2_decap_8 FILLER_4_788 ();
 sg13g2_decap_8 FILLER_4_795 ();
 sg13g2_decap_8 FILLER_4_802 ();
 sg13g2_decap_8 FILLER_4_809 ();
 sg13g2_decap_8 FILLER_4_816 ();
 sg13g2_decap_8 FILLER_4_823 ();
 sg13g2_decap_8 FILLER_4_830 ();
 sg13g2_decap_8 FILLER_4_837 ();
 sg13g2_decap_8 FILLER_4_844 ();
 sg13g2_decap_8 FILLER_4_851 ();
 sg13g2_decap_8 FILLER_4_858 ();
 sg13g2_decap_8 FILLER_4_865 ();
 sg13g2_decap_8 FILLER_4_872 ();
 sg13g2_decap_8 FILLER_4_879 ();
 sg13g2_decap_8 FILLER_4_886 ();
 sg13g2_decap_8 FILLER_4_893 ();
 sg13g2_decap_8 FILLER_4_900 ();
 sg13g2_decap_8 FILLER_4_907 ();
 sg13g2_decap_8 FILLER_4_914 ();
 sg13g2_decap_4 FILLER_4_921 ();
 sg13g2_decap_8 FILLER_5_4 ();
 sg13g2_decap_8 FILLER_5_11 ();
 sg13g2_decap_8 FILLER_5_18 ();
 sg13g2_decap_8 FILLER_5_25 ();
 sg13g2_decap_8 FILLER_5_32 ();
 sg13g2_decap_8 FILLER_5_39 ();
 sg13g2_decap_8 FILLER_5_46 ();
 sg13g2_decap_8 FILLER_5_53 ();
 sg13g2_decap_8 FILLER_5_60 ();
 sg13g2_decap_8 FILLER_5_67 ();
 sg13g2_decap_8 FILLER_5_74 ();
 sg13g2_decap_8 FILLER_5_81 ();
 sg13g2_decap_8 FILLER_5_88 ();
 sg13g2_decap_8 FILLER_5_95 ();
 sg13g2_decap_8 FILLER_5_102 ();
 sg13g2_decap_8 FILLER_5_109 ();
 sg13g2_decap_8 FILLER_5_116 ();
 sg13g2_decap_8 FILLER_5_123 ();
 sg13g2_decap_8 FILLER_5_130 ();
 sg13g2_decap_8 FILLER_5_137 ();
 sg13g2_decap_8 FILLER_5_144 ();
 sg13g2_decap_8 FILLER_5_151 ();
 sg13g2_decap_8 FILLER_5_158 ();
 sg13g2_decap_8 FILLER_5_165 ();
 sg13g2_decap_8 FILLER_5_172 ();
 sg13g2_decap_8 FILLER_5_179 ();
 sg13g2_decap_8 FILLER_5_186 ();
 sg13g2_decap_8 FILLER_5_193 ();
 sg13g2_decap_8 FILLER_5_200 ();
 sg13g2_decap_8 FILLER_5_207 ();
 sg13g2_decap_8 FILLER_5_214 ();
 sg13g2_decap_8 FILLER_5_221 ();
 sg13g2_decap_8 FILLER_5_228 ();
 sg13g2_decap_8 FILLER_5_235 ();
 sg13g2_decap_8 FILLER_5_242 ();
 sg13g2_decap_8 FILLER_5_249 ();
 sg13g2_decap_8 FILLER_5_256 ();
 sg13g2_decap_8 FILLER_5_263 ();
 sg13g2_decap_8 FILLER_5_270 ();
 sg13g2_decap_8 FILLER_5_277 ();
 sg13g2_decap_8 FILLER_5_284 ();
 sg13g2_decap_8 FILLER_5_291 ();
 sg13g2_decap_8 FILLER_5_298 ();
 sg13g2_decap_8 FILLER_5_305 ();
 sg13g2_decap_8 FILLER_5_312 ();
 sg13g2_decap_8 FILLER_5_319 ();
 sg13g2_decap_8 FILLER_5_326 ();
 sg13g2_decap_8 FILLER_5_333 ();
 sg13g2_decap_8 FILLER_5_340 ();
 sg13g2_decap_8 FILLER_5_347 ();
 sg13g2_decap_8 FILLER_5_354 ();
 sg13g2_decap_8 FILLER_5_361 ();
 sg13g2_decap_8 FILLER_5_368 ();
 sg13g2_decap_8 FILLER_5_375 ();
 sg13g2_decap_8 FILLER_5_382 ();
 sg13g2_decap_8 FILLER_5_389 ();
 sg13g2_decap_8 FILLER_5_396 ();
 sg13g2_decap_8 FILLER_5_403 ();
 sg13g2_decap_8 FILLER_5_410 ();
 sg13g2_decap_8 FILLER_5_417 ();
 sg13g2_decap_8 FILLER_5_424 ();
 sg13g2_decap_8 FILLER_5_431 ();
 sg13g2_decap_8 FILLER_5_438 ();
 sg13g2_decap_8 FILLER_5_445 ();
 sg13g2_decap_8 FILLER_5_452 ();
 sg13g2_decap_8 FILLER_5_459 ();
 sg13g2_decap_8 FILLER_5_466 ();
 sg13g2_decap_8 FILLER_5_473 ();
 sg13g2_decap_8 FILLER_5_480 ();
 sg13g2_decap_8 FILLER_5_487 ();
 sg13g2_decap_8 FILLER_5_494 ();
 sg13g2_decap_8 FILLER_5_501 ();
 sg13g2_decap_8 FILLER_5_508 ();
 sg13g2_decap_8 FILLER_5_515 ();
 sg13g2_decap_8 FILLER_5_522 ();
 sg13g2_decap_8 FILLER_5_529 ();
 sg13g2_decap_8 FILLER_5_536 ();
 sg13g2_decap_8 FILLER_5_543 ();
 sg13g2_decap_8 FILLER_5_550 ();
 sg13g2_decap_8 FILLER_5_557 ();
 sg13g2_decap_8 FILLER_5_564 ();
 sg13g2_decap_8 FILLER_5_571 ();
 sg13g2_decap_8 FILLER_5_578 ();
 sg13g2_decap_8 FILLER_5_585 ();
 sg13g2_decap_8 FILLER_5_592 ();
 sg13g2_decap_8 FILLER_5_599 ();
 sg13g2_decap_8 FILLER_5_606 ();
 sg13g2_decap_8 FILLER_5_613 ();
 sg13g2_decap_8 FILLER_5_620 ();
 sg13g2_decap_8 FILLER_5_627 ();
 sg13g2_decap_8 FILLER_5_634 ();
 sg13g2_decap_8 FILLER_5_641 ();
 sg13g2_decap_8 FILLER_5_648 ();
 sg13g2_decap_8 FILLER_5_655 ();
 sg13g2_decap_8 FILLER_5_662 ();
 sg13g2_decap_8 FILLER_5_669 ();
 sg13g2_decap_8 FILLER_5_676 ();
 sg13g2_decap_8 FILLER_5_683 ();
 sg13g2_decap_8 FILLER_5_690 ();
 sg13g2_decap_8 FILLER_5_697 ();
 sg13g2_decap_8 FILLER_5_704 ();
 sg13g2_decap_8 FILLER_5_711 ();
 sg13g2_decap_8 FILLER_5_718 ();
 sg13g2_decap_8 FILLER_5_725 ();
 sg13g2_decap_8 FILLER_5_732 ();
 sg13g2_decap_8 FILLER_5_739 ();
 sg13g2_decap_8 FILLER_5_746 ();
 sg13g2_decap_8 FILLER_5_753 ();
 sg13g2_decap_8 FILLER_5_760 ();
 sg13g2_decap_8 FILLER_5_767 ();
 sg13g2_decap_8 FILLER_5_774 ();
 sg13g2_decap_8 FILLER_5_781 ();
 sg13g2_decap_8 FILLER_5_788 ();
 sg13g2_decap_8 FILLER_5_795 ();
 sg13g2_decap_8 FILLER_5_802 ();
 sg13g2_decap_8 FILLER_5_809 ();
 sg13g2_decap_8 FILLER_5_816 ();
 sg13g2_decap_8 FILLER_5_823 ();
 sg13g2_decap_8 FILLER_5_830 ();
 sg13g2_decap_8 FILLER_5_837 ();
 sg13g2_decap_8 FILLER_5_844 ();
 sg13g2_decap_8 FILLER_5_851 ();
 sg13g2_decap_8 FILLER_5_858 ();
 sg13g2_decap_8 FILLER_5_865 ();
 sg13g2_decap_8 FILLER_5_872 ();
 sg13g2_decap_8 FILLER_5_879 ();
 sg13g2_decap_8 FILLER_5_886 ();
 sg13g2_decap_8 FILLER_5_893 ();
 sg13g2_decap_8 FILLER_5_900 ();
 sg13g2_decap_8 FILLER_5_907 ();
 sg13g2_decap_8 FILLER_5_914 ();
 sg13g2_decap_4 FILLER_5_921 ();
 sg13g2_decap_8 FILLER_6_4 ();
 sg13g2_decap_8 FILLER_6_11 ();
 sg13g2_decap_8 FILLER_6_18 ();
 sg13g2_decap_8 FILLER_6_25 ();
 sg13g2_decap_8 FILLER_6_32 ();
 sg13g2_decap_8 FILLER_6_39 ();
 sg13g2_decap_8 FILLER_6_46 ();
 sg13g2_decap_8 FILLER_6_53 ();
 sg13g2_decap_8 FILLER_6_60 ();
 sg13g2_decap_8 FILLER_6_67 ();
 sg13g2_decap_8 FILLER_6_74 ();
 sg13g2_decap_8 FILLER_6_81 ();
 sg13g2_decap_8 FILLER_6_88 ();
 sg13g2_decap_8 FILLER_6_95 ();
 sg13g2_decap_8 FILLER_6_102 ();
 sg13g2_decap_8 FILLER_6_109 ();
 sg13g2_decap_8 FILLER_6_116 ();
 sg13g2_decap_8 FILLER_6_123 ();
 sg13g2_decap_8 FILLER_6_130 ();
 sg13g2_decap_8 FILLER_6_137 ();
 sg13g2_decap_8 FILLER_6_144 ();
 sg13g2_decap_8 FILLER_6_151 ();
 sg13g2_decap_8 FILLER_6_158 ();
 sg13g2_decap_8 FILLER_6_165 ();
 sg13g2_decap_8 FILLER_6_172 ();
 sg13g2_decap_8 FILLER_6_179 ();
 sg13g2_decap_8 FILLER_6_186 ();
 sg13g2_decap_8 FILLER_6_193 ();
 sg13g2_decap_8 FILLER_6_200 ();
 sg13g2_decap_8 FILLER_6_207 ();
 sg13g2_decap_8 FILLER_6_214 ();
 sg13g2_decap_8 FILLER_6_221 ();
 sg13g2_decap_8 FILLER_6_228 ();
 sg13g2_decap_8 FILLER_6_235 ();
 sg13g2_decap_8 FILLER_6_242 ();
 sg13g2_decap_8 FILLER_6_249 ();
 sg13g2_decap_8 FILLER_6_256 ();
 sg13g2_decap_8 FILLER_6_263 ();
 sg13g2_decap_8 FILLER_6_270 ();
 sg13g2_decap_8 FILLER_6_277 ();
 sg13g2_decap_8 FILLER_6_284 ();
 sg13g2_decap_8 FILLER_6_291 ();
 sg13g2_decap_8 FILLER_6_298 ();
 sg13g2_decap_8 FILLER_6_305 ();
 sg13g2_decap_8 FILLER_6_312 ();
 sg13g2_decap_8 FILLER_6_319 ();
 sg13g2_decap_8 FILLER_6_326 ();
 sg13g2_decap_8 FILLER_6_333 ();
 sg13g2_decap_8 FILLER_6_340 ();
 sg13g2_decap_8 FILLER_6_347 ();
 sg13g2_decap_8 FILLER_6_354 ();
 sg13g2_decap_8 FILLER_6_361 ();
 sg13g2_decap_8 FILLER_6_368 ();
 sg13g2_decap_8 FILLER_6_375 ();
 sg13g2_decap_8 FILLER_6_382 ();
 sg13g2_decap_8 FILLER_6_389 ();
 sg13g2_decap_8 FILLER_6_396 ();
 sg13g2_decap_8 FILLER_6_403 ();
 sg13g2_decap_8 FILLER_6_410 ();
 sg13g2_decap_8 FILLER_6_417 ();
 sg13g2_decap_8 FILLER_6_424 ();
 sg13g2_decap_8 FILLER_6_431 ();
 sg13g2_decap_8 FILLER_6_438 ();
 sg13g2_decap_8 FILLER_6_445 ();
 sg13g2_decap_8 FILLER_6_452 ();
 sg13g2_decap_8 FILLER_6_459 ();
 sg13g2_decap_8 FILLER_6_466 ();
 sg13g2_decap_8 FILLER_6_473 ();
 sg13g2_decap_8 FILLER_6_480 ();
 sg13g2_decap_8 FILLER_6_487 ();
 sg13g2_decap_8 FILLER_6_494 ();
 sg13g2_decap_8 FILLER_6_501 ();
 sg13g2_decap_8 FILLER_6_508 ();
 sg13g2_decap_8 FILLER_6_515 ();
 sg13g2_decap_8 FILLER_6_522 ();
 sg13g2_decap_8 FILLER_6_529 ();
 sg13g2_decap_8 FILLER_6_536 ();
 sg13g2_decap_8 FILLER_6_543 ();
 sg13g2_decap_8 FILLER_6_550 ();
 sg13g2_decap_8 FILLER_6_557 ();
 sg13g2_decap_8 FILLER_6_564 ();
 sg13g2_decap_8 FILLER_6_571 ();
 sg13g2_decap_8 FILLER_6_578 ();
 sg13g2_decap_8 FILLER_6_585 ();
 sg13g2_decap_8 FILLER_6_592 ();
 sg13g2_decap_8 FILLER_6_599 ();
 sg13g2_decap_8 FILLER_6_606 ();
 sg13g2_decap_8 FILLER_6_613 ();
 sg13g2_decap_8 FILLER_6_620 ();
 sg13g2_decap_8 FILLER_6_627 ();
 sg13g2_decap_8 FILLER_6_634 ();
 sg13g2_decap_8 FILLER_6_641 ();
 sg13g2_decap_8 FILLER_6_648 ();
 sg13g2_decap_8 FILLER_6_655 ();
 sg13g2_decap_8 FILLER_6_662 ();
 sg13g2_decap_8 FILLER_6_669 ();
 sg13g2_decap_8 FILLER_6_676 ();
 sg13g2_decap_8 FILLER_6_683 ();
 sg13g2_decap_8 FILLER_6_690 ();
 sg13g2_decap_8 FILLER_6_697 ();
 sg13g2_decap_8 FILLER_6_704 ();
 sg13g2_decap_8 FILLER_6_711 ();
 sg13g2_decap_8 FILLER_6_718 ();
 sg13g2_decap_8 FILLER_6_725 ();
 sg13g2_decap_8 FILLER_6_732 ();
 sg13g2_decap_8 FILLER_6_739 ();
 sg13g2_decap_8 FILLER_6_746 ();
 sg13g2_decap_8 FILLER_6_753 ();
 sg13g2_decap_8 FILLER_6_760 ();
 sg13g2_decap_8 FILLER_6_767 ();
 sg13g2_decap_8 FILLER_6_774 ();
 sg13g2_decap_8 FILLER_6_781 ();
 sg13g2_decap_8 FILLER_6_788 ();
 sg13g2_decap_8 FILLER_6_795 ();
 sg13g2_decap_8 FILLER_6_802 ();
 sg13g2_decap_8 FILLER_6_809 ();
 sg13g2_decap_8 FILLER_6_816 ();
 sg13g2_decap_8 FILLER_6_823 ();
 sg13g2_decap_8 FILLER_6_830 ();
 sg13g2_decap_8 FILLER_6_837 ();
 sg13g2_decap_8 FILLER_6_844 ();
 sg13g2_decap_8 FILLER_6_851 ();
 sg13g2_decap_8 FILLER_6_858 ();
 sg13g2_decap_8 FILLER_6_865 ();
 sg13g2_decap_8 FILLER_6_872 ();
 sg13g2_decap_8 FILLER_6_879 ();
 sg13g2_decap_8 FILLER_6_886 ();
 sg13g2_decap_8 FILLER_6_893 ();
 sg13g2_decap_8 FILLER_6_900 ();
 sg13g2_decap_8 FILLER_6_907 ();
 sg13g2_decap_8 FILLER_6_914 ();
 sg13g2_decap_4 FILLER_6_921 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_133 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_decap_8 FILLER_7_154 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_8 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_175 ();
 sg13g2_decap_8 FILLER_7_182 ();
 sg13g2_decap_8 FILLER_7_189 ();
 sg13g2_decap_8 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_8 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_224 ();
 sg13g2_decap_8 FILLER_7_231 ();
 sg13g2_decap_8 FILLER_7_238 ();
 sg13g2_decap_8 FILLER_7_245 ();
 sg13g2_decap_8 FILLER_7_252 ();
 sg13g2_decap_8 FILLER_7_259 ();
 sg13g2_decap_8 FILLER_7_266 ();
 sg13g2_decap_8 FILLER_7_273 ();
 sg13g2_decap_8 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_287 ();
 sg13g2_decap_8 FILLER_7_294 ();
 sg13g2_decap_8 FILLER_7_301 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_decap_8 FILLER_7_448 ();
 sg13g2_decap_8 FILLER_7_455 ();
 sg13g2_decap_8 FILLER_7_462 ();
 sg13g2_decap_8 FILLER_7_469 ();
 sg13g2_decap_8 FILLER_7_476 ();
 sg13g2_decap_8 FILLER_7_483 ();
 sg13g2_decap_8 FILLER_7_490 ();
 sg13g2_decap_8 FILLER_7_497 ();
 sg13g2_decap_8 FILLER_7_504 ();
 sg13g2_decap_8 FILLER_7_511 ();
 sg13g2_decap_8 FILLER_7_518 ();
 sg13g2_decap_8 FILLER_7_525 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_553 ();
 sg13g2_decap_8 FILLER_7_560 ();
 sg13g2_decap_8 FILLER_7_567 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_8 FILLER_7_581 ();
 sg13g2_decap_8 FILLER_7_588 ();
 sg13g2_decap_8 FILLER_7_595 ();
 sg13g2_decap_8 FILLER_7_602 ();
 sg13g2_decap_8 FILLER_7_609 ();
 sg13g2_decap_8 FILLER_7_616 ();
 sg13g2_decap_8 FILLER_7_623 ();
 sg13g2_decap_8 FILLER_7_630 ();
 sg13g2_decap_8 FILLER_7_637 ();
 sg13g2_decap_8 FILLER_7_644 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_decap_8 FILLER_7_658 ();
 sg13g2_decap_8 FILLER_7_665 ();
 sg13g2_decap_8 FILLER_7_672 ();
 sg13g2_decap_8 FILLER_7_679 ();
 sg13g2_decap_8 FILLER_7_686 ();
 sg13g2_decap_8 FILLER_7_693 ();
 sg13g2_decap_8 FILLER_7_700 ();
 sg13g2_decap_8 FILLER_7_707 ();
 sg13g2_decap_8 FILLER_7_714 ();
 sg13g2_decap_8 FILLER_7_721 ();
 sg13g2_decap_8 FILLER_7_728 ();
 sg13g2_decap_8 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_742 ();
 sg13g2_decap_8 FILLER_7_749 ();
 sg13g2_decap_8 FILLER_7_756 ();
 sg13g2_decap_8 FILLER_7_763 ();
 sg13g2_decap_8 FILLER_7_770 ();
 sg13g2_decap_8 FILLER_7_777 ();
 sg13g2_decap_8 FILLER_7_784 ();
 sg13g2_decap_8 FILLER_7_791 ();
 sg13g2_decap_8 FILLER_7_798 ();
 sg13g2_decap_8 FILLER_7_805 ();
 sg13g2_decap_8 FILLER_7_812 ();
 sg13g2_decap_8 FILLER_7_819 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_decap_8 FILLER_7_833 ();
 sg13g2_decap_8 FILLER_7_840 ();
 sg13g2_decap_8 FILLER_7_847 ();
 sg13g2_decap_8 FILLER_7_854 ();
 sg13g2_decap_8 FILLER_7_861 ();
 sg13g2_decap_8 FILLER_7_868 ();
 sg13g2_decap_8 FILLER_7_875 ();
 sg13g2_decap_8 FILLER_7_882 ();
 sg13g2_decap_8 FILLER_7_889 ();
 sg13g2_decap_8 FILLER_7_896 ();
 sg13g2_decap_8 FILLER_7_903 ();
 sg13g2_decap_8 FILLER_7_910 ();
 sg13g2_decap_8 FILLER_7_917 ();
 sg13g2_fill_1 FILLER_7_924 ();
 sg13g2_decap_8 FILLER_8_4 ();
 sg13g2_decap_8 FILLER_8_11 ();
 sg13g2_decap_8 FILLER_8_18 ();
 sg13g2_decap_8 FILLER_8_25 ();
 sg13g2_decap_8 FILLER_8_32 ();
 sg13g2_decap_8 FILLER_8_39 ();
 sg13g2_decap_8 FILLER_8_46 ();
 sg13g2_decap_8 FILLER_8_53 ();
 sg13g2_decap_8 FILLER_8_60 ();
 sg13g2_decap_8 FILLER_8_67 ();
 sg13g2_decap_8 FILLER_8_74 ();
 sg13g2_decap_8 FILLER_8_81 ();
 sg13g2_decap_8 FILLER_8_88 ();
 sg13g2_decap_8 FILLER_8_95 ();
 sg13g2_decap_8 FILLER_8_102 ();
 sg13g2_decap_8 FILLER_8_109 ();
 sg13g2_decap_8 FILLER_8_116 ();
 sg13g2_decap_8 FILLER_8_123 ();
 sg13g2_decap_8 FILLER_8_130 ();
 sg13g2_decap_8 FILLER_8_137 ();
 sg13g2_decap_8 FILLER_8_144 ();
 sg13g2_decap_8 FILLER_8_151 ();
 sg13g2_decap_8 FILLER_8_158 ();
 sg13g2_decap_8 FILLER_8_165 ();
 sg13g2_decap_8 FILLER_8_172 ();
 sg13g2_decap_8 FILLER_8_179 ();
 sg13g2_decap_8 FILLER_8_186 ();
 sg13g2_decap_8 FILLER_8_193 ();
 sg13g2_decap_8 FILLER_8_200 ();
 sg13g2_decap_8 FILLER_8_207 ();
 sg13g2_decap_8 FILLER_8_214 ();
 sg13g2_decap_8 FILLER_8_221 ();
 sg13g2_decap_8 FILLER_8_228 ();
 sg13g2_decap_8 FILLER_8_235 ();
 sg13g2_decap_8 FILLER_8_242 ();
 sg13g2_decap_8 FILLER_8_249 ();
 sg13g2_decap_8 FILLER_8_256 ();
 sg13g2_decap_8 FILLER_8_263 ();
 sg13g2_decap_8 FILLER_8_270 ();
 sg13g2_decap_8 FILLER_8_277 ();
 sg13g2_decap_8 FILLER_8_284 ();
 sg13g2_decap_8 FILLER_8_291 ();
 sg13g2_decap_8 FILLER_8_298 ();
 sg13g2_decap_8 FILLER_8_305 ();
 sg13g2_decap_8 FILLER_8_312 ();
 sg13g2_decap_8 FILLER_8_319 ();
 sg13g2_decap_8 FILLER_8_326 ();
 sg13g2_decap_8 FILLER_8_333 ();
 sg13g2_decap_8 FILLER_8_340 ();
 sg13g2_decap_8 FILLER_8_347 ();
 sg13g2_decap_8 FILLER_8_354 ();
 sg13g2_decap_8 FILLER_8_361 ();
 sg13g2_decap_8 FILLER_8_368 ();
 sg13g2_decap_8 FILLER_8_375 ();
 sg13g2_decap_8 FILLER_8_382 ();
 sg13g2_decap_8 FILLER_8_389 ();
 sg13g2_decap_8 FILLER_8_396 ();
 sg13g2_decap_8 FILLER_8_403 ();
 sg13g2_decap_8 FILLER_8_410 ();
 sg13g2_decap_8 FILLER_8_417 ();
 sg13g2_decap_8 FILLER_8_424 ();
 sg13g2_decap_8 FILLER_8_431 ();
 sg13g2_decap_8 FILLER_8_438 ();
 sg13g2_decap_8 FILLER_8_445 ();
 sg13g2_decap_8 FILLER_8_452 ();
 sg13g2_decap_8 FILLER_8_459 ();
 sg13g2_decap_8 FILLER_8_466 ();
 sg13g2_decap_8 FILLER_8_473 ();
 sg13g2_decap_8 FILLER_8_480 ();
 sg13g2_decap_8 FILLER_8_487 ();
 sg13g2_decap_8 FILLER_8_494 ();
 sg13g2_decap_8 FILLER_8_501 ();
 sg13g2_decap_8 FILLER_8_508 ();
 sg13g2_decap_8 FILLER_8_515 ();
 sg13g2_decap_8 FILLER_8_522 ();
 sg13g2_decap_8 FILLER_8_529 ();
 sg13g2_decap_8 FILLER_8_536 ();
 sg13g2_decap_8 FILLER_8_543 ();
 sg13g2_decap_8 FILLER_8_550 ();
 sg13g2_decap_8 FILLER_8_557 ();
 sg13g2_decap_8 FILLER_8_564 ();
 sg13g2_decap_8 FILLER_8_571 ();
 sg13g2_decap_8 FILLER_8_578 ();
 sg13g2_decap_8 FILLER_8_585 ();
 sg13g2_decap_8 FILLER_8_592 ();
 sg13g2_decap_8 FILLER_8_599 ();
 sg13g2_decap_8 FILLER_8_606 ();
 sg13g2_decap_8 FILLER_8_613 ();
 sg13g2_decap_8 FILLER_8_620 ();
 sg13g2_decap_8 FILLER_8_627 ();
 sg13g2_decap_8 FILLER_8_634 ();
 sg13g2_decap_8 FILLER_8_641 ();
 sg13g2_decap_8 FILLER_8_648 ();
 sg13g2_decap_8 FILLER_8_655 ();
 sg13g2_decap_8 FILLER_8_662 ();
 sg13g2_decap_8 FILLER_8_669 ();
 sg13g2_decap_8 FILLER_8_676 ();
 sg13g2_decap_8 FILLER_8_683 ();
 sg13g2_decap_8 FILLER_8_690 ();
 sg13g2_decap_8 FILLER_8_697 ();
 sg13g2_decap_8 FILLER_8_704 ();
 sg13g2_decap_8 FILLER_8_711 ();
 sg13g2_decap_8 FILLER_8_718 ();
 sg13g2_decap_8 FILLER_8_725 ();
 sg13g2_decap_8 FILLER_8_732 ();
 sg13g2_decap_8 FILLER_8_739 ();
 sg13g2_decap_8 FILLER_8_746 ();
 sg13g2_decap_8 FILLER_8_753 ();
 sg13g2_decap_8 FILLER_8_760 ();
 sg13g2_decap_8 FILLER_8_767 ();
 sg13g2_decap_8 FILLER_8_774 ();
 sg13g2_decap_8 FILLER_8_781 ();
 sg13g2_decap_8 FILLER_8_788 ();
 sg13g2_decap_8 FILLER_8_795 ();
 sg13g2_decap_8 FILLER_8_802 ();
 sg13g2_decap_8 FILLER_8_809 ();
 sg13g2_decap_8 FILLER_8_816 ();
 sg13g2_decap_8 FILLER_8_823 ();
 sg13g2_decap_8 FILLER_8_830 ();
 sg13g2_decap_8 FILLER_8_837 ();
 sg13g2_decap_8 FILLER_8_844 ();
 sg13g2_decap_8 FILLER_8_851 ();
 sg13g2_decap_8 FILLER_8_858 ();
 sg13g2_decap_8 FILLER_8_865 ();
 sg13g2_decap_8 FILLER_8_872 ();
 sg13g2_decap_8 FILLER_8_879 ();
 sg13g2_decap_8 FILLER_8_886 ();
 sg13g2_decap_8 FILLER_8_893 ();
 sg13g2_decap_8 FILLER_8_900 ();
 sg13g2_decap_8 FILLER_8_907 ();
 sg13g2_decap_8 FILLER_8_914 ();
 sg13g2_decap_4 FILLER_8_921 ();
 sg13g2_decap_8 FILLER_9_4 ();
 sg13g2_decap_8 FILLER_9_11 ();
 sg13g2_decap_8 FILLER_9_18 ();
 sg13g2_decap_8 FILLER_9_25 ();
 sg13g2_decap_8 FILLER_9_32 ();
 sg13g2_decap_8 FILLER_9_39 ();
 sg13g2_decap_8 FILLER_9_46 ();
 sg13g2_decap_8 FILLER_9_53 ();
 sg13g2_decap_8 FILLER_9_60 ();
 sg13g2_decap_8 FILLER_9_67 ();
 sg13g2_decap_8 FILLER_9_74 ();
 sg13g2_decap_8 FILLER_9_81 ();
 sg13g2_decap_8 FILLER_9_88 ();
 sg13g2_decap_8 FILLER_9_95 ();
 sg13g2_decap_8 FILLER_9_102 ();
 sg13g2_decap_8 FILLER_9_109 ();
 sg13g2_decap_8 FILLER_9_116 ();
 sg13g2_decap_8 FILLER_9_123 ();
 sg13g2_decap_8 FILLER_9_130 ();
 sg13g2_decap_8 FILLER_9_137 ();
 sg13g2_decap_8 FILLER_9_144 ();
 sg13g2_decap_8 FILLER_9_151 ();
 sg13g2_decap_8 FILLER_9_158 ();
 sg13g2_decap_8 FILLER_9_165 ();
 sg13g2_decap_8 FILLER_9_172 ();
 sg13g2_decap_8 FILLER_9_179 ();
 sg13g2_decap_8 FILLER_9_186 ();
 sg13g2_decap_8 FILLER_9_193 ();
 sg13g2_decap_8 FILLER_9_200 ();
 sg13g2_decap_8 FILLER_9_207 ();
 sg13g2_decap_8 FILLER_9_214 ();
 sg13g2_decap_8 FILLER_9_221 ();
 sg13g2_decap_8 FILLER_9_228 ();
 sg13g2_decap_8 FILLER_9_235 ();
 sg13g2_decap_8 FILLER_9_242 ();
 sg13g2_decap_8 FILLER_9_249 ();
 sg13g2_decap_8 FILLER_9_256 ();
 sg13g2_decap_8 FILLER_9_263 ();
 sg13g2_decap_8 FILLER_9_270 ();
 sg13g2_decap_8 FILLER_9_277 ();
 sg13g2_decap_8 FILLER_9_284 ();
 sg13g2_decap_8 FILLER_9_291 ();
 sg13g2_decap_8 FILLER_9_298 ();
 sg13g2_decap_8 FILLER_9_305 ();
 sg13g2_decap_8 FILLER_9_312 ();
 sg13g2_decap_8 FILLER_9_319 ();
 sg13g2_decap_8 FILLER_9_326 ();
 sg13g2_decap_8 FILLER_9_333 ();
 sg13g2_decap_8 FILLER_9_340 ();
 sg13g2_decap_8 FILLER_9_347 ();
 sg13g2_decap_8 FILLER_9_354 ();
 sg13g2_decap_8 FILLER_9_361 ();
 sg13g2_decap_8 FILLER_9_368 ();
 sg13g2_decap_8 FILLER_9_375 ();
 sg13g2_decap_8 FILLER_9_382 ();
 sg13g2_decap_8 FILLER_9_389 ();
 sg13g2_decap_8 FILLER_9_396 ();
 sg13g2_decap_8 FILLER_9_403 ();
 sg13g2_decap_8 FILLER_9_410 ();
 sg13g2_decap_8 FILLER_9_417 ();
 sg13g2_decap_8 FILLER_9_424 ();
 sg13g2_decap_8 FILLER_9_431 ();
 sg13g2_decap_8 FILLER_9_438 ();
 sg13g2_decap_8 FILLER_9_445 ();
 sg13g2_decap_8 FILLER_9_452 ();
 sg13g2_decap_8 FILLER_9_459 ();
 sg13g2_decap_8 FILLER_9_466 ();
 sg13g2_decap_8 FILLER_9_473 ();
 sg13g2_decap_8 FILLER_9_480 ();
 sg13g2_decap_8 FILLER_9_487 ();
 sg13g2_decap_8 FILLER_9_494 ();
 sg13g2_decap_8 FILLER_9_501 ();
 sg13g2_decap_8 FILLER_9_508 ();
 sg13g2_decap_8 FILLER_9_515 ();
 sg13g2_decap_8 FILLER_9_522 ();
 sg13g2_decap_8 FILLER_9_529 ();
 sg13g2_decap_8 FILLER_9_536 ();
 sg13g2_decap_8 FILLER_9_543 ();
 sg13g2_decap_8 FILLER_9_550 ();
 sg13g2_decap_8 FILLER_9_557 ();
 sg13g2_decap_8 FILLER_9_564 ();
 sg13g2_decap_8 FILLER_9_571 ();
 sg13g2_decap_8 FILLER_9_578 ();
 sg13g2_decap_8 FILLER_9_585 ();
 sg13g2_decap_8 FILLER_9_592 ();
 sg13g2_decap_8 FILLER_9_599 ();
 sg13g2_decap_8 FILLER_9_606 ();
 sg13g2_decap_8 FILLER_9_613 ();
 sg13g2_decap_8 FILLER_9_620 ();
 sg13g2_decap_8 FILLER_9_627 ();
 sg13g2_decap_8 FILLER_9_634 ();
 sg13g2_decap_8 FILLER_9_641 ();
 sg13g2_decap_8 FILLER_9_648 ();
 sg13g2_decap_8 FILLER_9_655 ();
 sg13g2_decap_8 FILLER_9_662 ();
 sg13g2_decap_8 FILLER_9_669 ();
 sg13g2_decap_8 FILLER_9_676 ();
 sg13g2_decap_8 FILLER_9_683 ();
 sg13g2_decap_8 FILLER_9_690 ();
 sg13g2_decap_8 FILLER_9_697 ();
 sg13g2_decap_8 FILLER_9_704 ();
 sg13g2_decap_8 FILLER_9_711 ();
 sg13g2_decap_8 FILLER_9_718 ();
 sg13g2_decap_8 FILLER_9_725 ();
 sg13g2_decap_8 FILLER_9_732 ();
 sg13g2_decap_8 FILLER_9_739 ();
 sg13g2_decap_8 FILLER_9_746 ();
 sg13g2_decap_8 FILLER_9_753 ();
 sg13g2_decap_8 FILLER_9_760 ();
 sg13g2_decap_8 FILLER_9_767 ();
 sg13g2_decap_8 FILLER_9_774 ();
 sg13g2_decap_8 FILLER_9_781 ();
 sg13g2_decap_8 FILLER_9_788 ();
 sg13g2_decap_8 FILLER_9_795 ();
 sg13g2_decap_8 FILLER_9_802 ();
 sg13g2_decap_8 FILLER_9_809 ();
 sg13g2_decap_8 FILLER_9_816 ();
 sg13g2_decap_8 FILLER_9_823 ();
 sg13g2_decap_8 FILLER_9_830 ();
 sg13g2_decap_8 FILLER_9_837 ();
 sg13g2_decap_8 FILLER_9_844 ();
 sg13g2_decap_8 FILLER_9_851 ();
 sg13g2_decap_8 FILLER_9_858 ();
 sg13g2_decap_8 FILLER_9_865 ();
 sg13g2_decap_8 FILLER_9_872 ();
 sg13g2_decap_8 FILLER_9_879 ();
 sg13g2_decap_8 FILLER_9_886 ();
 sg13g2_decap_8 FILLER_9_893 ();
 sg13g2_decap_8 FILLER_9_900 ();
 sg13g2_decap_8 FILLER_9_907 ();
 sg13g2_decap_8 FILLER_9_914 ();
 sg13g2_decap_4 FILLER_9_921 ();
 sg13g2_decap_8 FILLER_10_4 ();
 sg13g2_decap_8 FILLER_10_11 ();
 sg13g2_decap_8 FILLER_10_18 ();
 sg13g2_decap_8 FILLER_10_25 ();
 sg13g2_decap_8 FILLER_10_32 ();
 sg13g2_decap_8 FILLER_10_39 ();
 sg13g2_decap_8 FILLER_10_46 ();
 sg13g2_decap_8 FILLER_10_53 ();
 sg13g2_decap_8 FILLER_10_60 ();
 sg13g2_decap_8 FILLER_10_67 ();
 sg13g2_decap_8 FILLER_10_74 ();
 sg13g2_decap_8 FILLER_10_81 ();
 sg13g2_decap_8 FILLER_10_88 ();
 sg13g2_decap_8 FILLER_10_95 ();
 sg13g2_decap_8 FILLER_10_102 ();
 sg13g2_decap_8 FILLER_10_109 ();
 sg13g2_decap_8 FILLER_10_116 ();
 sg13g2_decap_8 FILLER_10_123 ();
 sg13g2_decap_8 FILLER_10_130 ();
 sg13g2_decap_8 FILLER_10_137 ();
 sg13g2_decap_8 FILLER_10_144 ();
 sg13g2_decap_8 FILLER_10_151 ();
 sg13g2_decap_8 FILLER_10_158 ();
 sg13g2_decap_8 FILLER_10_165 ();
 sg13g2_decap_8 FILLER_10_172 ();
 sg13g2_decap_8 FILLER_10_179 ();
 sg13g2_decap_8 FILLER_10_186 ();
 sg13g2_decap_8 FILLER_10_193 ();
 sg13g2_decap_8 FILLER_10_200 ();
 sg13g2_decap_8 FILLER_10_207 ();
 sg13g2_decap_8 FILLER_10_214 ();
 sg13g2_decap_8 FILLER_10_221 ();
 sg13g2_decap_8 FILLER_10_228 ();
 sg13g2_decap_8 FILLER_10_235 ();
 sg13g2_decap_8 FILLER_10_242 ();
 sg13g2_decap_8 FILLER_10_249 ();
 sg13g2_decap_8 FILLER_10_256 ();
 sg13g2_decap_8 FILLER_10_263 ();
 sg13g2_decap_8 FILLER_10_270 ();
 sg13g2_decap_8 FILLER_10_277 ();
 sg13g2_decap_8 FILLER_10_284 ();
 sg13g2_decap_8 FILLER_10_291 ();
 sg13g2_decap_8 FILLER_10_298 ();
 sg13g2_decap_8 FILLER_10_305 ();
 sg13g2_decap_8 FILLER_10_312 ();
 sg13g2_decap_8 FILLER_10_319 ();
 sg13g2_decap_8 FILLER_10_326 ();
 sg13g2_decap_8 FILLER_10_333 ();
 sg13g2_decap_8 FILLER_10_340 ();
 sg13g2_decap_8 FILLER_10_347 ();
 sg13g2_decap_8 FILLER_10_354 ();
 sg13g2_decap_8 FILLER_10_361 ();
 sg13g2_decap_8 FILLER_10_368 ();
 sg13g2_decap_8 FILLER_10_375 ();
 sg13g2_decap_8 FILLER_10_382 ();
 sg13g2_decap_8 FILLER_10_389 ();
 sg13g2_decap_8 FILLER_10_396 ();
 sg13g2_decap_8 FILLER_10_403 ();
 sg13g2_decap_8 FILLER_10_410 ();
 sg13g2_decap_8 FILLER_10_417 ();
 sg13g2_decap_8 FILLER_10_424 ();
 sg13g2_decap_8 FILLER_10_431 ();
 sg13g2_decap_8 FILLER_10_438 ();
 sg13g2_decap_8 FILLER_10_445 ();
 sg13g2_decap_8 FILLER_10_452 ();
 sg13g2_decap_8 FILLER_10_459 ();
 sg13g2_decap_8 FILLER_10_466 ();
 sg13g2_decap_8 FILLER_10_473 ();
 sg13g2_decap_8 FILLER_10_480 ();
 sg13g2_decap_8 FILLER_10_487 ();
 sg13g2_decap_8 FILLER_10_494 ();
 sg13g2_decap_8 FILLER_10_501 ();
 sg13g2_decap_8 FILLER_10_508 ();
 sg13g2_decap_8 FILLER_10_515 ();
 sg13g2_decap_8 FILLER_10_522 ();
 sg13g2_decap_8 FILLER_10_529 ();
 sg13g2_decap_8 FILLER_10_536 ();
 sg13g2_decap_8 FILLER_10_543 ();
 sg13g2_decap_8 FILLER_10_550 ();
 sg13g2_decap_8 FILLER_10_557 ();
 sg13g2_decap_8 FILLER_10_564 ();
 sg13g2_decap_8 FILLER_10_571 ();
 sg13g2_decap_8 FILLER_10_578 ();
 sg13g2_decap_8 FILLER_10_585 ();
 sg13g2_decap_8 FILLER_10_592 ();
 sg13g2_decap_8 FILLER_10_599 ();
 sg13g2_decap_8 FILLER_10_606 ();
 sg13g2_decap_8 FILLER_10_613 ();
 sg13g2_decap_8 FILLER_10_620 ();
 sg13g2_decap_8 FILLER_10_627 ();
 sg13g2_decap_8 FILLER_10_634 ();
 sg13g2_decap_8 FILLER_10_641 ();
 sg13g2_decap_8 FILLER_10_648 ();
 sg13g2_decap_8 FILLER_10_655 ();
 sg13g2_decap_8 FILLER_10_662 ();
 sg13g2_decap_8 FILLER_10_669 ();
 sg13g2_decap_8 FILLER_10_676 ();
 sg13g2_decap_8 FILLER_10_683 ();
 sg13g2_decap_8 FILLER_10_690 ();
 sg13g2_decap_8 FILLER_10_697 ();
 sg13g2_decap_8 FILLER_10_704 ();
 sg13g2_decap_8 FILLER_10_711 ();
 sg13g2_decap_8 FILLER_10_718 ();
 sg13g2_decap_8 FILLER_10_725 ();
 sg13g2_decap_8 FILLER_10_732 ();
 sg13g2_decap_8 FILLER_10_739 ();
 sg13g2_decap_8 FILLER_10_746 ();
 sg13g2_decap_8 FILLER_10_753 ();
 sg13g2_decap_8 FILLER_10_760 ();
 sg13g2_decap_8 FILLER_10_767 ();
 sg13g2_decap_8 FILLER_10_774 ();
 sg13g2_decap_8 FILLER_10_781 ();
 sg13g2_decap_8 FILLER_10_788 ();
 sg13g2_decap_8 FILLER_10_795 ();
 sg13g2_decap_8 FILLER_10_802 ();
 sg13g2_decap_8 FILLER_10_809 ();
 sg13g2_decap_8 FILLER_10_816 ();
 sg13g2_decap_8 FILLER_10_823 ();
 sg13g2_decap_8 FILLER_10_830 ();
 sg13g2_decap_8 FILLER_10_837 ();
 sg13g2_decap_8 FILLER_10_844 ();
 sg13g2_decap_8 FILLER_10_851 ();
 sg13g2_decap_8 FILLER_10_858 ();
 sg13g2_decap_8 FILLER_10_865 ();
 sg13g2_decap_8 FILLER_10_872 ();
 sg13g2_decap_8 FILLER_10_879 ();
 sg13g2_decap_8 FILLER_10_886 ();
 sg13g2_decap_8 FILLER_10_893 ();
 sg13g2_decap_8 FILLER_10_900 ();
 sg13g2_decap_8 FILLER_10_907 ();
 sg13g2_decap_8 FILLER_10_914 ();
 sg13g2_decap_4 FILLER_10_921 ();
 sg13g2_decap_8 FILLER_11_4 ();
 sg13g2_decap_8 FILLER_11_11 ();
 sg13g2_decap_8 FILLER_11_18 ();
 sg13g2_decap_8 FILLER_11_25 ();
 sg13g2_decap_8 FILLER_11_32 ();
 sg13g2_decap_8 FILLER_11_39 ();
 sg13g2_decap_8 FILLER_11_46 ();
 sg13g2_decap_8 FILLER_11_53 ();
 sg13g2_decap_8 FILLER_11_60 ();
 sg13g2_decap_8 FILLER_11_67 ();
 sg13g2_decap_8 FILLER_11_74 ();
 sg13g2_decap_8 FILLER_11_81 ();
 sg13g2_decap_8 FILLER_11_88 ();
 sg13g2_decap_8 FILLER_11_95 ();
 sg13g2_decap_8 FILLER_11_102 ();
 sg13g2_decap_8 FILLER_11_109 ();
 sg13g2_decap_8 FILLER_11_116 ();
 sg13g2_decap_8 FILLER_11_123 ();
 sg13g2_decap_8 FILLER_11_130 ();
 sg13g2_decap_8 FILLER_11_137 ();
 sg13g2_decap_8 FILLER_11_144 ();
 sg13g2_decap_8 FILLER_11_151 ();
 sg13g2_decap_8 FILLER_11_158 ();
 sg13g2_decap_8 FILLER_11_165 ();
 sg13g2_decap_8 FILLER_11_172 ();
 sg13g2_decap_8 FILLER_11_179 ();
 sg13g2_decap_8 FILLER_11_186 ();
 sg13g2_decap_8 FILLER_11_193 ();
 sg13g2_decap_8 FILLER_11_200 ();
 sg13g2_decap_8 FILLER_11_207 ();
 sg13g2_decap_8 FILLER_11_214 ();
 sg13g2_decap_8 FILLER_11_221 ();
 sg13g2_decap_8 FILLER_11_228 ();
 sg13g2_decap_8 FILLER_11_235 ();
 sg13g2_decap_8 FILLER_11_242 ();
 sg13g2_decap_8 FILLER_11_249 ();
 sg13g2_decap_8 FILLER_11_256 ();
 sg13g2_decap_8 FILLER_11_263 ();
 sg13g2_decap_8 FILLER_11_270 ();
 sg13g2_decap_8 FILLER_11_277 ();
 sg13g2_decap_8 FILLER_11_284 ();
 sg13g2_decap_8 FILLER_11_291 ();
 sg13g2_decap_8 FILLER_11_298 ();
 sg13g2_decap_8 FILLER_11_305 ();
 sg13g2_decap_8 FILLER_11_312 ();
 sg13g2_decap_8 FILLER_11_319 ();
 sg13g2_decap_8 FILLER_11_326 ();
 sg13g2_decap_8 FILLER_11_333 ();
 sg13g2_decap_8 FILLER_11_340 ();
 sg13g2_decap_8 FILLER_11_347 ();
 sg13g2_decap_8 FILLER_11_354 ();
 sg13g2_decap_8 FILLER_11_361 ();
 sg13g2_decap_8 FILLER_11_368 ();
 sg13g2_decap_8 FILLER_11_375 ();
 sg13g2_decap_8 FILLER_11_382 ();
 sg13g2_decap_8 FILLER_11_389 ();
 sg13g2_decap_8 FILLER_11_396 ();
 sg13g2_decap_8 FILLER_11_403 ();
 sg13g2_decap_8 FILLER_11_410 ();
 sg13g2_decap_8 FILLER_11_417 ();
 sg13g2_decap_8 FILLER_11_424 ();
 sg13g2_decap_8 FILLER_11_431 ();
 sg13g2_decap_8 FILLER_11_438 ();
 sg13g2_decap_8 FILLER_11_445 ();
 sg13g2_decap_8 FILLER_11_452 ();
 sg13g2_decap_8 FILLER_11_459 ();
 sg13g2_decap_8 FILLER_11_466 ();
 sg13g2_decap_8 FILLER_11_473 ();
 sg13g2_decap_8 FILLER_11_480 ();
 sg13g2_decap_8 FILLER_11_487 ();
 sg13g2_decap_8 FILLER_11_494 ();
 sg13g2_decap_8 FILLER_11_501 ();
 sg13g2_decap_8 FILLER_11_508 ();
 sg13g2_decap_8 FILLER_11_515 ();
 sg13g2_decap_8 FILLER_11_522 ();
 sg13g2_decap_8 FILLER_11_529 ();
 sg13g2_decap_8 FILLER_11_536 ();
 sg13g2_decap_8 FILLER_11_543 ();
 sg13g2_decap_8 FILLER_11_550 ();
 sg13g2_decap_8 FILLER_11_557 ();
 sg13g2_decap_8 FILLER_11_564 ();
 sg13g2_decap_8 FILLER_11_571 ();
 sg13g2_decap_8 FILLER_11_578 ();
 sg13g2_decap_8 FILLER_11_585 ();
 sg13g2_decap_8 FILLER_11_592 ();
 sg13g2_decap_8 FILLER_11_599 ();
 sg13g2_decap_8 FILLER_11_606 ();
 sg13g2_decap_8 FILLER_11_613 ();
 sg13g2_decap_8 FILLER_11_620 ();
 sg13g2_decap_8 FILLER_11_627 ();
 sg13g2_decap_8 FILLER_11_634 ();
 sg13g2_decap_8 FILLER_11_641 ();
 sg13g2_decap_8 FILLER_11_648 ();
 sg13g2_decap_8 FILLER_11_655 ();
 sg13g2_decap_8 FILLER_11_662 ();
 sg13g2_decap_8 FILLER_11_669 ();
 sg13g2_decap_8 FILLER_11_676 ();
 sg13g2_decap_8 FILLER_11_683 ();
 sg13g2_decap_8 FILLER_11_690 ();
 sg13g2_decap_8 FILLER_11_697 ();
 sg13g2_decap_8 FILLER_11_704 ();
 sg13g2_decap_8 FILLER_11_711 ();
 sg13g2_decap_8 FILLER_11_718 ();
 sg13g2_decap_8 FILLER_11_725 ();
 sg13g2_decap_8 FILLER_11_732 ();
 sg13g2_decap_8 FILLER_11_739 ();
 sg13g2_decap_8 FILLER_11_746 ();
 sg13g2_decap_8 FILLER_11_753 ();
 sg13g2_decap_8 FILLER_11_760 ();
 sg13g2_decap_8 FILLER_11_767 ();
 sg13g2_decap_8 FILLER_11_774 ();
 sg13g2_decap_8 FILLER_11_781 ();
 sg13g2_decap_8 FILLER_11_788 ();
 sg13g2_decap_8 FILLER_11_795 ();
 sg13g2_decap_8 FILLER_11_802 ();
 sg13g2_decap_8 FILLER_11_809 ();
 sg13g2_decap_8 FILLER_11_816 ();
 sg13g2_decap_8 FILLER_11_823 ();
 sg13g2_decap_8 FILLER_11_830 ();
 sg13g2_decap_8 FILLER_11_837 ();
 sg13g2_decap_8 FILLER_11_844 ();
 sg13g2_decap_8 FILLER_11_851 ();
 sg13g2_decap_8 FILLER_11_858 ();
 sg13g2_decap_8 FILLER_11_865 ();
 sg13g2_decap_8 FILLER_11_872 ();
 sg13g2_decap_8 FILLER_11_879 ();
 sg13g2_decap_8 FILLER_11_886 ();
 sg13g2_decap_8 FILLER_11_893 ();
 sg13g2_decap_8 FILLER_11_900 ();
 sg13g2_decap_8 FILLER_11_907 ();
 sg13g2_decap_8 FILLER_11_914 ();
 sg13g2_decap_4 FILLER_11_921 ();
 sg13g2_decap_8 FILLER_12_4 ();
 sg13g2_decap_8 FILLER_12_11 ();
 sg13g2_decap_8 FILLER_12_18 ();
 sg13g2_decap_8 FILLER_12_25 ();
 sg13g2_decap_8 FILLER_12_32 ();
 sg13g2_decap_8 FILLER_12_39 ();
 sg13g2_decap_8 FILLER_12_46 ();
 sg13g2_decap_8 FILLER_12_53 ();
 sg13g2_decap_8 FILLER_12_60 ();
 sg13g2_decap_8 FILLER_12_67 ();
 sg13g2_decap_8 FILLER_12_74 ();
 sg13g2_decap_8 FILLER_12_81 ();
 sg13g2_decap_8 FILLER_12_88 ();
 sg13g2_decap_8 FILLER_12_95 ();
 sg13g2_decap_8 FILLER_12_102 ();
 sg13g2_decap_8 FILLER_12_109 ();
 sg13g2_decap_8 FILLER_12_116 ();
 sg13g2_decap_8 FILLER_12_123 ();
 sg13g2_decap_8 FILLER_12_130 ();
 sg13g2_decap_8 FILLER_12_137 ();
 sg13g2_decap_8 FILLER_12_144 ();
 sg13g2_decap_8 FILLER_12_151 ();
 sg13g2_decap_8 FILLER_12_158 ();
 sg13g2_decap_8 FILLER_12_165 ();
 sg13g2_decap_8 FILLER_12_172 ();
 sg13g2_decap_8 FILLER_12_179 ();
 sg13g2_decap_8 FILLER_12_186 ();
 sg13g2_decap_8 FILLER_12_193 ();
 sg13g2_decap_8 FILLER_12_200 ();
 sg13g2_decap_8 FILLER_12_207 ();
 sg13g2_decap_8 FILLER_12_214 ();
 sg13g2_decap_8 FILLER_12_221 ();
 sg13g2_decap_8 FILLER_12_228 ();
 sg13g2_decap_8 FILLER_12_235 ();
 sg13g2_decap_8 FILLER_12_242 ();
 sg13g2_decap_8 FILLER_12_249 ();
 sg13g2_decap_8 FILLER_12_256 ();
 sg13g2_decap_8 FILLER_12_263 ();
 sg13g2_decap_8 FILLER_12_270 ();
 sg13g2_decap_8 FILLER_12_277 ();
 sg13g2_decap_8 FILLER_12_284 ();
 sg13g2_decap_8 FILLER_12_291 ();
 sg13g2_decap_8 FILLER_12_298 ();
 sg13g2_decap_8 FILLER_12_305 ();
 sg13g2_decap_8 FILLER_12_312 ();
 sg13g2_decap_8 FILLER_12_319 ();
 sg13g2_decap_8 FILLER_12_326 ();
 sg13g2_decap_8 FILLER_12_333 ();
 sg13g2_decap_8 FILLER_12_340 ();
 sg13g2_decap_8 FILLER_12_347 ();
 sg13g2_decap_8 FILLER_12_354 ();
 sg13g2_decap_8 FILLER_12_361 ();
 sg13g2_decap_8 FILLER_12_368 ();
 sg13g2_decap_8 FILLER_12_375 ();
 sg13g2_decap_8 FILLER_12_382 ();
 sg13g2_decap_8 FILLER_12_389 ();
 sg13g2_decap_8 FILLER_12_396 ();
 sg13g2_decap_8 FILLER_12_403 ();
 sg13g2_decap_8 FILLER_12_410 ();
 sg13g2_decap_8 FILLER_12_417 ();
 sg13g2_decap_8 FILLER_12_424 ();
 sg13g2_decap_8 FILLER_12_431 ();
 sg13g2_decap_8 FILLER_12_438 ();
 sg13g2_decap_8 FILLER_12_445 ();
 sg13g2_decap_8 FILLER_12_452 ();
 sg13g2_decap_8 FILLER_12_459 ();
 sg13g2_decap_8 FILLER_12_466 ();
 sg13g2_decap_8 FILLER_12_473 ();
 sg13g2_decap_8 FILLER_12_480 ();
 sg13g2_decap_8 FILLER_12_487 ();
 sg13g2_decap_8 FILLER_12_494 ();
 sg13g2_decap_8 FILLER_12_501 ();
 sg13g2_decap_8 FILLER_12_508 ();
 sg13g2_decap_8 FILLER_12_515 ();
 sg13g2_decap_8 FILLER_12_522 ();
 sg13g2_decap_8 FILLER_12_529 ();
 sg13g2_decap_8 FILLER_12_536 ();
 sg13g2_decap_8 FILLER_12_543 ();
 sg13g2_decap_8 FILLER_12_550 ();
 sg13g2_decap_8 FILLER_12_557 ();
 sg13g2_decap_8 FILLER_12_564 ();
 sg13g2_decap_8 FILLER_12_571 ();
 sg13g2_decap_8 FILLER_12_578 ();
 sg13g2_decap_8 FILLER_12_585 ();
 sg13g2_decap_8 FILLER_12_592 ();
 sg13g2_decap_8 FILLER_12_599 ();
 sg13g2_decap_8 FILLER_12_606 ();
 sg13g2_decap_8 FILLER_12_613 ();
 sg13g2_decap_8 FILLER_12_620 ();
 sg13g2_decap_8 FILLER_12_627 ();
 sg13g2_decap_8 FILLER_12_634 ();
 sg13g2_decap_8 FILLER_12_641 ();
 sg13g2_decap_8 FILLER_12_648 ();
 sg13g2_decap_8 FILLER_12_655 ();
 sg13g2_decap_8 FILLER_12_662 ();
 sg13g2_decap_8 FILLER_12_669 ();
 sg13g2_decap_8 FILLER_12_676 ();
 sg13g2_decap_8 FILLER_12_683 ();
 sg13g2_decap_8 FILLER_12_690 ();
 sg13g2_decap_8 FILLER_12_697 ();
 sg13g2_decap_8 FILLER_12_704 ();
 sg13g2_decap_8 FILLER_12_711 ();
 sg13g2_decap_8 FILLER_12_718 ();
 sg13g2_decap_8 FILLER_12_725 ();
 sg13g2_decap_8 FILLER_12_732 ();
 sg13g2_decap_8 FILLER_12_739 ();
 sg13g2_decap_8 FILLER_12_746 ();
 sg13g2_decap_8 FILLER_12_753 ();
 sg13g2_decap_8 FILLER_12_760 ();
 sg13g2_decap_8 FILLER_12_767 ();
 sg13g2_decap_8 FILLER_12_774 ();
 sg13g2_decap_8 FILLER_12_781 ();
 sg13g2_decap_8 FILLER_12_788 ();
 sg13g2_decap_8 FILLER_12_795 ();
 sg13g2_decap_8 FILLER_12_802 ();
 sg13g2_decap_8 FILLER_12_809 ();
 sg13g2_decap_8 FILLER_12_816 ();
 sg13g2_decap_8 FILLER_12_823 ();
 sg13g2_decap_8 FILLER_12_830 ();
 sg13g2_decap_8 FILLER_12_837 ();
 sg13g2_decap_8 FILLER_12_844 ();
 sg13g2_decap_8 FILLER_12_851 ();
 sg13g2_decap_8 FILLER_12_858 ();
 sg13g2_decap_8 FILLER_12_865 ();
 sg13g2_decap_8 FILLER_12_872 ();
 sg13g2_decap_8 FILLER_12_879 ();
 sg13g2_decap_8 FILLER_12_886 ();
 sg13g2_decap_8 FILLER_12_893 ();
 sg13g2_decap_8 FILLER_12_900 ();
 sg13g2_decap_8 FILLER_12_907 ();
 sg13g2_decap_8 FILLER_12_914 ();
 sg13g2_decap_4 FILLER_12_921 ();
 sg13g2_decap_8 FILLER_13_4 ();
 sg13g2_decap_8 FILLER_13_11 ();
 sg13g2_decap_8 FILLER_13_18 ();
 sg13g2_decap_8 FILLER_13_25 ();
 sg13g2_decap_8 FILLER_13_32 ();
 sg13g2_decap_8 FILLER_13_39 ();
 sg13g2_decap_8 FILLER_13_46 ();
 sg13g2_decap_8 FILLER_13_53 ();
 sg13g2_decap_8 FILLER_13_60 ();
 sg13g2_decap_8 FILLER_13_67 ();
 sg13g2_decap_8 FILLER_13_74 ();
 sg13g2_decap_8 FILLER_13_81 ();
 sg13g2_decap_8 FILLER_13_88 ();
 sg13g2_decap_8 FILLER_13_95 ();
 sg13g2_decap_8 FILLER_13_102 ();
 sg13g2_decap_8 FILLER_13_109 ();
 sg13g2_decap_8 FILLER_13_116 ();
 sg13g2_decap_8 FILLER_13_123 ();
 sg13g2_decap_8 FILLER_13_130 ();
 sg13g2_decap_8 FILLER_13_137 ();
 sg13g2_decap_8 FILLER_13_144 ();
 sg13g2_decap_8 FILLER_13_151 ();
 sg13g2_decap_8 FILLER_13_158 ();
 sg13g2_decap_8 FILLER_13_165 ();
 sg13g2_decap_8 FILLER_13_172 ();
 sg13g2_decap_8 FILLER_13_179 ();
 sg13g2_decap_8 FILLER_13_186 ();
 sg13g2_decap_8 FILLER_13_193 ();
 sg13g2_decap_8 FILLER_13_200 ();
 sg13g2_decap_8 FILLER_13_207 ();
 sg13g2_decap_8 FILLER_13_214 ();
 sg13g2_decap_8 FILLER_13_221 ();
 sg13g2_decap_8 FILLER_13_228 ();
 sg13g2_decap_8 FILLER_13_235 ();
 sg13g2_decap_8 FILLER_13_242 ();
 sg13g2_decap_8 FILLER_13_249 ();
 sg13g2_decap_8 FILLER_13_256 ();
 sg13g2_decap_8 FILLER_13_263 ();
 sg13g2_decap_8 FILLER_13_270 ();
 sg13g2_decap_8 FILLER_13_277 ();
 sg13g2_decap_8 FILLER_13_284 ();
 sg13g2_decap_8 FILLER_13_291 ();
 sg13g2_decap_8 FILLER_13_298 ();
 sg13g2_decap_8 FILLER_13_305 ();
 sg13g2_decap_8 FILLER_13_312 ();
 sg13g2_decap_8 FILLER_13_319 ();
 sg13g2_decap_8 FILLER_13_326 ();
 sg13g2_decap_8 FILLER_13_333 ();
 sg13g2_decap_8 FILLER_13_340 ();
 sg13g2_decap_8 FILLER_13_347 ();
 sg13g2_decap_8 FILLER_13_354 ();
 sg13g2_decap_8 FILLER_13_361 ();
 sg13g2_decap_8 FILLER_13_368 ();
 sg13g2_decap_8 FILLER_13_375 ();
 sg13g2_decap_8 FILLER_13_382 ();
 sg13g2_decap_8 FILLER_13_389 ();
 sg13g2_decap_8 FILLER_13_396 ();
 sg13g2_decap_8 FILLER_13_403 ();
 sg13g2_decap_8 FILLER_13_410 ();
 sg13g2_decap_8 FILLER_13_417 ();
 sg13g2_decap_8 FILLER_13_424 ();
 sg13g2_decap_8 FILLER_13_431 ();
 sg13g2_decap_8 FILLER_13_438 ();
 sg13g2_decap_8 FILLER_13_445 ();
 sg13g2_decap_8 FILLER_13_452 ();
 sg13g2_decap_8 FILLER_13_459 ();
 sg13g2_decap_8 FILLER_13_466 ();
 sg13g2_decap_8 FILLER_13_473 ();
 sg13g2_decap_8 FILLER_13_480 ();
 sg13g2_decap_8 FILLER_13_487 ();
 sg13g2_decap_8 FILLER_13_494 ();
 sg13g2_decap_8 FILLER_13_501 ();
 sg13g2_decap_8 FILLER_13_508 ();
 sg13g2_decap_8 FILLER_13_515 ();
 sg13g2_decap_8 FILLER_13_522 ();
 sg13g2_decap_8 FILLER_13_529 ();
 sg13g2_decap_8 FILLER_13_536 ();
 sg13g2_decap_8 FILLER_13_543 ();
 sg13g2_decap_8 FILLER_13_550 ();
 sg13g2_decap_8 FILLER_13_557 ();
 sg13g2_decap_8 FILLER_13_564 ();
 sg13g2_decap_8 FILLER_13_571 ();
 sg13g2_decap_8 FILLER_13_578 ();
 sg13g2_decap_8 FILLER_13_585 ();
 sg13g2_decap_8 FILLER_13_592 ();
 sg13g2_decap_8 FILLER_13_599 ();
 sg13g2_decap_8 FILLER_13_606 ();
 sg13g2_decap_8 FILLER_13_613 ();
 sg13g2_decap_8 FILLER_13_620 ();
 sg13g2_decap_8 FILLER_13_627 ();
 sg13g2_decap_8 FILLER_13_634 ();
 sg13g2_decap_8 FILLER_13_641 ();
 sg13g2_decap_8 FILLER_13_648 ();
 sg13g2_decap_8 FILLER_13_655 ();
 sg13g2_decap_8 FILLER_13_662 ();
 sg13g2_decap_8 FILLER_13_669 ();
 sg13g2_decap_8 FILLER_13_676 ();
 sg13g2_decap_8 FILLER_13_683 ();
 sg13g2_decap_8 FILLER_13_690 ();
 sg13g2_decap_8 FILLER_13_697 ();
 sg13g2_decap_8 FILLER_13_704 ();
 sg13g2_decap_8 FILLER_13_711 ();
 sg13g2_decap_8 FILLER_13_718 ();
 sg13g2_decap_8 FILLER_13_725 ();
 sg13g2_decap_8 FILLER_13_732 ();
 sg13g2_decap_8 FILLER_13_739 ();
 sg13g2_decap_8 FILLER_13_746 ();
 sg13g2_decap_8 FILLER_13_753 ();
 sg13g2_decap_8 FILLER_13_760 ();
 sg13g2_decap_8 FILLER_13_767 ();
 sg13g2_decap_8 FILLER_13_774 ();
 sg13g2_decap_8 FILLER_13_781 ();
 sg13g2_decap_8 FILLER_13_788 ();
 sg13g2_decap_8 FILLER_13_795 ();
 sg13g2_decap_8 FILLER_13_802 ();
 sg13g2_decap_8 FILLER_13_809 ();
 sg13g2_decap_8 FILLER_13_816 ();
 sg13g2_decap_8 FILLER_13_823 ();
 sg13g2_decap_8 FILLER_13_830 ();
 sg13g2_decap_8 FILLER_13_837 ();
 sg13g2_decap_8 FILLER_13_844 ();
 sg13g2_decap_8 FILLER_13_851 ();
 sg13g2_decap_8 FILLER_13_858 ();
 sg13g2_decap_8 FILLER_13_865 ();
 sg13g2_decap_8 FILLER_13_872 ();
 sg13g2_decap_8 FILLER_13_879 ();
 sg13g2_decap_8 FILLER_13_886 ();
 sg13g2_decap_8 FILLER_13_893 ();
 sg13g2_decap_8 FILLER_13_900 ();
 sg13g2_decap_8 FILLER_13_907 ();
 sg13g2_decap_8 FILLER_13_914 ();
 sg13g2_decap_4 FILLER_13_921 ();
 sg13g2_decap_8 FILLER_14_4 ();
 sg13g2_decap_8 FILLER_14_11 ();
 sg13g2_decap_8 FILLER_14_18 ();
 sg13g2_decap_8 FILLER_14_25 ();
 sg13g2_decap_8 FILLER_14_32 ();
 sg13g2_decap_8 FILLER_14_39 ();
 sg13g2_decap_8 FILLER_14_46 ();
 sg13g2_decap_8 FILLER_14_53 ();
 sg13g2_decap_8 FILLER_14_60 ();
 sg13g2_decap_8 FILLER_14_67 ();
 sg13g2_decap_8 FILLER_14_74 ();
 sg13g2_decap_8 FILLER_14_81 ();
 sg13g2_decap_8 FILLER_14_88 ();
 sg13g2_decap_8 FILLER_14_95 ();
 sg13g2_decap_8 FILLER_14_102 ();
 sg13g2_decap_8 FILLER_14_109 ();
 sg13g2_decap_8 FILLER_14_116 ();
 sg13g2_decap_8 FILLER_14_123 ();
 sg13g2_decap_8 FILLER_14_130 ();
 sg13g2_decap_8 FILLER_14_137 ();
 sg13g2_decap_8 FILLER_14_144 ();
 sg13g2_decap_8 FILLER_14_151 ();
 sg13g2_decap_8 FILLER_14_158 ();
 sg13g2_decap_8 FILLER_14_165 ();
 sg13g2_decap_8 FILLER_14_172 ();
 sg13g2_decap_8 FILLER_14_179 ();
 sg13g2_decap_8 FILLER_14_186 ();
 sg13g2_decap_8 FILLER_14_193 ();
 sg13g2_decap_8 FILLER_14_200 ();
 sg13g2_decap_8 FILLER_14_207 ();
 sg13g2_decap_8 FILLER_14_214 ();
 sg13g2_decap_8 FILLER_14_221 ();
 sg13g2_decap_8 FILLER_14_228 ();
 sg13g2_decap_8 FILLER_14_235 ();
 sg13g2_decap_8 FILLER_14_242 ();
 sg13g2_decap_8 FILLER_14_249 ();
 sg13g2_decap_8 FILLER_14_256 ();
 sg13g2_decap_8 FILLER_14_263 ();
 sg13g2_decap_8 FILLER_14_270 ();
 sg13g2_decap_8 FILLER_14_277 ();
 sg13g2_decap_8 FILLER_14_284 ();
 sg13g2_decap_8 FILLER_14_291 ();
 sg13g2_decap_8 FILLER_14_298 ();
 sg13g2_decap_8 FILLER_14_305 ();
 sg13g2_decap_8 FILLER_14_312 ();
 sg13g2_decap_8 FILLER_14_319 ();
 sg13g2_decap_8 FILLER_14_326 ();
 sg13g2_decap_8 FILLER_14_333 ();
 sg13g2_decap_8 FILLER_14_340 ();
 sg13g2_decap_8 FILLER_14_347 ();
 sg13g2_decap_8 FILLER_14_354 ();
 sg13g2_decap_8 FILLER_14_361 ();
 sg13g2_decap_8 FILLER_14_368 ();
 sg13g2_decap_8 FILLER_14_375 ();
 sg13g2_decap_8 FILLER_14_382 ();
 sg13g2_decap_8 FILLER_14_389 ();
 sg13g2_decap_8 FILLER_14_396 ();
 sg13g2_decap_8 FILLER_14_403 ();
 sg13g2_decap_8 FILLER_14_410 ();
 sg13g2_decap_8 FILLER_14_417 ();
 sg13g2_decap_8 FILLER_14_424 ();
 sg13g2_decap_8 FILLER_14_431 ();
 sg13g2_decap_8 FILLER_14_438 ();
 sg13g2_decap_8 FILLER_14_445 ();
 sg13g2_decap_8 FILLER_14_452 ();
 sg13g2_decap_8 FILLER_14_459 ();
 sg13g2_decap_8 FILLER_14_466 ();
 sg13g2_decap_8 FILLER_14_473 ();
 sg13g2_decap_8 FILLER_14_480 ();
 sg13g2_decap_8 FILLER_14_487 ();
 sg13g2_decap_8 FILLER_14_494 ();
 sg13g2_decap_8 FILLER_14_501 ();
 sg13g2_decap_8 FILLER_14_508 ();
 sg13g2_decap_8 FILLER_14_515 ();
 sg13g2_decap_8 FILLER_14_522 ();
 sg13g2_decap_8 FILLER_14_529 ();
 sg13g2_decap_8 FILLER_14_536 ();
 sg13g2_decap_8 FILLER_14_543 ();
 sg13g2_decap_8 FILLER_14_550 ();
 sg13g2_decap_8 FILLER_14_557 ();
 sg13g2_decap_8 FILLER_14_564 ();
 sg13g2_decap_8 FILLER_14_571 ();
 sg13g2_decap_8 FILLER_14_578 ();
 sg13g2_decap_8 FILLER_14_585 ();
 sg13g2_decap_8 FILLER_14_592 ();
 sg13g2_decap_8 FILLER_14_599 ();
 sg13g2_decap_8 FILLER_14_606 ();
 sg13g2_decap_8 FILLER_14_613 ();
 sg13g2_decap_8 FILLER_14_620 ();
 sg13g2_decap_8 FILLER_14_627 ();
 sg13g2_decap_8 FILLER_14_634 ();
 sg13g2_decap_8 FILLER_14_641 ();
 sg13g2_decap_8 FILLER_14_648 ();
 sg13g2_decap_8 FILLER_14_655 ();
 sg13g2_decap_8 FILLER_14_662 ();
 sg13g2_decap_8 FILLER_14_669 ();
 sg13g2_decap_8 FILLER_14_676 ();
 sg13g2_decap_8 FILLER_14_683 ();
 sg13g2_decap_8 FILLER_14_690 ();
 sg13g2_decap_8 FILLER_14_697 ();
 sg13g2_decap_8 FILLER_14_704 ();
 sg13g2_decap_8 FILLER_14_711 ();
 sg13g2_decap_8 FILLER_14_718 ();
 sg13g2_decap_8 FILLER_14_725 ();
 sg13g2_decap_8 FILLER_14_732 ();
 sg13g2_decap_8 FILLER_14_739 ();
 sg13g2_decap_8 FILLER_14_746 ();
 sg13g2_decap_8 FILLER_14_753 ();
 sg13g2_decap_8 FILLER_14_760 ();
 sg13g2_decap_8 FILLER_14_767 ();
 sg13g2_decap_8 FILLER_14_774 ();
 sg13g2_decap_8 FILLER_14_781 ();
 sg13g2_decap_8 FILLER_14_788 ();
 sg13g2_decap_8 FILLER_14_795 ();
 sg13g2_decap_8 FILLER_14_802 ();
 sg13g2_decap_8 FILLER_14_809 ();
 sg13g2_decap_8 FILLER_14_816 ();
 sg13g2_decap_8 FILLER_14_823 ();
 sg13g2_decap_8 FILLER_14_830 ();
 sg13g2_decap_8 FILLER_14_837 ();
 sg13g2_decap_8 FILLER_14_844 ();
 sg13g2_decap_8 FILLER_14_851 ();
 sg13g2_decap_8 FILLER_14_858 ();
 sg13g2_decap_8 FILLER_14_865 ();
 sg13g2_decap_8 FILLER_14_872 ();
 sg13g2_decap_8 FILLER_14_879 ();
 sg13g2_decap_8 FILLER_14_886 ();
 sg13g2_decap_8 FILLER_14_893 ();
 sg13g2_decap_8 FILLER_14_900 ();
 sg13g2_decap_8 FILLER_14_907 ();
 sg13g2_decap_8 FILLER_14_914 ();
 sg13g2_decap_4 FILLER_14_921 ();
 sg13g2_decap_8 FILLER_15_4 ();
 sg13g2_decap_8 FILLER_15_11 ();
 sg13g2_decap_8 FILLER_15_18 ();
 sg13g2_decap_8 FILLER_15_25 ();
 sg13g2_decap_8 FILLER_15_32 ();
 sg13g2_decap_8 FILLER_15_39 ();
 sg13g2_decap_8 FILLER_15_46 ();
 sg13g2_decap_8 FILLER_15_53 ();
 sg13g2_decap_8 FILLER_15_60 ();
 sg13g2_decap_8 FILLER_15_67 ();
 sg13g2_decap_8 FILLER_15_74 ();
 sg13g2_decap_8 FILLER_15_81 ();
 sg13g2_decap_8 FILLER_15_88 ();
 sg13g2_decap_8 FILLER_15_95 ();
 sg13g2_decap_8 FILLER_15_102 ();
 sg13g2_decap_8 FILLER_15_109 ();
 sg13g2_decap_8 FILLER_15_116 ();
 sg13g2_decap_8 FILLER_15_123 ();
 sg13g2_decap_8 FILLER_15_130 ();
 sg13g2_decap_8 FILLER_15_137 ();
 sg13g2_decap_8 FILLER_15_144 ();
 sg13g2_decap_8 FILLER_15_151 ();
 sg13g2_decap_8 FILLER_15_158 ();
 sg13g2_decap_8 FILLER_15_165 ();
 sg13g2_decap_8 FILLER_15_172 ();
 sg13g2_decap_8 FILLER_15_179 ();
 sg13g2_decap_8 FILLER_15_186 ();
 sg13g2_decap_8 FILLER_15_193 ();
 sg13g2_decap_8 FILLER_15_200 ();
 sg13g2_decap_8 FILLER_15_207 ();
 sg13g2_decap_8 FILLER_15_214 ();
 sg13g2_decap_8 FILLER_15_221 ();
 sg13g2_decap_8 FILLER_15_228 ();
 sg13g2_decap_8 FILLER_15_235 ();
 sg13g2_decap_8 FILLER_15_242 ();
 sg13g2_decap_8 FILLER_15_249 ();
 sg13g2_decap_8 FILLER_15_256 ();
 sg13g2_decap_8 FILLER_15_263 ();
 sg13g2_decap_8 FILLER_15_270 ();
 sg13g2_decap_8 FILLER_15_277 ();
 sg13g2_decap_8 FILLER_15_284 ();
 sg13g2_decap_8 FILLER_15_291 ();
 sg13g2_decap_8 FILLER_15_298 ();
 sg13g2_decap_8 FILLER_15_305 ();
 sg13g2_decap_8 FILLER_15_312 ();
 sg13g2_decap_8 FILLER_15_319 ();
 sg13g2_decap_8 FILLER_15_326 ();
 sg13g2_decap_8 FILLER_15_333 ();
 sg13g2_decap_8 FILLER_15_340 ();
 sg13g2_decap_8 FILLER_15_347 ();
 sg13g2_decap_8 FILLER_15_354 ();
 sg13g2_decap_8 FILLER_15_361 ();
 sg13g2_decap_8 FILLER_15_368 ();
 sg13g2_decap_8 FILLER_15_375 ();
 sg13g2_decap_8 FILLER_15_382 ();
 sg13g2_decap_8 FILLER_15_389 ();
 sg13g2_decap_8 FILLER_15_396 ();
 sg13g2_decap_8 FILLER_15_403 ();
 sg13g2_decap_8 FILLER_15_410 ();
 sg13g2_decap_8 FILLER_15_417 ();
 sg13g2_decap_8 FILLER_15_424 ();
 sg13g2_decap_8 FILLER_15_431 ();
 sg13g2_decap_8 FILLER_15_438 ();
 sg13g2_decap_8 FILLER_15_445 ();
 sg13g2_decap_8 FILLER_15_452 ();
 sg13g2_decap_8 FILLER_15_459 ();
 sg13g2_decap_8 FILLER_15_466 ();
 sg13g2_decap_8 FILLER_15_473 ();
 sg13g2_decap_8 FILLER_15_480 ();
 sg13g2_decap_8 FILLER_15_487 ();
 sg13g2_decap_8 FILLER_15_494 ();
 sg13g2_decap_8 FILLER_15_501 ();
 sg13g2_decap_8 FILLER_15_508 ();
 sg13g2_decap_8 FILLER_15_515 ();
 sg13g2_decap_8 FILLER_15_522 ();
 sg13g2_decap_8 FILLER_15_529 ();
 sg13g2_decap_8 FILLER_15_536 ();
 sg13g2_decap_8 FILLER_15_543 ();
 sg13g2_decap_8 FILLER_15_550 ();
 sg13g2_decap_8 FILLER_15_557 ();
 sg13g2_decap_8 FILLER_15_564 ();
 sg13g2_decap_8 FILLER_15_571 ();
 sg13g2_decap_8 FILLER_15_578 ();
 sg13g2_decap_8 FILLER_15_585 ();
 sg13g2_decap_8 FILLER_15_592 ();
 sg13g2_decap_8 FILLER_15_599 ();
 sg13g2_decap_8 FILLER_15_606 ();
 sg13g2_decap_8 FILLER_15_613 ();
 sg13g2_decap_8 FILLER_15_620 ();
 sg13g2_decap_8 FILLER_15_627 ();
 sg13g2_decap_8 FILLER_15_634 ();
 sg13g2_decap_8 FILLER_15_641 ();
 sg13g2_decap_8 FILLER_15_648 ();
 sg13g2_decap_8 FILLER_15_655 ();
 sg13g2_decap_8 FILLER_15_662 ();
 sg13g2_decap_8 FILLER_15_669 ();
 sg13g2_decap_8 FILLER_15_676 ();
 sg13g2_decap_8 FILLER_15_683 ();
 sg13g2_decap_8 FILLER_15_690 ();
 sg13g2_decap_8 FILLER_15_697 ();
 sg13g2_decap_8 FILLER_15_704 ();
 sg13g2_decap_8 FILLER_15_711 ();
 sg13g2_decap_8 FILLER_15_718 ();
 sg13g2_decap_8 FILLER_15_725 ();
 sg13g2_decap_8 FILLER_15_732 ();
 sg13g2_decap_8 FILLER_15_739 ();
 sg13g2_decap_8 FILLER_15_746 ();
 sg13g2_decap_8 FILLER_15_753 ();
 sg13g2_decap_8 FILLER_15_760 ();
 sg13g2_decap_8 FILLER_15_767 ();
 sg13g2_decap_8 FILLER_15_774 ();
 sg13g2_decap_8 FILLER_15_781 ();
 sg13g2_decap_8 FILLER_15_788 ();
 sg13g2_decap_8 FILLER_15_795 ();
 sg13g2_decap_8 FILLER_15_802 ();
 sg13g2_decap_8 FILLER_15_809 ();
 sg13g2_decap_8 FILLER_15_816 ();
 sg13g2_decap_8 FILLER_15_823 ();
 sg13g2_decap_8 FILLER_15_830 ();
 sg13g2_decap_8 FILLER_15_837 ();
 sg13g2_decap_8 FILLER_15_844 ();
 sg13g2_decap_8 FILLER_15_851 ();
 sg13g2_decap_8 FILLER_15_858 ();
 sg13g2_decap_8 FILLER_15_865 ();
 sg13g2_decap_8 FILLER_15_872 ();
 sg13g2_decap_8 FILLER_15_879 ();
 sg13g2_decap_8 FILLER_15_886 ();
 sg13g2_decap_8 FILLER_15_893 ();
 sg13g2_decap_8 FILLER_15_900 ();
 sg13g2_decap_8 FILLER_15_907 ();
 sg13g2_decap_8 FILLER_15_914 ();
 sg13g2_decap_4 FILLER_15_921 ();
 sg13g2_decap_8 FILLER_16_4 ();
 sg13g2_decap_8 FILLER_16_11 ();
 sg13g2_decap_8 FILLER_16_18 ();
 sg13g2_decap_8 FILLER_16_25 ();
 sg13g2_decap_8 FILLER_16_32 ();
 sg13g2_decap_8 FILLER_16_39 ();
 sg13g2_decap_8 FILLER_16_46 ();
 sg13g2_decap_8 FILLER_16_53 ();
 sg13g2_decap_8 FILLER_16_60 ();
 sg13g2_decap_8 FILLER_16_67 ();
 sg13g2_decap_8 FILLER_16_74 ();
 sg13g2_decap_8 FILLER_16_81 ();
 sg13g2_decap_8 FILLER_16_88 ();
 sg13g2_decap_8 FILLER_16_95 ();
 sg13g2_decap_8 FILLER_16_102 ();
 sg13g2_decap_8 FILLER_16_109 ();
 sg13g2_decap_8 FILLER_16_116 ();
 sg13g2_decap_8 FILLER_16_123 ();
 sg13g2_decap_8 FILLER_16_130 ();
 sg13g2_decap_8 FILLER_16_137 ();
 sg13g2_decap_8 FILLER_16_144 ();
 sg13g2_decap_8 FILLER_16_151 ();
 sg13g2_decap_8 FILLER_16_158 ();
 sg13g2_decap_8 FILLER_16_165 ();
 sg13g2_decap_8 FILLER_16_172 ();
 sg13g2_decap_8 FILLER_16_179 ();
 sg13g2_decap_8 FILLER_16_186 ();
 sg13g2_decap_8 FILLER_16_193 ();
 sg13g2_decap_8 FILLER_16_200 ();
 sg13g2_decap_8 FILLER_16_207 ();
 sg13g2_decap_8 FILLER_16_214 ();
 sg13g2_decap_8 FILLER_16_221 ();
 sg13g2_decap_8 FILLER_16_228 ();
 sg13g2_decap_8 FILLER_16_235 ();
 sg13g2_decap_8 FILLER_16_242 ();
 sg13g2_decap_8 FILLER_16_249 ();
 sg13g2_decap_8 FILLER_16_256 ();
 sg13g2_decap_8 FILLER_16_263 ();
 sg13g2_decap_8 FILLER_16_270 ();
 sg13g2_decap_8 FILLER_16_277 ();
 sg13g2_decap_8 FILLER_16_284 ();
 sg13g2_decap_8 FILLER_16_291 ();
 sg13g2_decap_8 FILLER_16_298 ();
 sg13g2_decap_8 FILLER_16_305 ();
 sg13g2_decap_8 FILLER_16_312 ();
 sg13g2_decap_8 FILLER_16_319 ();
 sg13g2_decap_8 FILLER_16_326 ();
 sg13g2_decap_8 FILLER_16_333 ();
 sg13g2_decap_8 FILLER_16_340 ();
 sg13g2_decap_8 FILLER_16_347 ();
 sg13g2_decap_8 FILLER_16_354 ();
 sg13g2_decap_8 FILLER_16_361 ();
 sg13g2_decap_8 FILLER_16_368 ();
 sg13g2_decap_8 FILLER_16_375 ();
 sg13g2_decap_8 FILLER_16_382 ();
 sg13g2_decap_8 FILLER_16_389 ();
 sg13g2_decap_8 FILLER_16_396 ();
 sg13g2_decap_8 FILLER_16_403 ();
 sg13g2_decap_8 FILLER_16_410 ();
 sg13g2_decap_8 FILLER_16_417 ();
 sg13g2_decap_8 FILLER_16_424 ();
 sg13g2_decap_8 FILLER_16_431 ();
 sg13g2_decap_8 FILLER_16_438 ();
 sg13g2_decap_8 FILLER_16_445 ();
 sg13g2_decap_8 FILLER_16_452 ();
 sg13g2_decap_8 FILLER_16_459 ();
 sg13g2_decap_8 FILLER_16_466 ();
 sg13g2_decap_8 FILLER_16_473 ();
 sg13g2_decap_8 FILLER_16_480 ();
 sg13g2_decap_8 FILLER_16_487 ();
 sg13g2_decap_8 FILLER_16_494 ();
 sg13g2_decap_8 FILLER_16_501 ();
 sg13g2_decap_8 FILLER_16_508 ();
 sg13g2_decap_8 FILLER_16_515 ();
 sg13g2_decap_8 FILLER_16_522 ();
 sg13g2_decap_8 FILLER_16_529 ();
 sg13g2_decap_8 FILLER_16_536 ();
 sg13g2_decap_8 FILLER_16_543 ();
 sg13g2_decap_8 FILLER_16_550 ();
 sg13g2_decap_8 FILLER_16_557 ();
 sg13g2_decap_8 FILLER_16_564 ();
 sg13g2_decap_8 FILLER_16_571 ();
 sg13g2_decap_8 FILLER_16_578 ();
 sg13g2_decap_8 FILLER_16_585 ();
 sg13g2_decap_8 FILLER_16_592 ();
 sg13g2_decap_8 FILLER_16_599 ();
 sg13g2_decap_8 FILLER_16_606 ();
 sg13g2_decap_8 FILLER_16_613 ();
 sg13g2_decap_8 FILLER_16_620 ();
 sg13g2_decap_8 FILLER_16_627 ();
 sg13g2_decap_8 FILLER_16_634 ();
 sg13g2_decap_8 FILLER_16_641 ();
 sg13g2_decap_8 FILLER_16_648 ();
 sg13g2_decap_8 FILLER_16_655 ();
 sg13g2_decap_8 FILLER_16_662 ();
 sg13g2_decap_8 FILLER_16_669 ();
 sg13g2_decap_8 FILLER_16_676 ();
 sg13g2_decap_8 FILLER_16_683 ();
 sg13g2_decap_8 FILLER_16_690 ();
 sg13g2_decap_8 FILLER_16_697 ();
 sg13g2_decap_8 FILLER_16_704 ();
 sg13g2_decap_8 FILLER_16_711 ();
 sg13g2_decap_8 FILLER_16_718 ();
 sg13g2_decap_8 FILLER_16_725 ();
 sg13g2_decap_8 FILLER_16_732 ();
 sg13g2_decap_8 FILLER_16_739 ();
 sg13g2_decap_8 FILLER_16_746 ();
 sg13g2_decap_8 FILLER_16_753 ();
 sg13g2_decap_8 FILLER_16_760 ();
 sg13g2_decap_8 FILLER_16_767 ();
 sg13g2_decap_8 FILLER_16_774 ();
 sg13g2_decap_8 FILLER_16_781 ();
 sg13g2_decap_8 FILLER_16_788 ();
 sg13g2_decap_8 FILLER_16_795 ();
 sg13g2_decap_8 FILLER_16_802 ();
 sg13g2_decap_8 FILLER_16_809 ();
 sg13g2_decap_8 FILLER_16_816 ();
 sg13g2_decap_8 FILLER_16_823 ();
 sg13g2_decap_8 FILLER_16_830 ();
 sg13g2_decap_8 FILLER_16_837 ();
 sg13g2_decap_8 FILLER_16_844 ();
 sg13g2_decap_8 FILLER_16_851 ();
 sg13g2_decap_8 FILLER_16_858 ();
 sg13g2_decap_8 FILLER_16_865 ();
 sg13g2_decap_8 FILLER_16_872 ();
 sg13g2_decap_8 FILLER_16_879 ();
 sg13g2_decap_8 FILLER_16_886 ();
 sg13g2_decap_8 FILLER_16_893 ();
 sg13g2_decap_8 FILLER_16_900 ();
 sg13g2_decap_8 FILLER_16_907 ();
 sg13g2_decap_8 FILLER_16_914 ();
 sg13g2_decap_4 FILLER_16_921 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_decap_8 FILLER_17_49 ();
 sg13g2_decap_8 FILLER_17_56 ();
 sg13g2_decap_8 FILLER_17_63 ();
 sg13g2_decap_8 FILLER_17_70 ();
 sg13g2_decap_8 FILLER_17_77 ();
 sg13g2_decap_8 FILLER_17_84 ();
 sg13g2_decap_8 FILLER_17_91 ();
 sg13g2_decap_8 FILLER_17_98 ();
 sg13g2_decap_8 FILLER_17_105 ();
 sg13g2_decap_8 FILLER_17_112 ();
 sg13g2_decap_8 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_133 ();
 sg13g2_decap_8 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_147 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_8 FILLER_17_161 ();
 sg13g2_decap_8 FILLER_17_168 ();
 sg13g2_decap_8 FILLER_17_175 ();
 sg13g2_decap_8 FILLER_17_182 ();
 sg13g2_decap_8 FILLER_17_189 ();
 sg13g2_decap_8 FILLER_17_196 ();
 sg13g2_decap_8 FILLER_17_203 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_decap_8 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_231 ();
 sg13g2_decap_8 FILLER_17_238 ();
 sg13g2_decap_8 FILLER_17_245 ();
 sg13g2_decap_8 FILLER_17_252 ();
 sg13g2_decap_8 FILLER_17_259 ();
 sg13g2_decap_8 FILLER_17_266 ();
 sg13g2_decap_8 FILLER_17_273 ();
 sg13g2_decap_8 FILLER_17_280 ();
 sg13g2_decap_8 FILLER_17_287 ();
 sg13g2_decap_8 FILLER_17_294 ();
 sg13g2_decap_8 FILLER_17_301 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_decap_8 FILLER_17_315 ();
 sg13g2_decap_8 FILLER_17_322 ();
 sg13g2_decap_8 FILLER_17_329 ();
 sg13g2_decap_8 FILLER_17_336 ();
 sg13g2_decap_8 FILLER_17_343 ();
 sg13g2_decap_8 FILLER_17_350 ();
 sg13g2_decap_8 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_8 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_378 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_decap_8 FILLER_17_427 ();
 sg13g2_decap_8 FILLER_17_434 ();
 sg13g2_decap_8 FILLER_17_441 ();
 sg13g2_decap_8 FILLER_17_448 ();
 sg13g2_decap_8 FILLER_17_455 ();
 sg13g2_decap_8 FILLER_17_462 ();
 sg13g2_decap_8 FILLER_17_469 ();
 sg13g2_decap_8 FILLER_17_476 ();
 sg13g2_decap_8 FILLER_17_483 ();
 sg13g2_decap_8 FILLER_17_490 ();
 sg13g2_decap_8 FILLER_17_497 ();
 sg13g2_decap_8 FILLER_17_504 ();
 sg13g2_decap_8 FILLER_17_511 ();
 sg13g2_decap_8 FILLER_17_518 ();
 sg13g2_decap_8 FILLER_17_525 ();
 sg13g2_decap_8 FILLER_17_532 ();
 sg13g2_decap_8 FILLER_17_539 ();
 sg13g2_decap_8 FILLER_17_546 ();
 sg13g2_decap_8 FILLER_17_553 ();
 sg13g2_decap_8 FILLER_17_560 ();
 sg13g2_decap_8 FILLER_17_567 ();
 sg13g2_decap_8 FILLER_17_574 ();
 sg13g2_decap_8 FILLER_17_581 ();
 sg13g2_decap_8 FILLER_17_588 ();
 sg13g2_decap_8 FILLER_17_595 ();
 sg13g2_decap_8 FILLER_17_602 ();
 sg13g2_decap_8 FILLER_17_609 ();
 sg13g2_decap_8 FILLER_17_616 ();
 sg13g2_decap_8 FILLER_17_623 ();
 sg13g2_decap_8 FILLER_17_630 ();
 sg13g2_decap_8 FILLER_17_637 ();
 sg13g2_decap_8 FILLER_17_644 ();
 sg13g2_decap_8 FILLER_17_651 ();
 sg13g2_decap_8 FILLER_17_658 ();
 sg13g2_decap_8 FILLER_17_665 ();
 sg13g2_decap_8 FILLER_17_672 ();
 sg13g2_decap_8 FILLER_17_679 ();
 sg13g2_decap_8 FILLER_17_686 ();
 sg13g2_decap_8 FILLER_17_693 ();
 sg13g2_decap_8 FILLER_17_700 ();
 sg13g2_decap_8 FILLER_17_707 ();
 sg13g2_decap_8 FILLER_17_714 ();
 sg13g2_decap_8 FILLER_17_721 ();
 sg13g2_decap_8 FILLER_17_728 ();
 sg13g2_decap_8 FILLER_17_735 ();
 sg13g2_decap_8 FILLER_17_742 ();
 sg13g2_decap_8 FILLER_17_749 ();
 sg13g2_decap_8 FILLER_17_756 ();
 sg13g2_decap_8 FILLER_17_763 ();
 sg13g2_decap_8 FILLER_17_770 ();
 sg13g2_decap_8 FILLER_17_777 ();
 sg13g2_decap_8 FILLER_17_784 ();
 sg13g2_decap_8 FILLER_17_791 ();
 sg13g2_decap_8 FILLER_17_798 ();
 sg13g2_decap_8 FILLER_17_805 ();
 sg13g2_decap_8 FILLER_17_812 ();
 sg13g2_decap_8 FILLER_17_819 ();
 sg13g2_decap_8 FILLER_17_826 ();
 sg13g2_decap_8 FILLER_17_833 ();
 sg13g2_decap_8 FILLER_17_840 ();
 sg13g2_decap_8 FILLER_17_847 ();
 sg13g2_decap_8 FILLER_17_854 ();
 sg13g2_decap_8 FILLER_17_861 ();
 sg13g2_decap_8 FILLER_17_868 ();
 sg13g2_decap_8 FILLER_17_875 ();
 sg13g2_decap_8 FILLER_17_882 ();
 sg13g2_decap_8 FILLER_17_889 ();
 sg13g2_decap_8 FILLER_17_896 ();
 sg13g2_decap_8 FILLER_17_903 ();
 sg13g2_decap_8 FILLER_17_910 ();
 sg13g2_decap_8 FILLER_17_917 ();
 sg13g2_fill_1 FILLER_17_924 ();
 sg13g2_decap_8 FILLER_18_4 ();
 sg13g2_decap_8 FILLER_18_11 ();
 sg13g2_decap_8 FILLER_18_18 ();
 sg13g2_decap_8 FILLER_18_25 ();
 sg13g2_decap_8 FILLER_18_32 ();
 sg13g2_decap_8 FILLER_18_39 ();
 sg13g2_decap_8 FILLER_18_46 ();
 sg13g2_decap_8 FILLER_18_53 ();
 sg13g2_decap_8 FILLER_18_60 ();
 sg13g2_decap_8 FILLER_18_67 ();
 sg13g2_decap_8 FILLER_18_74 ();
 sg13g2_decap_8 FILLER_18_81 ();
 sg13g2_decap_8 FILLER_18_88 ();
 sg13g2_decap_8 FILLER_18_95 ();
 sg13g2_decap_8 FILLER_18_102 ();
 sg13g2_decap_8 FILLER_18_109 ();
 sg13g2_decap_8 FILLER_18_116 ();
 sg13g2_decap_8 FILLER_18_123 ();
 sg13g2_decap_8 FILLER_18_130 ();
 sg13g2_decap_8 FILLER_18_137 ();
 sg13g2_decap_8 FILLER_18_144 ();
 sg13g2_decap_8 FILLER_18_151 ();
 sg13g2_decap_8 FILLER_18_158 ();
 sg13g2_decap_8 FILLER_18_165 ();
 sg13g2_decap_8 FILLER_18_172 ();
 sg13g2_decap_8 FILLER_18_179 ();
 sg13g2_decap_8 FILLER_18_186 ();
 sg13g2_decap_8 FILLER_18_193 ();
 sg13g2_decap_8 FILLER_18_200 ();
 sg13g2_decap_8 FILLER_18_207 ();
 sg13g2_decap_8 FILLER_18_214 ();
 sg13g2_decap_8 FILLER_18_221 ();
 sg13g2_decap_8 FILLER_18_228 ();
 sg13g2_decap_8 FILLER_18_235 ();
 sg13g2_decap_8 FILLER_18_242 ();
 sg13g2_decap_8 FILLER_18_249 ();
 sg13g2_decap_8 FILLER_18_256 ();
 sg13g2_decap_8 FILLER_18_263 ();
 sg13g2_decap_8 FILLER_18_270 ();
 sg13g2_decap_8 FILLER_18_277 ();
 sg13g2_decap_8 FILLER_18_284 ();
 sg13g2_decap_8 FILLER_18_291 ();
 sg13g2_decap_8 FILLER_18_298 ();
 sg13g2_decap_8 FILLER_18_305 ();
 sg13g2_decap_8 FILLER_18_312 ();
 sg13g2_decap_8 FILLER_18_319 ();
 sg13g2_decap_8 FILLER_18_326 ();
 sg13g2_decap_8 FILLER_18_333 ();
 sg13g2_decap_8 FILLER_18_340 ();
 sg13g2_decap_8 FILLER_18_347 ();
 sg13g2_decap_8 FILLER_18_354 ();
 sg13g2_decap_8 FILLER_18_361 ();
 sg13g2_decap_8 FILLER_18_368 ();
 sg13g2_decap_8 FILLER_18_375 ();
 sg13g2_decap_8 FILLER_18_382 ();
 sg13g2_decap_8 FILLER_18_389 ();
 sg13g2_decap_8 FILLER_18_396 ();
 sg13g2_decap_8 FILLER_18_403 ();
 sg13g2_decap_8 FILLER_18_410 ();
 sg13g2_decap_8 FILLER_18_417 ();
 sg13g2_decap_8 FILLER_18_424 ();
 sg13g2_decap_8 FILLER_18_431 ();
 sg13g2_decap_8 FILLER_18_438 ();
 sg13g2_decap_8 FILLER_18_445 ();
 sg13g2_decap_8 FILLER_18_452 ();
 sg13g2_decap_8 FILLER_18_459 ();
 sg13g2_decap_8 FILLER_18_466 ();
 sg13g2_decap_8 FILLER_18_473 ();
 sg13g2_decap_8 FILLER_18_480 ();
 sg13g2_decap_8 FILLER_18_487 ();
 sg13g2_decap_8 FILLER_18_494 ();
 sg13g2_decap_8 FILLER_18_501 ();
 sg13g2_decap_8 FILLER_18_508 ();
 sg13g2_decap_8 FILLER_18_515 ();
 sg13g2_decap_8 FILLER_18_522 ();
 sg13g2_decap_8 FILLER_18_529 ();
 sg13g2_decap_8 FILLER_18_536 ();
 sg13g2_decap_8 FILLER_18_543 ();
 sg13g2_decap_8 FILLER_18_550 ();
 sg13g2_decap_8 FILLER_18_557 ();
 sg13g2_decap_8 FILLER_18_564 ();
 sg13g2_decap_8 FILLER_18_571 ();
 sg13g2_decap_8 FILLER_18_578 ();
 sg13g2_decap_8 FILLER_18_585 ();
 sg13g2_decap_8 FILLER_18_592 ();
 sg13g2_decap_8 FILLER_18_599 ();
 sg13g2_decap_8 FILLER_18_606 ();
 sg13g2_decap_8 FILLER_18_613 ();
 sg13g2_decap_8 FILLER_18_620 ();
 sg13g2_decap_8 FILLER_18_627 ();
 sg13g2_decap_8 FILLER_18_634 ();
 sg13g2_decap_8 FILLER_18_641 ();
 sg13g2_decap_8 FILLER_18_648 ();
 sg13g2_decap_8 FILLER_18_655 ();
 sg13g2_decap_8 FILLER_18_662 ();
 sg13g2_decap_8 FILLER_18_669 ();
 sg13g2_decap_8 FILLER_18_676 ();
 sg13g2_decap_8 FILLER_18_683 ();
 sg13g2_decap_8 FILLER_18_690 ();
 sg13g2_decap_8 FILLER_18_697 ();
 sg13g2_decap_8 FILLER_18_704 ();
 sg13g2_decap_8 FILLER_18_711 ();
 sg13g2_decap_8 FILLER_18_718 ();
 sg13g2_decap_8 FILLER_18_725 ();
 sg13g2_decap_8 FILLER_18_732 ();
 sg13g2_decap_8 FILLER_18_739 ();
 sg13g2_decap_8 FILLER_18_746 ();
 sg13g2_decap_8 FILLER_18_753 ();
 sg13g2_decap_8 FILLER_18_760 ();
 sg13g2_decap_8 FILLER_18_767 ();
 sg13g2_decap_8 FILLER_18_774 ();
 sg13g2_decap_8 FILLER_18_781 ();
 sg13g2_decap_8 FILLER_18_788 ();
 sg13g2_decap_8 FILLER_18_795 ();
 sg13g2_decap_8 FILLER_18_802 ();
 sg13g2_decap_8 FILLER_18_809 ();
 sg13g2_decap_8 FILLER_18_816 ();
 sg13g2_decap_8 FILLER_18_823 ();
 sg13g2_decap_8 FILLER_18_830 ();
 sg13g2_decap_8 FILLER_18_837 ();
 sg13g2_decap_8 FILLER_18_844 ();
 sg13g2_decap_8 FILLER_18_851 ();
 sg13g2_decap_8 FILLER_18_858 ();
 sg13g2_decap_8 FILLER_18_865 ();
 sg13g2_decap_8 FILLER_18_872 ();
 sg13g2_decap_8 FILLER_18_879 ();
 sg13g2_decap_8 FILLER_18_886 ();
 sg13g2_decap_8 FILLER_18_893 ();
 sg13g2_decap_8 FILLER_18_900 ();
 sg13g2_decap_8 FILLER_18_907 ();
 sg13g2_decap_8 FILLER_18_914 ();
 sg13g2_decap_4 FILLER_18_921 ();
 sg13g2_decap_8 FILLER_19_4 ();
 sg13g2_decap_8 FILLER_19_11 ();
 sg13g2_decap_8 FILLER_19_18 ();
 sg13g2_decap_8 FILLER_19_25 ();
 sg13g2_decap_8 FILLER_19_32 ();
 sg13g2_decap_8 FILLER_19_39 ();
 sg13g2_decap_8 FILLER_19_46 ();
 sg13g2_decap_8 FILLER_19_53 ();
 sg13g2_decap_8 FILLER_19_60 ();
 sg13g2_decap_8 FILLER_19_67 ();
 sg13g2_decap_8 FILLER_19_74 ();
 sg13g2_decap_8 FILLER_19_81 ();
 sg13g2_decap_8 FILLER_19_88 ();
 sg13g2_decap_8 FILLER_19_95 ();
 sg13g2_decap_8 FILLER_19_102 ();
 sg13g2_decap_8 FILLER_19_109 ();
 sg13g2_decap_8 FILLER_19_116 ();
 sg13g2_decap_8 FILLER_19_123 ();
 sg13g2_decap_8 FILLER_19_130 ();
 sg13g2_decap_8 FILLER_19_137 ();
 sg13g2_decap_8 FILLER_19_144 ();
 sg13g2_decap_8 FILLER_19_151 ();
 sg13g2_decap_8 FILLER_19_158 ();
 sg13g2_decap_8 FILLER_19_165 ();
 sg13g2_decap_8 FILLER_19_172 ();
 sg13g2_decap_8 FILLER_19_179 ();
 sg13g2_decap_8 FILLER_19_186 ();
 sg13g2_decap_8 FILLER_19_193 ();
 sg13g2_decap_8 FILLER_19_200 ();
 sg13g2_decap_8 FILLER_19_207 ();
 sg13g2_decap_8 FILLER_19_214 ();
 sg13g2_decap_8 FILLER_19_221 ();
 sg13g2_decap_8 FILLER_19_228 ();
 sg13g2_decap_8 FILLER_19_235 ();
 sg13g2_decap_8 FILLER_19_242 ();
 sg13g2_decap_8 FILLER_19_249 ();
 sg13g2_decap_8 FILLER_19_256 ();
 sg13g2_decap_8 FILLER_19_263 ();
 sg13g2_decap_8 FILLER_19_270 ();
 sg13g2_decap_8 FILLER_19_277 ();
 sg13g2_decap_8 FILLER_19_284 ();
 sg13g2_decap_8 FILLER_19_291 ();
 sg13g2_decap_8 FILLER_19_298 ();
 sg13g2_decap_8 FILLER_19_305 ();
 sg13g2_decap_8 FILLER_19_312 ();
 sg13g2_decap_8 FILLER_19_319 ();
 sg13g2_decap_8 FILLER_19_326 ();
 sg13g2_decap_8 FILLER_19_333 ();
 sg13g2_decap_8 FILLER_19_340 ();
 sg13g2_decap_8 FILLER_19_347 ();
 sg13g2_decap_8 FILLER_19_354 ();
 sg13g2_decap_8 FILLER_19_361 ();
 sg13g2_decap_8 FILLER_19_368 ();
 sg13g2_decap_8 FILLER_19_375 ();
 sg13g2_decap_8 FILLER_19_382 ();
 sg13g2_decap_8 FILLER_19_389 ();
 sg13g2_decap_8 FILLER_19_396 ();
 sg13g2_decap_8 FILLER_19_403 ();
 sg13g2_decap_8 FILLER_19_410 ();
 sg13g2_decap_8 FILLER_19_417 ();
 sg13g2_decap_8 FILLER_19_424 ();
 sg13g2_decap_8 FILLER_19_431 ();
 sg13g2_decap_8 FILLER_19_438 ();
 sg13g2_decap_8 FILLER_19_445 ();
 sg13g2_decap_8 FILLER_19_452 ();
 sg13g2_decap_8 FILLER_19_459 ();
 sg13g2_decap_8 FILLER_19_466 ();
 sg13g2_decap_8 FILLER_19_473 ();
 sg13g2_decap_8 FILLER_19_480 ();
 sg13g2_decap_8 FILLER_19_487 ();
 sg13g2_decap_8 FILLER_19_494 ();
 sg13g2_decap_8 FILLER_19_501 ();
 sg13g2_decap_8 FILLER_19_508 ();
 sg13g2_decap_8 FILLER_19_515 ();
 sg13g2_decap_8 FILLER_19_522 ();
 sg13g2_decap_8 FILLER_19_529 ();
 sg13g2_decap_8 FILLER_19_536 ();
 sg13g2_decap_8 FILLER_19_543 ();
 sg13g2_decap_8 FILLER_19_550 ();
 sg13g2_decap_8 FILLER_19_557 ();
 sg13g2_decap_8 FILLER_19_564 ();
 sg13g2_decap_8 FILLER_19_571 ();
 sg13g2_decap_8 FILLER_19_578 ();
 sg13g2_decap_8 FILLER_19_585 ();
 sg13g2_decap_8 FILLER_19_592 ();
 sg13g2_decap_8 FILLER_19_599 ();
 sg13g2_decap_8 FILLER_19_606 ();
 sg13g2_decap_8 FILLER_19_613 ();
 sg13g2_decap_8 FILLER_19_620 ();
 sg13g2_decap_8 FILLER_19_627 ();
 sg13g2_decap_8 FILLER_19_634 ();
 sg13g2_decap_8 FILLER_19_641 ();
 sg13g2_decap_8 FILLER_19_648 ();
 sg13g2_decap_8 FILLER_19_655 ();
 sg13g2_decap_8 FILLER_19_662 ();
 sg13g2_decap_8 FILLER_19_669 ();
 sg13g2_decap_8 FILLER_19_676 ();
 sg13g2_decap_8 FILLER_19_683 ();
 sg13g2_decap_8 FILLER_19_690 ();
 sg13g2_decap_8 FILLER_19_697 ();
 sg13g2_decap_8 FILLER_19_704 ();
 sg13g2_decap_8 FILLER_19_711 ();
 sg13g2_decap_8 FILLER_19_718 ();
 sg13g2_decap_8 FILLER_19_725 ();
 sg13g2_decap_8 FILLER_19_732 ();
 sg13g2_decap_8 FILLER_19_739 ();
 sg13g2_decap_8 FILLER_19_746 ();
 sg13g2_decap_8 FILLER_19_753 ();
 sg13g2_decap_8 FILLER_19_760 ();
 sg13g2_decap_8 FILLER_19_767 ();
 sg13g2_decap_8 FILLER_19_774 ();
 sg13g2_decap_8 FILLER_19_781 ();
 sg13g2_decap_8 FILLER_19_788 ();
 sg13g2_decap_8 FILLER_19_795 ();
 sg13g2_decap_8 FILLER_19_802 ();
 sg13g2_decap_8 FILLER_19_809 ();
 sg13g2_decap_8 FILLER_19_816 ();
 sg13g2_decap_8 FILLER_19_823 ();
 sg13g2_decap_8 FILLER_19_830 ();
 sg13g2_decap_8 FILLER_19_837 ();
 sg13g2_decap_8 FILLER_19_844 ();
 sg13g2_decap_8 FILLER_19_851 ();
 sg13g2_decap_8 FILLER_19_858 ();
 sg13g2_decap_8 FILLER_19_865 ();
 sg13g2_decap_8 FILLER_19_872 ();
 sg13g2_decap_8 FILLER_19_879 ();
 sg13g2_decap_8 FILLER_19_886 ();
 sg13g2_decap_8 FILLER_19_893 ();
 sg13g2_decap_8 FILLER_19_900 ();
 sg13g2_decap_8 FILLER_19_907 ();
 sg13g2_decap_8 FILLER_19_914 ();
 sg13g2_decap_4 FILLER_19_921 ();
 sg13g2_decap_8 FILLER_20_4 ();
 sg13g2_decap_8 FILLER_20_11 ();
 sg13g2_decap_8 FILLER_20_18 ();
 sg13g2_decap_8 FILLER_20_25 ();
 sg13g2_decap_8 FILLER_20_32 ();
 sg13g2_decap_8 FILLER_20_39 ();
 sg13g2_decap_8 FILLER_20_46 ();
 sg13g2_decap_8 FILLER_20_53 ();
 sg13g2_decap_8 FILLER_20_60 ();
 sg13g2_decap_8 FILLER_20_67 ();
 sg13g2_decap_8 FILLER_20_74 ();
 sg13g2_decap_8 FILLER_20_81 ();
 sg13g2_decap_8 FILLER_20_88 ();
 sg13g2_decap_8 FILLER_20_95 ();
 sg13g2_decap_8 FILLER_20_102 ();
 sg13g2_decap_8 FILLER_20_109 ();
 sg13g2_decap_8 FILLER_20_116 ();
 sg13g2_decap_8 FILLER_20_123 ();
 sg13g2_decap_8 FILLER_20_130 ();
 sg13g2_decap_8 FILLER_20_137 ();
 sg13g2_decap_8 FILLER_20_144 ();
 sg13g2_decap_8 FILLER_20_151 ();
 sg13g2_decap_8 FILLER_20_158 ();
 sg13g2_decap_8 FILLER_20_165 ();
 sg13g2_decap_8 FILLER_20_172 ();
 sg13g2_decap_8 FILLER_20_179 ();
 sg13g2_decap_8 FILLER_20_186 ();
 sg13g2_decap_8 FILLER_20_193 ();
 sg13g2_decap_8 FILLER_20_200 ();
 sg13g2_decap_8 FILLER_20_207 ();
 sg13g2_decap_8 FILLER_20_214 ();
 sg13g2_decap_8 FILLER_20_221 ();
 sg13g2_decap_8 FILLER_20_228 ();
 sg13g2_decap_8 FILLER_20_235 ();
 sg13g2_decap_8 FILLER_20_242 ();
 sg13g2_decap_8 FILLER_20_249 ();
 sg13g2_decap_8 FILLER_20_256 ();
 sg13g2_decap_8 FILLER_20_263 ();
 sg13g2_decap_8 FILLER_20_270 ();
 sg13g2_decap_8 FILLER_20_277 ();
 sg13g2_decap_8 FILLER_20_284 ();
 sg13g2_decap_8 FILLER_20_291 ();
 sg13g2_decap_8 FILLER_20_298 ();
 sg13g2_decap_8 FILLER_20_305 ();
 sg13g2_decap_8 FILLER_20_312 ();
 sg13g2_decap_8 FILLER_20_319 ();
 sg13g2_decap_8 FILLER_20_326 ();
 sg13g2_decap_8 FILLER_20_333 ();
 sg13g2_decap_8 FILLER_20_340 ();
 sg13g2_decap_8 FILLER_20_347 ();
 sg13g2_decap_8 FILLER_20_354 ();
 sg13g2_decap_8 FILLER_20_361 ();
 sg13g2_decap_8 FILLER_20_368 ();
 sg13g2_decap_8 FILLER_20_375 ();
 sg13g2_decap_8 FILLER_20_382 ();
 sg13g2_decap_8 FILLER_20_389 ();
 sg13g2_decap_8 FILLER_20_396 ();
 sg13g2_decap_8 FILLER_20_403 ();
 sg13g2_decap_8 FILLER_20_410 ();
 sg13g2_decap_8 FILLER_20_417 ();
 sg13g2_decap_8 FILLER_20_424 ();
 sg13g2_decap_8 FILLER_20_431 ();
 sg13g2_decap_8 FILLER_20_438 ();
 sg13g2_decap_8 FILLER_20_445 ();
 sg13g2_decap_8 FILLER_20_452 ();
 sg13g2_decap_8 FILLER_20_459 ();
 sg13g2_decap_8 FILLER_20_466 ();
 sg13g2_decap_8 FILLER_20_473 ();
 sg13g2_decap_8 FILLER_20_480 ();
 sg13g2_decap_8 FILLER_20_487 ();
 sg13g2_decap_8 FILLER_20_494 ();
 sg13g2_decap_8 FILLER_20_501 ();
 sg13g2_decap_8 FILLER_20_508 ();
 sg13g2_decap_8 FILLER_20_515 ();
 sg13g2_decap_8 FILLER_20_522 ();
 sg13g2_decap_8 FILLER_20_529 ();
 sg13g2_decap_8 FILLER_20_536 ();
 sg13g2_decap_8 FILLER_20_543 ();
 sg13g2_decap_8 FILLER_20_550 ();
 sg13g2_decap_8 FILLER_20_557 ();
 sg13g2_decap_8 FILLER_20_564 ();
 sg13g2_decap_8 FILLER_20_571 ();
 sg13g2_decap_8 FILLER_20_578 ();
 sg13g2_decap_8 FILLER_20_585 ();
 sg13g2_decap_8 FILLER_20_592 ();
 sg13g2_decap_8 FILLER_20_599 ();
 sg13g2_decap_8 FILLER_20_606 ();
 sg13g2_decap_8 FILLER_20_613 ();
 sg13g2_decap_8 FILLER_20_620 ();
 sg13g2_decap_8 FILLER_20_627 ();
 sg13g2_decap_8 FILLER_20_634 ();
 sg13g2_decap_8 FILLER_20_641 ();
 sg13g2_decap_8 FILLER_20_648 ();
 sg13g2_decap_8 FILLER_20_655 ();
 sg13g2_decap_8 FILLER_20_662 ();
 sg13g2_decap_8 FILLER_20_669 ();
 sg13g2_decap_8 FILLER_20_676 ();
 sg13g2_decap_8 FILLER_20_683 ();
 sg13g2_decap_8 FILLER_20_690 ();
 sg13g2_decap_8 FILLER_20_697 ();
 sg13g2_decap_8 FILLER_20_704 ();
 sg13g2_decap_8 FILLER_20_711 ();
 sg13g2_decap_8 FILLER_20_718 ();
 sg13g2_decap_8 FILLER_20_725 ();
 sg13g2_decap_8 FILLER_20_732 ();
 sg13g2_decap_8 FILLER_20_739 ();
 sg13g2_decap_8 FILLER_20_746 ();
 sg13g2_decap_8 FILLER_20_753 ();
 sg13g2_decap_8 FILLER_20_760 ();
 sg13g2_decap_8 FILLER_20_767 ();
 sg13g2_decap_8 FILLER_20_774 ();
 sg13g2_decap_8 FILLER_20_781 ();
 sg13g2_decap_8 FILLER_20_788 ();
 sg13g2_decap_8 FILLER_20_795 ();
 sg13g2_decap_8 FILLER_20_802 ();
 sg13g2_decap_8 FILLER_20_809 ();
 sg13g2_decap_8 FILLER_20_816 ();
 sg13g2_decap_8 FILLER_20_823 ();
 sg13g2_decap_8 FILLER_20_830 ();
 sg13g2_decap_8 FILLER_20_837 ();
 sg13g2_decap_8 FILLER_20_844 ();
 sg13g2_decap_8 FILLER_20_851 ();
 sg13g2_decap_8 FILLER_20_858 ();
 sg13g2_decap_8 FILLER_20_865 ();
 sg13g2_decap_8 FILLER_20_872 ();
 sg13g2_decap_8 FILLER_20_879 ();
 sg13g2_decap_8 FILLER_20_886 ();
 sg13g2_decap_8 FILLER_20_893 ();
 sg13g2_decap_8 FILLER_20_900 ();
 sg13g2_decap_8 FILLER_20_907 ();
 sg13g2_decap_8 FILLER_20_914 ();
 sg13g2_decap_4 FILLER_20_921 ();
 sg13g2_decap_8 FILLER_21_4 ();
 sg13g2_decap_8 FILLER_21_11 ();
 sg13g2_decap_8 FILLER_21_18 ();
 sg13g2_decap_8 FILLER_21_25 ();
 sg13g2_decap_8 FILLER_21_32 ();
 sg13g2_decap_8 FILLER_21_39 ();
 sg13g2_decap_8 FILLER_21_46 ();
 sg13g2_decap_8 FILLER_21_53 ();
 sg13g2_decap_8 FILLER_21_60 ();
 sg13g2_decap_8 FILLER_21_67 ();
 sg13g2_decap_8 FILLER_21_74 ();
 sg13g2_decap_8 FILLER_21_81 ();
 sg13g2_decap_8 FILLER_21_88 ();
 sg13g2_decap_8 FILLER_21_95 ();
 sg13g2_decap_8 FILLER_21_102 ();
 sg13g2_decap_8 FILLER_21_109 ();
 sg13g2_decap_8 FILLER_21_116 ();
 sg13g2_decap_8 FILLER_21_123 ();
 sg13g2_decap_8 FILLER_21_130 ();
 sg13g2_decap_8 FILLER_21_137 ();
 sg13g2_decap_8 FILLER_21_144 ();
 sg13g2_decap_8 FILLER_21_151 ();
 sg13g2_decap_8 FILLER_21_158 ();
 sg13g2_decap_8 FILLER_21_165 ();
 sg13g2_decap_8 FILLER_21_172 ();
 sg13g2_decap_8 FILLER_21_179 ();
 sg13g2_decap_8 FILLER_21_186 ();
 sg13g2_decap_8 FILLER_21_193 ();
 sg13g2_decap_8 FILLER_21_200 ();
 sg13g2_decap_8 FILLER_21_207 ();
 sg13g2_decap_8 FILLER_21_214 ();
 sg13g2_decap_8 FILLER_21_221 ();
 sg13g2_decap_8 FILLER_21_228 ();
 sg13g2_decap_8 FILLER_21_235 ();
 sg13g2_decap_8 FILLER_21_242 ();
 sg13g2_decap_8 FILLER_21_249 ();
 sg13g2_decap_8 FILLER_21_256 ();
 sg13g2_decap_8 FILLER_21_263 ();
 sg13g2_decap_8 FILLER_21_270 ();
 sg13g2_decap_8 FILLER_21_277 ();
 sg13g2_decap_8 FILLER_21_284 ();
 sg13g2_decap_8 FILLER_21_291 ();
 sg13g2_decap_8 FILLER_21_298 ();
 sg13g2_decap_8 FILLER_21_305 ();
 sg13g2_decap_8 FILLER_21_312 ();
 sg13g2_decap_8 FILLER_21_319 ();
 sg13g2_decap_8 FILLER_21_326 ();
 sg13g2_decap_8 FILLER_21_333 ();
 sg13g2_decap_8 FILLER_21_340 ();
 sg13g2_decap_8 FILLER_21_347 ();
 sg13g2_decap_8 FILLER_21_354 ();
 sg13g2_decap_8 FILLER_21_361 ();
 sg13g2_decap_8 FILLER_21_368 ();
 sg13g2_decap_8 FILLER_21_375 ();
 sg13g2_decap_8 FILLER_21_382 ();
 sg13g2_decap_8 FILLER_21_389 ();
 sg13g2_decap_8 FILLER_21_396 ();
 sg13g2_decap_8 FILLER_21_403 ();
 sg13g2_decap_8 FILLER_21_410 ();
 sg13g2_decap_8 FILLER_21_417 ();
 sg13g2_decap_8 FILLER_21_424 ();
 sg13g2_decap_8 FILLER_21_431 ();
 sg13g2_decap_8 FILLER_21_438 ();
 sg13g2_decap_8 FILLER_21_445 ();
 sg13g2_decap_8 FILLER_21_452 ();
 sg13g2_decap_8 FILLER_21_459 ();
 sg13g2_decap_8 FILLER_21_466 ();
 sg13g2_decap_8 FILLER_21_473 ();
 sg13g2_decap_8 FILLER_21_480 ();
 sg13g2_decap_8 FILLER_21_487 ();
 sg13g2_decap_8 FILLER_21_494 ();
 sg13g2_decap_8 FILLER_21_501 ();
 sg13g2_decap_8 FILLER_21_508 ();
 sg13g2_decap_8 FILLER_21_515 ();
 sg13g2_decap_8 FILLER_21_522 ();
 sg13g2_decap_8 FILLER_21_529 ();
 sg13g2_decap_8 FILLER_21_536 ();
 sg13g2_decap_8 FILLER_21_543 ();
 sg13g2_decap_8 FILLER_21_550 ();
 sg13g2_decap_8 FILLER_21_557 ();
 sg13g2_decap_8 FILLER_21_564 ();
 sg13g2_decap_8 FILLER_21_571 ();
 sg13g2_decap_8 FILLER_21_578 ();
 sg13g2_decap_8 FILLER_21_585 ();
 sg13g2_decap_8 FILLER_21_592 ();
 sg13g2_decap_8 FILLER_21_599 ();
 sg13g2_decap_8 FILLER_21_606 ();
 sg13g2_decap_8 FILLER_21_613 ();
 sg13g2_decap_8 FILLER_21_620 ();
 sg13g2_decap_8 FILLER_21_627 ();
 sg13g2_decap_8 FILLER_21_634 ();
 sg13g2_decap_8 FILLER_21_641 ();
 sg13g2_decap_8 FILLER_21_648 ();
 sg13g2_decap_8 FILLER_21_655 ();
 sg13g2_decap_8 FILLER_21_662 ();
 sg13g2_decap_8 FILLER_21_669 ();
 sg13g2_decap_8 FILLER_21_676 ();
 sg13g2_decap_8 FILLER_21_683 ();
 sg13g2_decap_8 FILLER_21_690 ();
 sg13g2_decap_8 FILLER_21_697 ();
 sg13g2_decap_8 FILLER_21_704 ();
 sg13g2_decap_8 FILLER_21_711 ();
 sg13g2_decap_8 FILLER_21_718 ();
 sg13g2_decap_8 FILLER_21_725 ();
 sg13g2_decap_8 FILLER_21_732 ();
 sg13g2_decap_8 FILLER_21_739 ();
 sg13g2_decap_8 FILLER_21_746 ();
 sg13g2_decap_8 FILLER_21_753 ();
 sg13g2_decap_8 FILLER_21_760 ();
 sg13g2_decap_8 FILLER_21_767 ();
 sg13g2_decap_8 FILLER_21_774 ();
 sg13g2_decap_8 FILLER_21_781 ();
 sg13g2_decap_8 FILLER_21_788 ();
 sg13g2_decap_8 FILLER_21_795 ();
 sg13g2_decap_8 FILLER_21_802 ();
 sg13g2_decap_8 FILLER_21_809 ();
 sg13g2_decap_8 FILLER_21_816 ();
 sg13g2_decap_8 FILLER_21_823 ();
 sg13g2_decap_8 FILLER_21_830 ();
 sg13g2_decap_8 FILLER_21_837 ();
 sg13g2_decap_8 FILLER_21_844 ();
 sg13g2_decap_8 FILLER_21_851 ();
 sg13g2_decap_8 FILLER_21_858 ();
 sg13g2_decap_8 FILLER_21_865 ();
 sg13g2_decap_8 FILLER_21_872 ();
 sg13g2_decap_8 FILLER_21_879 ();
 sg13g2_decap_8 FILLER_21_886 ();
 sg13g2_decap_8 FILLER_21_893 ();
 sg13g2_decap_8 FILLER_21_900 ();
 sg13g2_decap_8 FILLER_21_907 ();
 sg13g2_decap_8 FILLER_21_914 ();
 sg13g2_decap_4 FILLER_21_921 ();
 sg13g2_decap_8 FILLER_22_4 ();
 sg13g2_decap_8 FILLER_22_11 ();
 sg13g2_decap_8 FILLER_22_18 ();
 sg13g2_decap_8 FILLER_22_25 ();
 sg13g2_decap_8 FILLER_22_32 ();
 sg13g2_decap_8 FILLER_22_39 ();
 sg13g2_decap_8 FILLER_22_46 ();
 sg13g2_decap_8 FILLER_22_53 ();
 sg13g2_decap_8 FILLER_22_60 ();
 sg13g2_decap_8 FILLER_22_67 ();
 sg13g2_decap_8 FILLER_22_74 ();
 sg13g2_decap_8 FILLER_22_81 ();
 sg13g2_decap_8 FILLER_22_88 ();
 sg13g2_decap_8 FILLER_22_95 ();
 sg13g2_decap_8 FILLER_22_102 ();
 sg13g2_decap_8 FILLER_22_109 ();
 sg13g2_decap_8 FILLER_22_116 ();
 sg13g2_decap_8 FILLER_22_123 ();
 sg13g2_decap_8 FILLER_22_130 ();
 sg13g2_decap_8 FILLER_22_137 ();
 sg13g2_decap_8 FILLER_22_144 ();
 sg13g2_decap_8 FILLER_22_151 ();
 sg13g2_decap_8 FILLER_22_158 ();
 sg13g2_decap_8 FILLER_22_165 ();
 sg13g2_decap_8 FILLER_22_172 ();
 sg13g2_decap_8 FILLER_22_179 ();
 sg13g2_decap_8 FILLER_22_186 ();
 sg13g2_decap_8 FILLER_22_193 ();
 sg13g2_decap_8 FILLER_22_200 ();
 sg13g2_decap_8 FILLER_22_207 ();
 sg13g2_decap_8 FILLER_22_214 ();
 sg13g2_decap_8 FILLER_22_221 ();
 sg13g2_decap_8 FILLER_22_228 ();
 sg13g2_decap_8 FILLER_22_235 ();
 sg13g2_decap_8 FILLER_22_242 ();
 sg13g2_decap_8 FILLER_22_249 ();
 sg13g2_decap_8 FILLER_22_256 ();
 sg13g2_decap_8 FILLER_22_263 ();
 sg13g2_decap_8 FILLER_22_270 ();
 sg13g2_decap_8 FILLER_22_277 ();
 sg13g2_decap_8 FILLER_22_284 ();
 sg13g2_decap_8 FILLER_22_291 ();
 sg13g2_decap_8 FILLER_22_298 ();
 sg13g2_decap_8 FILLER_22_305 ();
 sg13g2_decap_8 FILLER_22_312 ();
 sg13g2_decap_8 FILLER_22_319 ();
 sg13g2_decap_8 FILLER_22_326 ();
 sg13g2_decap_8 FILLER_22_333 ();
 sg13g2_decap_8 FILLER_22_340 ();
 sg13g2_decap_8 FILLER_22_347 ();
 sg13g2_decap_8 FILLER_22_354 ();
 sg13g2_decap_8 FILLER_22_361 ();
 sg13g2_decap_8 FILLER_22_368 ();
 sg13g2_decap_8 FILLER_22_375 ();
 sg13g2_decap_8 FILLER_22_382 ();
 sg13g2_decap_8 FILLER_22_389 ();
 sg13g2_decap_8 FILLER_22_396 ();
 sg13g2_decap_8 FILLER_22_403 ();
 sg13g2_decap_8 FILLER_22_410 ();
 sg13g2_decap_8 FILLER_22_417 ();
 sg13g2_decap_8 FILLER_22_424 ();
 sg13g2_decap_8 FILLER_22_431 ();
 sg13g2_decap_8 FILLER_22_438 ();
 sg13g2_decap_8 FILLER_22_445 ();
 sg13g2_decap_8 FILLER_22_452 ();
 sg13g2_decap_8 FILLER_22_459 ();
 sg13g2_decap_8 FILLER_22_466 ();
 sg13g2_decap_8 FILLER_22_473 ();
 sg13g2_decap_8 FILLER_22_480 ();
 sg13g2_decap_8 FILLER_22_487 ();
 sg13g2_decap_8 FILLER_22_494 ();
 sg13g2_decap_8 FILLER_22_501 ();
 sg13g2_decap_8 FILLER_22_508 ();
 sg13g2_decap_8 FILLER_22_515 ();
 sg13g2_decap_8 FILLER_22_522 ();
 sg13g2_decap_8 FILLER_22_529 ();
 sg13g2_decap_8 FILLER_22_536 ();
 sg13g2_decap_8 FILLER_22_543 ();
 sg13g2_decap_8 FILLER_22_550 ();
 sg13g2_decap_8 FILLER_22_557 ();
 sg13g2_decap_8 FILLER_22_564 ();
 sg13g2_decap_8 FILLER_22_571 ();
 sg13g2_decap_8 FILLER_22_578 ();
 sg13g2_decap_8 FILLER_22_585 ();
 sg13g2_decap_8 FILLER_22_592 ();
 sg13g2_decap_8 FILLER_22_599 ();
 sg13g2_decap_8 FILLER_22_606 ();
 sg13g2_decap_8 FILLER_22_613 ();
 sg13g2_decap_8 FILLER_22_620 ();
 sg13g2_decap_8 FILLER_22_627 ();
 sg13g2_decap_8 FILLER_22_634 ();
 sg13g2_decap_8 FILLER_22_641 ();
 sg13g2_decap_8 FILLER_22_648 ();
 sg13g2_decap_8 FILLER_22_655 ();
 sg13g2_decap_8 FILLER_22_662 ();
 sg13g2_decap_8 FILLER_22_669 ();
 sg13g2_decap_8 FILLER_22_676 ();
 sg13g2_decap_8 FILLER_22_683 ();
 sg13g2_decap_8 FILLER_22_690 ();
 sg13g2_decap_8 FILLER_22_697 ();
 sg13g2_decap_8 FILLER_22_704 ();
 sg13g2_decap_8 FILLER_22_711 ();
 sg13g2_decap_8 FILLER_22_718 ();
 sg13g2_decap_8 FILLER_22_725 ();
 sg13g2_decap_8 FILLER_22_732 ();
 sg13g2_decap_8 FILLER_22_739 ();
 sg13g2_decap_8 FILLER_22_746 ();
 sg13g2_decap_8 FILLER_22_753 ();
 sg13g2_decap_8 FILLER_22_760 ();
 sg13g2_decap_8 FILLER_22_767 ();
 sg13g2_decap_8 FILLER_22_774 ();
 sg13g2_decap_8 FILLER_22_781 ();
 sg13g2_decap_8 FILLER_22_788 ();
 sg13g2_decap_8 FILLER_22_795 ();
 sg13g2_decap_8 FILLER_22_802 ();
 sg13g2_decap_8 FILLER_22_809 ();
 sg13g2_decap_8 FILLER_22_816 ();
 sg13g2_decap_8 FILLER_22_823 ();
 sg13g2_decap_8 FILLER_22_830 ();
 sg13g2_decap_8 FILLER_22_837 ();
 sg13g2_decap_8 FILLER_22_844 ();
 sg13g2_decap_8 FILLER_22_851 ();
 sg13g2_decap_8 FILLER_22_858 ();
 sg13g2_decap_8 FILLER_22_865 ();
 sg13g2_decap_8 FILLER_22_872 ();
 sg13g2_decap_8 FILLER_22_879 ();
 sg13g2_decap_8 FILLER_22_886 ();
 sg13g2_decap_8 FILLER_22_893 ();
 sg13g2_decap_8 FILLER_22_900 ();
 sg13g2_decap_8 FILLER_22_907 ();
 sg13g2_decap_8 FILLER_22_914 ();
 sg13g2_decap_4 FILLER_22_921 ();
 sg13g2_decap_8 FILLER_23_4 ();
 sg13g2_decap_8 FILLER_23_11 ();
 sg13g2_decap_8 FILLER_23_18 ();
 sg13g2_decap_8 FILLER_23_25 ();
 sg13g2_decap_8 FILLER_23_32 ();
 sg13g2_decap_8 FILLER_23_39 ();
 sg13g2_decap_8 FILLER_23_46 ();
 sg13g2_decap_8 FILLER_23_53 ();
 sg13g2_decap_8 FILLER_23_60 ();
 sg13g2_decap_8 FILLER_23_67 ();
 sg13g2_decap_8 FILLER_23_74 ();
 sg13g2_decap_8 FILLER_23_81 ();
 sg13g2_decap_8 FILLER_23_88 ();
 sg13g2_decap_8 FILLER_23_95 ();
 sg13g2_decap_8 FILLER_23_102 ();
 sg13g2_decap_8 FILLER_23_109 ();
 sg13g2_decap_8 FILLER_23_116 ();
 sg13g2_decap_8 FILLER_23_123 ();
 sg13g2_decap_8 FILLER_23_130 ();
 sg13g2_decap_8 FILLER_23_137 ();
 sg13g2_decap_8 FILLER_23_144 ();
 sg13g2_decap_8 FILLER_23_151 ();
 sg13g2_decap_8 FILLER_23_158 ();
 sg13g2_decap_8 FILLER_23_165 ();
 sg13g2_decap_8 FILLER_23_172 ();
 sg13g2_decap_8 FILLER_23_179 ();
 sg13g2_decap_8 FILLER_23_186 ();
 sg13g2_decap_8 FILLER_23_193 ();
 sg13g2_decap_8 FILLER_23_200 ();
 sg13g2_decap_8 FILLER_23_207 ();
 sg13g2_decap_8 FILLER_23_214 ();
 sg13g2_decap_8 FILLER_23_221 ();
 sg13g2_decap_8 FILLER_23_228 ();
 sg13g2_decap_8 FILLER_23_235 ();
 sg13g2_decap_8 FILLER_23_242 ();
 sg13g2_decap_8 FILLER_23_249 ();
 sg13g2_decap_8 FILLER_23_256 ();
 sg13g2_decap_8 FILLER_23_263 ();
 sg13g2_decap_8 FILLER_23_270 ();
 sg13g2_decap_8 FILLER_23_277 ();
 sg13g2_decap_8 FILLER_23_284 ();
 sg13g2_decap_8 FILLER_23_291 ();
 sg13g2_decap_8 FILLER_23_298 ();
 sg13g2_decap_8 FILLER_23_305 ();
 sg13g2_decap_8 FILLER_23_312 ();
 sg13g2_decap_8 FILLER_23_319 ();
 sg13g2_decap_8 FILLER_23_326 ();
 sg13g2_decap_8 FILLER_23_333 ();
 sg13g2_decap_8 FILLER_23_340 ();
 sg13g2_decap_8 FILLER_23_347 ();
 sg13g2_decap_8 FILLER_23_354 ();
 sg13g2_decap_8 FILLER_23_361 ();
 sg13g2_decap_8 FILLER_23_368 ();
 sg13g2_decap_8 FILLER_23_375 ();
 sg13g2_decap_8 FILLER_23_382 ();
 sg13g2_decap_8 FILLER_23_389 ();
 sg13g2_decap_8 FILLER_23_396 ();
 sg13g2_decap_8 FILLER_23_403 ();
 sg13g2_decap_8 FILLER_23_410 ();
 sg13g2_decap_8 FILLER_23_417 ();
 sg13g2_decap_8 FILLER_23_424 ();
 sg13g2_decap_8 FILLER_23_431 ();
 sg13g2_decap_8 FILLER_23_438 ();
 sg13g2_decap_8 FILLER_23_445 ();
 sg13g2_decap_8 FILLER_23_452 ();
 sg13g2_decap_8 FILLER_23_459 ();
 sg13g2_decap_8 FILLER_23_466 ();
 sg13g2_decap_8 FILLER_23_473 ();
 sg13g2_decap_8 FILLER_23_480 ();
 sg13g2_decap_8 FILLER_23_487 ();
 sg13g2_decap_8 FILLER_23_494 ();
 sg13g2_decap_8 FILLER_23_501 ();
 sg13g2_decap_8 FILLER_23_508 ();
 sg13g2_decap_8 FILLER_23_515 ();
 sg13g2_decap_8 FILLER_23_522 ();
 sg13g2_decap_8 FILLER_23_529 ();
 sg13g2_decap_8 FILLER_23_536 ();
 sg13g2_decap_8 FILLER_23_543 ();
 sg13g2_decap_8 FILLER_23_550 ();
 sg13g2_decap_8 FILLER_23_557 ();
 sg13g2_decap_8 FILLER_23_564 ();
 sg13g2_decap_8 FILLER_23_571 ();
 sg13g2_decap_8 FILLER_23_578 ();
 sg13g2_decap_8 FILLER_23_585 ();
 sg13g2_decap_8 FILLER_23_592 ();
 sg13g2_decap_8 FILLER_23_599 ();
 sg13g2_decap_8 FILLER_23_606 ();
 sg13g2_decap_8 FILLER_23_613 ();
 sg13g2_decap_8 FILLER_23_620 ();
 sg13g2_decap_8 FILLER_23_627 ();
 sg13g2_decap_8 FILLER_23_634 ();
 sg13g2_decap_8 FILLER_23_641 ();
 sg13g2_decap_8 FILLER_23_648 ();
 sg13g2_decap_8 FILLER_23_655 ();
 sg13g2_decap_8 FILLER_23_662 ();
 sg13g2_decap_8 FILLER_23_669 ();
 sg13g2_decap_8 FILLER_23_676 ();
 sg13g2_decap_8 FILLER_23_683 ();
 sg13g2_decap_8 FILLER_23_690 ();
 sg13g2_decap_8 FILLER_23_697 ();
 sg13g2_decap_8 FILLER_23_704 ();
 sg13g2_decap_8 FILLER_23_711 ();
 sg13g2_decap_8 FILLER_23_718 ();
 sg13g2_decap_8 FILLER_23_725 ();
 sg13g2_decap_8 FILLER_23_732 ();
 sg13g2_decap_8 FILLER_23_739 ();
 sg13g2_decap_8 FILLER_23_746 ();
 sg13g2_decap_8 FILLER_23_753 ();
 sg13g2_decap_8 FILLER_23_760 ();
 sg13g2_decap_8 FILLER_23_767 ();
 sg13g2_decap_8 FILLER_23_774 ();
 sg13g2_decap_8 FILLER_23_781 ();
 sg13g2_decap_8 FILLER_23_788 ();
 sg13g2_decap_8 FILLER_23_795 ();
 sg13g2_decap_8 FILLER_23_802 ();
 sg13g2_decap_8 FILLER_23_809 ();
 sg13g2_decap_8 FILLER_23_816 ();
 sg13g2_decap_8 FILLER_23_823 ();
 sg13g2_decap_8 FILLER_23_830 ();
 sg13g2_decap_8 FILLER_23_837 ();
 sg13g2_decap_8 FILLER_23_844 ();
 sg13g2_decap_8 FILLER_23_851 ();
 sg13g2_decap_8 FILLER_23_858 ();
 sg13g2_decap_8 FILLER_23_865 ();
 sg13g2_decap_8 FILLER_23_872 ();
 sg13g2_decap_8 FILLER_23_879 ();
 sg13g2_decap_8 FILLER_23_886 ();
 sg13g2_decap_8 FILLER_23_893 ();
 sg13g2_decap_8 FILLER_23_900 ();
 sg13g2_decap_8 FILLER_23_907 ();
 sg13g2_decap_8 FILLER_23_914 ();
 sg13g2_decap_4 FILLER_23_921 ();
 sg13g2_decap_8 FILLER_24_4 ();
 sg13g2_decap_8 FILLER_24_11 ();
 sg13g2_decap_8 FILLER_24_18 ();
 sg13g2_decap_8 FILLER_24_25 ();
 sg13g2_decap_8 FILLER_24_32 ();
 sg13g2_decap_8 FILLER_24_39 ();
 sg13g2_decap_8 FILLER_24_46 ();
 sg13g2_decap_8 FILLER_24_53 ();
 sg13g2_decap_8 FILLER_24_60 ();
 sg13g2_decap_8 FILLER_24_67 ();
 sg13g2_fill_2 FILLER_24_74 ();
 sg13g2_fill_1 FILLER_24_76 ();
 sg13g2_decap_8 FILLER_24_82 ();
 sg13g2_decap_8 FILLER_24_89 ();
 sg13g2_decap_8 FILLER_24_96 ();
 sg13g2_decap_8 FILLER_24_103 ();
 sg13g2_decap_8 FILLER_24_110 ();
 sg13g2_decap_8 FILLER_24_117 ();
 sg13g2_decap_8 FILLER_24_124 ();
 sg13g2_decap_8 FILLER_24_131 ();
 sg13g2_decap_8 FILLER_24_138 ();
 sg13g2_decap_8 FILLER_24_145 ();
 sg13g2_decap_8 FILLER_24_152 ();
 sg13g2_decap_8 FILLER_24_159 ();
 sg13g2_decap_8 FILLER_24_166 ();
 sg13g2_decap_8 FILLER_24_173 ();
 sg13g2_decap_8 FILLER_24_180 ();
 sg13g2_decap_8 FILLER_24_187 ();
 sg13g2_decap_8 FILLER_24_194 ();
 sg13g2_decap_8 FILLER_24_201 ();
 sg13g2_decap_8 FILLER_24_208 ();
 sg13g2_decap_8 FILLER_24_215 ();
 sg13g2_decap_8 FILLER_24_222 ();
 sg13g2_decap_8 FILLER_24_229 ();
 sg13g2_decap_8 FILLER_24_236 ();
 sg13g2_decap_8 FILLER_24_243 ();
 sg13g2_decap_8 FILLER_24_250 ();
 sg13g2_decap_8 FILLER_24_257 ();
 sg13g2_decap_8 FILLER_24_264 ();
 sg13g2_decap_8 FILLER_24_271 ();
 sg13g2_decap_8 FILLER_24_278 ();
 sg13g2_decap_8 FILLER_24_285 ();
 sg13g2_decap_8 FILLER_24_292 ();
 sg13g2_decap_8 FILLER_24_299 ();
 sg13g2_decap_8 FILLER_24_306 ();
 sg13g2_decap_8 FILLER_24_313 ();
 sg13g2_decap_8 FILLER_24_320 ();
 sg13g2_decap_8 FILLER_24_327 ();
 sg13g2_decap_8 FILLER_24_334 ();
 sg13g2_decap_8 FILLER_24_341 ();
 sg13g2_decap_8 FILLER_24_348 ();
 sg13g2_decap_8 FILLER_24_355 ();
 sg13g2_decap_8 FILLER_24_362 ();
 sg13g2_decap_8 FILLER_24_369 ();
 sg13g2_decap_8 FILLER_24_376 ();
 sg13g2_decap_8 FILLER_24_383 ();
 sg13g2_decap_8 FILLER_24_390 ();
 sg13g2_decap_8 FILLER_24_397 ();
 sg13g2_decap_8 FILLER_24_404 ();
 sg13g2_decap_8 FILLER_24_411 ();
 sg13g2_decap_8 FILLER_24_418 ();
 sg13g2_decap_8 FILLER_24_425 ();
 sg13g2_decap_8 FILLER_24_432 ();
 sg13g2_decap_8 FILLER_24_439 ();
 sg13g2_decap_8 FILLER_24_446 ();
 sg13g2_decap_8 FILLER_24_453 ();
 sg13g2_decap_8 FILLER_24_460 ();
 sg13g2_decap_8 FILLER_24_467 ();
 sg13g2_decap_8 FILLER_24_474 ();
 sg13g2_decap_8 FILLER_24_481 ();
 sg13g2_decap_8 FILLER_24_488 ();
 sg13g2_decap_8 FILLER_24_495 ();
 sg13g2_decap_8 FILLER_24_502 ();
 sg13g2_decap_8 FILLER_24_509 ();
 sg13g2_decap_8 FILLER_24_516 ();
 sg13g2_decap_8 FILLER_24_523 ();
 sg13g2_decap_8 FILLER_24_530 ();
 sg13g2_decap_8 FILLER_24_537 ();
 sg13g2_decap_8 FILLER_24_544 ();
 sg13g2_decap_8 FILLER_24_551 ();
 sg13g2_decap_8 FILLER_24_558 ();
 sg13g2_decap_8 FILLER_24_565 ();
 sg13g2_decap_8 FILLER_24_572 ();
 sg13g2_decap_8 FILLER_24_579 ();
 sg13g2_decap_8 FILLER_24_586 ();
 sg13g2_decap_8 FILLER_24_593 ();
 sg13g2_decap_8 FILLER_24_600 ();
 sg13g2_decap_8 FILLER_24_607 ();
 sg13g2_decap_8 FILLER_24_614 ();
 sg13g2_decap_8 FILLER_24_621 ();
 sg13g2_decap_8 FILLER_24_628 ();
 sg13g2_decap_8 FILLER_24_635 ();
 sg13g2_decap_8 FILLER_24_642 ();
 sg13g2_decap_8 FILLER_24_649 ();
 sg13g2_decap_8 FILLER_24_656 ();
 sg13g2_decap_8 FILLER_24_663 ();
 sg13g2_decap_8 FILLER_24_670 ();
 sg13g2_decap_8 FILLER_24_677 ();
 sg13g2_decap_8 FILLER_24_684 ();
 sg13g2_decap_8 FILLER_24_691 ();
 sg13g2_decap_8 FILLER_24_698 ();
 sg13g2_decap_8 FILLER_24_705 ();
 sg13g2_decap_8 FILLER_24_712 ();
 sg13g2_decap_8 FILLER_24_719 ();
 sg13g2_decap_8 FILLER_24_726 ();
 sg13g2_decap_8 FILLER_24_733 ();
 sg13g2_decap_8 FILLER_24_740 ();
 sg13g2_decap_8 FILLER_24_747 ();
 sg13g2_decap_8 FILLER_24_754 ();
 sg13g2_decap_8 FILLER_24_761 ();
 sg13g2_decap_8 FILLER_24_768 ();
 sg13g2_decap_8 FILLER_24_775 ();
 sg13g2_decap_8 FILLER_24_782 ();
 sg13g2_decap_8 FILLER_24_789 ();
 sg13g2_decap_8 FILLER_24_796 ();
 sg13g2_decap_8 FILLER_24_803 ();
 sg13g2_decap_8 FILLER_24_810 ();
 sg13g2_decap_8 FILLER_24_817 ();
 sg13g2_decap_8 FILLER_24_824 ();
 sg13g2_decap_8 FILLER_24_831 ();
 sg13g2_decap_8 FILLER_24_838 ();
 sg13g2_decap_8 FILLER_24_845 ();
 sg13g2_decap_8 FILLER_24_852 ();
 sg13g2_decap_8 FILLER_24_859 ();
 sg13g2_decap_8 FILLER_24_866 ();
 sg13g2_decap_8 FILLER_24_873 ();
 sg13g2_decap_8 FILLER_24_880 ();
 sg13g2_decap_8 FILLER_24_887 ();
 sg13g2_decap_8 FILLER_24_894 ();
 sg13g2_decap_8 FILLER_24_901 ();
 sg13g2_decap_8 FILLER_24_908 ();
 sg13g2_decap_8 FILLER_24_915 ();
 sg13g2_fill_2 FILLER_24_922 ();
 sg13g2_fill_1 FILLER_24_924 ();
 sg13g2_decap_8 FILLER_25_4 ();
 sg13g2_decap_8 FILLER_25_11 ();
 sg13g2_decap_8 FILLER_25_18 ();
 sg13g2_decap_8 FILLER_25_25 ();
 sg13g2_decap_8 FILLER_25_32 ();
 sg13g2_decap_8 FILLER_25_39 ();
 sg13g2_decap_8 FILLER_25_46 ();
 sg13g2_decap_8 FILLER_25_53 ();
 sg13g2_decap_8 FILLER_25_60 ();
 sg13g2_decap_8 FILLER_25_67 ();
 sg13g2_decap_8 FILLER_25_90 ();
 sg13g2_decap_8 FILLER_25_97 ();
 sg13g2_decap_8 FILLER_25_104 ();
 sg13g2_decap_8 FILLER_25_111 ();
 sg13g2_decap_8 FILLER_25_118 ();
 sg13g2_decap_8 FILLER_25_125 ();
 sg13g2_decap_8 FILLER_25_132 ();
 sg13g2_decap_8 FILLER_25_139 ();
 sg13g2_decap_8 FILLER_25_146 ();
 sg13g2_decap_8 FILLER_25_153 ();
 sg13g2_decap_8 FILLER_25_160 ();
 sg13g2_decap_8 FILLER_25_167 ();
 sg13g2_decap_8 FILLER_25_174 ();
 sg13g2_decap_8 FILLER_25_181 ();
 sg13g2_decap_8 FILLER_25_188 ();
 sg13g2_decap_8 FILLER_25_195 ();
 sg13g2_decap_8 FILLER_25_202 ();
 sg13g2_decap_8 FILLER_25_209 ();
 sg13g2_decap_8 FILLER_25_216 ();
 sg13g2_decap_8 FILLER_25_223 ();
 sg13g2_decap_8 FILLER_25_230 ();
 sg13g2_decap_8 FILLER_25_237 ();
 sg13g2_decap_8 FILLER_25_244 ();
 sg13g2_decap_8 FILLER_25_251 ();
 sg13g2_decap_8 FILLER_25_258 ();
 sg13g2_decap_8 FILLER_25_265 ();
 sg13g2_decap_8 FILLER_25_272 ();
 sg13g2_decap_8 FILLER_25_279 ();
 sg13g2_decap_8 FILLER_25_286 ();
 sg13g2_decap_8 FILLER_25_293 ();
 sg13g2_decap_8 FILLER_25_300 ();
 sg13g2_decap_8 FILLER_25_307 ();
 sg13g2_decap_8 FILLER_25_314 ();
 sg13g2_decap_8 FILLER_25_321 ();
 sg13g2_decap_8 FILLER_25_328 ();
 sg13g2_decap_8 FILLER_25_335 ();
 sg13g2_decap_8 FILLER_25_342 ();
 sg13g2_decap_8 FILLER_25_349 ();
 sg13g2_decap_8 FILLER_25_356 ();
 sg13g2_decap_8 FILLER_25_363 ();
 sg13g2_decap_8 FILLER_25_370 ();
 sg13g2_decap_8 FILLER_25_377 ();
 sg13g2_decap_8 FILLER_25_384 ();
 sg13g2_decap_8 FILLER_25_391 ();
 sg13g2_decap_8 FILLER_25_398 ();
 sg13g2_decap_8 FILLER_25_405 ();
 sg13g2_decap_8 FILLER_25_412 ();
 sg13g2_decap_8 FILLER_25_419 ();
 sg13g2_decap_8 FILLER_25_426 ();
 sg13g2_decap_8 FILLER_25_433 ();
 sg13g2_decap_8 FILLER_25_440 ();
 sg13g2_decap_8 FILLER_25_447 ();
 sg13g2_decap_8 FILLER_25_454 ();
 sg13g2_decap_8 FILLER_25_461 ();
 sg13g2_decap_8 FILLER_25_468 ();
 sg13g2_decap_8 FILLER_25_475 ();
 sg13g2_decap_8 FILLER_25_482 ();
 sg13g2_decap_8 FILLER_25_489 ();
 sg13g2_decap_8 FILLER_25_496 ();
 sg13g2_decap_8 FILLER_25_503 ();
 sg13g2_decap_8 FILLER_25_510 ();
 sg13g2_decap_8 FILLER_25_517 ();
 sg13g2_decap_8 FILLER_25_524 ();
 sg13g2_decap_8 FILLER_25_531 ();
 sg13g2_decap_8 FILLER_25_538 ();
 sg13g2_decap_8 FILLER_25_545 ();
 sg13g2_decap_8 FILLER_25_552 ();
 sg13g2_decap_8 FILLER_25_559 ();
 sg13g2_decap_8 FILLER_25_566 ();
 sg13g2_decap_8 FILLER_25_573 ();
 sg13g2_decap_8 FILLER_25_580 ();
 sg13g2_decap_8 FILLER_25_587 ();
 sg13g2_decap_8 FILLER_25_594 ();
 sg13g2_decap_8 FILLER_25_601 ();
 sg13g2_decap_8 FILLER_25_608 ();
 sg13g2_decap_8 FILLER_25_615 ();
 sg13g2_decap_8 FILLER_25_622 ();
 sg13g2_decap_8 FILLER_25_629 ();
 sg13g2_decap_8 FILLER_25_636 ();
 sg13g2_decap_8 FILLER_25_643 ();
 sg13g2_decap_8 FILLER_25_650 ();
 sg13g2_decap_8 FILLER_25_657 ();
 sg13g2_decap_8 FILLER_25_664 ();
 sg13g2_decap_8 FILLER_25_671 ();
 sg13g2_decap_8 FILLER_25_678 ();
 sg13g2_decap_8 FILLER_25_685 ();
 sg13g2_decap_8 FILLER_25_692 ();
 sg13g2_decap_8 FILLER_25_699 ();
 sg13g2_decap_8 FILLER_25_706 ();
 sg13g2_decap_8 FILLER_25_713 ();
 sg13g2_decap_8 FILLER_25_720 ();
 sg13g2_decap_8 FILLER_25_727 ();
 sg13g2_decap_8 FILLER_25_734 ();
 sg13g2_decap_8 FILLER_25_741 ();
 sg13g2_decap_8 FILLER_25_748 ();
 sg13g2_decap_8 FILLER_25_755 ();
 sg13g2_decap_8 FILLER_25_762 ();
 sg13g2_decap_8 FILLER_25_769 ();
 sg13g2_decap_8 FILLER_25_776 ();
 sg13g2_decap_8 FILLER_25_783 ();
 sg13g2_decap_8 FILLER_25_790 ();
 sg13g2_decap_8 FILLER_25_797 ();
 sg13g2_decap_8 FILLER_25_804 ();
 sg13g2_decap_8 FILLER_25_811 ();
 sg13g2_decap_8 FILLER_25_818 ();
 sg13g2_decap_8 FILLER_25_825 ();
 sg13g2_decap_8 FILLER_25_832 ();
 sg13g2_decap_8 FILLER_25_839 ();
 sg13g2_decap_8 FILLER_25_846 ();
 sg13g2_decap_8 FILLER_25_853 ();
 sg13g2_decap_8 FILLER_25_860 ();
 sg13g2_decap_8 FILLER_25_867 ();
 sg13g2_decap_8 FILLER_25_874 ();
 sg13g2_decap_8 FILLER_25_881 ();
 sg13g2_decap_8 FILLER_25_888 ();
 sg13g2_decap_8 FILLER_25_895 ();
 sg13g2_decap_8 FILLER_25_902 ();
 sg13g2_decap_8 FILLER_25_909 ();
 sg13g2_decap_8 FILLER_25_916 ();
 sg13g2_fill_2 FILLER_25_923 ();
 sg13g2_decap_8 FILLER_26_4 ();
 sg13g2_decap_8 FILLER_26_11 ();
 sg13g2_decap_8 FILLER_26_18 ();
 sg13g2_fill_2 FILLER_26_25 ();
 sg13g2_decap_8 FILLER_26_40 ();
 sg13g2_decap_8 FILLER_26_47 ();
 sg13g2_decap_8 FILLER_26_54 ();
 sg13g2_decap_8 FILLER_26_61 ();
 sg13g2_decap_8 FILLER_26_68 ();
 sg13g2_decap_4 FILLER_26_75 ();
 sg13g2_fill_1 FILLER_26_79 ();
 sg13g2_decap_8 FILLER_26_88 ();
 sg13g2_decap_8 FILLER_26_95 ();
 sg13g2_decap_8 FILLER_26_102 ();
 sg13g2_decap_8 FILLER_26_109 ();
 sg13g2_decap_8 FILLER_26_116 ();
 sg13g2_decap_8 FILLER_26_123 ();
 sg13g2_decap_8 FILLER_26_130 ();
 sg13g2_decap_8 FILLER_26_137 ();
 sg13g2_decap_8 FILLER_26_144 ();
 sg13g2_decap_8 FILLER_26_151 ();
 sg13g2_decap_8 FILLER_26_158 ();
 sg13g2_decap_8 FILLER_26_165 ();
 sg13g2_decap_8 FILLER_26_172 ();
 sg13g2_decap_8 FILLER_26_179 ();
 sg13g2_decap_8 FILLER_26_186 ();
 sg13g2_decap_8 FILLER_26_193 ();
 sg13g2_decap_8 FILLER_26_200 ();
 sg13g2_decap_8 FILLER_26_207 ();
 sg13g2_decap_8 FILLER_26_214 ();
 sg13g2_decap_8 FILLER_26_221 ();
 sg13g2_decap_8 FILLER_26_228 ();
 sg13g2_decap_8 FILLER_26_235 ();
 sg13g2_decap_8 FILLER_26_242 ();
 sg13g2_decap_8 FILLER_26_249 ();
 sg13g2_decap_8 FILLER_26_256 ();
 sg13g2_decap_8 FILLER_26_263 ();
 sg13g2_decap_8 FILLER_26_270 ();
 sg13g2_decap_8 FILLER_26_277 ();
 sg13g2_decap_8 FILLER_26_284 ();
 sg13g2_decap_8 FILLER_26_291 ();
 sg13g2_decap_8 FILLER_26_298 ();
 sg13g2_decap_8 FILLER_26_305 ();
 sg13g2_decap_8 FILLER_26_312 ();
 sg13g2_decap_8 FILLER_26_319 ();
 sg13g2_decap_8 FILLER_26_326 ();
 sg13g2_decap_8 FILLER_26_333 ();
 sg13g2_decap_8 FILLER_26_340 ();
 sg13g2_decap_8 FILLER_26_347 ();
 sg13g2_decap_8 FILLER_26_354 ();
 sg13g2_decap_8 FILLER_26_361 ();
 sg13g2_decap_8 FILLER_26_368 ();
 sg13g2_decap_8 FILLER_26_375 ();
 sg13g2_decap_8 FILLER_26_382 ();
 sg13g2_decap_8 FILLER_26_389 ();
 sg13g2_decap_8 FILLER_26_396 ();
 sg13g2_decap_8 FILLER_26_403 ();
 sg13g2_decap_8 FILLER_26_410 ();
 sg13g2_decap_8 FILLER_26_417 ();
 sg13g2_decap_8 FILLER_26_424 ();
 sg13g2_decap_8 FILLER_26_431 ();
 sg13g2_decap_8 FILLER_26_438 ();
 sg13g2_decap_8 FILLER_26_445 ();
 sg13g2_decap_8 FILLER_26_452 ();
 sg13g2_decap_8 FILLER_26_459 ();
 sg13g2_decap_8 FILLER_26_466 ();
 sg13g2_decap_8 FILLER_26_473 ();
 sg13g2_decap_8 FILLER_26_480 ();
 sg13g2_decap_8 FILLER_26_487 ();
 sg13g2_decap_8 FILLER_26_494 ();
 sg13g2_decap_8 FILLER_26_501 ();
 sg13g2_decap_8 FILLER_26_508 ();
 sg13g2_decap_8 FILLER_26_515 ();
 sg13g2_decap_8 FILLER_26_522 ();
 sg13g2_decap_8 FILLER_26_529 ();
 sg13g2_decap_8 FILLER_26_536 ();
 sg13g2_decap_8 FILLER_26_543 ();
 sg13g2_decap_8 FILLER_26_550 ();
 sg13g2_decap_8 FILLER_26_557 ();
 sg13g2_decap_8 FILLER_26_564 ();
 sg13g2_decap_8 FILLER_26_571 ();
 sg13g2_decap_8 FILLER_26_578 ();
 sg13g2_decap_8 FILLER_26_585 ();
 sg13g2_decap_8 FILLER_26_592 ();
 sg13g2_decap_8 FILLER_26_599 ();
 sg13g2_decap_8 FILLER_26_606 ();
 sg13g2_decap_8 FILLER_26_613 ();
 sg13g2_decap_8 FILLER_26_620 ();
 sg13g2_decap_8 FILLER_26_627 ();
 sg13g2_decap_8 FILLER_26_634 ();
 sg13g2_decap_8 FILLER_26_641 ();
 sg13g2_decap_8 FILLER_26_648 ();
 sg13g2_decap_8 FILLER_26_655 ();
 sg13g2_decap_8 FILLER_26_662 ();
 sg13g2_decap_8 FILLER_26_669 ();
 sg13g2_decap_8 FILLER_26_676 ();
 sg13g2_decap_8 FILLER_26_683 ();
 sg13g2_decap_8 FILLER_26_690 ();
 sg13g2_decap_8 FILLER_26_697 ();
 sg13g2_decap_8 FILLER_26_704 ();
 sg13g2_decap_8 FILLER_26_711 ();
 sg13g2_decap_8 FILLER_26_718 ();
 sg13g2_decap_8 FILLER_26_725 ();
 sg13g2_decap_8 FILLER_26_732 ();
 sg13g2_decap_8 FILLER_26_739 ();
 sg13g2_decap_8 FILLER_26_746 ();
 sg13g2_decap_8 FILLER_26_753 ();
 sg13g2_decap_8 FILLER_26_760 ();
 sg13g2_decap_8 FILLER_26_767 ();
 sg13g2_decap_8 FILLER_26_774 ();
 sg13g2_decap_8 FILLER_26_781 ();
 sg13g2_decap_8 FILLER_26_788 ();
 sg13g2_decap_8 FILLER_26_795 ();
 sg13g2_decap_8 FILLER_26_802 ();
 sg13g2_decap_8 FILLER_26_809 ();
 sg13g2_decap_8 FILLER_26_816 ();
 sg13g2_decap_8 FILLER_26_823 ();
 sg13g2_decap_8 FILLER_26_830 ();
 sg13g2_decap_8 FILLER_26_837 ();
 sg13g2_decap_8 FILLER_26_844 ();
 sg13g2_decap_8 FILLER_26_851 ();
 sg13g2_decap_8 FILLER_26_858 ();
 sg13g2_decap_8 FILLER_26_865 ();
 sg13g2_decap_8 FILLER_26_872 ();
 sg13g2_decap_8 FILLER_26_879 ();
 sg13g2_decap_8 FILLER_26_886 ();
 sg13g2_decap_8 FILLER_26_893 ();
 sg13g2_decap_8 FILLER_26_900 ();
 sg13g2_decap_8 FILLER_26_907 ();
 sg13g2_decap_8 FILLER_26_914 ();
 sg13g2_decap_4 FILLER_26_921 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_8 FILLER_27_28 ();
 sg13g2_decap_8 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_42 ();
 sg13g2_decap_8 FILLER_27_49 ();
 sg13g2_decap_8 FILLER_27_56 ();
 sg13g2_decap_8 FILLER_27_63 ();
 sg13g2_decap_8 FILLER_27_70 ();
 sg13g2_decap_8 FILLER_27_77 ();
 sg13g2_decap_8 FILLER_27_84 ();
 sg13g2_decap_8 FILLER_27_91 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_decap_8 FILLER_27_126 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_decap_8 FILLER_27_168 ();
 sg13g2_decap_8 FILLER_27_175 ();
 sg13g2_decap_8 FILLER_27_182 ();
 sg13g2_decap_8 FILLER_27_189 ();
 sg13g2_decap_8 FILLER_27_196 ();
 sg13g2_decap_8 FILLER_27_203 ();
 sg13g2_decap_8 FILLER_27_210 ();
 sg13g2_decap_8 FILLER_27_217 ();
 sg13g2_decap_8 FILLER_27_224 ();
 sg13g2_decap_8 FILLER_27_231 ();
 sg13g2_decap_8 FILLER_27_238 ();
 sg13g2_decap_8 FILLER_27_245 ();
 sg13g2_decap_8 FILLER_27_252 ();
 sg13g2_decap_8 FILLER_27_259 ();
 sg13g2_decap_8 FILLER_27_266 ();
 sg13g2_decap_8 FILLER_27_273 ();
 sg13g2_decap_8 FILLER_27_280 ();
 sg13g2_decap_8 FILLER_27_287 ();
 sg13g2_decap_8 FILLER_27_294 ();
 sg13g2_decap_8 FILLER_27_301 ();
 sg13g2_decap_8 FILLER_27_308 ();
 sg13g2_decap_8 FILLER_27_315 ();
 sg13g2_decap_8 FILLER_27_322 ();
 sg13g2_decap_8 FILLER_27_329 ();
 sg13g2_decap_8 FILLER_27_336 ();
 sg13g2_decap_8 FILLER_27_343 ();
 sg13g2_decap_8 FILLER_27_350 ();
 sg13g2_decap_8 FILLER_27_357 ();
 sg13g2_decap_8 FILLER_27_364 ();
 sg13g2_decap_8 FILLER_27_371 ();
 sg13g2_decap_8 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_385 ();
 sg13g2_decap_8 FILLER_27_392 ();
 sg13g2_decap_8 FILLER_27_399 ();
 sg13g2_decap_8 FILLER_27_406 ();
 sg13g2_decap_8 FILLER_27_413 ();
 sg13g2_decap_8 FILLER_27_420 ();
 sg13g2_decap_8 FILLER_27_427 ();
 sg13g2_decap_8 FILLER_27_434 ();
 sg13g2_decap_8 FILLER_27_441 ();
 sg13g2_decap_8 FILLER_27_448 ();
 sg13g2_decap_8 FILLER_27_455 ();
 sg13g2_decap_8 FILLER_27_462 ();
 sg13g2_decap_8 FILLER_27_469 ();
 sg13g2_decap_8 FILLER_27_476 ();
 sg13g2_decap_8 FILLER_27_483 ();
 sg13g2_decap_8 FILLER_27_490 ();
 sg13g2_decap_8 FILLER_27_497 ();
 sg13g2_decap_8 FILLER_27_504 ();
 sg13g2_decap_8 FILLER_27_511 ();
 sg13g2_decap_8 FILLER_27_518 ();
 sg13g2_decap_8 FILLER_27_525 ();
 sg13g2_decap_8 FILLER_27_532 ();
 sg13g2_decap_8 FILLER_27_539 ();
 sg13g2_decap_8 FILLER_27_546 ();
 sg13g2_decap_8 FILLER_27_553 ();
 sg13g2_decap_8 FILLER_27_560 ();
 sg13g2_decap_8 FILLER_27_567 ();
 sg13g2_decap_8 FILLER_27_574 ();
 sg13g2_decap_8 FILLER_27_581 ();
 sg13g2_decap_8 FILLER_27_588 ();
 sg13g2_decap_8 FILLER_27_595 ();
 sg13g2_decap_8 FILLER_27_602 ();
 sg13g2_decap_8 FILLER_27_609 ();
 sg13g2_decap_8 FILLER_27_616 ();
 sg13g2_decap_8 FILLER_27_623 ();
 sg13g2_decap_8 FILLER_27_630 ();
 sg13g2_decap_8 FILLER_27_637 ();
 sg13g2_decap_8 FILLER_27_644 ();
 sg13g2_decap_8 FILLER_27_651 ();
 sg13g2_decap_8 FILLER_27_658 ();
 sg13g2_decap_8 FILLER_27_665 ();
 sg13g2_decap_8 FILLER_27_672 ();
 sg13g2_decap_8 FILLER_27_679 ();
 sg13g2_decap_8 FILLER_27_686 ();
 sg13g2_decap_8 FILLER_27_693 ();
 sg13g2_decap_8 FILLER_27_700 ();
 sg13g2_decap_8 FILLER_27_707 ();
 sg13g2_decap_8 FILLER_27_714 ();
 sg13g2_decap_8 FILLER_27_721 ();
 sg13g2_decap_8 FILLER_27_728 ();
 sg13g2_decap_8 FILLER_27_735 ();
 sg13g2_decap_8 FILLER_27_742 ();
 sg13g2_decap_8 FILLER_27_749 ();
 sg13g2_decap_8 FILLER_27_756 ();
 sg13g2_decap_8 FILLER_27_763 ();
 sg13g2_decap_8 FILLER_27_770 ();
 sg13g2_decap_8 FILLER_27_777 ();
 sg13g2_decap_8 FILLER_27_784 ();
 sg13g2_decap_8 FILLER_27_791 ();
 sg13g2_decap_8 FILLER_27_798 ();
 sg13g2_decap_8 FILLER_27_805 ();
 sg13g2_decap_8 FILLER_27_812 ();
 sg13g2_decap_8 FILLER_27_819 ();
 sg13g2_decap_8 FILLER_27_826 ();
 sg13g2_decap_8 FILLER_27_833 ();
 sg13g2_decap_8 FILLER_27_840 ();
 sg13g2_decap_8 FILLER_27_847 ();
 sg13g2_decap_8 FILLER_27_854 ();
 sg13g2_decap_8 FILLER_27_861 ();
 sg13g2_decap_8 FILLER_27_868 ();
 sg13g2_decap_8 FILLER_27_875 ();
 sg13g2_decap_8 FILLER_27_882 ();
 sg13g2_decap_8 FILLER_27_889 ();
 sg13g2_decap_8 FILLER_27_896 ();
 sg13g2_decap_8 FILLER_27_903 ();
 sg13g2_decap_8 FILLER_27_910 ();
 sg13g2_decap_8 FILLER_27_917 ();
 sg13g2_fill_1 FILLER_27_924 ();
 sg13g2_decap_8 FILLER_28_4 ();
 sg13g2_decap_8 FILLER_28_11 ();
 sg13g2_decap_8 FILLER_28_18 ();
 sg13g2_decap_8 FILLER_28_25 ();
 sg13g2_decap_8 FILLER_28_32 ();
 sg13g2_decap_8 FILLER_28_39 ();
 sg13g2_decap_8 FILLER_28_46 ();
 sg13g2_decap_8 FILLER_28_53 ();
 sg13g2_decap_8 FILLER_28_60 ();
 sg13g2_decap_8 FILLER_28_67 ();
 sg13g2_decap_8 FILLER_28_74 ();
 sg13g2_decap_8 FILLER_28_81 ();
 sg13g2_decap_8 FILLER_28_88 ();
 sg13g2_decap_8 FILLER_28_95 ();
 sg13g2_decap_4 FILLER_28_102 ();
 sg13g2_fill_2 FILLER_28_106 ();
 sg13g2_fill_1 FILLER_28_116 ();
 sg13g2_decap_8 FILLER_28_125 ();
 sg13g2_decap_8 FILLER_28_132 ();
 sg13g2_decap_8 FILLER_28_139 ();
 sg13g2_decap_8 FILLER_28_146 ();
 sg13g2_decap_8 FILLER_28_153 ();
 sg13g2_decap_8 FILLER_28_160 ();
 sg13g2_decap_8 FILLER_28_167 ();
 sg13g2_decap_8 FILLER_28_174 ();
 sg13g2_decap_8 FILLER_28_181 ();
 sg13g2_decap_8 FILLER_28_188 ();
 sg13g2_decap_8 FILLER_28_195 ();
 sg13g2_decap_8 FILLER_28_202 ();
 sg13g2_decap_8 FILLER_28_209 ();
 sg13g2_decap_8 FILLER_28_216 ();
 sg13g2_decap_8 FILLER_28_223 ();
 sg13g2_decap_8 FILLER_28_230 ();
 sg13g2_decap_8 FILLER_28_237 ();
 sg13g2_decap_8 FILLER_28_244 ();
 sg13g2_decap_8 FILLER_28_251 ();
 sg13g2_decap_8 FILLER_28_258 ();
 sg13g2_decap_8 FILLER_28_265 ();
 sg13g2_decap_8 FILLER_28_272 ();
 sg13g2_decap_8 FILLER_28_279 ();
 sg13g2_decap_8 FILLER_28_286 ();
 sg13g2_decap_8 FILLER_28_293 ();
 sg13g2_decap_8 FILLER_28_300 ();
 sg13g2_decap_8 FILLER_28_307 ();
 sg13g2_decap_8 FILLER_28_314 ();
 sg13g2_decap_8 FILLER_28_321 ();
 sg13g2_decap_8 FILLER_28_328 ();
 sg13g2_decap_8 FILLER_28_335 ();
 sg13g2_decap_8 FILLER_28_342 ();
 sg13g2_decap_8 FILLER_28_349 ();
 sg13g2_decap_8 FILLER_28_356 ();
 sg13g2_decap_8 FILLER_28_363 ();
 sg13g2_decap_8 FILLER_28_370 ();
 sg13g2_decap_8 FILLER_28_377 ();
 sg13g2_decap_8 FILLER_28_384 ();
 sg13g2_decap_8 FILLER_28_391 ();
 sg13g2_decap_8 FILLER_28_398 ();
 sg13g2_decap_8 FILLER_28_405 ();
 sg13g2_decap_8 FILLER_28_412 ();
 sg13g2_decap_8 FILLER_28_419 ();
 sg13g2_decap_8 FILLER_28_426 ();
 sg13g2_decap_8 FILLER_28_433 ();
 sg13g2_decap_8 FILLER_28_440 ();
 sg13g2_decap_8 FILLER_28_447 ();
 sg13g2_decap_8 FILLER_28_454 ();
 sg13g2_decap_8 FILLER_28_461 ();
 sg13g2_decap_8 FILLER_28_468 ();
 sg13g2_decap_8 FILLER_28_475 ();
 sg13g2_decap_8 FILLER_28_482 ();
 sg13g2_decap_8 FILLER_28_489 ();
 sg13g2_decap_8 FILLER_28_496 ();
 sg13g2_decap_8 FILLER_28_503 ();
 sg13g2_decap_8 FILLER_28_510 ();
 sg13g2_decap_8 FILLER_28_517 ();
 sg13g2_decap_8 FILLER_28_524 ();
 sg13g2_decap_8 FILLER_28_531 ();
 sg13g2_decap_8 FILLER_28_538 ();
 sg13g2_decap_8 FILLER_28_545 ();
 sg13g2_decap_8 FILLER_28_552 ();
 sg13g2_decap_8 FILLER_28_559 ();
 sg13g2_decap_8 FILLER_28_566 ();
 sg13g2_decap_8 FILLER_28_573 ();
 sg13g2_decap_8 FILLER_28_580 ();
 sg13g2_decap_8 FILLER_28_587 ();
 sg13g2_decap_8 FILLER_28_594 ();
 sg13g2_decap_8 FILLER_28_601 ();
 sg13g2_decap_8 FILLER_28_608 ();
 sg13g2_decap_8 FILLER_28_615 ();
 sg13g2_decap_8 FILLER_28_622 ();
 sg13g2_decap_8 FILLER_28_629 ();
 sg13g2_decap_8 FILLER_28_636 ();
 sg13g2_decap_8 FILLER_28_643 ();
 sg13g2_decap_8 FILLER_28_650 ();
 sg13g2_decap_8 FILLER_28_657 ();
 sg13g2_decap_8 FILLER_28_664 ();
 sg13g2_decap_8 FILLER_28_671 ();
 sg13g2_decap_8 FILLER_28_678 ();
 sg13g2_decap_8 FILLER_28_685 ();
 sg13g2_decap_8 FILLER_28_692 ();
 sg13g2_decap_8 FILLER_28_699 ();
 sg13g2_decap_8 FILLER_28_706 ();
 sg13g2_decap_8 FILLER_28_713 ();
 sg13g2_decap_8 FILLER_28_720 ();
 sg13g2_decap_8 FILLER_28_727 ();
 sg13g2_decap_8 FILLER_28_734 ();
 sg13g2_decap_8 FILLER_28_741 ();
 sg13g2_decap_8 FILLER_28_748 ();
 sg13g2_decap_8 FILLER_28_755 ();
 sg13g2_decap_8 FILLER_28_762 ();
 sg13g2_decap_8 FILLER_28_769 ();
 sg13g2_decap_8 FILLER_28_776 ();
 sg13g2_decap_8 FILLER_28_783 ();
 sg13g2_decap_8 FILLER_28_790 ();
 sg13g2_decap_8 FILLER_28_797 ();
 sg13g2_decap_8 FILLER_28_804 ();
 sg13g2_decap_8 FILLER_28_811 ();
 sg13g2_decap_8 FILLER_28_818 ();
 sg13g2_decap_8 FILLER_28_825 ();
 sg13g2_decap_8 FILLER_28_832 ();
 sg13g2_decap_8 FILLER_28_839 ();
 sg13g2_decap_8 FILLER_28_846 ();
 sg13g2_decap_8 FILLER_28_853 ();
 sg13g2_decap_8 FILLER_28_860 ();
 sg13g2_decap_8 FILLER_28_867 ();
 sg13g2_decap_8 FILLER_28_874 ();
 sg13g2_decap_8 FILLER_28_881 ();
 sg13g2_decap_8 FILLER_28_888 ();
 sg13g2_decap_8 FILLER_28_895 ();
 sg13g2_decap_8 FILLER_28_902 ();
 sg13g2_decap_8 FILLER_28_909 ();
 sg13g2_decap_8 FILLER_28_916 ();
 sg13g2_fill_2 FILLER_28_923 ();
 sg13g2_decap_8 FILLER_29_4 ();
 sg13g2_decap_8 FILLER_29_11 ();
 sg13g2_decap_8 FILLER_29_18 ();
 sg13g2_decap_8 FILLER_29_25 ();
 sg13g2_decap_8 FILLER_29_32 ();
 sg13g2_decap_8 FILLER_29_39 ();
 sg13g2_decap_8 FILLER_29_46 ();
 sg13g2_decap_8 FILLER_29_53 ();
 sg13g2_decap_8 FILLER_29_60 ();
 sg13g2_decap_8 FILLER_29_67 ();
 sg13g2_decap_8 FILLER_29_74 ();
 sg13g2_decap_8 FILLER_29_81 ();
 sg13g2_decap_8 FILLER_29_88 ();
 sg13g2_decap_8 FILLER_29_95 ();
 sg13g2_decap_8 FILLER_29_102 ();
 sg13g2_decap_8 FILLER_29_109 ();
 sg13g2_fill_2 FILLER_29_116 ();
 sg13g2_fill_1 FILLER_29_118 ();
 sg13g2_decap_8 FILLER_29_124 ();
 sg13g2_decap_8 FILLER_29_131 ();
 sg13g2_decap_8 FILLER_29_138 ();
 sg13g2_decap_8 FILLER_29_145 ();
 sg13g2_decap_8 FILLER_29_152 ();
 sg13g2_decap_8 FILLER_29_159 ();
 sg13g2_decap_8 FILLER_29_166 ();
 sg13g2_decap_8 FILLER_29_173 ();
 sg13g2_decap_8 FILLER_29_180 ();
 sg13g2_decap_8 FILLER_29_187 ();
 sg13g2_decap_8 FILLER_29_194 ();
 sg13g2_decap_8 FILLER_29_201 ();
 sg13g2_decap_8 FILLER_29_208 ();
 sg13g2_decap_8 FILLER_29_215 ();
 sg13g2_decap_8 FILLER_29_222 ();
 sg13g2_decap_8 FILLER_29_229 ();
 sg13g2_decap_8 FILLER_29_236 ();
 sg13g2_decap_8 FILLER_29_243 ();
 sg13g2_decap_8 FILLER_29_250 ();
 sg13g2_decap_8 FILLER_29_257 ();
 sg13g2_decap_8 FILLER_29_264 ();
 sg13g2_decap_8 FILLER_29_271 ();
 sg13g2_decap_8 FILLER_29_278 ();
 sg13g2_decap_8 FILLER_29_285 ();
 sg13g2_decap_8 FILLER_29_292 ();
 sg13g2_decap_8 FILLER_29_299 ();
 sg13g2_decap_8 FILLER_29_306 ();
 sg13g2_decap_8 FILLER_29_313 ();
 sg13g2_decap_8 FILLER_29_320 ();
 sg13g2_decap_8 FILLER_29_327 ();
 sg13g2_decap_8 FILLER_29_334 ();
 sg13g2_decap_8 FILLER_29_341 ();
 sg13g2_decap_8 FILLER_29_348 ();
 sg13g2_decap_8 FILLER_29_355 ();
 sg13g2_decap_8 FILLER_29_362 ();
 sg13g2_decap_8 FILLER_29_369 ();
 sg13g2_decap_8 FILLER_29_376 ();
 sg13g2_decap_8 FILLER_29_383 ();
 sg13g2_decap_8 FILLER_29_390 ();
 sg13g2_decap_8 FILLER_29_397 ();
 sg13g2_decap_8 FILLER_29_404 ();
 sg13g2_decap_8 FILLER_29_411 ();
 sg13g2_decap_8 FILLER_29_418 ();
 sg13g2_decap_8 FILLER_29_425 ();
 sg13g2_decap_8 FILLER_29_432 ();
 sg13g2_decap_8 FILLER_29_439 ();
 sg13g2_decap_8 FILLER_29_446 ();
 sg13g2_decap_8 FILLER_29_453 ();
 sg13g2_decap_8 FILLER_29_460 ();
 sg13g2_decap_8 FILLER_29_467 ();
 sg13g2_decap_8 FILLER_29_474 ();
 sg13g2_decap_8 FILLER_29_481 ();
 sg13g2_decap_8 FILLER_29_488 ();
 sg13g2_decap_8 FILLER_29_495 ();
 sg13g2_decap_8 FILLER_29_502 ();
 sg13g2_decap_8 FILLER_29_509 ();
 sg13g2_decap_8 FILLER_29_516 ();
 sg13g2_decap_8 FILLER_29_523 ();
 sg13g2_decap_8 FILLER_29_530 ();
 sg13g2_decap_8 FILLER_29_537 ();
 sg13g2_decap_8 FILLER_29_544 ();
 sg13g2_decap_8 FILLER_29_551 ();
 sg13g2_decap_8 FILLER_29_558 ();
 sg13g2_decap_8 FILLER_29_565 ();
 sg13g2_decap_8 FILLER_29_572 ();
 sg13g2_decap_8 FILLER_29_579 ();
 sg13g2_decap_8 FILLER_29_586 ();
 sg13g2_decap_8 FILLER_29_593 ();
 sg13g2_decap_8 FILLER_29_600 ();
 sg13g2_decap_8 FILLER_29_607 ();
 sg13g2_decap_8 FILLER_29_614 ();
 sg13g2_decap_8 FILLER_29_621 ();
 sg13g2_decap_8 FILLER_29_628 ();
 sg13g2_decap_8 FILLER_29_635 ();
 sg13g2_decap_8 FILLER_29_642 ();
 sg13g2_decap_8 FILLER_29_649 ();
 sg13g2_decap_8 FILLER_29_656 ();
 sg13g2_decap_8 FILLER_29_663 ();
 sg13g2_decap_8 FILLER_29_670 ();
 sg13g2_decap_8 FILLER_29_677 ();
 sg13g2_decap_8 FILLER_29_684 ();
 sg13g2_decap_8 FILLER_29_691 ();
 sg13g2_decap_8 FILLER_29_698 ();
 sg13g2_decap_8 FILLER_29_705 ();
 sg13g2_decap_8 FILLER_29_712 ();
 sg13g2_decap_8 FILLER_29_719 ();
 sg13g2_decap_8 FILLER_29_726 ();
 sg13g2_decap_8 FILLER_29_733 ();
 sg13g2_decap_8 FILLER_29_740 ();
 sg13g2_decap_8 FILLER_29_747 ();
 sg13g2_decap_8 FILLER_29_754 ();
 sg13g2_decap_8 FILLER_29_761 ();
 sg13g2_decap_8 FILLER_29_768 ();
 sg13g2_decap_8 FILLER_29_775 ();
 sg13g2_decap_8 FILLER_29_782 ();
 sg13g2_decap_8 FILLER_29_789 ();
 sg13g2_decap_8 FILLER_29_796 ();
 sg13g2_decap_8 FILLER_29_803 ();
 sg13g2_decap_8 FILLER_29_810 ();
 sg13g2_decap_8 FILLER_29_817 ();
 sg13g2_decap_8 FILLER_29_824 ();
 sg13g2_decap_8 FILLER_29_831 ();
 sg13g2_decap_8 FILLER_29_838 ();
 sg13g2_decap_8 FILLER_29_845 ();
 sg13g2_decap_8 FILLER_29_852 ();
 sg13g2_decap_8 FILLER_29_859 ();
 sg13g2_decap_8 FILLER_29_866 ();
 sg13g2_decap_8 FILLER_29_873 ();
 sg13g2_decap_8 FILLER_29_880 ();
 sg13g2_decap_8 FILLER_29_887 ();
 sg13g2_decap_8 FILLER_29_894 ();
 sg13g2_decap_8 FILLER_29_901 ();
 sg13g2_decap_8 FILLER_29_908 ();
 sg13g2_decap_8 FILLER_29_915 ();
 sg13g2_fill_2 FILLER_29_922 ();
 sg13g2_fill_1 FILLER_29_924 ();
 sg13g2_decap_8 FILLER_30_4 ();
 sg13g2_fill_1 FILLER_30_11 ();
 sg13g2_decap_8 FILLER_30_24 ();
 sg13g2_decap_4 FILLER_30_31 ();
 sg13g2_fill_1 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_40 ();
 sg13g2_decap_8 FILLER_30_47 ();
 sg13g2_decap_8 FILLER_30_54 ();
 sg13g2_decap_8 FILLER_30_61 ();
 sg13g2_decap_8 FILLER_30_68 ();
 sg13g2_decap_8 FILLER_30_75 ();
 sg13g2_decap_8 FILLER_30_82 ();
 sg13g2_decap_8 FILLER_30_89 ();
 sg13g2_decap_8 FILLER_30_96 ();
 sg13g2_decap_8 FILLER_30_103 ();
 sg13g2_decap_8 FILLER_30_114 ();
 sg13g2_decap_8 FILLER_30_121 ();
 sg13g2_decap_8 FILLER_30_128 ();
 sg13g2_decap_8 FILLER_30_135 ();
 sg13g2_decap_8 FILLER_30_142 ();
 sg13g2_decap_8 FILLER_30_149 ();
 sg13g2_decap_8 FILLER_30_156 ();
 sg13g2_decap_8 FILLER_30_163 ();
 sg13g2_decap_8 FILLER_30_170 ();
 sg13g2_decap_8 FILLER_30_177 ();
 sg13g2_decap_8 FILLER_30_184 ();
 sg13g2_decap_8 FILLER_30_191 ();
 sg13g2_decap_8 FILLER_30_198 ();
 sg13g2_decap_8 FILLER_30_205 ();
 sg13g2_decap_8 FILLER_30_212 ();
 sg13g2_decap_8 FILLER_30_219 ();
 sg13g2_decap_8 FILLER_30_226 ();
 sg13g2_decap_8 FILLER_30_233 ();
 sg13g2_decap_8 FILLER_30_240 ();
 sg13g2_decap_8 FILLER_30_247 ();
 sg13g2_decap_8 FILLER_30_254 ();
 sg13g2_decap_8 FILLER_30_261 ();
 sg13g2_decap_8 FILLER_30_268 ();
 sg13g2_decap_8 FILLER_30_275 ();
 sg13g2_decap_8 FILLER_30_282 ();
 sg13g2_decap_8 FILLER_30_289 ();
 sg13g2_decap_8 FILLER_30_296 ();
 sg13g2_decap_8 FILLER_30_303 ();
 sg13g2_decap_8 FILLER_30_310 ();
 sg13g2_decap_8 FILLER_30_317 ();
 sg13g2_decap_8 FILLER_30_324 ();
 sg13g2_decap_8 FILLER_30_331 ();
 sg13g2_decap_8 FILLER_30_338 ();
 sg13g2_decap_8 FILLER_30_345 ();
 sg13g2_decap_8 FILLER_30_352 ();
 sg13g2_decap_8 FILLER_30_359 ();
 sg13g2_decap_8 FILLER_30_366 ();
 sg13g2_decap_8 FILLER_30_373 ();
 sg13g2_decap_8 FILLER_30_380 ();
 sg13g2_decap_8 FILLER_30_387 ();
 sg13g2_decap_8 FILLER_30_394 ();
 sg13g2_decap_8 FILLER_30_401 ();
 sg13g2_decap_8 FILLER_30_408 ();
 sg13g2_decap_8 FILLER_30_415 ();
 sg13g2_decap_8 FILLER_30_422 ();
 sg13g2_decap_8 FILLER_30_429 ();
 sg13g2_decap_8 FILLER_30_436 ();
 sg13g2_decap_8 FILLER_30_443 ();
 sg13g2_decap_8 FILLER_30_450 ();
 sg13g2_decap_8 FILLER_30_457 ();
 sg13g2_decap_8 FILLER_30_464 ();
 sg13g2_decap_8 FILLER_30_471 ();
 sg13g2_decap_8 FILLER_30_478 ();
 sg13g2_decap_8 FILLER_30_485 ();
 sg13g2_decap_8 FILLER_30_492 ();
 sg13g2_decap_8 FILLER_30_499 ();
 sg13g2_decap_8 FILLER_30_506 ();
 sg13g2_decap_8 FILLER_30_513 ();
 sg13g2_decap_8 FILLER_30_520 ();
 sg13g2_decap_8 FILLER_30_527 ();
 sg13g2_decap_8 FILLER_30_534 ();
 sg13g2_decap_8 FILLER_30_541 ();
 sg13g2_decap_8 FILLER_30_548 ();
 sg13g2_decap_8 FILLER_30_555 ();
 sg13g2_decap_8 FILLER_30_562 ();
 sg13g2_decap_8 FILLER_30_569 ();
 sg13g2_decap_8 FILLER_30_576 ();
 sg13g2_decap_8 FILLER_30_583 ();
 sg13g2_decap_8 FILLER_30_590 ();
 sg13g2_decap_8 FILLER_30_597 ();
 sg13g2_decap_8 FILLER_30_604 ();
 sg13g2_decap_8 FILLER_30_611 ();
 sg13g2_decap_8 FILLER_30_618 ();
 sg13g2_decap_8 FILLER_30_625 ();
 sg13g2_decap_8 FILLER_30_632 ();
 sg13g2_decap_8 FILLER_30_639 ();
 sg13g2_decap_8 FILLER_30_646 ();
 sg13g2_decap_8 FILLER_30_653 ();
 sg13g2_decap_8 FILLER_30_660 ();
 sg13g2_decap_8 FILLER_30_667 ();
 sg13g2_decap_8 FILLER_30_674 ();
 sg13g2_decap_8 FILLER_30_681 ();
 sg13g2_decap_8 FILLER_30_688 ();
 sg13g2_decap_8 FILLER_30_695 ();
 sg13g2_decap_8 FILLER_30_702 ();
 sg13g2_decap_8 FILLER_30_709 ();
 sg13g2_decap_8 FILLER_30_716 ();
 sg13g2_decap_8 FILLER_30_723 ();
 sg13g2_decap_8 FILLER_30_730 ();
 sg13g2_decap_8 FILLER_30_737 ();
 sg13g2_decap_8 FILLER_30_744 ();
 sg13g2_decap_8 FILLER_30_751 ();
 sg13g2_decap_8 FILLER_30_758 ();
 sg13g2_decap_8 FILLER_30_765 ();
 sg13g2_decap_8 FILLER_30_772 ();
 sg13g2_decap_8 FILLER_30_779 ();
 sg13g2_decap_8 FILLER_30_786 ();
 sg13g2_decap_8 FILLER_30_793 ();
 sg13g2_decap_8 FILLER_30_800 ();
 sg13g2_decap_8 FILLER_30_807 ();
 sg13g2_decap_8 FILLER_30_814 ();
 sg13g2_decap_8 FILLER_30_821 ();
 sg13g2_decap_8 FILLER_30_828 ();
 sg13g2_decap_8 FILLER_30_835 ();
 sg13g2_decap_8 FILLER_30_842 ();
 sg13g2_decap_8 FILLER_30_849 ();
 sg13g2_decap_8 FILLER_30_856 ();
 sg13g2_decap_8 FILLER_30_863 ();
 sg13g2_decap_8 FILLER_30_870 ();
 sg13g2_decap_8 FILLER_30_877 ();
 sg13g2_decap_8 FILLER_30_884 ();
 sg13g2_decap_8 FILLER_30_891 ();
 sg13g2_decap_8 FILLER_30_898 ();
 sg13g2_decap_8 FILLER_30_905 ();
 sg13g2_decap_8 FILLER_30_912 ();
 sg13g2_decap_4 FILLER_30_919 ();
 sg13g2_fill_2 FILLER_30_923 ();
 sg13g2_decap_8 FILLER_31_4 ();
 sg13g2_decap_8 FILLER_31_11 ();
 sg13g2_decap_8 FILLER_31_18 ();
 sg13g2_decap_8 FILLER_31_25 ();
 sg13g2_decap_4 FILLER_31_32 ();
 sg13g2_fill_2 FILLER_31_40 ();
 sg13g2_fill_2 FILLER_31_45 ();
 sg13g2_fill_1 FILLER_31_47 ();
 sg13g2_fill_2 FILLER_31_56 ();
 sg13g2_fill_1 FILLER_31_58 ();
 sg13g2_decap_8 FILLER_31_67 ();
 sg13g2_decap_8 FILLER_31_74 ();
 sg13g2_decap_8 FILLER_31_81 ();
 sg13g2_decap_8 FILLER_31_88 ();
 sg13g2_decap_4 FILLER_31_100 ();
 sg13g2_fill_2 FILLER_31_104 ();
 sg13g2_decap_8 FILLER_31_111 ();
 sg13g2_decap_8 FILLER_31_122 ();
 sg13g2_decap_8 FILLER_31_129 ();
 sg13g2_decap_8 FILLER_31_136 ();
 sg13g2_decap_8 FILLER_31_143 ();
 sg13g2_decap_8 FILLER_31_150 ();
 sg13g2_decap_8 FILLER_31_157 ();
 sg13g2_decap_8 FILLER_31_164 ();
 sg13g2_decap_8 FILLER_31_171 ();
 sg13g2_decap_8 FILLER_31_178 ();
 sg13g2_decap_8 FILLER_31_185 ();
 sg13g2_decap_8 FILLER_31_192 ();
 sg13g2_decap_8 FILLER_31_199 ();
 sg13g2_decap_8 FILLER_31_206 ();
 sg13g2_decap_8 FILLER_31_213 ();
 sg13g2_decap_8 FILLER_31_220 ();
 sg13g2_decap_8 FILLER_31_227 ();
 sg13g2_decap_8 FILLER_31_234 ();
 sg13g2_decap_8 FILLER_31_241 ();
 sg13g2_decap_8 FILLER_31_248 ();
 sg13g2_decap_8 FILLER_31_255 ();
 sg13g2_decap_8 FILLER_31_262 ();
 sg13g2_decap_8 FILLER_31_269 ();
 sg13g2_decap_8 FILLER_31_276 ();
 sg13g2_decap_8 FILLER_31_283 ();
 sg13g2_decap_8 FILLER_31_290 ();
 sg13g2_decap_8 FILLER_31_297 ();
 sg13g2_decap_8 FILLER_31_304 ();
 sg13g2_decap_8 FILLER_31_311 ();
 sg13g2_decap_8 FILLER_31_318 ();
 sg13g2_decap_8 FILLER_31_325 ();
 sg13g2_decap_8 FILLER_31_332 ();
 sg13g2_decap_8 FILLER_31_339 ();
 sg13g2_decap_8 FILLER_31_346 ();
 sg13g2_decap_8 FILLER_31_353 ();
 sg13g2_decap_8 FILLER_31_360 ();
 sg13g2_decap_8 FILLER_31_367 ();
 sg13g2_decap_8 FILLER_31_374 ();
 sg13g2_decap_8 FILLER_31_381 ();
 sg13g2_decap_8 FILLER_31_388 ();
 sg13g2_decap_8 FILLER_31_395 ();
 sg13g2_decap_8 FILLER_31_402 ();
 sg13g2_decap_8 FILLER_31_409 ();
 sg13g2_decap_8 FILLER_31_416 ();
 sg13g2_decap_8 FILLER_31_423 ();
 sg13g2_decap_8 FILLER_31_430 ();
 sg13g2_decap_8 FILLER_31_437 ();
 sg13g2_decap_8 FILLER_31_444 ();
 sg13g2_decap_8 FILLER_31_451 ();
 sg13g2_decap_8 FILLER_31_458 ();
 sg13g2_decap_8 FILLER_31_465 ();
 sg13g2_decap_8 FILLER_31_472 ();
 sg13g2_decap_8 FILLER_31_479 ();
 sg13g2_decap_8 FILLER_31_486 ();
 sg13g2_decap_8 FILLER_31_493 ();
 sg13g2_decap_8 FILLER_31_500 ();
 sg13g2_decap_8 FILLER_31_507 ();
 sg13g2_decap_8 FILLER_31_514 ();
 sg13g2_decap_8 FILLER_31_521 ();
 sg13g2_decap_8 FILLER_31_528 ();
 sg13g2_decap_8 FILLER_31_535 ();
 sg13g2_decap_8 FILLER_31_542 ();
 sg13g2_decap_8 FILLER_31_549 ();
 sg13g2_decap_8 FILLER_31_556 ();
 sg13g2_decap_8 FILLER_31_563 ();
 sg13g2_decap_8 FILLER_31_570 ();
 sg13g2_decap_8 FILLER_31_577 ();
 sg13g2_decap_8 FILLER_31_584 ();
 sg13g2_decap_8 FILLER_31_591 ();
 sg13g2_decap_8 FILLER_31_598 ();
 sg13g2_decap_8 FILLER_31_605 ();
 sg13g2_decap_8 FILLER_31_612 ();
 sg13g2_decap_8 FILLER_31_619 ();
 sg13g2_decap_8 FILLER_31_626 ();
 sg13g2_decap_8 FILLER_31_633 ();
 sg13g2_decap_8 FILLER_31_640 ();
 sg13g2_decap_8 FILLER_31_647 ();
 sg13g2_decap_8 FILLER_31_654 ();
 sg13g2_decap_8 FILLER_31_661 ();
 sg13g2_decap_8 FILLER_31_668 ();
 sg13g2_decap_8 FILLER_31_675 ();
 sg13g2_decap_8 FILLER_31_682 ();
 sg13g2_decap_8 FILLER_31_689 ();
 sg13g2_decap_8 FILLER_31_696 ();
 sg13g2_decap_8 FILLER_31_703 ();
 sg13g2_decap_8 FILLER_31_710 ();
 sg13g2_decap_8 FILLER_31_717 ();
 sg13g2_decap_8 FILLER_31_724 ();
 sg13g2_decap_8 FILLER_31_731 ();
 sg13g2_decap_8 FILLER_31_738 ();
 sg13g2_decap_8 FILLER_31_745 ();
 sg13g2_decap_8 FILLER_31_752 ();
 sg13g2_decap_8 FILLER_31_759 ();
 sg13g2_decap_8 FILLER_31_766 ();
 sg13g2_decap_8 FILLER_31_773 ();
 sg13g2_decap_8 FILLER_31_780 ();
 sg13g2_decap_8 FILLER_31_787 ();
 sg13g2_decap_8 FILLER_31_794 ();
 sg13g2_decap_8 FILLER_31_801 ();
 sg13g2_decap_8 FILLER_31_808 ();
 sg13g2_decap_8 FILLER_31_815 ();
 sg13g2_decap_8 FILLER_31_822 ();
 sg13g2_decap_8 FILLER_31_829 ();
 sg13g2_decap_8 FILLER_31_836 ();
 sg13g2_decap_8 FILLER_31_843 ();
 sg13g2_decap_8 FILLER_31_850 ();
 sg13g2_decap_8 FILLER_31_857 ();
 sg13g2_decap_8 FILLER_31_864 ();
 sg13g2_decap_8 FILLER_31_871 ();
 sg13g2_decap_8 FILLER_31_878 ();
 sg13g2_decap_8 FILLER_31_885 ();
 sg13g2_decap_8 FILLER_31_892 ();
 sg13g2_decap_8 FILLER_31_899 ();
 sg13g2_decap_8 FILLER_31_906 ();
 sg13g2_decap_8 FILLER_31_913 ();
 sg13g2_decap_4 FILLER_31_920 ();
 sg13g2_fill_1 FILLER_31_924 ();
 sg13g2_decap_8 FILLER_32_4 ();
 sg13g2_decap_8 FILLER_32_11 ();
 sg13g2_decap_8 FILLER_32_18 ();
 sg13g2_decap_8 FILLER_32_25 ();
 sg13g2_decap_8 FILLER_32_32 ();
 sg13g2_decap_8 FILLER_32_39 ();
 sg13g2_decap_8 FILLER_32_46 ();
 sg13g2_decap_8 FILLER_32_53 ();
 sg13g2_decap_8 FILLER_32_60 ();
 sg13g2_decap_8 FILLER_32_67 ();
 sg13g2_decap_8 FILLER_32_74 ();
 sg13g2_decap_8 FILLER_32_81 ();
 sg13g2_decap_8 FILLER_32_88 ();
 sg13g2_decap_8 FILLER_32_95 ();
 sg13g2_decap_8 FILLER_32_102 ();
 sg13g2_decap_8 FILLER_32_109 ();
 sg13g2_decap_4 FILLER_32_116 ();
 sg13g2_fill_2 FILLER_32_120 ();
 sg13g2_decap_8 FILLER_32_130 ();
 sg13g2_decap_8 FILLER_32_137 ();
 sg13g2_decap_8 FILLER_32_144 ();
 sg13g2_decap_8 FILLER_32_151 ();
 sg13g2_decap_8 FILLER_32_158 ();
 sg13g2_decap_8 FILLER_32_165 ();
 sg13g2_decap_8 FILLER_32_172 ();
 sg13g2_decap_8 FILLER_32_179 ();
 sg13g2_decap_8 FILLER_32_186 ();
 sg13g2_decap_8 FILLER_32_193 ();
 sg13g2_decap_8 FILLER_32_200 ();
 sg13g2_decap_8 FILLER_32_207 ();
 sg13g2_decap_8 FILLER_32_214 ();
 sg13g2_decap_8 FILLER_32_221 ();
 sg13g2_decap_8 FILLER_32_228 ();
 sg13g2_decap_8 FILLER_32_235 ();
 sg13g2_decap_8 FILLER_32_242 ();
 sg13g2_decap_8 FILLER_32_249 ();
 sg13g2_decap_8 FILLER_32_256 ();
 sg13g2_decap_8 FILLER_32_263 ();
 sg13g2_decap_8 FILLER_32_270 ();
 sg13g2_decap_8 FILLER_32_277 ();
 sg13g2_decap_8 FILLER_32_284 ();
 sg13g2_decap_8 FILLER_32_291 ();
 sg13g2_decap_8 FILLER_32_298 ();
 sg13g2_decap_8 FILLER_32_305 ();
 sg13g2_decap_8 FILLER_32_312 ();
 sg13g2_decap_8 FILLER_32_319 ();
 sg13g2_decap_8 FILLER_32_326 ();
 sg13g2_decap_8 FILLER_32_333 ();
 sg13g2_decap_8 FILLER_32_340 ();
 sg13g2_decap_8 FILLER_32_347 ();
 sg13g2_decap_8 FILLER_32_354 ();
 sg13g2_decap_8 FILLER_32_361 ();
 sg13g2_decap_8 FILLER_32_368 ();
 sg13g2_decap_8 FILLER_32_375 ();
 sg13g2_decap_8 FILLER_32_382 ();
 sg13g2_decap_8 FILLER_32_389 ();
 sg13g2_decap_8 FILLER_32_396 ();
 sg13g2_decap_8 FILLER_32_403 ();
 sg13g2_decap_8 FILLER_32_410 ();
 sg13g2_decap_8 FILLER_32_417 ();
 sg13g2_decap_8 FILLER_32_424 ();
 sg13g2_decap_8 FILLER_32_431 ();
 sg13g2_decap_8 FILLER_32_438 ();
 sg13g2_decap_8 FILLER_32_445 ();
 sg13g2_decap_8 FILLER_32_452 ();
 sg13g2_decap_8 FILLER_32_459 ();
 sg13g2_decap_8 FILLER_32_466 ();
 sg13g2_decap_8 FILLER_32_473 ();
 sg13g2_decap_8 FILLER_32_480 ();
 sg13g2_decap_8 FILLER_32_487 ();
 sg13g2_decap_8 FILLER_32_494 ();
 sg13g2_decap_8 FILLER_32_501 ();
 sg13g2_decap_8 FILLER_32_508 ();
 sg13g2_decap_8 FILLER_32_515 ();
 sg13g2_decap_8 FILLER_32_522 ();
 sg13g2_decap_8 FILLER_32_529 ();
 sg13g2_decap_8 FILLER_32_536 ();
 sg13g2_decap_8 FILLER_32_543 ();
 sg13g2_decap_8 FILLER_32_550 ();
 sg13g2_decap_8 FILLER_32_557 ();
 sg13g2_decap_8 FILLER_32_564 ();
 sg13g2_decap_8 FILLER_32_571 ();
 sg13g2_decap_8 FILLER_32_578 ();
 sg13g2_decap_8 FILLER_32_585 ();
 sg13g2_decap_8 FILLER_32_592 ();
 sg13g2_decap_8 FILLER_32_599 ();
 sg13g2_decap_8 FILLER_32_606 ();
 sg13g2_decap_8 FILLER_32_613 ();
 sg13g2_decap_8 FILLER_32_620 ();
 sg13g2_decap_8 FILLER_32_627 ();
 sg13g2_decap_8 FILLER_32_634 ();
 sg13g2_decap_8 FILLER_32_641 ();
 sg13g2_decap_8 FILLER_32_648 ();
 sg13g2_decap_8 FILLER_32_655 ();
 sg13g2_decap_8 FILLER_32_662 ();
 sg13g2_decap_8 FILLER_32_669 ();
 sg13g2_decap_8 FILLER_32_676 ();
 sg13g2_decap_8 FILLER_32_683 ();
 sg13g2_decap_8 FILLER_32_690 ();
 sg13g2_decap_8 FILLER_32_697 ();
 sg13g2_decap_8 FILLER_32_704 ();
 sg13g2_decap_8 FILLER_32_711 ();
 sg13g2_decap_8 FILLER_32_718 ();
 sg13g2_decap_8 FILLER_32_725 ();
 sg13g2_decap_8 FILLER_32_732 ();
 sg13g2_decap_8 FILLER_32_739 ();
 sg13g2_decap_8 FILLER_32_746 ();
 sg13g2_decap_8 FILLER_32_753 ();
 sg13g2_decap_8 FILLER_32_760 ();
 sg13g2_decap_8 FILLER_32_767 ();
 sg13g2_decap_8 FILLER_32_774 ();
 sg13g2_decap_8 FILLER_32_781 ();
 sg13g2_decap_8 FILLER_32_788 ();
 sg13g2_decap_8 FILLER_32_795 ();
 sg13g2_decap_8 FILLER_32_802 ();
 sg13g2_decap_8 FILLER_32_809 ();
 sg13g2_decap_8 FILLER_32_816 ();
 sg13g2_decap_8 FILLER_32_823 ();
 sg13g2_decap_8 FILLER_32_830 ();
 sg13g2_decap_8 FILLER_32_837 ();
 sg13g2_decap_8 FILLER_32_844 ();
 sg13g2_decap_8 FILLER_32_851 ();
 sg13g2_decap_8 FILLER_32_858 ();
 sg13g2_decap_8 FILLER_32_865 ();
 sg13g2_decap_8 FILLER_32_872 ();
 sg13g2_decap_8 FILLER_32_879 ();
 sg13g2_decap_8 FILLER_32_886 ();
 sg13g2_decap_8 FILLER_32_893 ();
 sg13g2_decap_8 FILLER_32_900 ();
 sg13g2_decap_8 FILLER_32_907 ();
 sg13g2_decap_8 FILLER_32_914 ();
 sg13g2_decap_4 FILLER_32_921 ();
 sg13g2_decap_8 FILLER_33_4 ();
 sg13g2_decap_8 FILLER_33_11 ();
 sg13g2_decap_8 FILLER_33_18 ();
 sg13g2_decap_4 FILLER_33_25 ();
 sg13g2_decap_8 FILLER_33_33 ();
 sg13g2_decap_8 FILLER_33_40 ();
 sg13g2_decap_8 FILLER_33_51 ();
 sg13g2_decap_8 FILLER_33_58 ();
 sg13g2_decap_8 FILLER_33_65 ();
 sg13g2_decap_8 FILLER_33_72 ();
 sg13g2_decap_8 FILLER_33_79 ();
 sg13g2_decap_8 FILLER_33_86 ();
 sg13g2_decap_8 FILLER_33_93 ();
 sg13g2_decap_8 FILLER_33_100 ();
 sg13g2_fill_2 FILLER_33_107 ();
 sg13g2_decap_8 FILLER_33_114 ();
 sg13g2_decap_8 FILLER_33_121 ();
 sg13g2_decap_8 FILLER_33_128 ();
 sg13g2_decap_8 FILLER_33_135 ();
 sg13g2_decap_8 FILLER_33_142 ();
 sg13g2_decap_8 FILLER_33_149 ();
 sg13g2_decap_8 FILLER_33_156 ();
 sg13g2_decap_8 FILLER_33_163 ();
 sg13g2_decap_8 FILLER_33_170 ();
 sg13g2_decap_8 FILLER_33_177 ();
 sg13g2_decap_8 FILLER_33_184 ();
 sg13g2_decap_8 FILLER_33_191 ();
 sg13g2_decap_8 FILLER_33_198 ();
 sg13g2_decap_8 FILLER_33_205 ();
 sg13g2_decap_8 FILLER_33_212 ();
 sg13g2_decap_8 FILLER_33_219 ();
 sg13g2_decap_8 FILLER_33_226 ();
 sg13g2_decap_8 FILLER_33_233 ();
 sg13g2_decap_8 FILLER_33_240 ();
 sg13g2_decap_8 FILLER_33_247 ();
 sg13g2_decap_8 FILLER_33_254 ();
 sg13g2_decap_8 FILLER_33_261 ();
 sg13g2_decap_8 FILLER_33_268 ();
 sg13g2_decap_8 FILLER_33_275 ();
 sg13g2_decap_8 FILLER_33_282 ();
 sg13g2_decap_8 FILLER_33_289 ();
 sg13g2_decap_8 FILLER_33_296 ();
 sg13g2_decap_8 FILLER_33_303 ();
 sg13g2_decap_8 FILLER_33_310 ();
 sg13g2_decap_8 FILLER_33_317 ();
 sg13g2_decap_8 FILLER_33_324 ();
 sg13g2_decap_8 FILLER_33_331 ();
 sg13g2_decap_8 FILLER_33_338 ();
 sg13g2_decap_8 FILLER_33_345 ();
 sg13g2_decap_8 FILLER_33_352 ();
 sg13g2_decap_8 FILLER_33_359 ();
 sg13g2_decap_8 FILLER_33_366 ();
 sg13g2_decap_8 FILLER_33_373 ();
 sg13g2_decap_8 FILLER_33_380 ();
 sg13g2_decap_8 FILLER_33_387 ();
 sg13g2_decap_8 FILLER_33_394 ();
 sg13g2_decap_8 FILLER_33_401 ();
 sg13g2_decap_8 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_33_415 ();
 sg13g2_decap_8 FILLER_33_422 ();
 sg13g2_decap_8 FILLER_33_429 ();
 sg13g2_decap_8 FILLER_33_436 ();
 sg13g2_decap_8 FILLER_33_443 ();
 sg13g2_decap_8 FILLER_33_450 ();
 sg13g2_decap_8 FILLER_33_457 ();
 sg13g2_decap_8 FILLER_33_464 ();
 sg13g2_decap_8 FILLER_33_471 ();
 sg13g2_decap_8 FILLER_33_478 ();
 sg13g2_decap_8 FILLER_33_485 ();
 sg13g2_decap_8 FILLER_33_492 ();
 sg13g2_decap_8 FILLER_33_499 ();
 sg13g2_decap_8 FILLER_33_506 ();
 sg13g2_decap_8 FILLER_33_513 ();
 sg13g2_decap_8 FILLER_33_520 ();
 sg13g2_decap_8 FILLER_33_527 ();
 sg13g2_decap_8 FILLER_33_534 ();
 sg13g2_decap_8 FILLER_33_541 ();
 sg13g2_decap_8 FILLER_33_548 ();
 sg13g2_decap_8 FILLER_33_555 ();
 sg13g2_decap_8 FILLER_33_562 ();
 sg13g2_decap_8 FILLER_33_569 ();
 sg13g2_decap_8 FILLER_33_576 ();
 sg13g2_decap_8 FILLER_33_583 ();
 sg13g2_decap_8 FILLER_33_590 ();
 sg13g2_decap_8 FILLER_33_597 ();
 sg13g2_decap_8 FILLER_33_604 ();
 sg13g2_decap_8 FILLER_33_611 ();
 sg13g2_decap_8 FILLER_33_618 ();
 sg13g2_decap_8 FILLER_33_625 ();
 sg13g2_decap_8 FILLER_33_632 ();
 sg13g2_decap_8 FILLER_33_639 ();
 sg13g2_decap_8 FILLER_33_646 ();
 sg13g2_decap_8 FILLER_33_653 ();
 sg13g2_decap_8 FILLER_33_660 ();
 sg13g2_decap_8 FILLER_33_667 ();
 sg13g2_decap_8 FILLER_33_674 ();
 sg13g2_decap_8 FILLER_33_681 ();
 sg13g2_decap_8 FILLER_33_688 ();
 sg13g2_decap_8 FILLER_33_695 ();
 sg13g2_decap_8 FILLER_33_702 ();
 sg13g2_decap_8 FILLER_33_709 ();
 sg13g2_decap_8 FILLER_33_716 ();
 sg13g2_decap_8 FILLER_33_723 ();
 sg13g2_decap_8 FILLER_33_730 ();
 sg13g2_decap_8 FILLER_33_737 ();
 sg13g2_decap_8 FILLER_33_744 ();
 sg13g2_decap_8 FILLER_33_751 ();
 sg13g2_decap_8 FILLER_33_758 ();
 sg13g2_decap_8 FILLER_33_765 ();
 sg13g2_decap_8 FILLER_33_772 ();
 sg13g2_decap_8 FILLER_33_779 ();
 sg13g2_decap_8 FILLER_33_786 ();
 sg13g2_decap_8 FILLER_33_793 ();
 sg13g2_decap_8 FILLER_33_800 ();
 sg13g2_decap_8 FILLER_33_807 ();
 sg13g2_decap_8 FILLER_33_814 ();
 sg13g2_decap_8 FILLER_33_821 ();
 sg13g2_decap_8 FILLER_33_828 ();
 sg13g2_decap_8 FILLER_33_835 ();
 sg13g2_decap_8 FILLER_33_842 ();
 sg13g2_decap_8 FILLER_33_849 ();
 sg13g2_decap_8 FILLER_33_856 ();
 sg13g2_decap_8 FILLER_33_863 ();
 sg13g2_decap_8 FILLER_33_870 ();
 sg13g2_decap_8 FILLER_33_877 ();
 sg13g2_decap_8 FILLER_33_884 ();
 sg13g2_decap_8 FILLER_33_891 ();
 sg13g2_decap_8 FILLER_33_898 ();
 sg13g2_decap_8 FILLER_33_905 ();
 sg13g2_decap_8 FILLER_33_912 ();
 sg13g2_decap_4 FILLER_33_919 ();
 sg13g2_fill_2 FILLER_33_923 ();
 sg13g2_decap_8 FILLER_34_4 ();
 sg13g2_decap_8 FILLER_34_11 ();
 sg13g2_decap_8 FILLER_34_18 ();
 sg13g2_decap_4 FILLER_34_25 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_118 ();
 sg13g2_decap_8 FILLER_34_125 ();
 sg13g2_decap_8 FILLER_34_132 ();
 sg13g2_decap_8 FILLER_34_139 ();
 sg13g2_decap_8 FILLER_34_146 ();
 sg13g2_decap_8 FILLER_34_153 ();
 sg13g2_decap_8 FILLER_34_160 ();
 sg13g2_decap_8 FILLER_34_167 ();
 sg13g2_decap_8 FILLER_34_174 ();
 sg13g2_decap_8 FILLER_34_181 ();
 sg13g2_decap_8 FILLER_34_188 ();
 sg13g2_decap_8 FILLER_34_195 ();
 sg13g2_decap_8 FILLER_34_202 ();
 sg13g2_decap_8 FILLER_34_209 ();
 sg13g2_decap_8 FILLER_34_216 ();
 sg13g2_decap_8 FILLER_34_223 ();
 sg13g2_decap_8 FILLER_34_230 ();
 sg13g2_decap_8 FILLER_34_237 ();
 sg13g2_decap_8 FILLER_34_244 ();
 sg13g2_decap_8 FILLER_34_251 ();
 sg13g2_decap_8 FILLER_34_258 ();
 sg13g2_decap_8 FILLER_34_265 ();
 sg13g2_decap_8 FILLER_34_272 ();
 sg13g2_decap_8 FILLER_34_279 ();
 sg13g2_decap_8 FILLER_34_286 ();
 sg13g2_decap_8 FILLER_34_293 ();
 sg13g2_decap_8 FILLER_34_300 ();
 sg13g2_decap_8 FILLER_34_307 ();
 sg13g2_decap_8 FILLER_34_314 ();
 sg13g2_decap_8 FILLER_34_321 ();
 sg13g2_decap_8 FILLER_34_328 ();
 sg13g2_decap_8 FILLER_34_335 ();
 sg13g2_decap_8 FILLER_34_342 ();
 sg13g2_decap_8 FILLER_34_349 ();
 sg13g2_decap_8 FILLER_34_356 ();
 sg13g2_decap_8 FILLER_34_363 ();
 sg13g2_decap_8 FILLER_34_370 ();
 sg13g2_decap_8 FILLER_34_377 ();
 sg13g2_decap_8 FILLER_34_384 ();
 sg13g2_decap_8 FILLER_34_391 ();
 sg13g2_decap_8 FILLER_34_398 ();
 sg13g2_decap_8 FILLER_34_405 ();
 sg13g2_decap_8 FILLER_34_412 ();
 sg13g2_decap_8 FILLER_34_419 ();
 sg13g2_decap_8 FILLER_34_426 ();
 sg13g2_decap_8 FILLER_34_433 ();
 sg13g2_decap_8 FILLER_34_440 ();
 sg13g2_decap_8 FILLER_34_447 ();
 sg13g2_decap_8 FILLER_34_454 ();
 sg13g2_decap_8 FILLER_34_461 ();
 sg13g2_decap_8 FILLER_34_468 ();
 sg13g2_decap_8 FILLER_34_475 ();
 sg13g2_decap_8 FILLER_34_482 ();
 sg13g2_decap_8 FILLER_34_489 ();
 sg13g2_decap_8 FILLER_34_496 ();
 sg13g2_decap_8 FILLER_34_503 ();
 sg13g2_decap_8 FILLER_34_510 ();
 sg13g2_decap_8 FILLER_34_517 ();
 sg13g2_decap_8 FILLER_34_524 ();
 sg13g2_decap_8 FILLER_34_531 ();
 sg13g2_decap_8 FILLER_34_538 ();
 sg13g2_decap_8 FILLER_34_545 ();
 sg13g2_decap_8 FILLER_34_552 ();
 sg13g2_decap_8 FILLER_34_559 ();
 sg13g2_decap_8 FILLER_34_566 ();
 sg13g2_decap_8 FILLER_34_573 ();
 sg13g2_decap_8 FILLER_34_580 ();
 sg13g2_decap_8 FILLER_34_587 ();
 sg13g2_decap_8 FILLER_34_594 ();
 sg13g2_decap_8 FILLER_34_601 ();
 sg13g2_decap_8 FILLER_34_608 ();
 sg13g2_decap_8 FILLER_34_615 ();
 sg13g2_decap_8 FILLER_34_622 ();
 sg13g2_decap_8 FILLER_34_629 ();
 sg13g2_decap_8 FILLER_34_636 ();
 sg13g2_decap_8 FILLER_34_643 ();
 sg13g2_decap_8 FILLER_34_650 ();
 sg13g2_decap_8 FILLER_34_657 ();
 sg13g2_decap_8 FILLER_34_664 ();
 sg13g2_decap_8 FILLER_34_671 ();
 sg13g2_decap_8 FILLER_34_678 ();
 sg13g2_decap_8 FILLER_34_685 ();
 sg13g2_decap_8 FILLER_34_692 ();
 sg13g2_decap_8 FILLER_34_699 ();
 sg13g2_decap_8 FILLER_34_706 ();
 sg13g2_decap_8 FILLER_34_713 ();
 sg13g2_decap_8 FILLER_34_720 ();
 sg13g2_decap_8 FILLER_34_727 ();
 sg13g2_decap_8 FILLER_34_734 ();
 sg13g2_decap_8 FILLER_34_741 ();
 sg13g2_decap_8 FILLER_34_748 ();
 sg13g2_decap_8 FILLER_34_755 ();
 sg13g2_decap_8 FILLER_34_762 ();
 sg13g2_decap_8 FILLER_34_769 ();
 sg13g2_decap_8 FILLER_34_776 ();
 sg13g2_decap_8 FILLER_34_783 ();
 sg13g2_decap_8 FILLER_34_790 ();
 sg13g2_decap_8 FILLER_34_797 ();
 sg13g2_decap_8 FILLER_34_804 ();
 sg13g2_decap_8 FILLER_34_811 ();
 sg13g2_decap_8 FILLER_34_818 ();
 sg13g2_decap_8 FILLER_34_825 ();
 sg13g2_decap_8 FILLER_34_832 ();
 sg13g2_decap_8 FILLER_34_839 ();
 sg13g2_decap_8 FILLER_34_846 ();
 sg13g2_decap_8 FILLER_34_853 ();
 sg13g2_decap_8 FILLER_34_860 ();
 sg13g2_decap_8 FILLER_34_867 ();
 sg13g2_decap_8 FILLER_34_874 ();
 sg13g2_decap_8 FILLER_34_881 ();
 sg13g2_decap_8 FILLER_34_888 ();
 sg13g2_decap_8 FILLER_34_895 ();
 sg13g2_decap_8 FILLER_34_902 ();
 sg13g2_decap_8 FILLER_34_909 ();
 sg13g2_decap_8 FILLER_34_916 ();
 sg13g2_fill_2 FILLER_34_923 ();
 sg13g2_decap_8 FILLER_35_4 ();
 sg13g2_decap_8 FILLER_35_11 ();
 sg13g2_decap_8 FILLER_35_18 ();
 sg13g2_decap_8 FILLER_35_25 ();
 sg13g2_decap_8 FILLER_35_32 ();
 sg13g2_decap_8 FILLER_35_39 ();
 sg13g2_decap_8 FILLER_35_46 ();
 sg13g2_decap_8 FILLER_35_53 ();
 sg13g2_decap_8 FILLER_35_60 ();
 sg13g2_decap_8 FILLER_35_67 ();
 sg13g2_decap_8 FILLER_35_74 ();
 sg13g2_decap_8 FILLER_35_81 ();
 sg13g2_decap_8 FILLER_35_88 ();
 sg13g2_decap_8 FILLER_35_95 ();
 sg13g2_decap_8 FILLER_35_102 ();
 sg13g2_decap_8 FILLER_35_114 ();
 sg13g2_decap_8 FILLER_35_121 ();
 sg13g2_decap_8 FILLER_35_128 ();
 sg13g2_decap_8 FILLER_35_135 ();
 sg13g2_decap_8 FILLER_35_142 ();
 sg13g2_decap_8 FILLER_35_149 ();
 sg13g2_decap_8 FILLER_35_156 ();
 sg13g2_decap_8 FILLER_35_163 ();
 sg13g2_decap_8 FILLER_35_170 ();
 sg13g2_decap_8 FILLER_35_177 ();
 sg13g2_decap_8 FILLER_35_184 ();
 sg13g2_decap_8 FILLER_35_191 ();
 sg13g2_decap_8 FILLER_35_198 ();
 sg13g2_decap_8 FILLER_35_205 ();
 sg13g2_decap_8 FILLER_35_212 ();
 sg13g2_decap_8 FILLER_35_219 ();
 sg13g2_decap_8 FILLER_35_226 ();
 sg13g2_decap_8 FILLER_35_233 ();
 sg13g2_decap_8 FILLER_35_240 ();
 sg13g2_decap_8 FILLER_35_247 ();
 sg13g2_decap_8 FILLER_35_254 ();
 sg13g2_decap_8 FILLER_35_261 ();
 sg13g2_decap_8 FILLER_35_268 ();
 sg13g2_decap_8 FILLER_35_275 ();
 sg13g2_decap_8 FILLER_35_282 ();
 sg13g2_decap_8 FILLER_35_289 ();
 sg13g2_decap_8 FILLER_35_296 ();
 sg13g2_decap_8 FILLER_35_303 ();
 sg13g2_decap_8 FILLER_35_310 ();
 sg13g2_decap_8 FILLER_35_317 ();
 sg13g2_decap_8 FILLER_35_324 ();
 sg13g2_decap_8 FILLER_35_331 ();
 sg13g2_decap_8 FILLER_35_338 ();
 sg13g2_decap_8 FILLER_35_345 ();
 sg13g2_decap_8 FILLER_35_352 ();
 sg13g2_decap_8 FILLER_35_359 ();
 sg13g2_decap_8 FILLER_35_366 ();
 sg13g2_decap_8 FILLER_35_373 ();
 sg13g2_decap_8 FILLER_35_380 ();
 sg13g2_decap_8 FILLER_35_387 ();
 sg13g2_decap_8 FILLER_35_394 ();
 sg13g2_decap_8 FILLER_35_401 ();
 sg13g2_decap_8 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_35_415 ();
 sg13g2_decap_8 FILLER_35_422 ();
 sg13g2_decap_8 FILLER_35_429 ();
 sg13g2_decap_8 FILLER_35_436 ();
 sg13g2_decap_8 FILLER_35_443 ();
 sg13g2_decap_8 FILLER_35_450 ();
 sg13g2_decap_8 FILLER_35_457 ();
 sg13g2_decap_8 FILLER_35_464 ();
 sg13g2_decap_8 FILLER_35_471 ();
 sg13g2_decap_8 FILLER_35_478 ();
 sg13g2_decap_8 FILLER_35_485 ();
 sg13g2_decap_8 FILLER_35_492 ();
 sg13g2_decap_8 FILLER_35_499 ();
 sg13g2_decap_8 FILLER_35_506 ();
 sg13g2_decap_8 FILLER_35_513 ();
 sg13g2_decap_8 FILLER_35_520 ();
 sg13g2_decap_8 FILLER_35_527 ();
 sg13g2_decap_8 FILLER_35_534 ();
 sg13g2_decap_8 FILLER_35_541 ();
 sg13g2_decap_8 FILLER_35_548 ();
 sg13g2_decap_8 FILLER_35_555 ();
 sg13g2_decap_8 FILLER_35_562 ();
 sg13g2_decap_8 FILLER_35_569 ();
 sg13g2_decap_8 FILLER_35_576 ();
 sg13g2_decap_8 FILLER_35_583 ();
 sg13g2_decap_8 FILLER_35_590 ();
 sg13g2_decap_8 FILLER_35_597 ();
 sg13g2_decap_8 FILLER_35_604 ();
 sg13g2_decap_8 FILLER_35_611 ();
 sg13g2_decap_8 FILLER_35_618 ();
 sg13g2_decap_8 FILLER_35_625 ();
 sg13g2_decap_8 FILLER_35_632 ();
 sg13g2_decap_8 FILLER_35_639 ();
 sg13g2_decap_8 FILLER_35_646 ();
 sg13g2_decap_8 FILLER_35_653 ();
 sg13g2_decap_8 FILLER_35_660 ();
 sg13g2_decap_8 FILLER_35_667 ();
 sg13g2_decap_8 FILLER_35_674 ();
 sg13g2_decap_8 FILLER_35_681 ();
 sg13g2_decap_8 FILLER_35_688 ();
 sg13g2_decap_8 FILLER_35_695 ();
 sg13g2_decap_8 FILLER_35_702 ();
 sg13g2_decap_8 FILLER_35_709 ();
 sg13g2_decap_8 FILLER_35_716 ();
 sg13g2_decap_8 FILLER_35_723 ();
 sg13g2_decap_8 FILLER_35_730 ();
 sg13g2_decap_8 FILLER_35_737 ();
 sg13g2_decap_8 FILLER_35_744 ();
 sg13g2_decap_8 FILLER_35_751 ();
 sg13g2_decap_8 FILLER_35_758 ();
 sg13g2_decap_8 FILLER_35_765 ();
 sg13g2_decap_8 FILLER_35_772 ();
 sg13g2_decap_8 FILLER_35_779 ();
 sg13g2_decap_8 FILLER_35_786 ();
 sg13g2_decap_8 FILLER_35_793 ();
 sg13g2_decap_8 FILLER_35_800 ();
 sg13g2_decap_8 FILLER_35_807 ();
 sg13g2_decap_8 FILLER_35_814 ();
 sg13g2_decap_8 FILLER_35_821 ();
 sg13g2_decap_8 FILLER_35_828 ();
 sg13g2_decap_8 FILLER_35_835 ();
 sg13g2_decap_8 FILLER_35_842 ();
 sg13g2_decap_8 FILLER_35_849 ();
 sg13g2_decap_8 FILLER_35_856 ();
 sg13g2_decap_8 FILLER_35_863 ();
 sg13g2_decap_8 FILLER_35_870 ();
 sg13g2_decap_8 FILLER_35_877 ();
 sg13g2_decap_8 FILLER_35_884 ();
 sg13g2_decap_8 FILLER_35_891 ();
 sg13g2_decap_8 FILLER_35_898 ();
 sg13g2_decap_8 FILLER_35_905 ();
 sg13g2_decap_8 FILLER_35_912 ();
 sg13g2_decap_4 FILLER_35_919 ();
 sg13g2_fill_2 FILLER_35_923 ();
 sg13g2_decap_8 FILLER_36_4 ();
 sg13g2_decap_8 FILLER_36_11 ();
 sg13g2_decap_8 FILLER_36_18 ();
 sg13g2_decap_8 FILLER_36_25 ();
 sg13g2_decap_8 FILLER_36_32 ();
 sg13g2_decap_8 FILLER_36_39 ();
 sg13g2_decap_8 FILLER_36_46 ();
 sg13g2_decap_8 FILLER_36_53 ();
 sg13g2_decap_8 FILLER_36_60 ();
 sg13g2_decap_8 FILLER_36_67 ();
 sg13g2_decap_8 FILLER_36_74 ();
 sg13g2_decap_8 FILLER_36_81 ();
 sg13g2_decap_8 FILLER_36_88 ();
 sg13g2_decap_8 FILLER_36_95 ();
 sg13g2_decap_8 FILLER_36_102 ();
 sg13g2_decap_8 FILLER_36_109 ();
 sg13g2_decap_8 FILLER_36_116 ();
 sg13g2_decap_8 FILLER_36_123 ();
 sg13g2_decap_8 FILLER_36_130 ();
 sg13g2_decap_8 FILLER_36_137 ();
 sg13g2_decap_8 FILLER_36_144 ();
 sg13g2_decap_8 FILLER_36_151 ();
 sg13g2_decap_8 FILLER_36_158 ();
 sg13g2_decap_8 FILLER_36_165 ();
 sg13g2_decap_8 FILLER_36_172 ();
 sg13g2_decap_8 FILLER_36_179 ();
 sg13g2_decap_8 FILLER_36_186 ();
 sg13g2_decap_8 FILLER_36_193 ();
 sg13g2_decap_8 FILLER_36_200 ();
 sg13g2_decap_8 FILLER_36_207 ();
 sg13g2_decap_8 FILLER_36_214 ();
 sg13g2_decap_8 FILLER_36_221 ();
 sg13g2_decap_8 FILLER_36_228 ();
 sg13g2_decap_8 FILLER_36_235 ();
 sg13g2_decap_8 FILLER_36_242 ();
 sg13g2_decap_8 FILLER_36_249 ();
 sg13g2_decap_8 FILLER_36_256 ();
 sg13g2_decap_8 FILLER_36_263 ();
 sg13g2_decap_8 FILLER_36_270 ();
 sg13g2_decap_8 FILLER_36_277 ();
 sg13g2_decap_8 FILLER_36_284 ();
 sg13g2_decap_8 FILLER_36_291 ();
 sg13g2_decap_8 FILLER_36_298 ();
 sg13g2_decap_8 FILLER_36_305 ();
 sg13g2_decap_8 FILLER_36_312 ();
 sg13g2_decap_8 FILLER_36_319 ();
 sg13g2_decap_8 FILLER_36_326 ();
 sg13g2_decap_8 FILLER_36_333 ();
 sg13g2_decap_8 FILLER_36_340 ();
 sg13g2_decap_8 FILLER_36_347 ();
 sg13g2_decap_8 FILLER_36_354 ();
 sg13g2_decap_8 FILLER_36_361 ();
 sg13g2_decap_8 FILLER_36_368 ();
 sg13g2_decap_8 FILLER_36_375 ();
 sg13g2_decap_8 FILLER_36_382 ();
 sg13g2_decap_8 FILLER_36_389 ();
 sg13g2_decap_8 FILLER_36_396 ();
 sg13g2_decap_8 FILLER_36_403 ();
 sg13g2_decap_8 FILLER_36_410 ();
 sg13g2_decap_8 FILLER_36_417 ();
 sg13g2_decap_8 FILLER_36_424 ();
 sg13g2_decap_8 FILLER_36_431 ();
 sg13g2_decap_8 FILLER_36_438 ();
 sg13g2_decap_8 FILLER_36_445 ();
 sg13g2_decap_8 FILLER_36_452 ();
 sg13g2_decap_8 FILLER_36_459 ();
 sg13g2_decap_8 FILLER_36_466 ();
 sg13g2_decap_8 FILLER_36_473 ();
 sg13g2_decap_8 FILLER_36_480 ();
 sg13g2_decap_8 FILLER_36_487 ();
 sg13g2_decap_8 FILLER_36_494 ();
 sg13g2_decap_8 FILLER_36_501 ();
 sg13g2_decap_8 FILLER_36_508 ();
 sg13g2_decap_8 FILLER_36_515 ();
 sg13g2_decap_8 FILLER_36_522 ();
 sg13g2_decap_8 FILLER_36_529 ();
 sg13g2_decap_8 FILLER_36_536 ();
 sg13g2_decap_8 FILLER_36_543 ();
 sg13g2_decap_8 FILLER_36_550 ();
 sg13g2_decap_8 FILLER_36_557 ();
 sg13g2_decap_8 FILLER_36_564 ();
 sg13g2_decap_8 FILLER_36_571 ();
 sg13g2_decap_8 FILLER_36_578 ();
 sg13g2_decap_8 FILLER_36_585 ();
 sg13g2_decap_8 FILLER_36_592 ();
 sg13g2_decap_8 FILLER_36_599 ();
 sg13g2_decap_8 FILLER_36_606 ();
 sg13g2_decap_8 FILLER_36_613 ();
 sg13g2_decap_8 FILLER_36_620 ();
 sg13g2_decap_8 FILLER_36_627 ();
 sg13g2_decap_8 FILLER_36_634 ();
 sg13g2_decap_8 FILLER_36_641 ();
 sg13g2_decap_8 FILLER_36_648 ();
 sg13g2_decap_8 FILLER_36_655 ();
 sg13g2_decap_8 FILLER_36_662 ();
 sg13g2_decap_8 FILLER_36_669 ();
 sg13g2_decap_8 FILLER_36_676 ();
 sg13g2_decap_8 FILLER_36_683 ();
 sg13g2_decap_8 FILLER_36_690 ();
 sg13g2_decap_8 FILLER_36_697 ();
 sg13g2_decap_8 FILLER_36_704 ();
 sg13g2_decap_8 FILLER_36_711 ();
 sg13g2_decap_8 FILLER_36_718 ();
 sg13g2_decap_8 FILLER_36_725 ();
 sg13g2_decap_8 FILLER_36_732 ();
 sg13g2_decap_8 FILLER_36_739 ();
 sg13g2_decap_8 FILLER_36_746 ();
 sg13g2_decap_8 FILLER_36_753 ();
 sg13g2_decap_8 FILLER_36_760 ();
 sg13g2_decap_8 FILLER_36_767 ();
 sg13g2_decap_8 FILLER_36_774 ();
 sg13g2_decap_8 FILLER_36_781 ();
 sg13g2_decap_8 FILLER_36_788 ();
 sg13g2_decap_8 FILLER_36_795 ();
 sg13g2_decap_8 FILLER_36_802 ();
 sg13g2_decap_8 FILLER_36_809 ();
 sg13g2_decap_8 FILLER_36_816 ();
 sg13g2_decap_8 FILLER_36_823 ();
 sg13g2_decap_8 FILLER_36_830 ();
 sg13g2_decap_8 FILLER_36_837 ();
 sg13g2_decap_8 FILLER_36_844 ();
 sg13g2_decap_8 FILLER_36_851 ();
 sg13g2_decap_8 FILLER_36_858 ();
 sg13g2_decap_8 FILLER_36_865 ();
 sg13g2_decap_8 FILLER_36_872 ();
 sg13g2_decap_8 FILLER_36_879 ();
 sg13g2_decap_8 FILLER_36_886 ();
 sg13g2_decap_8 FILLER_36_893 ();
 sg13g2_decap_8 FILLER_36_900 ();
 sg13g2_decap_8 FILLER_36_907 ();
 sg13g2_decap_8 FILLER_36_914 ();
 sg13g2_decap_4 FILLER_36_921 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_decap_8 FILLER_37_91 ();
 sg13g2_decap_8 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_105 ();
 sg13g2_decap_8 FILLER_37_112 ();
 sg13g2_decap_8 FILLER_37_119 ();
 sg13g2_decap_8 FILLER_37_126 ();
 sg13g2_decap_8 FILLER_37_133 ();
 sg13g2_decap_8 FILLER_37_140 ();
 sg13g2_decap_8 FILLER_37_147 ();
 sg13g2_decap_8 FILLER_37_154 ();
 sg13g2_decap_8 FILLER_37_161 ();
 sg13g2_decap_8 FILLER_37_168 ();
 sg13g2_decap_8 FILLER_37_175 ();
 sg13g2_decap_8 FILLER_37_182 ();
 sg13g2_decap_8 FILLER_37_189 ();
 sg13g2_decap_8 FILLER_37_196 ();
 sg13g2_decap_8 FILLER_37_203 ();
 sg13g2_decap_8 FILLER_37_210 ();
 sg13g2_decap_8 FILLER_37_217 ();
 sg13g2_decap_8 FILLER_37_224 ();
 sg13g2_decap_8 FILLER_37_231 ();
 sg13g2_decap_8 FILLER_37_238 ();
 sg13g2_decap_8 FILLER_37_245 ();
 sg13g2_decap_8 FILLER_37_252 ();
 sg13g2_decap_8 FILLER_37_259 ();
 sg13g2_decap_8 FILLER_37_266 ();
 sg13g2_decap_8 FILLER_37_273 ();
 sg13g2_decap_8 FILLER_37_280 ();
 sg13g2_decap_8 FILLER_37_287 ();
 sg13g2_decap_8 FILLER_37_294 ();
 sg13g2_decap_8 FILLER_37_301 ();
 sg13g2_decap_8 FILLER_37_308 ();
 sg13g2_decap_8 FILLER_37_315 ();
 sg13g2_decap_8 FILLER_37_322 ();
 sg13g2_decap_8 FILLER_37_329 ();
 sg13g2_decap_8 FILLER_37_336 ();
 sg13g2_decap_8 FILLER_37_343 ();
 sg13g2_decap_8 FILLER_37_350 ();
 sg13g2_decap_8 FILLER_37_357 ();
 sg13g2_decap_8 FILLER_37_364 ();
 sg13g2_decap_8 FILLER_37_371 ();
 sg13g2_decap_8 FILLER_37_378 ();
 sg13g2_decap_8 FILLER_37_385 ();
 sg13g2_decap_8 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_399 ();
 sg13g2_decap_8 FILLER_37_406 ();
 sg13g2_decap_8 FILLER_37_413 ();
 sg13g2_decap_8 FILLER_37_420 ();
 sg13g2_decap_8 FILLER_37_427 ();
 sg13g2_decap_8 FILLER_37_434 ();
 sg13g2_decap_8 FILLER_37_441 ();
 sg13g2_decap_8 FILLER_37_448 ();
 sg13g2_decap_8 FILLER_37_455 ();
 sg13g2_decap_8 FILLER_37_462 ();
 sg13g2_decap_8 FILLER_37_469 ();
 sg13g2_decap_8 FILLER_37_476 ();
 sg13g2_decap_8 FILLER_37_483 ();
 sg13g2_decap_8 FILLER_37_490 ();
 sg13g2_decap_8 FILLER_37_497 ();
 sg13g2_decap_8 FILLER_37_504 ();
 sg13g2_decap_8 FILLER_37_511 ();
 sg13g2_decap_8 FILLER_37_518 ();
 sg13g2_decap_8 FILLER_37_525 ();
 sg13g2_decap_8 FILLER_37_532 ();
 sg13g2_decap_8 FILLER_37_539 ();
 sg13g2_decap_8 FILLER_37_546 ();
 sg13g2_decap_8 FILLER_37_553 ();
 sg13g2_decap_8 FILLER_37_560 ();
 sg13g2_decap_8 FILLER_37_567 ();
 sg13g2_decap_8 FILLER_37_574 ();
 sg13g2_decap_8 FILLER_37_581 ();
 sg13g2_decap_8 FILLER_37_588 ();
 sg13g2_decap_8 FILLER_37_595 ();
 sg13g2_decap_8 FILLER_37_602 ();
 sg13g2_decap_8 FILLER_37_609 ();
 sg13g2_decap_8 FILLER_37_616 ();
 sg13g2_decap_8 FILLER_37_623 ();
 sg13g2_decap_8 FILLER_37_630 ();
 sg13g2_decap_8 FILLER_37_637 ();
 sg13g2_decap_8 FILLER_37_644 ();
 sg13g2_decap_8 FILLER_37_651 ();
 sg13g2_decap_8 FILLER_37_658 ();
 sg13g2_decap_8 FILLER_37_665 ();
 sg13g2_decap_8 FILLER_37_672 ();
 sg13g2_decap_8 FILLER_37_679 ();
 sg13g2_decap_8 FILLER_37_686 ();
 sg13g2_decap_8 FILLER_37_693 ();
 sg13g2_decap_8 FILLER_37_700 ();
 sg13g2_decap_8 FILLER_37_707 ();
 sg13g2_decap_8 FILLER_37_714 ();
 sg13g2_decap_8 FILLER_37_721 ();
 sg13g2_decap_8 FILLER_37_728 ();
 sg13g2_decap_8 FILLER_37_735 ();
 sg13g2_decap_8 FILLER_37_742 ();
 sg13g2_decap_8 FILLER_37_749 ();
 sg13g2_decap_8 FILLER_37_756 ();
 sg13g2_decap_8 FILLER_37_763 ();
 sg13g2_decap_8 FILLER_37_770 ();
 sg13g2_decap_8 FILLER_37_777 ();
 sg13g2_decap_8 FILLER_37_784 ();
 sg13g2_decap_8 FILLER_37_791 ();
 sg13g2_decap_8 FILLER_37_798 ();
 sg13g2_decap_8 FILLER_37_805 ();
 sg13g2_decap_8 FILLER_37_812 ();
 sg13g2_decap_8 FILLER_37_819 ();
 sg13g2_decap_8 FILLER_37_826 ();
 sg13g2_decap_8 FILLER_37_833 ();
 sg13g2_decap_8 FILLER_37_840 ();
 sg13g2_decap_8 FILLER_37_847 ();
 sg13g2_decap_8 FILLER_37_854 ();
 sg13g2_decap_8 FILLER_37_861 ();
 sg13g2_decap_8 FILLER_37_868 ();
 sg13g2_decap_8 FILLER_37_875 ();
 sg13g2_decap_8 FILLER_37_882 ();
 sg13g2_decap_8 FILLER_37_889 ();
 sg13g2_decap_8 FILLER_37_896 ();
 sg13g2_decap_8 FILLER_37_903 ();
 sg13g2_decap_8 FILLER_37_910 ();
 sg13g2_decap_8 FILLER_37_917 ();
 sg13g2_fill_1 FILLER_37_924 ();
 sg13g2_decap_8 FILLER_38_4 ();
 sg13g2_decap_4 FILLER_38_11 ();
 sg13g2_fill_2 FILLER_38_15 ();
 sg13g2_decap_8 FILLER_38_33 ();
 sg13g2_decap_8 FILLER_38_40 ();
 sg13g2_decap_8 FILLER_38_47 ();
 sg13g2_decap_8 FILLER_38_54 ();
 sg13g2_decap_8 FILLER_38_61 ();
 sg13g2_decap_8 FILLER_38_68 ();
 sg13g2_decap_8 FILLER_38_75 ();
 sg13g2_decap_8 FILLER_38_82 ();
 sg13g2_decap_8 FILLER_38_89 ();
 sg13g2_decap_8 FILLER_38_96 ();
 sg13g2_decap_8 FILLER_38_103 ();
 sg13g2_decap_8 FILLER_38_110 ();
 sg13g2_decap_8 FILLER_38_117 ();
 sg13g2_decap_8 FILLER_38_124 ();
 sg13g2_decap_8 FILLER_38_131 ();
 sg13g2_decap_8 FILLER_38_138 ();
 sg13g2_decap_8 FILLER_38_145 ();
 sg13g2_decap_8 FILLER_38_152 ();
 sg13g2_decap_8 FILLER_38_159 ();
 sg13g2_decap_8 FILLER_38_166 ();
 sg13g2_decap_8 FILLER_38_173 ();
 sg13g2_decap_8 FILLER_38_180 ();
 sg13g2_decap_8 FILLER_38_187 ();
 sg13g2_decap_8 FILLER_38_194 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_decap_8 FILLER_38_208 ();
 sg13g2_decap_8 FILLER_38_215 ();
 sg13g2_decap_8 FILLER_38_222 ();
 sg13g2_decap_8 FILLER_38_229 ();
 sg13g2_decap_8 FILLER_38_236 ();
 sg13g2_decap_8 FILLER_38_243 ();
 sg13g2_decap_8 FILLER_38_250 ();
 sg13g2_decap_8 FILLER_38_257 ();
 sg13g2_decap_8 FILLER_38_264 ();
 sg13g2_decap_8 FILLER_38_271 ();
 sg13g2_decap_8 FILLER_38_278 ();
 sg13g2_decap_8 FILLER_38_285 ();
 sg13g2_decap_8 FILLER_38_292 ();
 sg13g2_decap_8 FILLER_38_299 ();
 sg13g2_decap_8 FILLER_38_306 ();
 sg13g2_decap_8 FILLER_38_313 ();
 sg13g2_decap_8 FILLER_38_320 ();
 sg13g2_decap_8 FILLER_38_327 ();
 sg13g2_decap_8 FILLER_38_334 ();
 sg13g2_decap_8 FILLER_38_341 ();
 sg13g2_decap_8 FILLER_38_348 ();
 sg13g2_decap_8 FILLER_38_355 ();
 sg13g2_decap_8 FILLER_38_362 ();
 sg13g2_decap_8 FILLER_38_369 ();
 sg13g2_decap_8 FILLER_38_376 ();
 sg13g2_decap_8 FILLER_38_383 ();
 sg13g2_decap_8 FILLER_38_390 ();
 sg13g2_decap_8 FILLER_38_397 ();
 sg13g2_decap_8 FILLER_38_404 ();
 sg13g2_decap_8 FILLER_38_411 ();
 sg13g2_decap_8 FILLER_38_418 ();
 sg13g2_decap_8 FILLER_38_425 ();
 sg13g2_decap_8 FILLER_38_432 ();
 sg13g2_decap_8 FILLER_38_439 ();
 sg13g2_decap_8 FILLER_38_446 ();
 sg13g2_decap_8 FILLER_38_453 ();
 sg13g2_decap_8 FILLER_38_460 ();
 sg13g2_decap_8 FILLER_38_467 ();
 sg13g2_decap_8 FILLER_38_474 ();
 sg13g2_decap_8 FILLER_38_481 ();
 sg13g2_decap_8 FILLER_38_488 ();
 sg13g2_decap_8 FILLER_38_495 ();
 sg13g2_decap_8 FILLER_38_502 ();
 sg13g2_decap_8 FILLER_38_509 ();
 sg13g2_decap_8 FILLER_38_516 ();
 sg13g2_decap_8 FILLER_38_523 ();
 sg13g2_decap_8 FILLER_38_530 ();
 sg13g2_decap_8 FILLER_38_537 ();
 sg13g2_decap_8 FILLER_38_544 ();
 sg13g2_decap_8 FILLER_38_551 ();
 sg13g2_decap_8 FILLER_38_558 ();
 sg13g2_decap_8 FILLER_38_565 ();
 sg13g2_decap_8 FILLER_38_572 ();
 sg13g2_decap_8 FILLER_38_579 ();
 sg13g2_decap_8 FILLER_38_586 ();
 sg13g2_decap_8 FILLER_38_593 ();
 sg13g2_decap_8 FILLER_38_600 ();
 sg13g2_decap_8 FILLER_38_607 ();
 sg13g2_decap_8 FILLER_38_614 ();
 sg13g2_decap_8 FILLER_38_621 ();
 sg13g2_decap_8 FILLER_38_628 ();
 sg13g2_decap_8 FILLER_38_635 ();
 sg13g2_decap_8 FILLER_38_642 ();
 sg13g2_decap_8 FILLER_38_649 ();
 sg13g2_decap_8 FILLER_38_656 ();
 sg13g2_decap_8 FILLER_38_663 ();
 sg13g2_decap_8 FILLER_38_670 ();
 sg13g2_decap_8 FILLER_38_677 ();
 sg13g2_decap_8 FILLER_38_684 ();
 sg13g2_decap_8 FILLER_38_691 ();
 sg13g2_decap_8 FILLER_38_698 ();
 sg13g2_decap_8 FILLER_38_705 ();
 sg13g2_decap_8 FILLER_38_712 ();
 sg13g2_decap_8 FILLER_38_719 ();
 sg13g2_decap_8 FILLER_38_726 ();
 sg13g2_decap_8 FILLER_38_733 ();
 sg13g2_decap_8 FILLER_38_740 ();
 sg13g2_decap_8 FILLER_38_747 ();
 sg13g2_decap_8 FILLER_38_754 ();
 sg13g2_decap_8 FILLER_38_761 ();
 sg13g2_decap_8 FILLER_38_768 ();
 sg13g2_decap_8 FILLER_38_775 ();
 sg13g2_decap_8 FILLER_38_782 ();
 sg13g2_decap_8 FILLER_38_789 ();
 sg13g2_decap_8 FILLER_38_796 ();
 sg13g2_decap_8 FILLER_38_803 ();
 sg13g2_decap_8 FILLER_38_810 ();
 sg13g2_decap_8 FILLER_38_817 ();
 sg13g2_decap_8 FILLER_38_824 ();
 sg13g2_decap_8 FILLER_38_831 ();
 sg13g2_decap_8 FILLER_38_838 ();
 sg13g2_decap_8 FILLER_38_845 ();
 sg13g2_decap_8 FILLER_38_852 ();
 sg13g2_decap_8 FILLER_38_859 ();
 sg13g2_decap_8 FILLER_38_866 ();
 sg13g2_decap_8 FILLER_38_873 ();
 sg13g2_decap_8 FILLER_38_880 ();
 sg13g2_decap_8 FILLER_38_887 ();
 sg13g2_decap_8 FILLER_38_894 ();
 sg13g2_decap_8 FILLER_38_901 ();
 sg13g2_decap_8 FILLER_38_908 ();
 sg13g2_decap_8 FILLER_38_915 ();
 sg13g2_fill_2 FILLER_38_922 ();
 sg13g2_fill_1 FILLER_38_924 ();
 sg13g2_decap_8 FILLER_39_4 ();
 sg13g2_decap_8 FILLER_39_11 ();
 sg13g2_fill_2 FILLER_39_18 ();
 sg13g2_fill_1 FILLER_39_20 ();
 sg13g2_fill_1 FILLER_39_29 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_decap_8 FILLER_39_77 ();
 sg13g2_decap_8 FILLER_39_84 ();
 sg13g2_decap_8 FILLER_39_91 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_119 ();
 sg13g2_decap_8 FILLER_39_126 ();
 sg13g2_decap_8 FILLER_39_133 ();
 sg13g2_decap_8 FILLER_39_140 ();
 sg13g2_decap_8 FILLER_39_147 ();
 sg13g2_decap_8 FILLER_39_154 ();
 sg13g2_decap_8 FILLER_39_161 ();
 sg13g2_decap_8 FILLER_39_168 ();
 sg13g2_decap_8 FILLER_39_175 ();
 sg13g2_decap_8 FILLER_39_182 ();
 sg13g2_decap_8 FILLER_39_189 ();
 sg13g2_decap_8 FILLER_39_196 ();
 sg13g2_decap_8 FILLER_39_203 ();
 sg13g2_decap_8 FILLER_39_210 ();
 sg13g2_decap_8 FILLER_39_217 ();
 sg13g2_decap_8 FILLER_39_224 ();
 sg13g2_decap_8 FILLER_39_231 ();
 sg13g2_decap_8 FILLER_39_238 ();
 sg13g2_decap_8 FILLER_39_245 ();
 sg13g2_decap_8 FILLER_39_252 ();
 sg13g2_decap_8 FILLER_39_259 ();
 sg13g2_decap_8 FILLER_39_266 ();
 sg13g2_decap_8 FILLER_39_273 ();
 sg13g2_decap_8 FILLER_39_280 ();
 sg13g2_decap_8 FILLER_39_287 ();
 sg13g2_decap_8 FILLER_39_294 ();
 sg13g2_decap_8 FILLER_39_301 ();
 sg13g2_decap_8 FILLER_39_308 ();
 sg13g2_decap_8 FILLER_39_315 ();
 sg13g2_decap_8 FILLER_39_322 ();
 sg13g2_decap_8 FILLER_39_329 ();
 sg13g2_decap_8 FILLER_39_336 ();
 sg13g2_decap_8 FILLER_39_343 ();
 sg13g2_decap_8 FILLER_39_350 ();
 sg13g2_decap_8 FILLER_39_357 ();
 sg13g2_decap_8 FILLER_39_364 ();
 sg13g2_decap_8 FILLER_39_371 ();
 sg13g2_decap_8 FILLER_39_378 ();
 sg13g2_decap_8 FILLER_39_385 ();
 sg13g2_decap_8 FILLER_39_392 ();
 sg13g2_decap_8 FILLER_39_399 ();
 sg13g2_decap_8 FILLER_39_406 ();
 sg13g2_decap_8 FILLER_39_413 ();
 sg13g2_decap_8 FILLER_39_420 ();
 sg13g2_decap_8 FILLER_39_427 ();
 sg13g2_decap_8 FILLER_39_434 ();
 sg13g2_decap_8 FILLER_39_441 ();
 sg13g2_decap_8 FILLER_39_448 ();
 sg13g2_decap_8 FILLER_39_455 ();
 sg13g2_decap_8 FILLER_39_462 ();
 sg13g2_decap_8 FILLER_39_469 ();
 sg13g2_decap_8 FILLER_39_476 ();
 sg13g2_decap_8 FILLER_39_483 ();
 sg13g2_decap_8 FILLER_39_490 ();
 sg13g2_decap_8 FILLER_39_497 ();
 sg13g2_decap_8 FILLER_39_504 ();
 sg13g2_decap_8 FILLER_39_511 ();
 sg13g2_decap_8 FILLER_39_518 ();
 sg13g2_decap_8 FILLER_39_525 ();
 sg13g2_decap_8 FILLER_39_532 ();
 sg13g2_decap_8 FILLER_39_539 ();
 sg13g2_decap_8 FILLER_39_546 ();
 sg13g2_decap_8 FILLER_39_553 ();
 sg13g2_decap_8 FILLER_39_560 ();
 sg13g2_decap_8 FILLER_39_567 ();
 sg13g2_decap_8 FILLER_39_574 ();
 sg13g2_decap_8 FILLER_39_581 ();
 sg13g2_decap_8 FILLER_39_588 ();
 sg13g2_decap_8 FILLER_39_595 ();
 sg13g2_decap_8 FILLER_39_602 ();
 sg13g2_decap_8 FILLER_39_609 ();
 sg13g2_decap_8 FILLER_39_616 ();
 sg13g2_decap_8 FILLER_39_623 ();
 sg13g2_decap_8 FILLER_39_630 ();
 sg13g2_decap_8 FILLER_39_637 ();
 sg13g2_decap_8 FILLER_39_644 ();
 sg13g2_decap_8 FILLER_39_651 ();
 sg13g2_decap_8 FILLER_39_658 ();
 sg13g2_decap_8 FILLER_39_665 ();
 sg13g2_decap_8 FILLER_39_672 ();
 sg13g2_decap_8 FILLER_39_679 ();
 sg13g2_decap_8 FILLER_39_686 ();
 sg13g2_decap_8 FILLER_39_693 ();
 sg13g2_decap_8 FILLER_39_700 ();
 sg13g2_decap_8 FILLER_39_707 ();
 sg13g2_decap_8 FILLER_39_714 ();
 sg13g2_decap_8 FILLER_39_721 ();
 sg13g2_decap_8 FILLER_39_728 ();
 sg13g2_decap_8 FILLER_39_735 ();
 sg13g2_decap_8 FILLER_39_742 ();
 sg13g2_decap_8 FILLER_39_749 ();
 sg13g2_decap_8 FILLER_39_756 ();
 sg13g2_decap_8 FILLER_39_763 ();
 sg13g2_decap_8 FILLER_39_770 ();
 sg13g2_decap_8 FILLER_39_777 ();
 sg13g2_decap_8 FILLER_39_784 ();
 sg13g2_decap_8 FILLER_39_791 ();
 sg13g2_decap_8 FILLER_39_798 ();
 sg13g2_decap_8 FILLER_39_805 ();
 sg13g2_decap_8 FILLER_39_812 ();
 sg13g2_decap_8 FILLER_39_819 ();
 sg13g2_decap_8 FILLER_39_826 ();
 sg13g2_decap_8 FILLER_39_833 ();
 sg13g2_decap_8 FILLER_39_840 ();
 sg13g2_decap_8 FILLER_39_847 ();
 sg13g2_decap_8 FILLER_39_854 ();
 sg13g2_decap_8 FILLER_39_861 ();
 sg13g2_decap_8 FILLER_39_868 ();
 sg13g2_decap_8 FILLER_39_875 ();
 sg13g2_decap_8 FILLER_39_882 ();
 sg13g2_decap_8 FILLER_39_889 ();
 sg13g2_decap_8 FILLER_39_896 ();
 sg13g2_decap_8 FILLER_39_903 ();
 sg13g2_decap_8 FILLER_39_910 ();
 sg13g2_decap_8 FILLER_39_917 ();
 sg13g2_fill_1 FILLER_39_924 ();
 sg13g2_decap_8 FILLER_40_4 ();
 sg13g2_decap_8 FILLER_40_11 ();
 sg13g2_decap_8 FILLER_40_18 ();
 sg13g2_decap_8 FILLER_40_25 ();
 sg13g2_decap_8 FILLER_40_32 ();
 sg13g2_decap_8 FILLER_40_39 ();
 sg13g2_decap_8 FILLER_40_46 ();
 sg13g2_decap_8 FILLER_40_53 ();
 sg13g2_decap_8 FILLER_40_60 ();
 sg13g2_decap_8 FILLER_40_67 ();
 sg13g2_decap_8 FILLER_40_74 ();
 sg13g2_decap_8 FILLER_40_81 ();
 sg13g2_decap_8 FILLER_40_88 ();
 sg13g2_decap_8 FILLER_40_95 ();
 sg13g2_decap_8 FILLER_40_102 ();
 sg13g2_decap_8 FILLER_40_109 ();
 sg13g2_decap_8 FILLER_40_116 ();
 sg13g2_decap_8 FILLER_40_123 ();
 sg13g2_decap_8 FILLER_40_130 ();
 sg13g2_decap_8 FILLER_40_137 ();
 sg13g2_decap_8 FILLER_40_144 ();
 sg13g2_decap_8 FILLER_40_151 ();
 sg13g2_decap_8 FILLER_40_158 ();
 sg13g2_decap_8 FILLER_40_165 ();
 sg13g2_decap_8 FILLER_40_172 ();
 sg13g2_decap_8 FILLER_40_179 ();
 sg13g2_decap_8 FILLER_40_186 ();
 sg13g2_decap_8 FILLER_40_193 ();
 sg13g2_decap_8 FILLER_40_200 ();
 sg13g2_decap_8 FILLER_40_207 ();
 sg13g2_decap_8 FILLER_40_214 ();
 sg13g2_decap_8 FILLER_40_221 ();
 sg13g2_decap_8 FILLER_40_228 ();
 sg13g2_decap_8 FILLER_40_235 ();
 sg13g2_decap_8 FILLER_40_242 ();
 sg13g2_decap_8 FILLER_40_249 ();
 sg13g2_decap_8 FILLER_40_256 ();
 sg13g2_decap_8 FILLER_40_263 ();
 sg13g2_decap_8 FILLER_40_270 ();
 sg13g2_decap_8 FILLER_40_277 ();
 sg13g2_decap_8 FILLER_40_284 ();
 sg13g2_decap_8 FILLER_40_291 ();
 sg13g2_decap_8 FILLER_40_298 ();
 sg13g2_decap_8 FILLER_40_305 ();
 sg13g2_decap_8 FILLER_40_312 ();
 sg13g2_decap_8 FILLER_40_319 ();
 sg13g2_decap_8 FILLER_40_326 ();
 sg13g2_decap_8 FILLER_40_333 ();
 sg13g2_decap_8 FILLER_40_340 ();
 sg13g2_decap_8 FILLER_40_347 ();
 sg13g2_decap_8 FILLER_40_354 ();
 sg13g2_decap_8 FILLER_40_361 ();
 sg13g2_decap_8 FILLER_40_368 ();
 sg13g2_decap_8 FILLER_40_375 ();
 sg13g2_decap_8 FILLER_40_382 ();
 sg13g2_decap_8 FILLER_40_389 ();
 sg13g2_decap_8 FILLER_40_396 ();
 sg13g2_decap_8 FILLER_40_403 ();
 sg13g2_decap_8 FILLER_40_410 ();
 sg13g2_decap_8 FILLER_40_417 ();
 sg13g2_decap_8 FILLER_40_424 ();
 sg13g2_decap_8 FILLER_40_431 ();
 sg13g2_decap_8 FILLER_40_438 ();
 sg13g2_decap_8 FILLER_40_445 ();
 sg13g2_decap_8 FILLER_40_452 ();
 sg13g2_decap_8 FILLER_40_459 ();
 sg13g2_decap_8 FILLER_40_466 ();
 sg13g2_decap_8 FILLER_40_473 ();
 sg13g2_decap_8 FILLER_40_480 ();
 sg13g2_decap_8 FILLER_40_487 ();
 sg13g2_decap_8 FILLER_40_494 ();
 sg13g2_decap_8 FILLER_40_501 ();
 sg13g2_decap_8 FILLER_40_508 ();
 sg13g2_decap_8 FILLER_40_515 ();
 sg13g2_decap_8 FILLER_40_522 ();
 sg13g2_decap_8 FILLER_40_529 ();
 sg13g2_decap_8 FILLER_40_536 ();
 sg13g2_decap_8 FILLER_40_543 ();
 sg13g2_decap_8 FILLER_40_550 ();
 sg13g2_decap_8 FILLER_40_557 ();
 sg13g2_decap_8 FILLER_40_564 ();
 sg13g2_decap_8 FILLER_40_571 ();
 sg13g2_decap_8 FILLER_40_578 ();
 sg13g2_decap_8 FILLER_40_585 ();
 sg13g2_decap_8 FILLER_40_592 ();
 sg13g2_decap_8 FILLER_40_599 ();
 sg13g2_decap_8 FILLER_40_606 ();
 sg13g2_decap_8 FILLER_40_613 ();
 sg13g2_decap_8 FILLER_40_620 ();
 sg13g2_decap_8 FILLER_40_627 ();
 sg13g2_decap_8 FILLER_40_634 ();
 sg13g2_decap_8 FILLER_40_641 ();
 sg13g2_decap_8 FILLER_40_648 ();
 sg13g2_decap_8 FILLER_40_655 ();
 sg13g2_decap_8 FILLER_40_662 ();
 sg13g2_decap_8 FILLER_40_669 ();
 sg13g2_decap_8 FILLER_40_676 ();
 sg13g2_decap_8 FILLER_40_683 ();
 sg13g2_decap_8 FILLER_40_690 ();
 sg13g2_decap_8 FILLER_40_697 ();
 sg13g2_decap_8 FILLER_40_704 ();
 sg13g2_decap_8 FILLER_40_711 ();
 sg13g2_decap_8 FILLER_40_718 ();
 sg13g2_decap_8 FILLER_40_725 ();
 sg13g2_decap_8 FILLER_40_732 ();
 sg13g2_decap_8 FILLER_40_739 ();
 sg13g2_decap_8 FILLER_40_746 ();
 sg13g2_decap_8 FILLER_40_753 ();
 sg13g2_decap_8 FILLER_40_760 ();
 sg13g2_decap_8 FILLER_40_767 ();
 sg13g2_decap_8 FILLER_40_774 ();
 sg13g2_decap_8 FILLER_40_781 ();
 sg13g2_decap_8 FILLER_40_788 ();
 sg13g2_decap_8 FILLER_40_795 ();
 sg13g2_decap_8 FILLER_40_802 ();
 sg13g2_decap_8 FILLER_40_809 ();
 sg13g2_decap_8 FILLER_40_816 ();
 sg13g2_decap_8 FILLER_40_823 ();
 sg13g2_decap_8 FILLER_40_830 ();
 sg13g2_decap_8 FILLER_40_837 ();
 sg13g2_decap_8 FILLER_40_844 ();
 sg13g2_decap_8 FILLER_40_851 ();
 sg13g2_decap_8 FILLER_40_858 ();
 sg13g2_decap_8 FILLER_40_865 ();
 sg13g2_decap_8 FILLER_40_872 ();
 sg13g2_decap_8 FILLER_40_879 ();
 sg13g2_decap_8 FILLER_40_886 ();
 sg13g2_decap_8 FILLER_40_893 ();
 sg13g2_decap_8 FILLER_40_900 ();
 sg13g2_decap_8 FILLER_40_907 ();
 sg13g2_decap_8 FILLER_40_914 ();
 sg13g2_decap_4 FILLER_40_921 ();
 sg13g2_decap_8 FILLER_41_4 ();
 sg13g2_decap_8 FILLER_41_11 ();
 sg13g2_decap_8 FILLER_41_18 ();
 sg13g2_decap_8 FILLER_41_25 ();
 sg13g2_decap_4 FILLER_41_32 ();
 sg13g2_decap_8 FILLER_41_44 ();
 sg13g2_decap_8 FILLER_41_51 ();
 sg13g2_decap_8 FILLER_41_58 ();
 sg13g2_decap_8 FILLER_41_65 ();
 sg13g2_decap_8 FILLER_41_72 ();
 sg13g2_decap_8 FILLER_41_79 ();
 sg13g2_decap_8 FILLER_41_86 ();
 sg13g2_decap_8 FILLER_41_93 ();
 sg13g2_decap_8 FILLER_41_100 ();
 sg13g2_decap_8 FILLER_41_107 ();
 sg13g2_decap_8 FILLER_41_114 ();
 sg13g2_decap_8 FILLER_41_121 ();
 sg13g2_decap_8 FILLER_41_128 ();
 sg13g2_decap_8 FILLER_41_135 ();
 sg13g2_decap_8 FILLER_41_142 ();
 sg13g2_decap_8 FILLER_41_149 ();
 sg13g2_decap_8 FILLER_41_156 ();
 sg13g2_decap_8 FILLER_41_163 ();
 sg13g2_decap_8 FILLER_41_170 ();
 sg13g2_decap_8 FILLER_41_177 ();
 sg13g2_decap_8 FILLER_41_184 ();
 sg13g2_decap_8 FILLER_41_191 ();
 sg13g2_decap_8 FILLER_41_198 ();
 sg13g2_decap_8 FILLER_41_205 ();
 sg13g2_decap_8 FILLER_41_212 ();
 sg13g2_decap_8 FILLER_41_219 ();
 sg13g2_decap_8 FILLER_41_226 ();
 sg13g2_decap_8 FILLER_41_233 ();
 sg13g2_decap_8 FILLER_41_240 ();
 sg13g2_decap_8 FILLER_41_247 ();
 sg13g2_decap_8 FILLER_41_254 ();
 sg13g2_decap_8 FILLER_41_261 ();
 sg13g2_decap_8 FILLER_41_268 ();
 sg13g2_decap_8 FILLER_41_275 ();
 sg13g2_decap_8 FILLER_41_282 ();
 sg13g2_decap_8 FILLER_41_289 ();
 sg13g2_decap_8 FILLER_41_296 ();
 sg13g2_decap_8 FILLER_41_303 ();
 sg13g2_decap_8 FILLER_41_310 ();
 sg13g2_decap_8 FILLER_41_317 ();
 sg13g2_decap_8 FILLER_41_324 ();
 sg13g2_decap_8 FILLER_41_331 ();
 sg13g2_decap_8 FILLER_41_338 ();
 sg13g2_decap_8 FILLER_41_345 ();
 sg13g2_decap_8 FILLER_41_352 ();
 sg13g2_decap_8 FILLER_41_359 ();
 sg13g2_decap_8 FILLER_41_366 ();
 sg13g2_decap_8 FILLER_41_373 ();
 sg13g2_decap_8 FILLER_41_380 ();
 sg13g2_decap_8 FILLER_41_387 ();
 sg13g2_decap_8 FILLER_41_394 ();
 sg13g2_decap_8 FILLER_41_401 ();
 sg13g2_decap_8 FILLER_41_408 ();
 sg13g2_decap_8 FILLER_41_415 ();
 sg13g2_decap_8 FILLER_41_422 ();
 sg13g2_decap_8 FILLER_41_429 ();
 sg13g2_decap_8 FILLER_41_436 ();
 sg13g2_decap_8 FILLER_41_443 ();
 sg13g2_decap_8 FILLER_41_450 ();
 sg13g2_decap_8 FILLER_41_457 ();
 sg13g2_decap_8 FILLER_41_464 ();
 sg13g2_decap_8 FILLER_41_471 ();
 sg13g2_decap_8 FILLER_41_478 ();
 sg13g2_decap_8 FILLER_41_485 ();
 sg13g2_decap_8 FILLER_41_492 ();
 sg13g2_decap_8 FILLER_41_499 ();
 sg13g2_decap_8 FILLER_41_506 ();
 sg13g2_decap_8 FILLER_41_513 ();
 sg13g2_decap_8 FILLER_41_520 ();
 sg13g2_decap_8 FILLER_41_527 ();
 sg13g2_decap_8 FILLER_41_534 ();
 sg13g2_decap_8 FILLER_41_541 ();
 sg13g2_decap_8 FILLER_41_548 ();
 sg13g2_decap_8 FILLER_41_555 ();
 sg13g2_decap_8 FILLER_41_562 ();
 sg13g2_decap_8 FILLER_41_569 ();
 sg13g2_decap_8 FILLER_41_576 ();
 sg13g2_decap_8 FILLER_41_583 ();
 sg13g2_decap_8 FILLER_41_590 ();
 sg13g2_decap_8 FILLER_41_597 ();
 sg13g2_decap_8 FILLER_41_604 ();
 sg13g2_decap_8 FILLER_41_611 ();
 sg13g2_decap_8 FILLER_41_618 ();
 sg13g2_decap_8 FILLER_41_625 ();
 sg13g2_decap_8 FILLER_41_632 ();
 sg13g2_decap_8 FILLER_41_639 ();
 sg13g2_decap_8 FILLER_41_646 ();
 sg13g2_decap_8 FILLER_41_653 ();
 sg13g2_decap_8 FILLER_41_660 ();
 sg13g2_decap_8 FILLER_41_667 ();
 sg13g2_decap_8 FILLER_41_674 ();
 sg13g2_decap_8 FILLER_41_681 ();
 sg13g2_decap_8 FILLER_41_688 ();
 sg13g2_decap_8 FILLER_41_695 ();
 sg13g2_decap_8 FILLER_41_702 ();
 sg13g2_decap_8 FILLER_41_709 ();
 sg13g2_decap_8 FILLER_41_716 ();
 sg13g2_decap_8 FILLER_41_723 ();
 sg13g2_decap_8 FILLER_41_730 ();
 sg13g2_decap_8 FILLER_41_737 ();
 sg13g2_decap_8 FILLER_41_744 ();
 sg13g2_decap_8 FILLER_41_751 ();
 sg13g2_decap_8 FILLER_41_758 ();
 sg13g2_decap_8 FILLER_41_765 ();
 sg13g2_decap_8 FILLER_41_772 ();
 sg13g2_decap_8 FILLER_41_779 ();
 sg13g2_decap_8 FILLER_41_786 ();
 sg13g2_decap_8 FILLER_41_793 ();
 sg13g2_decap_8 FILLER_41_800 ();
 sg13g2_decap_8 FILLER_41_807 ();
 sg13g2_decap_8 FILLER_41_814 ();
 sg13g2_decap_8 FILLER_41_821 ();
 sg13g2_decap_8 FILLER_41_828 ();
 sg13g2_decap_8 FILLER_41_835 ();
 sg13g2_decap_8 FILLER_41_842 ();
 sg13g2_decap_8 FILLER_41_849 ();
 sg13g2_decap_8 FILLER_41_856 ();
 sg13g2_decap_8 FILLER_41_863 ();
 sg13g2_decap_8 FILLER_41_870 ();
 sg13g2_decap_8 FILLER_41_877 ();
 sg13g2_decap_8 FILLER_41_884 ();
 sg13g2_decap_8 FILLER_41_891 ();
 sg13g2_decap_8 FILLER_41_898 ();
 sg13g2_decap_8 FILLER_41_905 ();
 sg13g2_decap_8 FILLER_41_912 ();
 sg13g2_decap_4 FILLER_41_919 ();
 sg13g2_fill_2 FILLER_41_923 ();
 sg13g2_decap_8 FILLER_42_4 ();
 sg13g2_decap_8 FILLER_42_11 ();
 sg13g2_decap_8 FILLER_42_18 ();
 sg13g2_decap_8 FILLER_42_25 ();
 sg13g2_fill_2 FILLER_42_32 ();
 sg13g2_fill_1 FILLER_42_34 ();
 sg13g2_decap_8 FILLER_42_43 ();
 sg13g2_decap_8 FILLER_42_50 ();
 sg13g2_decap_8 FILLER_42_57 ();
 sg13g2_decap_8 FILLER_42_64 ();
 sg13g2_decap_8 FILLER_42_71 ();
 sg13g2_decap_8 FILLER_42_78 ();
 sg13g2_decap_8 FILLER_42_85 ();
 sg13g2_decap_8 FILLER_42_92 ();
 sg13g2_decap_8 FILLER_42_99 ();
 sg13g2_decap_8 FILLER_42_106 ();
 sg13g2_decap_8 FILLER_42_113 ();
 sg13g2_decap_8 FILLER_42_120 ();
 sg13g2_decap_8 FILLER_42_127 ();
 sg13g2_decap_8 FILLER_42_134 ();
 sg13g2_decap_8 FILLER_42_141 ();
 sg13g2_decap_8 FILLER_42_148 ();
 sg13g2_decap_8 FILLER_42_155 ();
 sg13g2_decap_8 FILLER_42_162 ();
 sg13g2_decap_8 FILLER_42_169 ();
 sg13g2_decap_8 FILLER_42_176 ();
 sg13g2_decap_8 FILLER_42_183 ();
 sg13g2_decap_8 FILLER_42_190 ();
 sg13g2_decap_8 FILLER_42_197 ();
 sg13g2_decap_8 FILLER_42_204 ();
 sg13g2_decap_8 FILLER_42_211 ();
 sg13g2_decap_8 FILLER_42_218 ();
 sg13g2_decap_8 FILLER_42_225 ();
 sg13g2_decap_8 FILLER_42_232 ();
 sg13g2_decap_8 FILLER_42_239 ();
 sg13g2_decap_8 FILLER_42_246 ();
 sg13g2_decap_8 FILLER_42_253 ();
 sg13g2_decap_8 FILLER_42_260 ();
 sg13g2_decap_8 FILLER_42_267 ();
 sg13g2_decap_8 FILLER_42_274 ();
 sg13g2_decap_8 FILLER_42_281 ();
 sg13g2_decap_8 FILLER_42_288 ();
 sg13g2_decap_8 FILLER_42_295 ();
 sg13g2_decap_8 FILLER_42_302 ();
 sg13g2_decap_8 FILLER_42_309 ();
 sg13g2_decap_8 FILLER_42_316 ();
 sg13g2_decap_8 FILLER_42_323 ();
 sg13g2_decap_8 FILLER_42_330 ();
 sg13g2_decap_8 FILLER_42_337 ();
 sg13g2_decap_8 FILLER_42_344 ();
 sg13g2_decap_8 FILLER_42_351 ();
 sg13g2_decap_8 FILLER_42_358 ();
 sg13g2_decap_8 FILLER_42_365 ();
 sg13g2_decap_8 FILLER_42_372 ();
 sg13g2_decap_8 FILLER_42_379 ();
 sg13g2_decap_8 FILLER_42_386 ();
 sg13g2_decap_8 FILLER_42_393 ();
 sg13g2_decap_8 FILLER_42_400 ();
 sg13g2_decap_8 FILLER_42_407 ();
 sg13g2_decap_8 FILLER_42_414 ();
 sg13g2_decap_8 FILLER_42_421 ();
 sg13g2_decap_8 FILLER_42_428 ();
 sg13g2_decap_8 FILLER_42_435 ();
 sg13g2_decap_8 FILLER_42_442 ();
 sg13g2_decap_8 FILLER_42_449 ();
 sg13g2_decap_8 FILLER_42_456 ();
 sg13g2_decap_8 FILLER_42_463 ();
 sg13g2_decap_8 FILLER_42_470 ();
 sg13g2_decap_8 FILLER_42_477 ();
 sg13g2_decap_8 FILLER_42_484 ();
 sg13g2_decap_8 FILLER_42_491 ();
 sg13g2_decap_8 FILLER_42_498 ();
 sg13g2_decap_8 FILLER_42_505 ();
 sg13g2_decap_8 FILLER_42_512 ();
 sg13g2_decap_8 FILLER_42_519 ();
 sg13g2_decap_8 FILLER_42_526 ();
 sg13g2_decap_8 FILLER_42_533 ();
 sg13g2_decap_8 FILLER_42_540 ();
 sg13g2_decap_8 FILLER_42_547 ();
 sg13g2_decap_8 FILLER_42_554 ();
 sg13g2_decap_8 FILLER_42_561 ();
 sg13g2_decap_8 FILLER_42_568 ();
 sg13g2_decap_8 FILLER_42_575 ();
 sg13g2_decap_8 FILLER_42_582 ();
 sg13g2_decap_8 FILLER_42_589 ();
 sg13g2_decap_8 FILLER_42_596 ();
 sg13g2_decap_8 FILLER_42_603 ();
 sg13g2_decap_8 FILLER_42_610 ();
 sg13g2_decap_8 FILLER_42_617 ();
 sg13g2_decap_8 FILLER_42_624 ();
 sg13g2_decap_8 FILLER_42_631 ();
 sg13g2_decap_8 FILLER_42_638 ();
 sg13g2_decap_8 FILLER_42_645 ();
 sg13g2_decap_8 FILLER_42_652 ();
 sg13g2_decap_8 FILLER_42_659 ();
 sg13g2_decap_8 FILLER_42_666 ();
 sg13g2_decap_8 FILLER_42_673 ();
 sg13g2_decap_8 FILLER_42_680 ();
 sg13g2_decap_8 FILLER_42_687 ();
 sg13g2_decap_8 FILLER_42_694 ();
 sg13g2_decap_8 FILLER_42_701 ();
 sg13g2_decap_8 FILLER_42_708 ();
 sg13g2_decap_8 FILLER_42_715 ();
 sg13g2_decap_8 FILLER_42_722 ();
 sg13g2_decap_8 FILLER_42_729 ();
 sg13g2_decap_8 FILLER_42_736 ();
 sg13g2_decap_8 FILLER_42_743 ();
 sg13g2_decap_8 FILLER_42_750 ();
 sg13g2_decap_8 FILLER_42_757 ();
 sg13g2_decap_8 FILLER_42_764 ();
 sg13g2_decap_8 FILLER_42_771 ();
 sg13g2_decap_8 FILLER_42_778 ();
 sg13g2_decap_8 FILLER_42_785 ();
 sg13g2_decap_8 FILLER_42_792 ();
 sg13g2_decap_8 FILLER_42_799 ();
 sg13g2_decap_8 FILLER_42_806 ();
 sg13g2_decap_8 FILLER_42_813 ();
 sg13g2_decap_8 FILLER_42_820 ();
 sg13g2_decap_8 FILLER_42_827 ();
 sg13g2_decap_8 FILLER_42_834 ();
 sg13g2_decap_8 FILLER_42_841 ();
 sg13g2_decap_8 FILLER_42_848 ();
 sg13g2_decap_8 FILLER_42_855 ();
 sg13g2_decap_8 FILLER_42_862 ();
 sg13g2_decap_8 FILLER_42_869 ();
 sg13g2_decap_8 FILLER_42_876 ();
 sg13g2_decap_8 FILLER_42_883 ();
 sg13g2_decap_8 FILLER_42_890 ();
 sg13g2_decap_8 FILLER_42_897 ();
 sg13g2_decap_8 FILLER_42_904 ();
 sg13g2_decap_8 FILLER_42_911 ();
 sg13g2_decap_8 FILLER_42_918 ();
 sg13g2_decap_8 FILLER_43_4 ();
 sg13g2_decap_8 FILLER_43_11 ();
 sg13g2_decap_8 FILLER_43_18 ();
 sg13g2_decap_8 FILLER_43_25 ();
 sg13g2_decap_8 FILLER_43_32 ();
 sg13g2_decap_8 FILLER_43_39 ();
 sg13g2_decap_8 FILLER_43_46 ();
 sg13g2_decap_8 FILLER_43_53 ();
 sg13g2_decap_8 FILLER_43_60 ();
 sg13g2_decap_8 FILLER_43_67 ();
 sg13g2_decap_8 FILLER_43_74 ();
 sg13g2_decap_8 FILLER_43_81 ();
 sg13g2_decap_8 FILLER_43_88 ();
 sg13g2_decap_8 FILLER_43_95 ();
 sg13g2_decap_8 FILLER_43_102 ();
 sg13g2_decap_8 FILLER_43_109 ();
 sg13g2_decap_8 FILLER_43_116 ();
 sg13g2_decap_8 FILLER_43_123 ();
 sg13g2_decap_8 FILLER_43_130 ();
 sg13g2_decap_8 FILLER_43_137 ();
 sg13g2_decap_8 FILLER_43_144 ();
 sg13g2_decap_8 FILLER_43_151 ();
 sg13g2_decap_8 FILLER_43_158 ();
 sg13g2_decap_8 FILLER_43_165 ();
 sg13g2_decap_8 FILLER_43_172 ();
 sg13g2_decap_8 FILLER_43_179 ();
 sg13g2_decap_8 FILLER_43_186 ();
 sg13g2_decap_8 FILLER_43_193 ();
 sg13g2_decap_8 FILLER_43_200 ();
 sg13g2_decap_8 FILLER_43_207 ();
 sg13g2_decap_8 FILLER_43_214 ();
 sg13g2_decap_8 FILLER_43_221 ();
 sg13g2_decap_8 FILLER_43_228 ();
 sg13g2_decap_8 FILLER_43_235 ();
 sg13g2_decap_8 FILLER_43_242 ();
 sg13g2_decap_8 FILLER_43_249 ();
 sg13g2_decap_8 FILLER_43_256 ();
 sg13g2_decap_8 FILLER_43_263 ();
 sg13g2_decap_8 FILLER_43_270 ();
 sg13g2_decap_8 FILLER_43_277 ();
 sg13g2_decap_8 FILLER_43_284 ();
 sg13g2_decap_8 FILLER_43_291 ();
 sg13g2_decap_8 FILLER_43_298 ();
 sg13g2_decap_8 FILLER_43_305 ();
 sg13g2_decap_8 FILLER_43_312 ();
 sg13g2_decap_8 FILLER_43_319 ();
 sg13g2_decap_8 FILLER_43_326 ();
 sg13g2_decap_8 FILLER_43_333 ();
 sg13g2_decap_8 FILLER_43_340 ();
 sg13g2_decap_8 FILLER_43_347 ();
 sg13g2_decap_8 FILLER_43_354 ();
 sg13g2_decap_8 FILLER_43_361 ();
 sg13g2_decap_8 FILLER_43_368 ();
 sg13g2_decap_8 FILLER_43_375 ();
 sg13g2_decap_8 FILLER_43_382 ();
 sg13g2_decap_8 FILLER_43_389 ();
 sg13g2_decap_8 FILLER_43_396 ();
 sg13g2_decap_8 FILLER_43_403 ();
 sg13g2_decap_8 FILLER_43_410 ();
 sg13g2_decap_8 FILLER_43_417 ();
 sg13g2_decap_8 FILLER_43_424 ();
 sg13g2_decap_8 FILLER_43_431 ();
 sg13g2_decap_8 FILLER_43_438 ();
 sg13g2_decap_8 FILLER_43_445 ();
 sg13g2_decap_8 FILLER_43_452 ();
 sg13g2_decap_8 FILLER_43_459 ();
 sg13g2_decap_8 FILLER_43_466 ();
 sg13g2_decap_8 FILLER_43_473 ();
 sg13g2_decap_8 FILLER_43_480 ();
 sg13g2_decap_8 FILLER_43_487 ();
 sg13g2_decap_8 FILLER_43_494 ();
 sg13g2_decap_8 FILLER_43_501 ();
 sg13g2_decap_8 FILLER_43_508 ();
 sg13g2_decap_8 FILLER_43_515 ();
 sg13g2_decap_8 FILLER_43_522 ();
 sg13g2_decap_8 FILLER_43_529 ();
 sg13g2_decap_8 FILLER_43_536 ();
 sg13g2_decap_8 FILLER_43_543 ();
 sg13g2_decap_8 FILLER_43_550 ();
 sg13g2_decap_8 FILLER_43_557 ();
 sg13g2_decap_8 FILLER_43_564 ();
 sg13g2_decap_8 FILLER_43_571 ();
 sg13g2_decap_8 FILLER_43_578 ();
 sg13g2_decap_8 FILLER_43_585 ();
 sg13g2_decap_8 FILLER_43_592 ();
 sg13g2_decap_8 FILLER_43_599 ();
 sg13g2_decap_8 FILLER_43_606 ();
 sg13g2_decap_8 FILLER_43_613 ();
 sg13g2_decap_8 FILLER_43_620 ();
 sg13g2_decap_8 FILLER_43_627 ();
 sg13g2_decap_8 FILLER_43_634 ();
 sg13g2_decap_8 FILLER_43_641 ();
 sg13g2_decap_8 FILLER_43_648 ();
 sg13g2_decap_8 FILLER_43_655 ();
 sg13g2_decap_8 FILLER_43_662 ();
 sg13g2_decap_8 FILLER_43_669 ();
 sg13g2_decap_8 FILLER_43_676 ();
 sg13g2_decap_8 FILLER_43_683 ();
 sg13g2_decap_8 FILLER_43_690 ();
 sg13g2_decap_8 FILLER_43_697 ();
 sg13g2_decap_8 FILLER_43_704 ();
 sg13g2_decap_8 FILLER_43_711 ();
 sg13g2_decap_8 FILLER_43_718 ();
 sg13g2_decap_8 FILLER_43_725 ();
 sg13g2_decap_8 FILLER_43_732 ();
 sg13g2_decap_8 FILLER_43_739 ();
 sg13g2_decap_8 FILLER_43_746 ();
 sg13g2_decap_8 FILLER_43_753 ();
 sg13g2_decap_8 FILLER_43_760 ();
 sg13g2_decap_8 FILLER_43_767 ();
 sg13g2_decap_8 FILLER_43_774 ();
 sg13g2_decap_8 FILLER_43_781 ();
 sg13g2_decap_8 FILLER_43_788 ();
 sg13g2_decap_8 FILLER_43_795 ();
 sg13g2_decap_8 FILLER_43_802 ();
 sg13g2_decap_8 FILLER_43_809 ();
 sg13g2_decap_8 FILLER_43_816 ();
 sg13g2_decap_8 FILLER_43_823 ();
 sg13g2_decap_8 FILLER_43_830 ();
 sg13g2_decap_8 FILLER_43_837 ();
 sg13g2_decap_8 FILLER_43_844 ();
 sg13g2_decap_8 FILLER_43_851 ();
 sg13g2_decap_8 FILLER_43_858 ();
 sg13g2_decap_8 FILLER_43_865 ();
 sg13g2_decap_8 FILLER_43_872 ();
 sg13g2_decap_8 FILLER_43_879 ();
 sg13g2_decap_8 FILLER_43_886 ();
 sg13g2_decap_8 FILLER_43_893 ();
 sg13g2_decap_8 FILLER_43_900 ();
 sg13g2_decap_8 FILLER_43_907 ();
 sg13g2_decap_8 FILLER_43_914 ();
 sg13g2_decap_4 FILLER_43_921 ();
 sg13g2_decap_8 FILLER_44_4 ();
 sg13g2_decap_8 FILLER_44_11 ();
 sg13g2_decap_8 FILLER_44_18 ();
 sg13g2_decap_8 FILLER_44_25 ();
 sg13g2_decap_8 FILLER_44_32 ();
 sg13g2_decap_8 FILLER_44_39 ();
 sg13g2_decap_8 FILLER_44_46 ();
 sg13g2_decap_8 FILLER_44_53 ();
 sg13g2_decap_8 FILLER_44_60 ();
 sg13g2_decap_8 FILLER_44_67 ();
 sg13g2_decap_8 FILLER_44_74 ();
 sg13g2_decap_8 FILLER_44_81 ();
 sg13g2_decap_8 FILLER_44_88 ();
 sg13g2_decap_8 FILLER_44_95 ();
 sg13g2_decap_8 FILLER_44_102 ();
 sg13g2_decap_8 FILLER_44_109 ();
 sg13g2_decap_8 FILLER_44_116 ();
 sg13g2_decap_8 FILLER_44_123 ();
 sg13g2_decap_8 FILLER_44_130 ();
 sg13g2_decap_8 FILLER_44_137 ();
 sg13g2_decap_8 FILLER_44_144 ();
 sg13g2_decap_8 FILLER_44_151 ();
 sg13g2_decap_8 FILLER_44_158 ();
 sg13g2_decap_8 FILLER_44_165 ();
 sg13g2_decap_8 FILLER_44_172 ();
 sg13g2_decap_8 FILLER_44_179 ();
 sg13g2_decap_8 FILLER_44_186 ();
 sg13g2_decap_8 FILLER_44_193 ();
 sg13g2_decap_8 FILLER_44_200 ();
 sg13g2_decap_8 FILLER_44_207 ();
 sg13g2_decap_8 FILLER_44_214 ();
 sg13g2_decap_8 FILLER_44_221 ();
 sg13g2_decap_8 FILLER_44_228 ();
 sg13g2_decap_8 FILLER_44_235 ();
 sg13g2_decap_8 FILLER_44_242 ();
 sg13g2_decap_8 FILLER_44_249 ();
 sg13g2_decap_8 FILLER_44_256 ();
 sg13g2_decap_8 FILLER_44_263 ();
 sg13g2_decap_8 FILLER_44_270 ();
 sg13g2_decap_8 FILLER_44_277 ();
 sg13g2_decap_8 FILLER_44_284 ();
 sg13g2_decap_8 FILLER_44_291 ();
 sg13g2_decap_8 FILLER_44_298 ();
 sg13g2_decap_8 FILLER_44_305 ();
 sg13g2_decap_8 FILLER_44_312 ();
 sg13g2_decap_8 FILLER_44_319 ();
 sg13g2_decap_8 FILLER_44_326 ();
 sg13g2_decap_8 FILLER_44_333 ();
 sg13g2_decap_8 FILLER_44_340 ();
 sg13g2_decap_8 FILLER_44_347 ();
 sg13g2_decap_8 FILLER_44_354 ();
 sg13g2_decap_8 FILLER_44_361 ();
 sg13g2_decap_8 FILLER_44_368 ();
 sg13g2_decap_8 FILLER_44_375 ();
 sg13g2_decap_8 FILLER_44_382 ();
 sg13g2_decap_8 FILLER_44_389 ();
 sg13g2_decap_8 FILLER_44_396 ();
 sg13g2_decap_8 FILLER_44_403 ();
 sg13g2_decap_8 FILLER_44_410 ();
 sg13g2_decap_8 FILLER_44_417 ();
 sg13g2_decap_8 FILLER_44_424 ();
 sg13g2_decap_8 FILLER_44_431 ();
 sg13g2_decap_8 FILLER_44_438 ();
 sg13g2_decap_8 FILLER_44_445 ();
 sg13g2_decap_8 FILLER_44_452 ();
 sg13g2_decap_8 FILLER_44_459 ();
 sg13g2_decap_8 FILLER_44_466 ();
 sg13g2_decap_8 FILLER_44_473 ();
 sg13g2_decap_8 FILLER_44_480 ();
 sg13g2_decap_8 FILLER_44_487 ();
 sg13g2_decap_8 FILLER_44_494 ();
 sg13g2_decap_8 FILLER_44_501 ();
 sg13g2_decap_8 FILLER_44_508 ();
 sg13g2_decap_8 FILLER_44_515 ();
 sg13g2_decap_8 FILLER_44_522 ();
 sg13g2_decap_8 FILLER_44_529 ();
 sg13g2_decap_8 FILLER_44_536 ();
 sg13g2_decap_8 FILLER_44_543 ();
 sg13g2_decap_8 FILLER_44_550 ();
 sg13g2_decap_8 FILLER_44_557 ();
 sg13g2_decap_8 FILLER_44_564 ();
 sg13g2_decap_8 FILLER_44_571 ();
 sg13g2_decap_8 FILLER_44_578 ();
 sg13g2_decap_8 FILLER_44_585 ();
 sg13g2_decap_8 FILLER_44_592 ();
 sg13g2_decap_8 FILLER_44_599 ();
 sg13g2_decap_8 FILLER_44_606 ();
 sg13g2_decap_8 FILLER_44_613 ();
 sg13g2_decap_8 FILLER_44_620 ();
 sg13g2_decap_8 FILLER_44_627 ();
 sg13g2_decap_8 FILLER_44_634 ();
 sg13g2_decap_8 FILLER_44_641 ();
 sg13g2_decap_8 FILLER_44_648 ();
 sg13g2_decap_8 FILLER_44_655 ();
 sg13g2_decap_8 FILLER_44_662 ();
 sg13g2_decap_8 FILLER_44_669 ();
 sg13g2_decap_8 FILLER_44_676 ();
 sg13g2_decap_8 FILLER_44_683 ();
 sg13g2_decap_8 FILLER_44_690 ();
 sg13g2_decap_8 FILLER_44_697 ();
 sg13g2_decap_8 FILLER_44_704 ();
 sg13g2_decap_8 FILLER_44_711 ();
 sg13g2_decap_8 FILLER_44_718 ();
 sg13g2_decap_8 FILLER_44_725 ();
 sg13g2_decap_8 FILLER_44_732 ();
 sg13g2_decap_8 FILLER_44_739 ();
 sg13g2_decap_8 FILLER_44_746 ();
 sg13g2_decap_8 FILLER_44_753 ();
 sg13g2_decap_8 FILLER_44_760 ();
 sg13g2_decap_8 FILLER_44_767 ();
 sg13g2_decap_8 FILLER_44_774 ();
 sg13g2_decap_8 FILLER_44_781 ();
 sg13g2_decap_8 FILLER_44_788 ();
 sg13g2_decap_8 FILLER_44_795 ();
 sg13g2_decap_8 FILLER_44_802 ();
 sg13g2_decap_8 FILLER_44_809 ();
 sg13g2_decap_8 FILLER_44_816 ();
 sg13g2_decap_8 FILLER_44_823 ();
 sg13g2_decap_8 FILLER_44_830 ();
 sg13g2_decap_8 FILLER_44_837 ();
 sg13g2_decap_8 FILLER_44_844 ();
 sg13g2_decap_8 FILLER_44_851 ();
 sg13g2_decap_8 FILLER_44_858 ();
 sg13g2_decap_8 FILLER_44_865 ();
 sg13g2_decap_8 FILLER_44_872 ();
 sg13g2_decap_8 FILLER_44_879 ();
 sg13g2_decap_8 FILLER_44_886 ();
 sg13g2_decap_8 FILLER_44_893 ();
 sg13g2_decap_8 FILLER_44_900 ();
 sg13g2_decap_8 FILLER_44_907 ();
 sg13g2_decap_8 FILLER_44_914 ();
 sg13g2_decap_4 FILLER_44_921 ();
 sg13g2_decap_8 FILLER_45_4 ();
 sg13g2_decap_8 FILLER_45_11 ();
 sg13g2_decap_8 FILLER_45_18 ();
 sg13g2_decap_8 FILLER_45_25 ();
 sg13g2_decap_8 FILLER_45_32 ();
 sg13g2_decap_8 FILLER_45_39 ();
 sg13g2_decap_8 FILLER_45_46 ();
 sg13g2_decap_8 FILLER_45_53 ();
 sg13g2_decap_8 FILLER_45_60 ();
 sg13g2_decap_8 FILLER_45_67 ();
 sg13g2_decap_8 FILLER_45_74 ();
 sg13g2_decap_8 FILLER_45_81 ();
 sg13g2_decap_8 FILLER_45_88 ();
 sg13g2_decap_8 FILLER_45_95 ();
 sg13g2_decap_8 FILLER_45_102 ();
 sg13g2_decap_8 FILLER_45_109 ();
 sg13g2_decap_8 FILLER_45_116 ();
 sg13g2_decap_8 FILLER_45_123 ();
 sg13g2_decap_8 FILLER_45_130 ();
 sg13g2_decap_8 FILLER_45_137 ();
 sg13g2_decap_8 FILLER_45_144 ();
 sg13g2_decap_8 FILLER_45_151 ();
 sg13g2_decap_8 FILLER_45_158 ();
 sg13g2_decap_8 FILLER_45_165 ();
 sg13g2_decap_8 FILLER_45_172 ();
 sg13g2_decap_8 FILLER_45_179 ();
 sg13g2_decap_8 FILLER_45_186 ();
 sg13g2_decap_8 FILLER_45_193 ();
 sg13g2_decap_8 FILLER_45_200 ();
 sg13g2_decap_8 FILLER_45_207 ();
 sg13g2_decap_8 FILLER_45_214 ();
 sg13g2_decap_8 FILLER_45_221 ();
 sg13g2_decap_8 FILLER_45_228 ();
 sg13g2_decap_8 FILLER_45_235 ();
 sg13g2_decap_8 FILLER_45_242 ();
 sg13g2_decap_8 FILLER_45_249 ();
 sg13g2_decap_8 FILLER_45_256 ();
 sg13g2_decap_8 FILLER_45_263 ();
 sg13g2_decap_8 FILLER_45_270 ();
 sg13g2_decap_8 FILLER_45_277 ();
 sg13g2_decap_8 FILLER_45_284 ();
 sg13g2_decap_8 FILLER_45_291 ();
 sg13g2_decap_8 FILLER_45_298 ();
 sg13g2_decap_8 FILLER_45_305 ();
 sg13g2_decap_8 FILLER_45_312 ();
 sg13g2_decap_8 FILLER_45_319 ();
 sg13g2_decap_8 FILLER_45_326 ();
 sg13g2_decap_8 FILLER_45_333 ();
 sg13g2_decap_8 FILLER_45_340 ();
 sg13g2_decap_8 FILLER_45_347 ();
 sg13g2_decap_8 FILLER_45_354 ();
 sg13g2_decap_8 FILLER_45_361 ();
 sg13g2_decap_8 FILLER_45_368 ();
 sg13g2_decap_8 FILLER_45_375 ();
 sg13g2_decap_8 FILLER_45_382 ();
 sg13g2_decap_8 FILLER_45_389 ();
 sg13g2_decap_8 FILLER_45_396 ();
 sg13g2_decap_8 FILLER_45_403 ();
 sg13g2_decap_8 FILLER_45_410 ();
 sg13g2_decap_8 FILLER_45_417 ();
 sg13g2_decap_8 FILLER_45_424 ();
 sg13g2_decap_8 FILLER_45_431 ();
 sg13g2_decap_8 FILLER_45_438 ();
 sg13g2_decap_8 FILLER_45_445 ();
 sg13g2_decap_8 FILLER_45_452 ();
 sg13g2_decap_8 FILLER_45_459 ();
 sg13g2_decap_8 FILLER_45_466 ();
 sg13g2_decap_8 FILLER_45_473 ();
 sg13g2_decap_8 FILLER_45_480 ();
 sg13g2_decap_8 FILLER_45_487 ();
 sg13g2_decap_8 FILLER_45_494 ();
 sg13g2_decap_8 FILLER_45_501 ();
 sg13g2_decap_8 FILLER_45_508 ();
 sg13g2_decap_8 FILLER_45_515 ();
 sg13g2_decap_8 FILLER_45_522 ();
 sg13g2_decap_8 FILLER_45_529 ();
 sg13g2_decap_8 FILLER_45_536 ();
 sg13g2_decap_8 FILLER_45_543 ();
 sg13g2_decap_8 FILLER_45_550 ();
 sg13g2_decap_8 FILLER_45_557 ();
 sg13g2_decap_8 FILLER_45_564 ();
 sg13g2_decap_8 FILLER_45_571 ();
 sg13g2_decap_8 FILLER_45_578 ();
 sg13g2_decap_8 FILLER_45_585 ();
 sg13g2_decap_8 FILLER_45_592 ();
 sg13g2_decap_8 FILLER_45_599 ();
 sg13g2_decap_8 FILLER_45_606 ();
 sg13g2_decap_8 FILLER_45_613 ();
 sg13g2_decap_8 FILLER_45_620 ();
 sg13g2_decap_8 FILLER_45_627 ();
 sg13g2_decap_8 FILLER_45_634 ();
 sg13g2_decap_8 FILLER_45_641 ();
 sg13g2_decap_8 FILLER_45_648 ();
 sg13g2_decap_8 FILLER_45_655 ();
 sg13g2_decap_8 FILLER_45_662 ();
 sg13g2_decap_8 FILLER_45_669 ();
 sg13g2_decap_8 FILLER_45_676 ();
 sg13g2_decap_8 FILLER_45_683 ();
 sg13g2_decap_8 FILLER_45_690 ();
 sg13g2_decap_8 FILLER_45_697 ();
 sg13g2_decap_8 FILLER_45_704 ();
 sg13g2_decap_8 FILLER_45_711 ();
 sg13g2_decap_8 FILLER_45_718 ();
 sg13g2_decap_8 FILLER_45_725 ();
 sg13g2_decap_8 FILLER_45_732 ();
 sg13g2_decap_8 FILLER_45_739 ();
 sg13g2_decap_8 FILLER_45_746 ();
 sg13g2_decap_8 FILLER_45_753 ();
 sg13g2_decap_8 FILLER_45_760 ();
 sg13g2_decap_8 FILLER_45_767 ();
 sg13g2_decap_8 FILLER_45_774 ();
 sg13g2_decap_8 FILLER_45_781 ();
 sg13g2_decap_8 FILLER_45_788 ();
 sg13g2_decap_8 FILLER_45_795 ();
 sg13g2_decap_8 FILLER_45_802 ();
 sg13g2_decap_8 FILLER_45_809 ();
 sg13g2_decap_8 FILLER_45_816 ();
 sg13g2_decap_8 FILLER_45_823 ();
 sg13g2_decap_8 FILLER_45_830 ();
 sg13g2_decap_8 FILLER_45_837 ();
 sg13g2_decap_8 FILLER_45_844 ();
 sg13g2_decap_8 FILLER_45_851 ();
 sg13g2_decap_8 FILLER_45_858 ();
 sg13g2_decap_8 FILLER_45_865 ();
 sg13g2_decap_8 FILLER_45_872 ();
 sg13g2_decap_8 FILLER_45_879 ();
 sg13g2_decap_8 FILLER_45_886 ();
 sg13g2_decap_8 FILLER_45_893 ();
 sg13g2_decap_8 FILLER_45_900 ();
 sg13g2_decap_8 FILLER_45_907 ();
 sg13g2_decap_8 FILLER_45_914 ();
 sg13g2_decap_4 FILLER_45_921 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_decap_8 FILLER_46_42 ();
 sg13g2_decap_8 FILLER_46_49 ();
 sg13g2_decap_8 FILLER_46_56 ();
 sg13g2_decap_8 FILLER_46_63 ();
 sg13g2_decap_8 FILLER_46_70 ();
 sg13g2_decap_8 FILLER_46_77 ();
 sg13g2_decap_8 FILLER_46_84 ();
 sg13g2_decap_8 FILLER_46_91 ();
 sg13g2_decap_8 FILLER_46_98 ();
 sg13g2_decap_8 FILLER_46_105 ();
 sg13g2_decap_8 FILLER_46_112 ();
 sg13g2_decap_8 FILLER_46_119 ();
 sg13g2_decap_8 FILLER_46_126 ();
 sg13g2_decap_8 FILLER_46_133 ();
 sg13g2_decap_8 FILLER_46_140 ();
 sg13g2_decap_8 FILLER_46_147 ();
 sg13g2_decap_8 FILLER_46_154 ();
 sg13g2_decap_8 FILLER_46_161 ();
 sg13g2_decap_8 FILLER_46_168 ();
 sg13g2_decap_8 FILLER_46_175 ();
 sg13g2_decap_8 FILLER_46_182 ();
 sg13g2_decap_8 FILLER_46_189 ();
 sg13g2_decap_8 FILLER_46_196 ();
 sg13g2_decap_8 FILLER_46_203 ();
 sg13g2_decap_8 FILLER_46_210 ();
 sg13g2_decap_8 FILLER_46_217 ();
 sg13g2_decap_8 FILLER_46_224 ();
 sg13g2_decap_8 FILLER_46_231 ();
 sg13g2_decap_8 FILLER_46_238 ();
 sg13g2_decap_8 FILLER_46_245 ();
 sg13g2_decap_8 FILLER_46_252 ();
 sg13g2_decap_8 FILLER_46_259 ();
 sg13g2_decap_8 FILLER_46_266 ();
 sg13g2_decap_8 FILLER_46_273 ();
 sg13g2_decap_8 FILLER_46_280 ();
 sg13g2_decap_8 FILLER_46_287 ();
 sg13g2_decap_8 FILLER_46_294 ();
 sg13g2_decap_8 FILLER_46_301 ();
 sg13g2_decap_8 FILLER_46_308 ();
 sg13g2_decap_8 FILLER_46_315 ();
 sg13g2_decap_8 FILLER_46_322 ();
 sg13g2_decap_8 FILLER_46_329 ();
 sg13g2_decap_8 FILLER_46_336 ();
 sg13g2_decap_8 FILLER_46_343 ();
 sg13g2_decap_8 FILLER_46_350 ();
 sg13g2_decap_8 FILLER_46_357 ();
 sg13g2_decap_8 FILLER_46_364 ();
 sg13g2_decap_8 FILLER_46_371 ();
 sg13g2_decap_8 FILLER_46_378 ();
 sg13g2_decap_8 FILLER_46_385 ();
 sg13g2_decap_8 FILLER_46_392 ();
 sg13g2_decap_8 FILLER_46_399 ();
 sg13g2_decap_8 FILLER_46_406 ();
 sg13g2_decap_8 FILLER_46_413 ();
 sg13g2_decap_8 FILLER_46_420 ();
 sg13g2_decap_8 FILLER_46_427 ();
 sg13g2_decap_8 FILLER_46_434 ();
 sg13g2_decap_8 FILLER_46_441 ();
 sg13g2_decap_8 FILLER_46_448 ();
 sg13g2_decap_8 FILLER_46_455 ();
 sg13g2_decap_8 FILLER_46_462 ();
 sg13g2_decap_8 FILLER_46_469 ();
 sg13g2_decap_8 FILLER_46_476 ();
 sg13g2_decap_8 FILLER_46_483 ();
 sg13g2_decap_8 FILLER_46_490 ();
 sg13g2_decap_8 FILLER_46_497 ();
 sg13g2_decap_8 FILLER_46_504 ();
 sg13g2_decap_8 FILLER_46_511 ();
 sg13g2_decap_8 FILLER_46_518 ();
 sg13g2_decap_8 FILLER_46_525 ();
 sg13g2_decap_8 FILLER_46_532 ();
 sg13g2_decap_8 FILLER_46_539 ();
 sg13g2_decap_8 FILLER_46_546 ();
 sg13g2_decap_8 FILLER_46_553 ();
 sg13g2_decap_8 FILLER_46_560 ();
 sg13g2_decap_8 FILLER_46_567 ();
 sg13g2_decap_8 FILLER_46_574 ();
 sg13g2_decap_8 FILLER_46_581 ();
 sg13g2_decap_8 FILLER_46_588 ();
 sg13g2_decap_8 FILLER_46_595 ();
 sg13g2_decap_8 FILLER_46_602 ();
 sg13g2_decap_8 FILLER_46_609 ();
 sg13g2_decap_8 FILLER_46_616 ();
 sg13g2_decap_8 FILLER_46_623 ();
 sg13g2_decap_8 FILLER_46_630 ();
 sg13g2_decap_8 FILLER_46_637 ();
 sg13g2_decap_8 FILLER_46_644 ();
 sg13g2_decap_8 FILLER_46_651 ();
 sg13g2_decap_8 FILLER_46_658 ();
 sg13g2_decap_8 FILLER_46_665 ();
 sg13g2_decap_8 FILLER_46_672 ();
 sg13g2_decap_8 FILLER_46_679 ();
 sg13g2_decap_8 FILLER_46_686 ();
 sg13g2_decap_8 FILLER_46_693 ();
 sg13g2_decap_8 FILLER_46_700 ();
 sg13g2_decap_8 FILLER_46_707 ();
 sg13g2_decap_8 FILLER_46_714 ();
 sg13g2_decap_8 FILLER_46_721 ();
 sg13g2_decap_8 FILLER_46_728 ();
 sg13g2_decap_8 FILLER_46_735 ();
 sg13g2_decap_8 FILLER_46_742 ();
 sg13g2_decap_8 FILLER_46_749 ();
 sg13g2_decap_8 FILLER_46_756 ();
 sg13g2_decap_8 FILLER_46_763 ();
 sg13g2_decap_8 FILLER_46_770 ();
 sg13g2_decap_8 FILLER_46_777 ();
 sg13g2_decap_8 FILLER_46_784 ();
 sg13g2_decap_8 FILLER_46_791 ();
 sg13g2_decap_8 FILLER_46_798 ();
 sg13g2_decap_8 FILLER_46_805 ();
 sg13g2_decap_8 FILLER_46_812 ();
 sg13g2_decap_8 FILLER_46_819 ();
 sg13g2_decap_8 FILLER_46_826 ();
 sg13g2_decap_8 FILLER_46_833 ();
 sg13g2_decap_8 FILLER_46_840 ();
 sg13g2_decap_8 FILLER_46_847 ();
 sg13g2_decap_8 FILLER_46_854 ();
 sg13g2_decap_8 FILLER_46_861 ();
 sg13g2_decap_8 FILLER_46_868 ();
 sg13g2_decap_8 FILLER_46_875 ();
 sg13g2_decap_8 FILLER_46_882 ();
 sg13g2_decap_8 FILLER_46_889 ();
 sg13g2_decap_8 FILLER_46_896 ();
 sg13g2_decap_8 FILLER_46_903 ();
 sg13g2_decap_8 FILLER_46_910 ();
 sg13g2_decap_8 FILLER_46_917 ();
 sg13g2_fill_1 FILLER_46_924 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_decap_8 FILLER_47_119 ();
 sg13g2_decap_8 FILLER_47_126 ();
 sg13g2_decap_8 FILLER_47_133 ();
 sg13g2_decap_8 FILLER_47_140 ();
 sg13g2_decap_8 FILLER_47_147 ();
 sg13g2_decap_8 FILLER_47_154 ();
 sg13g2_decap_8 FILLER_47_161 ();
 sg13g2_decap_8 FILLER_47_168 ();
 sg13g2_decap_8 FILLER_47_175 ();
 sg13g2_decap_8 FILLER_47_182 ();
 sg13g2_decap_8 FILLER_47_189 ();
 sg13g2_decap_8 FILLER_47_196 ();
 sg13g2_decap_8 FILLER_47_203 ();
 sg13g2_decap_8 FILLER_47_210 ();
 sg13g2_decap_8 FILLER_47_217 ();
 sg13g2_decap_8 FILLER_47_224 ();
 sg13g2_decap_8 FILLER_47_231 ();
 sg13g2_decap_8 FILLER_47_238 ();
 sg13g2_decap_8 FILLER_47_245 ();
 sg13g2_decap_8 FILLER_47_252 ();
 sg13g2_decap_8 FILLER_47_259 ();
 sg13g2_decap_8 FILLER_47_266 ();
 sg13g2_decap_8 FILLER_47_273 ();
 sg13g2_decap_8 FILLER_47_280 ();
 sg13g2_decap_8 FILLER_47_287 ();
 sg13g2_decap_8 FILLER_47_294 ();
 sg13g2_decap_8 FILLER_47_301 ();
 sg13g2_decap_8 FILLER_47_308 ();
 sg13g2_decap_8 FILLER_47_315 ();
 sg13g2_decap_8 FILLER_47_322 ();
 sg13g2_decap_8 FILLER_47_329 ();
 sg13g2_decap_8 FILLER_47_336 ();
 sg13g2_decap_8 FILLER_47_343 ();
 sg13g2_decap_8 FILLER_47_350 ();
 sg13g2_decap_8 FILLER_47_357 ();
 sg13g2_decap_8 FILLER_47_364 ();
 sg13g2_decap_8 FILLER_47_371 ();
 sg13g2_decap_8 FILLER_47_378 ();
 sg13g2_decap_8 FILLER_47_385 ();
 sg13g2_decap_8 FILLER_47_392 ();
 sg13g2_decap_8 FILLER_47_399 ();
 sg13g2_decap_8 FILLER_47_406 ();
 sg13g2_decap_8 FILLER_47_413 ();
 sg13g2_decap_8 FILLER_47_420 ();
 sg13g2_decap_8 FILLER_47_427 ();
 sg13g2_decap_8 FILLER_47_434 ();
 sg13g2_decap_8 FILLER_47_441 ();
 sg13g2_decap_8 FILLER_47_448 ();
 sg13g2_decap_8 FILLER_47_455 ();
 sg13g2_decap_8 FILLER_47_462 ();
 sg13g2_decap_8 FILLER_47_469 ();
 sg13g2_decap_8 FILLER_47_476 ();
 sg13g2_decap_8 FILLER_47_483 ();
 sg13g2_decap_8 FILLER_47_490 ();
 sg13g2_decap_8 FILLER_47_497 ();
 sg13g2_decap_8 FILLER_47_504 ();
 sg13g2_decap_8 FILLER_47_511 ();
 sg13g2_decap_8 FILLER_47_518 ();
 sg13g2_decap_8 FILLER_47_525 ();
 sg13g2_decap_8 FILLER_47_532 ();
 sg13g2_decap_8 FILLER_47_539 ();
 sg13g2_decap_8 FILLER_47_546 ();
 sg13g2_decap_8 FILLER_47_553 ();
 sg13g2_decap_8 FILLER_47_560 ();
 sg13g2_decap_8 FILLER_47_567 ();
 sg13g2_decap_8 FILLER_47_574 ();
 sg13g2_decap_8 FILLER_47_581 ();
 sg13g2_decap_8 FILLER_47_588 ();
 sg13g2_decap_8 FILLER_47_595 ();
 sg13g2_decap_8 FILLER_47_602 ();
 sg13g2_decap_8 FILLER_47_609 ();
 sg13g2_decap_8 FILLER_47_616 ();
 sg13g2_decap_8 FILLER_47_623 ();
 sg13g2_decap_8 FILLER_47_630 ();
 sg13g2_decap_8 FILLER_47_637 ();
 sg13g2_decap_8 FILLER_47_644 ();
 sg13g2_decap_8 FILLER_47_651 ();
 sg13g2_decap_8 FILLER_47_658 ();
 sg13g2_decap_8 FILLER_47_665 ();
 sg13g2_decap_8 FILLER_47_672 ();
 sg13g2_decap_8 FILLER_47_679 ();
 sg13g2_decap_8 FILLER_47_686 ();
 sg13g2_decap_8 FILLER_47_693 ();
 sg13g2_decap_8 FILLER_47_700 ();
 sg13g2_decap_8 FILLER_47_707 ();
 sg13g2_decap_8 FILLER_47_714 ();
 sg13g2_decap_8 FILLER_47_721 ();
 sg13g2_decap_8 FILLER_47_728 ();
 sg13g2_decap_8 FILLER_47_735 ();
 sg13g2_decap_8 FILLER_47_742 ();
 sg13g2_decap_8 FILLER_47_749 ();
 sg13g2_decap_8 FILLER_47_756 ();
 sg13g2_decap_8 FILLER_47_763 ();
 sg13g2_decap_8 FILLER_47_770 ();
 sg13g2_decap_8 FILLER_47_777 ();
 sg13g2_decap_8 FILLER_47_784 ();
 sg13g2_decap_8 FILLER_47_791 ();
 sg13g2_decap_8 FILLER_47_798 ();
 sg13g2_decap_8 FILLER_47_805 ();
 sg13g2_decap_8 FILLER_47_812 ();
 sg13g2_decap_8 FILLER_47_819 ();
 sg13g2_decap_8 FILLER_47_826 ();
 sg13g2_decap_8 FILLER_47_833 ();
 sg13g2_decap_8 FILLER_47_840 ();
 sg13g2_decap_8 FILLER_47_847 ();
 sg13g2_decap_8 FILLER_47_854 ();
 sg13g2_decap_8 FILLER_47_861 ();
 sg13g2_decap_8 FILLER_47_868 ();
 sg13g2_decap_8 FILLER_47_875 ();
 sg13g2_decap_8 FILLER_47_882 ();
 sg13g2_decap_8 FILLER_47_889 ();
 sg13g2_decap_8 FILLER_47_896 ();
 sg13g2_decap_8 FILLER_47_903 ();
 sg13g2_decap_8 FILLER_47_910 ();
 sg13g2_decap_8 FILLER_47_917 ();
 sg13g2_fill_1 FILLER_47_924 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_119 ();
 sg13g2_decap_8 FILLER_48_126 ();
 sg13g2_decap_8 FILLER_48_133 ();
 sg13g2_decap_8 FILLER_48_140 ();
 sg13g2_decap_8 FILLER_48_147 ();
 sg13g2_decap_8 FILLER_48_154 ();
 sg13g2_decap_8 FILLER_48_161 ();
 sg13g2_decap_8 FILLER_48_168 ();
 sg13g2_decap_8 FILLER_48_175 ();
 sg13g2_decap_8 FILLER_48_182 ();
 sg13g2_decap_8 FILLER_48_189 ();
 sg13g2_decap_8 FILLER_48_196 ();
 sg13g2_decap_8 FILLER_48_203 ();
 sg13g2_decap_8 FILLER_48_210 ();
 sg13g2_decap_8 FILLER_48_217 ();
 sg13g2_decap_8 FILLER_48_224 ();
 sg13g2_decap_8 FILLER_48_231 ();
 sg13g2_decap_8 FILLER_48_238 ();
 sg13g2_decap_8 FILLER_48_245 ();
 sg13g2_decap_8 FILLER_48_252 ();
 sg13g2_decap_8 FILLER_48_259 ();
 sg13g2_decap_8 FILLER_48_266 ();
 sg13g2_decap_8 FILLER_48_273 ();
 sg13g2_decap_8 FILLER_48_280 ();
 sg13g2_decap_8 FILLER_48_287 ();
 sg13g2_decap_8 FILLER_48_294 ();
 sg13g2_decap_8 FILLER_48_301 ();
 sg13g2_decap_8 FILLER_48_308 ();
 sg13g2_decap_8 FILLER_48_315 ();
 sg13g2_decap_8 FILLER_48_322 ();
 sg13g2_decap_8 FILLER_48_329 ();
 sg13g2_decap_8 FILLER_48_336 ();
 sg13g2_decap_8 FILLER_48_343 ();
 sg13g2_decap_8 FILLER_48_350 ();
 sg13g2_decap_8 FILLER_48_357 ();
 sg13g2_decap_8 FILLER_48_364 ();
 sg13g2_decap_8 FILLER_48_371 ();
 sg13g2_decap_8 FILLER_48_378 ();
 sg13g2_decap_8 FILLER_48_385 ();
 sg13g2_decap_8 FILLER_48_392 ();
 sg13g2_decap_8 FILLER_48_399 ();
 sg13g2_decap_8 FILLER_48_406 ();
 sg13g2_decap_8 FILLER_48_413 ();
 sg13g2_decap_8 FILLER_48_420 ();
 sg13g2_decap_8 FILLER_48_427 ();
 sg13g2_decap_8 FILLER_48_434 ();
 sg13g2_decap_8 FILLER_48_441 ();
 sg13g2_decap_8 FILLER_48_448 ();
 sg13g2_decap_8 FILLER_48_455 ();
 sg13g2_decap_8 FILLER_48_462 ();
 sg13g2_decap_8 FILLER_48_469 ();
 sg13g2_decap_8 FILLER_48_476 ();
 sg13g2_decap_8 FILLER_48_483 ();
 sg13g2_decap_8 FILLER_48_490 ();
 sg13g2_decap_8 FILLER_48_497 ();
 sg13g2_decap_8 FILLER_48_504 ();
 sg13g2_decap_8 FILLER_48_511 ();
 sg13g2_decap_8 FILLER_48_518 ();
 sg13g2_decap_8 FILLER_48_525 ();
 sg13g2_decap_8 FILLER_48_532 ();
 sg13g2_decap_8 FILLER_48_539 ();
 sg13g2_decap_8 FILLER_48_546 ();
 sg13g2_decap_8 FILLER_48_553 ();
 sg13g2_decap_8 FILLER_48_560 ();
 sg13g2_decap_8 FILLER_48_567 ();
 sg13g2_decap_8 FILLER_48_574 ();
 sg13g2_decap_8 FILLER_48_581 ();
 sg13g2_decap_8 FILLER_48_588 ();
 sg13g2_decap_8 FILLER_48_595 ();
 sg13g2_decap_8 FILLER_48_602 ();
 sg13g2_decap_8 FILLER_48_609 ();
 sg13g2_decap_8 FILLER_48_616 ();
 sg13g2_decap_8 FILLER_48_623 ();
 sg13g2_decap_8 FILLER_48_630 ();
 sg13g2_decap_8 FILLER_48_637 ();
 sg13g2_decap_8 FILLER_48_644 ();
 sg13g2_decap_8 FILLER_48_651 ();
 sg13g2_decap_8 FILLER_48_658 ();
 sg13g2_decap_8 FILLER_48_665 ();
 sg13g2_decap_8 FILLER_48_672 ();
 sg13g2_decap_8 FILLER_48_679 ();
 sg13g2_decap_8 FILLER_48_686 ();
 sg13g2_decap_8 FILLER_48_693 ();
 sg13g2_decap_8 FILLER_48_700 ();
 sg13g2_decap_8 FILLER_48_707 ();
 sg13g2_decap_8 FILLER_48_714 ();
 sg13g2_decap_8 FILLER_48_721 ();
 sg13g2_decap_8 FILLER_48_728 ();
 sg13g2_decap_8 FILLER_48_735 ();
 sg13g2_decap_8 FILLER_48_742 ();
 sg13g2_decap_8 FILLER_48_749 ();
 sg13g2_decap_8 FILLER_48_756 ();
 sg13g2_decap_8 FILLER_48_763 ();
 sg13g2_decap_8 FILLER_48_770 ();
 sg13g2_decap_8 FILLER_48_777 ();
 sg13g2_decap_8 FILLER_48_784 ();
 sg13g2_decap_8 FILLER_48_791 ();
 sg13g2_decap_8 FILLER_48_798 ();
 sg13g2_decap_8 FILLER_48_805 ();
 sg13g2_decap_8 FILLER_48_812 ();
 sg13g2_decap_8 FILLER_48_819 ();
 sg13g2_decap_8 FILLER_48_826 ();
 sg13g2_decap_8 FILLER_48_833 ();
 sg13g2_decap_8 FILLER_48_840 ();
 sg13g2_decap_8 FILLER_48_847 ();
 sg13g2_decap_8 FILLER_48_854 ();
 sg13g2_decap_8 FILLER_48_861 ();
 sg13g2_decap_8 FILLER_48_868 ();
 sg13g2_decap_8 FILLER_48_875 ();
 sg13g2_decap_8 FILLER_48_882 ();
 sg13g2_decap_8 FILLER_48_889 ();
 sg13g2_decap_8 FILLER_48_896 ();
 sg13g2_decap_8 FILLER_48_903 ();
 sg13g2_decap_8 FILLER_48_910 ();
 sg13g2_decap_8 FILLER_48_917 ();
 sg13g2_fill_1 FILLER_48_924 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_8 FILLER_49_42 ();
 sg13g2_decap_8 FILLER_49_49 ();
 sg13g2_decap_8 FILLER_49_56 ();
 sg13g2_decap_8 FILLER_49_63 ();
 sg13g2_decap_8 FILLER_49_70 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_84 ();
 sg13g2_decap_8 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_decap_8 FILLER_49_105 ();
 sg13g2_decap_8 FILLER_49_112 ();
 sg13g2_decap_8 FILLER_49_119 ();
 sg13g2_decap_8 FILLER_49_126 ();
 sg13g2_decap_8 FILLER_49_133 ();
 sg13g2_decap_8 FILLER_49_140 ();
 sg13g2_decap_8 FILLER_49_147 ();
 sg13g2_decap_8 FILLER_49_154 ();
 sg13g2_decap_8 FILLER_49_161 ();
 sg13g2_decap_8 FILLER_49_168 ();
 sg13g2_decap_8 FILLER_49_175 ();
 sg13g2_decap_8 FILLER_49_182 ();
 sg13g2_decap_8 FILLER_49_189 ();
 sg13g2_decap_8 FILLER_49_196 ();
 sg13g2_decap_8 FILLER_49_203 ();
 sg13g2_decap_8 FILLER_49_210 ();
 sg13g2_decap_8 FILLER_49_217 ();
 sg13g2_decap_8 FILLER_49_224 ();
 sg13g2_decap_8 FILLER_49_231 ();
 sg13g2_decap_8 FILLER_49_238 ();
 sg13g2_decap_8 FILLER_49_245 ();
 sg13g2_decap_8 FILLER_49_252 ();
 sg13g2_decap_8 FILLER_49_259 ();
 sg13g2_decap_8 FILLER_49_266 ();
 sg13g2_decap_8 FILLER_49_273 ();
 sg13g2_decap_8 FILLER_49_280 ();
 sg13g2_decap_8 FILLER_49_287 ();
 sg13g2_decap_8 FILLER_49_294 ();
 sg13g2_decap_8 FILLER_49_301 ();
 sg13g2_decap_8 FILLER_49_308 ();
 sg13g2_decap_8 FILLER_49_315 ();
 sg13g2_decap_8 FILLER_49_322 ();
 sg13g2_decap_8 FILLER_49_329 ();
 sg13g2_decap_8 FILLER_49_336 ();
 sg13g2_decap_8 FILLER_49_343 ();
 sg13g2_decap_8 FILLER_49_350 ();
 sg13g2_decap_8 FILLER_49_357 ();
 sg13g2_decap_8 FILLER_49_364 ();
 sg13g2_decap_8 FILLER_49_371 ();
 sg13g2_decap_8 FILLER_49_378 ();
 sg13g2_decap_8 FILLER_49_385 ();
 sg13g2_decap_8 FILLER_49_392 ();
 sg13g2_decap_8 FILLER_49_399 ();
 sg13g2_decap_8 FILLER_49_406 ();
 sg13g2_decap_8 FILLER_49_413 ();
 sg13g2_decap_8 FILLER_49_420 ();
 sg13g2_decap_8 FILLER_49_427 ();
 sg13g2_decap_8 FILLER_49_434 ();
 sg13g2_decap_8 FILLER_49_441 ();
 sg13g2_decap_8 FILLER_49_448 ();
 sg13g2_decap_8 FILLER_49_455 ();
 sg13g2_decap_8 FILLER_49_462 ();
 sg13g2_decap_8 FILLER_49_469 ();
 sg13g2_decap_8 FILLER_49_476 ();
 sg13g2_decap_8 FILLER_49_483 ();
 sg13g2_decap_8 FILLER_49_490 ();
 sg13g2_decap_8 FILLER_49_497 ();
 sg13g2_decap_8 FILLER_49_504 ();
 sg13g2_decap_8 FILLER_49_511 ();
 sg13g2_decap_8 FILLER_49_518 ();
 sg13g2_decap_8 FILLER_49_525 ();
 sg13g2_decap_8 FILLER_49_532 ();
 sg13g2_decap_8 FILLER_49_539 ();
 sg13g2_decap_8 FILLER_49_546 ();
 sg13g2_decap_8 FILLER_49_553 ();
 sg13g2_decap_8 FILLER_49_560 ();
 sg13g2_decap_8 FILLER_49_567 ();
 sg13g2_decap_8 FILLER_49_574 ();
 sg13g2_decap_8 FILLER_49_581 ();
 sg13g2_decap_8 FILLER_49_588 ();
 sg13g2_decap_8 FILLER_49_595 ();
 sg13g2_decap_8 FILLER_49_602 ();
 sg13g2_decap_8 FILLER_49_609 ();
 sg13g2_decap_8 FILLER_49_616 ();
 sg13g2_decap_8 FILLER_49_623 ();
 sg13g2_decap_8 FILLER_49_630 ();
 sg13g2_decap_8 FILLER_49_637 ();
 sg13g2_decap_8 FILLER_49_644 ();
 sg13g2_decap_8 FILLER_49_651 ();
 sg13g2_decap_8 FILLER_49_658 ();
 sg13g2_decap_8 FILLER_49_665 ();
 sg13g2_decap_8 FILLER_49_672 ();
 sg13g2_decap_8 FILLER_49_679 ();
 sg13g2_decap_8 FILLER_49_686 ();
 sg13g2_decap_8 FILLER_49_693 ();
 sg13g2_decap_8 FILLER_49_700 ();
 sg13g2_decap_8 FILLER_49_707 ();
 sg13g2_decap_8 FILLER_49_714 ();
 sg13g2_decap_8 FILLER_49_721 ();
 sg13g2_decap_8 FILLER_49_728 ();
 sg13g2_decap_8 FILLER_49_735 ();
 sg13g2_decap_8 FILLER_49_742 ();
 sg13g2_decap_8 FILLER_49_749 ();
 sg13g2_decap_8 FILLER_49_756 ();
 sg13g2_decap_8 FILLER_49_763 ();
 sg13g2_decap_8 FILLER_49_770 ();
 sg13g2_decap_8 FILLER_49_777 ();
 sg13g2_decap_8 FILLER_49_784 ();
 sg13g2_decap_8 FILLER_49_791 ();
 sg13g2_decap_8 FILLER_49_798 ();
 sg13g2_decap_8 FILLER_49_805 ();
 sg13g2_decap_8 FILLER_49_812 ();
 sg13g2_decap_8 FILLER_49_819 ();
 sg13g2_decap_8 FILLER_49_826 ();
 sg13g2_decap_8 FILLER_49_833 ();
 sg13g2_decap_8 FILLER_49_840 ();
 sg13g2_decap_8 FILLER_49_847 ();
 sg13g2_decap_8 FILLER_49_854 ();
 sg13g2_decap_8 FILLER_49_861 ();
 sg13g2_decap_8 FILLER_49_868 ();
 sg13g2_decap_8 FILLER_49_875 ();
 sg13g2_decap_8 FILLER_49_882 ();
 sg13g2_decap_8 FILLER_49_889 ();
 sg13g2_decap_8 FILLER_49_896 ();
 sg13g2_decap_8 FILLER_49_903 ();
 sg13g2_decap_8 FILLER_49_910 ();
 sg13g2_decap_8 FILLER_49_917 ();
 sg13g2_fill_1 FILLER_49_924 ();
 assign uio_oe[0] = net25;
 assign uio_oe[1] = net26;
 assign uio_oe[2] = net27;
 assign uio_oe[3] = net28;
 assign uio_oe[4] = net29;
 assign uio_oe[5] = net30;
 assign uio_oe[6] = net31;
 assign uio_oe[7] = net32;
 assign uio_out[0] = net33;
 assign uio_out[1] = net34;
 assign uio_out[2] = net35;
 assign uio_out[3] = net36;
 assign uio_out[4] = net37;
 assign uio_out[5] = net38;
 assign uio_out[6] = net39;
 assign uio_out[7] = net40;
endmodule
