* NGSPICE file created from E_TT_IF.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_dlhq_1 abstract view
.subckt sg13g2_dlhq_1 D GATE Q VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_mux4_1 abstract view
.subckt sg13g2_mux4_1 S0 A0 A1 A2 A3 S1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_antennanp abstract view
.subckt sg13g2_antennanp VDD VSS A
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

.subckt E_TT_IF CLK_TT_PROJECT E1END[0] E1END[1] E1END[2] E1END[3] E2END[0] E2END[1]
+ E2END[2] E2END[3] E2END[4] E2END[5] E2END[6] E2END[7] E2MID[0] E2MID[1] E2MID[2]
+ E2MID[3] E2MID[4] E2MID[5] E2MID[6] E2MID[7] E6END[0] E6END[10] E6END[11] E6END[1]
+ E6END[2] E6END[3] E6END[4] E6END[5] E6END[6] E6END[7] E6END[8] E6END[9] EE4END[0]
+ EE4END[10] EE4END[11] EE4END[12] EE4END[13] EE4END[14] EE4END[15] EE4END[1] EE4END[2]
+ EE4END[3] EE4END[4] EE4END[5] EE4END[6] EE4END[7] EE4END[8] EE4END[9] ENA_TT_PROJECT
+ FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13] FrameData[14]
+ FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19] FrameData[1]
+ FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24] FrameData[25]
+ FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2] FrameData[30]
+ FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6] FrameData[7] FrameData[8]
+ FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11] FrameData_O[12] FrameData_O[13]
+ FrameData_O[14] FrameData_O[15] FrameData_O[16] FrameData_O[17] FrameData_O[18]
+ FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21] FrameData_O[22] FrameData_O[23]
+ FrameData_O[24] FrameData_O[25] FrameData_O[26] FrameData_O[27] FrameData_O[28]
+ FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31] FrameData_O[3] FrameData_O[4]
+ FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8] FrameData_O[9] FrameStrobe[0]
+ FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13] FrameStrobe[14]
+ FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18] FrameStrobe[19]
+ FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5] FrameStrobe[6]
+ FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1] N1BEG[2] N1BEG[3]
+ N1END[0] N1END[1] N1END[2] N1END[3] N2BEG[0] N2BEG[1] N2BEG[2] N2BEG[3] N2BEG[4]
+ N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0] N2BEGb[1] N2BEGb[2] N2BEGb[3] N2BEGb[4] N2BEGb[5]
+ N2BEGb[6] N2BEGb[7] N2END[0] N2END[1] N2END[2] N2END[3] N2END[4] N2END[5] N2END[6]
+ N2END[7] N2MID[0] N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5] N2MID[6] N2MID[7]
+ N4BEG[0] N4BEG[10] N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2]
+ N4BEG[3] N4BEG[4] N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9] N4END[0] N4END[10]
+ N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2] N4END[3] N4END[4]
+ N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] RST_N_TT_PROJECT S1BEG[0] S1BEG[1]
+ S1BEG[2] S1BEG[3] S1END[0] S1END[1] S1END[2] S1END[3] S2BEG[0] S2BEG[1] S2BEG[2]
+ S2BEG[3] S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7] S2BEGb[0] S2BEGb[1] S2BEGb[2] S2BEGb[3]
+ S2BEGb[4] S2BEGb[5] S2BEGb[6] S2BEGb[7] S2END[0] S2END[1] S2END[2] S2END[3] S2END[4]
+ S2END[5] S2END[6] S2END[7] S2MID[0] S2MID[1] S2MID[2] S2MID[3] S2MID[4] S2MID[5]
+ S2MID[6] S2MID[7] S4BEG[0] S4BEG[10] S4BEG[11] S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15]
+ S4BEG[1] S4BEG[2] S4BEG[3] S4BEG[4] S4BEG[5] S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9]
+ S4END[0] S4END[10] S4END[11] S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2]
+ S4END[3] S4END[4] S4END[5] S4END[6] S4END[7] S4END[8] S4END[9] UIO_IN_TT_PROJECT0
+ UIO_IN_TT_PROJECT1 UIO_IN_TT_PROJECT2 UIO_IN_TT_PROJECT3 UIO_IN_TT_PROJECT4 UIO_IN_TT_PROJECT5
+ UIO_IN_TT_PROJECT6 UIO_IN_TT_PROJECT7 UIO_OE_TT_PROJECT0 UIO_OE_TT_PROJECT1 UIO_OE_TT_PROJECT2
+ UIO_OE_TT_PROJECT3 UIO_OE_TT_PROJECT4 UIO_OE_TT_PROJECT5 UIO_OE_TT_PROJECT6 UIO_OE_TT_PROJECT7
+ UIO_OUT_TT_PROJECT0 UIO_OUT_TT_PROJECT1 UIO_OUT_TT_PROJECT2 UIO_OUT_TT_PROJECT3
+ UIO_OUT_TT_PROJECT4 UIO_OUT_TT_PROJECT5 UIO_OUT_TT_PROJECT6 UIO_OUT_TT_PROJECT7
+ UI_IN_TT_PROJECT0 UI_IN_TT_PROJECT1 UI_IN_TT_PROJECT2 UI_IN_TT_PROJECT3 UI_IN_TT_PROJECT4
+ UI_IN_TT_PROJECT5 UI_IN_TT_PROJECT6 UI_IN_TT_PROJECT7 UO_OUT_TT_PROJECT0 UO_OUT_TT_PROJECT1
+ UO_OUT_TT_PROJECT2 UO_OUT_TT_PROJECT3 UO_OUT_TT_PROJECT4 UO_OUT_TT_PROJECT5 UO_OUT_TT_PROJECT6
+ UO_OUT_TT_PROJECT7 UserCLK UserCLKo VGND VPWR W1BEG[0] W1BEG[1] W1BEG[2] W1BEG[3]
+ W2BEG[0] W2BEG[1] W2BEG[2] W2BEG[3] W2BEG[4] W2BEG[5] W2BEG[6] W2BEG[7] W2BEGb[0]
+ W2BEGb[1] W2BEGb[2] W2BEGb[3] W2BEGb[4] W2BEGb[5] W2BEGb[6] W2BEGb[7] W6BEG[0] W6BEG[10]
+ W6BEG[11] W6BEG[1] W6BEG[2] W6BEG[3] W6BEG[4] W6BEG[5] W6BEG[6] W6BEG[7] W6BEG[8]
+ W6BEG[9] WW4BEG[0] WW4BEG[10] WW4BEG[11] WW4BEG[12] WW4BEG[13] WW4BEG[14] WW4BEG[15]
+ WW4BEG[1] WW4BEG[2] WW4BEG[3] WW4BEG[4] WW4BEG[5] WW4BEG[6] WW4BEG[7] WW4BEG[8]
+ WW4BEG[9]
X_1270_ S4END[7] S4BEG[3] VPWR VGND sg13g2_buf_1
X_0419_ VPWR _0038_ _0037_ VGND sg13g2_inv_1
X_0985_ FrameData[19] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit19.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_5_4 VPWR VGND sg13g2_fill_1
XFILLER_52_6 VPWR VGND sg13g2_fill_1
X_1184_ FrameData[25] FrameData_O[25] VPWR VGND sg13g2_buf_1
X_0770_ _0348_ _0347_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit19.Q Inst_E_TT_IF_switch_matrix.S4BEG0
+ VPWR VGND sg13g2_mux2_1
X_0968_ FrameData[2] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit2.Q VPWR
+ VGND sg13g2_dlhq_1
X_1322_ Inst_E_TT_IF_switch_matrix.WW4BEG6 WW4BEG[6] VPWR VGND sg13g2_buf_1
X_1253_ Inst_E_TT_IF_switch_matrix.S2BEG2 S2BEG[2] VPWR VGND sg13g2_buf_1
X_0899_ FrameData[29] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit29.Q VPWR
+ VGND sg13g2_dlhq_1
X_0753_ VGND VPWR _0332_ _0334_ Inst_E_TT_IF_switch_matrix.S4BEG3 _0330_ sg13g2_a21oi_1
X_0684_ _0079_ _0274_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit22.Q _0275_ VPWR VGND
+ sg13g2_mux2_1
X_0822_ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit21.Q UO_OUT_TT_PROJECT1 _0155_ UIO_OUT_TT_PROJECT5
+ _0096_ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit20.Q Inst_E_TT_IF_switch_matrix.WW4BEG13
+ VPWR VGND sg13g2_mux4_1
X_1236_ N4END[9] N4BEG[5] VPWR VGND sg13g2_buf_1
X_1098_ FrameData[4] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit4.Q VPWR
+ VGND sg13g2_dlhq_1
X_1167_ FrameData[8] FrameData_O[8] VPWR VGND sg13g2_buf_1
X_1305_ Inst_E_TT_IF_switch_matrix.W6BEG1 W6BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_38_128 VPWR VGND sg13g2_fill_2
X_1219_ Inst_E_TT_IF_switch_matrix.N2BEG4 N2BEG[4] VPWR VGND sg13g2_buf_1
X_0805_ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit2.Q VPWR _0379_ VGND E2MID[6] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit3.Q
+ sg13g2_o21ai_1
X_0736_ _0320_ _0319_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit6.Q Inst_E_TT_IF_switch_matrix.W1BEG2
+ VPWR VGND sg13g2_mux2_1
X_0667_ _0134_ _0096_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit25.Q _0259_ VPWR VGND
+ sg13g2_mux2_1
X_0598_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit18.Q E2END[2] UIO_OUT_TT_PROJECT5 UIO_OUT_TT_PROJECT2
+ UIO_OUT_TT_PROJECT6 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit17.Q _0198_ VPWR VGND
+ sg13g2_mux4_1
X_1021_ FrameData[23] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit23.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_29_74 VPWR VGND sg13g2_fill_2
X_0521_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit5.Q _0015_ _0130_ VPWR VGND sg13g2_nor2_1
X_0452_ UIO_IN_TT_PROJECT6 _0068_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit28.Q _0066_
+ _0063_ VPWR VGND sg13g2_a22oi_1
X_0383_ VPWR _0002_ S1END[3] VGND sg13g2_inv_1
XANTENNA_5 VPWR VGND Inst_E_TT_IF_switch_matrix.S4BEG2 sg13g2_antennanp
X_1004_ FrameData[6] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit6.Q VPWR
+ VGND sg13g2_dlhq_1
X_0719_ Inst_E_TT_IF_switch_matrix.W2BEG1 _0304_ _0306_ _0302_ _0298_ VPWR VGND sg13g2_a22oi_1
X_0504_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit11.Q _0014_ _0115_ VPWR VGND sg13g2_nor2_1
X_0435_ VPWR _0053_ _0052_ VGND sg13g2_inv_1
XFILLER_42_85 VPWR VGND sg13g2_fill_2
X_0418_ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit4.Q E2MID[3] E2MID[6] E2END[1] E2END[2]
+ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit5.Q _0037_ VPWR VGND sg13g2_mux4_1
X_0984_ FrameData[18] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit18.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_10_104 VPWR VGND sg13g2_fill_1
X_1183_ FrameData[24] FrameData_O[24] VPWR VGND sg13g2_buf_1
X_1252_ Inst_E_TT_IF_switch_matrix.S2BEG1 S2BEG[1] VPWR VGND sg13g2_buf_1
X_1321_ Inst_E_TT_IF_switch_matrix.WW4BEG5 WW4BEG[5] VPWR VGND sg13g2_buf_1
X_0898_ FrameData[28] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit28.Q VPWR
+ VGND sg13g2_dlhq_1
X_0967_ FrameData[1] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit1.Q VPWR
+ VGND sg13g2_dlhq_1
X_0752_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame7_bit27.Q _0333_ _0334_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit28.Q
+ sg13g2_a21oi_1
XFILLER_0_36 VPWR VGND sg13g2_fill_1
X_0821_ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit23.Q UO_OUT_TT_PROJECT2 _0162_ UIO_OUT_TT_PROJECT6
+ _0104_ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit22.Q Inst_E_TT_IF_switch_matrix.WW4BEG14
+ VPWR VGND sg13g2_mux4_1
XFILLER_49_170 VPWR VGND sg13g2_fill_1
X_1235_ N4END[8] N4BEG[4] VPWR VGND sg13g2_buf_1
X_0683_ VPWR VGND Inst_E_TT_IF_ConfigMem.Inst_frame0_bit30.Q _0273_ _0272_ _0002_
+ _0274_ Inst_E_TT_IF_ConfigMem.Inst_frame0_bit31.Q sg13g2_a221oi_1
X_1166_ FrameData[7] FrameData_O[7] VPWR VGND sg13g2_buf_1
X_1097_ FrameData[3] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit3.Q VPWR
+ VGND sg13g2_dlhq_1
X_1304_ Inst_E_TT_IF_switch_matrix.W6BEG0 W6BEG[0] VPWR VGND sg13g2_buf_1
XFILLER_18_43 VPWR VGND sg13g2_fill_1
XFILLER_18_21 VPWR VGND sg13g2_fill_1
X_0804_ _0376_ _0378_ Inst_E_TT_IF_switch_matrix.N4BEG0 VPWR VGND sg13g2_nor2_1
X_0666_ Inst_E_TT_IF_switch_matrix.W2BEG6 _0256_ _0258_ _0254_ _0253_ VPWR VGND sg13g2_a22oi_1
X_0735_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit4.Q N1END[2] S1END[2] UO_OUT_TT_PROJECT0
+ UO_OUT_TT_PROJECT5 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit5.Q _0320_ VPWR VGND sg13g2_mux4_1
X_0597_ _0193_ _0196_ _0197_ VPWR VGND sg13g2_nor2_1
X_1020_ FrameData[22] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit22.Q VPWR
+ VGND sg13g2_dlhq_1
X_1149_ FrameData[23] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit23.Q VPWR
+ VGND sg13g2_dlhq_1
X_1218_ Inst_E_TT_IF_switch_matrix.N2BEG3 N2BEG[3] VPWR VGND sg13g2_buf_1
XFILLER_20_88 VPWR VGND sg13g2_fill_2
XFILLER_43_198 VPWR VGND sg13g2_fill_2
X_0520_ E2MID[6] EE4END[6] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit5.Q _0129_ VPWR VGND
+ sg13g2_mux2_1
X_0451_ _0068_ _0067_ _0006_ _0065_ _0060_ VPWR VGND sg13g2_a22oi_1
XANTENNA_6 VPWR VGND N2END[0] sg13g2_antennanp
X_0382_ VPWR _0001_ E1END[3] VGND sg13g2_inv_1
X_1003_ FrameData[5] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit5.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_25_198 VPWR VGND sg13g2_fill_2
X_0649_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit31.Q _0120_ _0112_ _0052_ _0242_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit0.Q
+ _0243_ VPWR VGND sg13g2_mux4_1
X_0718_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame6_bit14.Q _0305_ _0306_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit15.Q
+ sg13g2_a21oi_1
XFILLER_16_165 VPWR VGND sg13g2_fill_1
X_0434_ Inst_E_TT_IF_ConfigMem.Inst_frame0_bit22.Q N2MID[7] N2END[7] S2MID[7] S2END[7]
+ Inst_E_TT_IF_ConfigMem.Inst_frame0_bit23.Q _0052_ VPWR VGND sg13g2_mux4_1
X_0503_ E2MID[0] EE4END[0] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit11.Q _0114_ VPWR
+ VGND sg13g2_mux2_1
XFILLER_42_97 VPWR VGND sg13g2_fill_1
X_0983_ FrameData[17] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit17.Q VPWR
+ VGND sg13g2_dlhq_1
X_0417_ VPWR _0036_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit16.Q VGND sg13g2_inv_1
XFILLER_53_96 VPWR VGND sg13g2_fill_2
X_1182_ FrameData[23] FrameData_O[23] VPWR VGND sg13g2_buf_1
X_1251_ Inst_E_TT_IF_switch_matrix.S2BEG0 S2BEG[0] VPWR VGND sg13g2_buf_1
X_1320_ Inst_E_TT_IF_switch_matrix.WW4BEG4 WW4BEG[4] VPWR VGND sg13g2_buf_1
XFILLER_5_197 VPWR VGND sg13g2_fill_2
X_0897_ FrameData[27] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit27.Q VPWR
+ VGND sg13g2_dlhq_1
X_0966_ FrameData[0] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit0.Q VPWR
+ VGND sg13g2_dlhq_1
X_1234_ N4END[7] N4BEG[3] VPWR VGND sg13g2_buf_1
X_0682_ N1END[3] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit30.Q Inst_E_TT_IF_ConfigMem.Inst_frame0_bit31.Q
+ _0273_ VPWR VGND sg13g2_nor3_1
X_1165_ FrameData[6] FrameData_O[6] VPWR VGND sg13g2_buf_1
X_0751_ EE4END[15] _0087_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit29.Q _0333_ VPWR VGND
+ sg13g2_mux2_1
X_1096_ FrameData[2] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit2.Q VPWR
+ VGND sg13g2_dlhq_1
X_0820_ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit25.Q UO_OUT_TT_PROJECT3 _0169_ UIO_OUT_TT_PROJECT7
+ _0112_ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit24.Q Inst_E_TT_IF_switch_matrix.WW4BEG15
+ VPWR VGND sg13g2_mux4_1
X_1303_ Inst_E_TT_IF_switch_matrix.W2BEGb7 W2BEGb[7] VPWR VGND sg13g2_buf_1
X_0949_ FrameData[15] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit15.Q VPWR
+ VGND sg13g2_dlhq_1
X_0803_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit15.Q _0377_ _0378_ VPWR VGND sg13g2_nor2_1
X_0665_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame6_bit29.Q _0257_ _0258_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit30.Q
+ sg13g2_a21oi_1
X_0734_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit4.Q UIO_OE_TT_PROJECT2 UIO_OE_TT_PROJECT3
+ UIO_OE_TT_PROJECT4 UIO_OE_TT_PROJECT5 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit5.Q
+ _0319_ VPWR VGND sg13g2_mux4_1
XFILLER_52_199 VPWR VGND sg13g2_fill_1
XFILLER_52_111 VPWR VGND sg13g2_fill_2
X_1079_ FrameData[17] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit17.Q VPWR
+ VGND sg13g2_dlhq_1
X_1217_ Inst_E_TT_IF_switch_matrix.N2BEG2 N2BEG[2] VPWR VGND sg13g2_buf_1
X_1148_ FrameData[22] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit22.Q VPWR
+ VGND sg13g2_dlhq_1
X_0596_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit19.Q VPWR _0196_ VGND Inst_E_TT_IF_ConfigMem.Inst_frame5_bit18.Q
+ _0195_ sg13g2_o21ai_1
XANTENNA_7 VPWR VGND N4END[10] sg13g2_antennanp
X_0381_ VPWR _0000_ E2END[3] VGND sg13g2_inv_1
X_0450_ E2MID[6] EE4END[6] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit29.Q _0067_ VPWR
+ VGND sg13g2_mux2_1
XFILLER_28_141 VPWR VGND sg13g2_fill_1
XFILLER_34_199 VPWR VGND sg13g2_fill_1
X_0648_ VPWR VGND Inst_E_TT_IF_ConfigMem.Inst_frame0_bit24.Q _0240_ _0241_ _0009_
+ _0242_ Inst_E_TT_IF_ConfigMem.Inst_frame0_bit25.Q sg13g2_a221oi_1
X_1002_ FrameData[4] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit4.Q VPWR
+ VGND sg13g2_dlhq_1
X_0579_ _0177_ _0180_ _0181_ VPWR VGND sg13g2_nor2_1
X_0717_ UIO_OUT_TT_PROJECT1 UIO_OE_TT_PROJECT6 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit13.Q
+ _0305_ VPWR VGND sg13g2_mux2_1
XFILLER_25_111 VPWR VGND sg13g2_fill_2
XFILLER_16_111 VPWR VGND sg13g2_fill_1
X_0433_ Inst_E_TT_IF_ConfigMem.Inst_frame0_bit6.Q N1END[3] N4END[3] S1END[3] S4END[3]
+ Inst_E_TT_IF_ConfigMem.Inst_frame0_bit7.Q _0051_ VPWR VGND sg13g2_mux4_1
X_0502_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit12.Q _0112_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit11.Q
+ _0113_ VPWR VGND sg13g2_nand3_1
XFILLER_22_147 VPWR VGND sg13g2_fill_2
XFILLER_26_77 VPWR VGND sg13g2_decap_8
X_0982_ FrameData[16] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit16.Q VPWR
+ VGND sg13g2_dlhq_1
X_0416_ VPWR _0035_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit19.Q VGND sg13g2_inv_1
X_1181_ FrameData[22] FrameData_O[22] VPWR VGND sg13g2_buf_1
X_0896_ FrameData[26] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit26.Q VPWR
+ VGND sg13g2_dlhq_1
X_1250_ Inst_E_TT_IF_switch_matrix.S1BEG3 S1BEG[3] VPWR VGND sg13g2_buf_1
X_0965_ FrameData[31] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit31.Q VPWR
+ VGND sg13g2_dlhq_1
X_1233_ N4END[6] N4BEG[2] VPWR VGND sg13g2_buf_1
X_0681_ _0272_ E6END[3] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit31.Q VPWR VGND sg13g2_nand2b_1
X_0750_ _0331_ VPWR _0332_ VGND _0031_ _0120_ sg13g2_o21ai_1
X_1164_ FrameData[5] FrameData_O[5] VPWR VGND sg13g2_buf_1
X_1095_ FrameData[1] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit1.Q VPWR
+ VGND sg13g2_dlhq_1
X_1302_ Inst_E_TT_IF_switch_matrix.W2BEGb6 W2BEGb[6] VPWR VGND sg13g2_buf_1
X_0879_ FrameData[9] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit9.Q VPWR
+ VGND sg13g2_dlhq_1
X_0948_ FrameData[14] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit14.Q VPWR
+ VGND sg13g2_dlhq_1
X_0802_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit14.Q E1END[0] EE4END[0] _0141_ _0111_
+ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit16.Q _0377_ VPWR VGND sg13g2_mux4_1
X_1147_ FrameData[21] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit21.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_52_178 VPWR VGND sg13g2_fill_1
X_1078_ FrameData[16] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit16.Q VPWR
+ VGND sg13g2_dlhq_1
X_1216_ Inst_E_TT_IF_switch_matrix.N2BEG1 N2BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_37_164 VPWR VGND sg13g2_fill_1
X_0664_ UIO_OUT_TT_PROJECT6 UIO_OE_TT_PROJECT1 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit28.Q
+ _0257_ VPWR VGND sg13g2_mux2_1
X_0733_ _0318_ _0317_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit9.Q Inst_E_TT_IF_switch_matrix.W1BEG3
+ VPWR VGND sg13g2_mux2_1
X_0595_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame5_bit17.Q _0069_ _0195_ _0194_
+ sg13g2_a21oi_1
XFILLER_29_55 VPWR VGND sg13g2_fill_2
XANTENNA_8 VPWR VGND N4END[4] sg13g2_antennanp
X_0716_ _0303_ VPWR _0304_ VGND UO_OUT_TT_PROJECT1 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit13.Q
+ sg13g2_o21ai_1
X_1001_ FrameData[3] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit3.Q VPWR
+ VGND sg13g2_dlhq_1
X_0647_ _0241_ E6END[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit25.Q VPWR VGND sg13g2_nand2b_1
X_0578_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit25.Q VPWR _0180_ VGND Inst_E_TT_IF_ConfigMem.Inst_frame5_bit24.Q
+ _0179_ sg13g2_o21ai_1
XFILLER_40_126 VPWR VGND sg13g2_fill_1
X_0501_ Inst_E_TT_IF_ConfigMem.Inst_frame0_bit8.Q N2MID[0] N2END[0] S2MID[0] S2END[0]
+ Inst_E_TT_IF_ConfigMem.Inst_frame0_bit9.Q _0112_ VPWR VGND sg13g2_mux4_1
X_0432_ _0042_ VPWR RST_N_TT_PROJECT VGND _0049_ _0050_ sg13g2_o21ai_1
XFILLER_31_115 VPWR VGND sg13g2_decap_8
XFILLER_26_23 VPWR VGND sg13g2_fill_1
X_0981_ FrameData[15] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit15.Q VPWR
+ VGND sg13g2_dlhq_1
X_0415_ VPWR _0034_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit22.Q VGND sg13g2_inv_1
X_1180_ FrameData[21] FrameData_O[21] VPWR VGND sg13g2_buf_1
X_0895_ FrameData[25] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit25.Q VPWR
+ VGND sg13g2_dlhq_1
X_0964_ FrameData[30] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit30.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_5_199 VPWR VGND sg13g2_fill_1
X_1232_ N4END[5] N4BEG[1] VPWR VGND sg13g2_buf_1
X_1301_ Inst_E_TT_IF_switch_matrix.W2BEGb5 W2BEGb[5] VPWR VGND sg13g2_buf_1
X_0680_ _0271_ _0270_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit23.Q VPWR VGND sg13g2_nand2b_1
X_0878_ FrameData[8] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit8.Q VPWR
+ VGND sg13g2_dlhq_1
X_1094_ FrameData[0] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit0.Q VPWR
+ VGND sg13g2_dlhq_1
X_1163_ FrameData[4] FrameData_O[4] VPWR VGND sg13g2_buf_1
X_0947_ FrameData[13] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit13.Q VPWR
+ VGND sg13g2_dlhq_1
X_1146_ FrameData[20] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit20.Q VPWR
+ VGND sg13g2_dlhq_1
X_1215_ Inst_E_TT_IF_switch_matrix.N2BEG0 N2BEG[0] VPWR VGND sg13g2_buf_1
X_1077_ FrameData[15] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit15.Q VPWR
+ VGND sg13g2_dlhq_1
X_0801_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame8_bit14.Q _0372_ _0376_ _0375_
+ sg13g2_a21oi_1
X_0663_ _0255_ VPWR _0256_ VGND UO_OUT_TT_PROJECT5 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit28.Q
+ sg13g2_o21ai_1
X_0732_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit7.Q N1END[3] S1END[3] UO_OUT_TT_PROJECT1
+ UO_OUT_TT_PROJECT4 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit8.Q _0318_ VPWR VGND sg13g2_mux4_1
X_0594_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit17.Q UIO_OE_TT_PROJECT5 _0194_ VPWR
+ VGND sg13g2_nor2b_1
XFILLER_28_132 VPWR VGND sg13g2_decap_8
XANTENNA_9 VPWR VGND N4END[7] sg13g2_antennanp
X_1000_ FrameData[2] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit2.Q VPWR
+ VGND sg13g2_dlhq_1
X_0715_ VGND VPWR _0028_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit13.Q _0303_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit14.Q
+ sg13g2_a21oi_1
X_1129_ FrameData[3] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit3.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_25_113 VPWR VGND sg13g2_fill_1
X_0646_ N1END[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit24.Q Inst_E_TT_IF_ConfigMem.Inst_frame0_bit25.Q
+ _0240_ VPWR VGND sg13g2_nor3_1
X_0577_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame5_bit23.Q _0051_ _0179_ _0178_
+ sg13g2_a21oi_1
X_0431_ _0050_ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit7.Q _0045_ VPWR VGND sg13g2_nand2_1
X_0500_ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit24.Q N1END[0] N4END[0] S1END[0] S4END[0]
+ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit25.Q _0111_ VPWR VGND sg13g2_mux4_1
X_0629_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame5_bit5.Q _0062_ _0225_ _0224_ sg13g2_a21oi_1
XFILLER_22_149 VPWR VGND sg13g2_fill_1
XFILLER_21_160 VPWR VGND sg13g2_fill_2
X_0414_ VPWR _0033_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit25.Q VGND sg13g2_inv_1
X_0980_ FrameData[14] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit14.Q VPWR
+ VGND sg13g2_dlhq_1
X_0894_ FrameData[24] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit24.Q VPWR
+ VGND sg13g2_dlhq_1
X_0963_ FrameData[29] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit29.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_13_91 VPWR VGND sg13g2_fill_1
XFILLER_49_163 VPWR VGND sg13g2_fill_2
X_1231_ N4END[4] N4BEG[0] VPWR VGND sg13g2_buf_1
X_0877_ FrameData[7] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit7.Q VPWR
+ VGND sg13g2_dlhq_1
X_1093_ FrameData[31] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit31.Q VPWR
+ VGND sg13g2_dlhq_1
X_1162_ FrameData[3] FrameData_O[3] VPWR VGND sg13g2_buf_1
X_0946_ FrameData[12] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit12.Q VPWR
+ VGND sg13g2_dlhq_1
X_1300_ Inst_E_TT_IF_switch_matrix.W2BEGb4 W2BEGb[4] VPWR VGND sg13g2_buf_1
X_1145_ FrameData[19] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit19.Q VPWR
+ VGND sg13g2_dlhq_1
X_1214_ Inst_E_TT_IF_switch_matrix.N1BEG3 N1BEG[3] VPWR VGND sg13g2_buf_1
XFILLER_37_199 VPWR VGND sg13g2_fill_1
X_0800_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit15.Q VPWR _0375_ VGND Inst_E_TT_IF_ConfigMem.Inst_frame8_bit14.Q
+ _0374_ sg13g2_o21ai_1
X_0662_ VGND VPWR _0023_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit28.Q _0255_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit29.Q
+ sg13g2_a21oi_1
X_0731_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit7.Q UIO_OE_TT_PROJECT1 UIO_OE_TT_PROJECT3
+ UIO_OE_TT_PROJECT4 UIO_OE_TT_PROJECT7 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit8.Q
+ _0317_ VPWR VGND sg13g2_mux4_1
X_0593_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame5_bit17.Q _0071_ _0193_ _0192_
+ sg13g2_a21oi_1
X_0929_ FrameData[27] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit27.Q VPWR
+ VGND sg13g2_dlhq_1
X_1076_ FrameData[14] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit14.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_19_111 VPWR VGND sg13g2_fill_1
X_1059_ FrameData[29] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit29.Q VPWR
+ VGND sg13g2_dlhq_1
X_1128_ FrameData[2] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit2.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_25_169 VPWR VGND sg13g2_fill_2
X_0714_ _0301_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit15.Q _0302_ VPWR VGND sg13g2_nor2b_1
X_0576_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit23.Q UIO_OE_TT_PROJECT7 _0178_ VPWR
+ VGND sg13g2_nor2b_1
X_0645_ _0237_ _0239_ Inst_E_TT_IF_switch_matrix.W2BEGb0 VPWR VGND sg13g2_nor2_1
X_0430_ VGND VPWR _0047_ _0048_ _0049_ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit4.Q sg13g2_a21oi_1
X_0628_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit6.Q VPWR _0224_ VGND Inst_E_TT_IF_ConfigMem.Inst_frame5_bit5.Q
+ _0104_ sg13g2_o21ai_1
X_0559_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit23.Q _0104_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit22.Q
+ _0163_ VPWR VGND sg13g2_nand3_1
X_0413_ VPWR _0032_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit26.Q VGND sg13g2_inv_1
XFILLER_27_90 VPWR VGND sg13g2_fill_1
X_0893_ FrameData[23] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit23.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_23_48 VPWR VGND sg13g2_fill_2
X_0962_ FrameData[28] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit28.Q VPWR
+ VGND sg13g2_dlhq_1
X_0876_ FrameData[6] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit6.Q VPWR
+ VGND sg13g2_dlhq_1
X_1230_ N2MID[7] N2BEGb[7] VPWR VGND sg13g2_buf_1
X_1092_ FrameData[30] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit30.Q VPWR
+ VGND sg13g2_dlhq_1
X_1161_ FrameData[2] FrameData_O[2] VPWR VGND sg13g2_buf_1
X_0945_ FrameData[11] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit11.Q VPWR
+ VGND sg13g2_dlhq_1
X_1213_ Inst_E_TT_IF_switch_matrix.N1BEG2 N1BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_24_80 VPWR VGND sg13g2_fill_1
X_0661_ _0247_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit30.Q _0254_ VPWR VGND sg13g2_nor2b_1
X_0730_ Inst_E_TT_IF_switch_matrix.W2BEG0 _0314_ _0316_ _0312_ _0311_ VPWR VGND sg13g2_a22oi_1
X_0592_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit18.Q VPWR _0192_ VGND Inst_E_TT_IF_ConfigMem.Inst_frame5_bit17.Q
+ _0096_ sg13g2_o21ai_1
X_1144_ FrameData[18] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit18.Q VPWR
+ VGND sg13g2_dlhq_1
X_0928_ FrameData[26] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit26.Q VPWR
+ VGND sg13g2_dlhq_1
X_1075_ FrameData[13] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit13.Q VPWR
+ VGND sg13g2_dlhq_1
X_0859_ Inst_E_TT_IF_ConfigMem.Inst_frame9_bit22.Q E1END[0] E6END[4] _0078_ _0242_
+ Inst_E_TT_IF_ConfigMem.Inst_frame9_bit23.Q Inst_E_TT_IF_switch_matrix.N1BEG0 VPWR
+ VGND sg13g2_mux4_1
XFILLER_19_167 VPWR VGND sg13g2_fill_1
X_1058_ FrameData[28] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit28.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_25_104 VPWR VGND sg13g2_decap_8
X_1127_ FrameData[1] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit1.Q VPWR
+ VGND sg13g2_dlhq_1
X_0644_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit4.Q _0238_ _0239_ VPWR VGND sg13g2_nor2_1
X_0713_ VGND VPWR _0299_ _0300_ _0301_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit14.Q
+ sg13g2_a21oi_1
X_0575_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame5_bit23.Q _0053_ _0177_ _0176_
+ sg13g2_a21oi_1
X_0489_ _0102_ _0101_ _0012_ _0099_ _0095_ VPWR VGND sg13g2_a22oi_1
X_0558_ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit10.Q N1END[1] N4END[1] S1END[1] S4END[1]
+ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit11.Q _0162_ VPWR VGND sg13g2_mux4_1
X_0627_ _0221_ _0223_ Inst_E_TT_IF_switch_matrix.W2BEGb2 VPWR VGND sg13g2_nor2_1
X_0412_ VPWR _0031_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit29.Q VGND sg13g2_inv_1
X_0892_ FrameData[22] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit22.Q VPWR
+ VGND sg13g2_dlhq_1
X_0961_ FrameData[27] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit27.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_48_79 VPWR VGND sg13g2_fill_1
X_1091_ FrameData[29] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit29.Q VPWR
+ VGND sg13g2_dlhq_1
X_1160_ FrameData[1] FrameData_O[1] VPWR VGND sg13g2_buf_1
XFILLER_1_172 VPWR VGND sg13g2_fill_2
X_0944_ FrameData[10] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit10.Q VPWR
+ VGND sg13g2_dlhq_1
X_0875_ FrameData[5] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit5.Q VPWR
+ VGND sg13g2_dlhq_1
X_1289_ Inst_E_TT_IF_switch_matrix.W2BEG1 W2BEG[1] VPWR VGND sg13g2_buf_1
X_0591_ _0189_ _0191_ Inst_E_TT_IF_switch_matrix.W2BEGb6 VPWR VGND sg13g2_nor2_1
X_0660_ _0251_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit28.Q _0252_ _0253_ VPWR VGND
+ sg13g2_a21o_1
X_1143_ FrameData[17] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit17.Q VPWR
+ VGND sg13g2_dlhq_1
X_0927_ FrameData[25] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit25.Q VPWR
+ VGND sg13g2_dlhq_1
X_1212_ Inst_E_TT_IF_switch_matrix.N1BEG1 N1BEG[1] VPWR VGND sg13g2_buf_1
X_0789_ _0104_ _0162_ _0035_ _0365_ VPWR VGND sg13g2_mux2_1
XFILLER_37_146 VPWR VGND sg13g2_fill_2
X_0858_ Inst_E_TT_IF_ConfigMem.Inst_frame9_bit24.Q E1END[1] E6END[5] _0069_ _0250_
+ Inst_E_TT_IF_ConfigMem.Inst_frame9_bit25.Q Inst_E_TT_IF_switch_matrix.N1BEG1 VPWR
+ VGND sg13g2_mux4_1
X_1074_ FrameData[12] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit12.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_29_37 VPWR VGND sg13g2_fill_1
X_1126_ FrameData[0] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit0.Q VPWR
+ VGND sg13g2_dlhq_1
X_0574_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit24.Q VPWR _0176_ VGND Inst_E_TT_IF_ConfigMem.Inst_frame5_bit23.Q
+ _0112_ sg13g2_o21ai_1
X_0643_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit2.Q E2END[7] UIO_OUT_TT_PROJECT0 UIO_OUT_TT_PROJECT3
+ UIO_OUT_TT_PROJECT7 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit3.Q _0238_ VPWR VGND sg13g2_mux4_1
X_0712_ _0300_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit13.Q _0104_ VPWR VGND sg13g2_nand2_1
X_1057_ FrameData[27] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit27.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_21_93 VPWR VGND sg13g2_decap_8
X_0488_ E2END[2] EE4END[10] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit17.Q _0101_ VPWR
+ VGND sg13g2_mux2_1
X_0557_ UI_IN_TT_PROJECT2 _0161_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit24.Q _0159_
+ _0156_ VPWR VGND sg13g2_a22oi_1
X_1109_ FrameData[15] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit15.Q VPWR
+ VGND sg13g2_dlhq_1
X_0626_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit10.Q _0222_ _0223_ VPWR VGND sg13g2_nor2_1
XFILLER_16_71 VPWR VGND sg13g2_fill_1
X_0411_ VPWR _0030_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit10.Q VGND sg13g2_inv_1
X_0609_ _0205_ _0207_ Inst_E_TT_IF_switch_matrix.W2BEGb4 VPWR VGND sg13g2_nor2_1
X_0891_ FrameData[21] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit21.Q VPWR
+ VGND sg13g2_dlhq_1
X_0960_ FrameData[26] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit26.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_48_58 VPWR VGND sg13g2_fill_1
XFILLER_49_188 VPWR VGND sg13g2_fill_2
X_1090_ FrameData[28] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit28.Q VPWR
+ VGND sg13g2_dlhq_1
X_0874_ FrameData[4] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit4.Q VPWR
+ VGND sg13g2_dlhq_1
X_1288_ Inst_E_TT_IF_switch_matrix.W2BEG0 W2BEG[0] VPWR VGND sg13g2_buf_1
X_0943_ FrameData[9] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit9.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_46_125 VPWR VGND sg13g2_fill_1
XFILLER_24_71 VPWR VGND sg13g2_decap_8
X_0857_ Inst_E_TT_IF_ConfigMem.Inst_frame9_bit26.Q E1END[2] E6END[6] _0060_ _0263_
+ Inst_E_TT_IF_ConfigMem.Inst_frame9_bit27.Q Inst_E_TT_IF_switch_matrix.N1BEG2 VPWR
+ VGND sg13g2_mux4_1
X_0926_ FrameData[24] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit24.Q VPWR
+ VGND sg13g2_dlhq_1
X_1211_ Inst_E_TT_IF_switch_matrix.N1BEG0 N1BEG[0] VPWR VGND sg13g2_buf_1
X_1142_ FrameData[16] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit16.Q VPWR
+ VGND sg13g2_dlhq_1
X_0590_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit22.Q _0190_ _0191_ VPWR VGND sg13g2_nor2_1
X_1073_ FrameData[11] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit11.Q VPWR
+ VGND sg13g2_dlhq_1
X_0788_ VGND VPWR _0362_ _0364_ Inst_E_TT_IF_switch_matrix.N4BEG2 _0360_ sg13g2_a21oi_1
X_0573_ UI_IN_TT_PROJECT0 _0175_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit18.Q _0173_
+ _0170_ VPWR VGND sg13g2_a22oi_1
XFILLER_19_147 VPWR VGND sg13g2_fill_2
XFILLER_19_93 VPWR VGND sg13g2_fill_1
X_0642_ _0233_ _0236_ _0237_ VPWR VGND sg13g2_nor2_1
X_0711_ _0299_ _0162_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit13.Q VPWR VGND sg13g2_nand2b_1
X_1056_ FrameData[26] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit26.Q VPWR
+ VGND sg13g2_dlhq_1
X_0909_ FrameData[7] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit7.Q VPWR
+ VGND sg13g2_dlhq_1
X_1125_ FrameData[31] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit31.Q VPWR
+ VGND sg13g2_dlhq_1
X_0487_ VPWR VGND E6END[10] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit16.Q _0099_ _0012_
+ _0100_ _0098_ sg13g2_a221oi_1
X_0556_ _0161_ _0160_ _0019_ _0158_ _0155_ VPWR VGND sg13g2_a22oi_1
XFILLER_30_0 VPWR VGND sg13g2_fill_2
X_0625_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit8.Q E2END[5] UIO_OUT_TT_PROJECT1 UIO_OUT_TT_PROJECT2
+ UIO_OUT_TT_PROJECT5 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit9.Q _0222_ VPWR VGND sg13g2_mux4_1
X_1039_ FrameData[9] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit9.Q VPWR
+ VGND sg13g2_dlhq_1
X_1108_ FrameData[14] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit14.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_21_175 VPWR VGND sg13g2_fill_1
XFILLER_8_113 VPWR VGND sg13g2_fill_1
XFILLER_8_135 VPWR VGND sg13g2_fill_1
XFILLER_8_179 VPWR VGND sg13g2_fill_2
X_0410_ VPWR _0029_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit18.Q VGND sg13g2_inv_1
X_0539_ E2END[4] EE4END[12] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit31.Q _0146_ VPWR
+ VGND sg13g2_mux2_1
X_0608_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit16.Q _0206_ _0207_ VPWR VGND sg13g2_nor2_1
X_0890_ FrameData[20] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit20.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_8_0 VPWR VGND sg13g2_fill_1
X_0873_ FrameData[3] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit3.Q VPWR
+ VGND sg13g2_dlhq_1
X_0942_ FrameData[8] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit8.Q VPWR
+ VGND sg13g2_dlhq_1
X_1287_ Inst_E_TT_IF_switch_matrix.W1BEG3 W1BEG[3] VPWR VGND sg13g2_buf_1
XFILLER_34_17 VPWR VGND sg13g2_fill_2
X_1141_ FrameData[15] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit15.Q VPWR
+ VGND sg13g2_dlhq_1
X_1210_ FrameStrobe[19] FrameStrobe_O[19] VPWR VGND sg13g2_buf_1
X_1072_ FrameData[10] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit10.Q VPWR
+ VGND sg13g2_dlhq_1
X_0787_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame8_bit20.Q _0363_ _0364_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit21.Q
+ sg13g2_a21oi_1
Xclkbuf_1_1__f_UserCLK clknet_0_UserCLK clknet_1_1__leaf_UserCLK VPWR VGND sg13g2_buf_8
X_0856_ Inst_E_TT_IF_ConfigMem.Inst_frame9_bit28.Q E1END[3] E6END[7] _0051_ _0274_
+ Inst_E_TT_IF_ConfigMem.Inst_frame9_bit29.Q Inst_E_TT_IF_switch_matrix.N1BEG3 VPWR
+ VGND sg13g2_mux4_1
X_0925_ FrameData[23] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit23.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_28_159 VPWR VGND sg13g2_fill_2
XFILLER_34_129 VPWR VGND sg13g2_fill_1
XFILLER_19_72 VPWR VGND sg13g2_fill_1
X_0641_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit4.Q VPWR _0236_ VGND Inst_E_TT_IF_ConfigMem.Inst_frame5_bit3.Q
+ _0235_ sg13g2_o21ai_1
X_0710_ _0251_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit13.Q _0297_ _0298_ VPWR VGND
+ sg13g2_a21o_1
X_1055_ FrameData[25] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit25.Q VPWR
+ VGND sg13g2_dlhq_1
X_0572_ _0175_ _0174_ _0021_ _0172_ _0169_ VPWR VGND sg13g2_a22oi_1
X_0908_ FrameData[6] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit6.Q VPWR
+ VGND sg13g2_dlhq_1
X_1124_ FrameData[30] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit30.Q VPWR
+ VGND sg13g2_dlhq_1
X_0839_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit11.Q E1END[0] E2END[3] E2MID[3] _0079_
+ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit10.Q Inst_E_TT_IF_switch_matrix.S2BEG4 VPWR
+ VGND sg13g2_mux4_1
X_0486_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit17.Q _0012_ _0099_ VPWR VGND sg13g2_nor2_1
X_0555_ E2END[2] EE4END[10] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit25.Q _0160_ VPWR
+ VGND sg13g2_mux2_1
X_0624_ _0217_ _0220_ _0221_ VPWR VGND sg13g2_nor2_1
X_1107_ FrameData[13] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit13.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_21_198 VPWR VGND sg13g2_fill_2
X_1038_ FrameData[8] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit8.Q VPWR
+ VGND sg13g2_dlhq_1
X_0538_ VPWR VGND E6END[4] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit30.Q _0144_ _0017_
+ _0145_ _0143_ sg13g2_a221oi_1
X_0469_ VPWR VGND EE4END[12] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit22.Q _0083_ _0010_
+ _0084_ _0082_ sg13g2_a221oi_1
X_0607_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit15.Q E2END[3] UIO_OUT_TT_PROJECT4 UIO_OUT_TT_PROJECT3
+ UIO_OUT_TT_PROJECT7 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit14.Q _0206_ VPWR VGND
+ sg13g2_mux4_1
X_0872_ FrameData[2] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit2.Q VPWR
+ VGND sg13g2_dlhq_1
X_0941_ FrameData[7] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit7.Q VPWR
+ VGND sg13g2_dlhq_1
X_1286_ Inst_E_TT_IF_switch_matrix.W1BEG2 W1BEG[2] VPWR VGND sg13g2_buf_1
X_1140_ FrameData[14] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit14.Q VPWR
+ VGND sg13g2_dlhq_1
X_1071_ FrameData[9] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit9.Q VPWR
+ VGND sg13g2_dlhq_1
X_1269_ S4END[6] S4BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_53_0 VPWR VGND sg13g2_fill_1
X_0786_ EE4END[2] _0095_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit22.Q _0363_ VPWR VGND
+ sg13g2_mux2_1
XFILLER_45_28 VPWR VGND sg13g2_fill_1
X_0924_ FrameData[22] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit22.Q VPWR
+ VGND sg13g2_dlhq_1
X_0855_ Inst_E_TT_IF_ConfigMem.Inst_frame9_bit30.Q E2MID[7] E2END[7] E6END[7] _0112_
+ Inst_E_TT_IF_ConfigMem.Inst_frame9_bit31.Q Inst_E_TT_IF_switch_matrix.N2BEG0 VPWR
+ VGND sg13g2_mux4_1
XFILLER_19_149 VPWR VGND sg13g2_fill_1
X_1123_ FrameData[29] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit29.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_51_71 VPWR VGND sg13g2_fill_2
X_1054_ FrameData[24] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit24.Q VPWR
+ VGND sg13g2_dlhq_1
X_0907_ FrameData[5] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit5.Q VPWR
+ VGND sg13g2_dlhq_1
X_0571_ E2END[0] EE4END[8] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit19.Q _0174_ VPWR
+ VGND sg13g2_mux2_1
XFILLER_18_171 VPWR VGND sg13g2_fill_1
X_0640_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame5_bit2.Q _0111_ _0235_ _0234_ sg13g2_a21oi_1
XANTENNA_70 VPWR VGND S2MID[6] sg13g2_antennanp
X_0769_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit18.Q E1END[0] EE4END[12] _0141_ _0111_
+ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit20.Q _0348_ VPWR VGND sg13g2_mux4_1
XFILLER_24_174 VPWR VGND sg13g2_fill_2
XFILLER_24_163 VPWR VGND sg13g2_fill_1
X_0838_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit12.Q E1END[1] E2MID[2] E2END[2] _0070_
+ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit13.Q Inst_E_TT_IF_switch_matrix.S2BEG5 VPWR
+ VGND sg13g2_mux4_1
X_0554_ VPWR VGND E6END[2] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit24.Q _0158_ _0019_
+ _0159_ _0157_ sg13g2_a221oi_1
XFILLER_30_133 VPWR VGND sg13g2_decap_4
X_0623_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit10.Q VPWR _0220_ VGND Inst_E_TT_IF_ConfigMem.Inst_frame5_bit9.Q
+ _0219_ sg13g2_o21ai_1
X_1106_ FrameData[12] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit12.Q VPWR
+ VGND sg13g2_dlhq_1
X_0485_ E2MID[2] EE4END[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit17.Q _0098_ VPWR
+ VGND sg13g2_mux2_1
XFILLER_21_100 VPWR VGND sg13g2_decap_8
X_1037_ FrameData[7] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit7.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_16_30 VPWR VGND sg13g2_fill_2
X_0399_ VPWR _0018_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit29.Q VGND sg13g2_inv_1
X_0537_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit31.Q _0017_ _0144_ VPWR VGND sg13g2_nor2_1
X_0468_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit23.Q _0010_ _0083_ VPWR VGND sg13g2_nor2_1
X_0606_ _0201_ _0204_ _0205_ VPWR VGND sg13g2_nor2_1
XFILLER_4_151 VPWR VGND sg13g2_fill_2
XFILLER_48_28 VPWR VGND sg13g2_fill_2
X_0871_ FrameData[1] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit1.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_38_83 VPWR VGND sg13g2_fill_2
X_0940_ FrameData[6] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit6.Q VPWR
+ VGND sg13g2_dlhq_1
X_1285_ Inst_E_TT_IF_switch_matrix.W1BEG1 W1BEG[1] VPWR VGND sg13g2_buf_1
X_1268_ S4END[5] S4BEG[1] VPWR VGND sg13g2_buf_1
X_0785_ _0361_ VPWR _0362_ VGND _0034_ _0127_ sg13g2_o21ai_1
X_0854_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit0.Q E2MID[6] E2END[6] E6END[6] _0104_
+ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit1.Q Inst_E_TT_IF_switch_matrix.N2BEG1 VPWR
+ VGND sg13g2_mux4_1
X_0923_ FrameData[21] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit21.Q VPWR
+ VGND sg13g2_dlhq_1
X_1070_ FrameData[8] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit8.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_28_139 VPWR VGND sg13g2_fill_2
XFILLER_1_34 VPWR VGND sg13g2_fill_2
XFILLER_51_153 VPWR VGND sg13g2_fill_1
X_1199_ FrameStrobe[8] FrameStrobe_O[8] VPWR VGND sg13g2_buf_1
X_1122_ FrameData[28] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit28.Q VPWR
+ VGND sg13g2_dlhq_1
X_1053_ FrameData[23] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit23.Q VPWR
+ VGND sg13g2_dlhq_1
X_0570_ VPWR VGND E6END[0] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit18.Q _0172_ _0021_
+ _0173_ _0171_ sg13g2_a221oi_1
X_0906_ FrameData[4] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit4.Q VPWR
+ VGND sg13g2_dlhq_1
X_0768_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit20.Q E6END[4] _0078_ _0169_ _0079_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit18.Q
+ _0347_ VPWR VGND sg13g2_mux4_1
X_0837_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit14.Q E1END[2] E2MID[1] E2END[1] _0061_
+ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit15.Q Inst_E_TT_IF_switch_matrix.S2BEG6 VPWR
+ VGND sg13g2_mux4_1
X_0699_ Inst_E_TT_IF_switch_matrix.W2BEG3 _0286_ _0288_ _0284_ _0283_ VPWR VGND sg13g2_a22oi_1
XANTENNA_60 VPWR VGND N2MID[5] sg13g2_antennanp
XANTENNA_71 VPWR VGND S2MID[6] sg13g2_antennanp
X_0484_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit18.Q _0096_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit17.Q
+ _0097_ VPWR VGND sg13g2_nand3_1
X_0553_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit25.Q _0019_ _0158_ VPWR VGND sg13g2_nor2_1
X_1105_ FrameData[11] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit11.Q VPWR
+ VGND sg13g2_dlhq_1
X_1036_ FrameData[6] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit6.Q VPWR
+ VGND sg13g2_dlhq_1
X_0622_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame5_bit8.Q _0095_ _0219_ _0218_ sg13g2_a21oi_1
X_0536_ E2MID[4] EE4END[4] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit31.Q _0143_ VPWR
+ VGND sg13g2_mux2_1
X_0467_ E1END[0] E2END[4] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit23.Q _0082_ VPWR VGND
+ sg13g2_mux2_1
X_0605_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit16.Q VPWR _0204_ VGND Inst_E_TT_IF_ConfigMem.Inst_frame5_bit15.Q
+ _0203_ sg13g2_o21ai_1
X_0398_ VPWR _0017_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit0.Q VGND sg13g2_inv_1
XFILLER_27_30 VPWR VGND sg13g2_fill_1
X_1019_ FrameData[21] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit21.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_4_78 VPWR VGND sg13g2_fill_1
X_0519_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit6.Q _0061_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit5.Q
+ _0128_ VPWR VGND sg13g2_nand3_1
X_0870_ FrameData[0] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit0.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_1_111 VPWR VGND sg13g2_fill_1
X_0999_ FrameData[1] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit1.Q VPWR
+ VGND sg13g2_dlhq_1
X_1284_ Inst_E_TT_IF_switch_matrix.W1BEG0 W1BEG[0] VPWR VGND sg13g2_buf_1
X_0784_ VGND VPWR _0004_ _0034_ _0361_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit20.Q
+ sg13g2_a21oi_1
X_0853_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit3.Q E2MID[5] E6END[5] E2END[5] _0096_
+ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit2.Q Inst_E_TT_IF_switch_matrix.N2BEG2 VPWR
+ VGND sg13g2_mux4_1
X_0922_ FrameData[20] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit20.Q VPWR
+ VGND sg13g2_dlhq_1
X_1267_ S4END[4] S4BEG[0] VPWR VGND sg13g2_buf_1
X_1198_ FrameStrobe[7] FrameStrobe_O[7] VPWR VGND sg13g2_buf_1
XFILLER_19_129 VPWR VGND sg13g2_fill_1
XFILLER_10_77 VPWR VGND sg13g2_fill_1
X_1052_ FrameData[22] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit22.Q VPWR
+ VGND sg13g2_dlhq_1
X_1121_ FrameData[27] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit27.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_18_140 VPWR VGND sg13g2_decap_8
X_0767_ _0346_ _0345_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit22.Q Inst_E_TT_IF_switch_matrix.S4BEG1
+ VPWR VGND sg13g2_mux2_1
X_0905_ FrameData[3] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit3.Q VPWR
+ VGND sg13g2_dlhq_1
X_1319_ Inst_E_TT_IF_switch_matrix.WW4BEG3 WW4BEG[3] VPWR VGND sg13g2_buf_1
X_0836_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit17.Q E1END[3] E2END[0] E2MID[0] _0052_
+ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit16.Q Inst_E_TT_IF_switch_matrix.S2BEG7 VPWR
+ VGND sg13g2_mux4_1
X_0698_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame6_bit20.Q _0287_ _0288_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit21.Q
+ sg13g2_a21oi_1
XANTENNA_72 VPWR VGND S2MID[6] sg13g2_antennanp
XANTENNA_61 VPWR VGND N4END[11] sg13g2_antennanp
Xclkbuf_1_0__f_UserCLK clknet_0_UserCLK clknet_1_0__leaf_UserCLK VPWR VGND sg13g2_buf_8
XANTENNA_50 VPWR VGND E6END[0] sg13g2_antennanp
XFILLER_24_176 VPWR VGND sg13g2_fill_1
X_0483_ Inst_E_TT_IF_ConfigMem.Inst_frame0_bit13.Q N2MID[2] S2MID[2] N2END[2] S2END[2]
+ Inst_E_TT_IF_ConfigMem.Inst_frame0_bit12.Q _0096_ VPWR VGND sg13g2_mux4_1
X_0552_ E2MID[2] EE4END[2] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit25.Q _0157_ VPWR
+ VGND sg13g2_mux2_1
X_1104_ FrameData[10] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit10.Q VPWR
+ VGND sg13g2_dlhq_1
X_1035_ FrameData[5] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit5.Q VPWR
+ VGND sg13g2_dlhq_1
X_0621_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit8.Q UIO_OE_TT_PROJECT2 _0218_ VPWR VGND
+ sg13g2_nor2b_1
X_0819_ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit26.Q N4END[0] S4END[0] _0087_ _0051_
+ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit27.Q Inst_E_TT_IF_switch_matrix.W6BEG0 VPWR
+ VGND sg13g2_mux4_1
XFILLER_7_183 VPWR VGND sg13g2_fill_2
X_0604_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame5_bit14.Q _0078_ _0203_ _0202_
+ sg13g2_a21oi_1
X_0397_ VPWR _0016_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit3.Q VGND sg13g2_inv_1
X_0535_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit0.Q _0079_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit31.Q
+ _0142_ VPWR VGND sg13g2_nand3_1
X_0466_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit24.Q _0079_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit23.Q
+ _0081_ VPWR VGND sg13g2_nand3_1
XFILLER_21_0 VPWR VGND sg13g2_fill_2
X_1018_ FrameData[20] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit20.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_4_197 VPWR VGND sg13g2_fill_2
X_0518_ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit20.Q N1END[2] N4END[2] S1END[2] S4END[2]
+ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit21.Q _0127_ VPWR VGND sg13g2_mux4_1
X_0449_ VPWR VGND EE4END[14] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit28.Q _0065_ _0006_
+ _0066_ _0064_ sg13g2_a221oi_1
X_1283_ clknet_1_1__leaf_UserCLK UserCLKo VPWR VGND sg13g2_buf_1
X_0998_ FrameData[0] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit0.Q VPWR
+ VGND sg13g2_dlhq_1
X_0783_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame8_bit20.Q _0356_ _0360_ _0359_
+ sg13g2_a21oi_1
X_0852_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit5.Q E2MID[4] E6END[4] E2END[4] _0088_
+ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit4.Q Inst_E_TT_IF_switch_matrix.N2BEG3 VPWR
+ VGND sg13g2_mux4_1
X_0921_ FrameData[19] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit19.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_51_199 VPWR VGND sg13g2_fill_1
X_1197_ FrameStrobe[6] FrameStrobe_O[6] VPWR VGND sg13g2_buf_1
X_1266_ S2MID[7] S2BEGb[7] VPWR VGND sg13g2_buf_1
XFILLER_42_199 VPWR VGND sg13g2_fill_1
XFILLER_51_0 VPWR VGND sg13g2_fill_2
X_1051_ FrameData[21] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit21.Q VPWR
+ VGND sg13g2_dlhq_1
X_0766_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit21.Q E1END[1] EE4END[13] _0134_ _0103_
+ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit23.Q _0346_ VPWR VGND sg13g2_mux4_1
XFILLER_33_199 VPWR VGND sg13g2_fill_1
X_1120_ FrameData[26] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit26.Q VPWR
+ VGND sg13g2_dlhq_1
X_0904_ FrameData[2] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit2.Q VPWR
+ VGND sg13g2_dlhq_1
X_0835_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit27.Q UO_OUT_TT_PROJECT0 _0051_ UIO_OE_TT_PROJECT4
+ _0052_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit26.Q Inst_E_TT_IF_switch_matrix.WW4BEG0
+ VPWR VGND sg13g2_mux4_1
X_0697_ UIO_OUT_TT_PROJECT3 UIO_OE_TT_PROJECT4 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit19.Q
+ _0287_ VPWR VGND sg13g2_mux2_1
X_1318_ Inst_E_TT_IF_switch_matrix.WW4BEG2 WW4BEG[2] VPWR VGND sg13g2_buf_1
XANTENNA_62 VPWR VGND N4END[12] sg13g2_antennanp
XANTENNA_40 VPWR VGND N2MID[2] sg13g2_antennanp
XFILLER_24_199 VPWR VGND sg13g2_fill_1
X_1249_ Inst_E_TT_IF_switch_matrix.S1BEG2 S1BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_2_90 VPWR VGND sg13g2_fill_1
XANTENNA_73 VPWR VGND S2MID[6] sg13g2_antennanp
XANTENNA_51 VPWR VGND E6END[0] sg13g2_antennanp
X_0482_ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit28.Q N1END[2] N4END[2] S1END[2] S4END[2]
+ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit29.Q _0095_ VPWR VGND sg13g2_mux4_1
X_0551_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit26.Q _0096_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit25.Q
+ _0156_ VPWR VGND sg13g2_nand3_1
X_1103_ FrameData[9] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit9.Q VPWR
+ VGND sg13g2_dlhq_1
X_0620_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame5_bit8.Q _0071_ _0217_ _0216_ sg13g2_a21oi_1
X_1034_ FrameData[4] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit4.Q VPWR
+ VGND sg13g2_dlhq_1
X_0749_ VGND VPWR _0001_ _0031_ _0331_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit27.Q
+ sg13g2_a21oi_1
X_0818_ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit28.Q N4END[1] S4END[1] _0095_ _0060_
+ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit29.Q Inst_E_TT_IF_switch_matrix.W6BEG1 VPWR
+ VGND sg13g2_mux4_1
XFILLER_32_54 VPWR VGND sg13g2_fill_2
X_0396_ VPWR _0015_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit6.Q VGND sg13g2_inv_1
X_0465_ VPWR _0080_ _0079_ VGND sg13g2_inv_1
X_0603_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit14.Q UIO_OE_TT_PROJECT4 _0202_ VPWR
+ VGND sg13g2_nor2b_1
X_0534_ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit16.Q N1END[0] N4END[0] S1END[0] S4END[0]
+ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit17.Q _0141_ VPWR VGND sg13g2_mux4_1
X_1017_ FrameData[19] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit19.Q VPWR
+ VGND sg13g2_dlhq_1
X_0517_ VGND VPWR _0122_ _0124_ UI_IN_TT_PROJECT7 _0126_ sg13g2_a21oi_1
X_0448_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit29.Q _0006_ _0065_ VPWR VGND sg13g2_nor2_1
X_1282_ Inst_E_TT_IF_switch_matrix.S4BEG3 S4BEG[15] VPWR VGND sg13g2_buf_1
X_0997_ FrameData[31] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit31.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_49_63 VPWR VGND sg13g2_fill_2
X_0920_ FrameData[18] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit18.Q VPWR
+ VGND sg13g2_dlhq_1
X_0782_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit21.Q VPWR _0359_ VGND Inst_E_TT_IF_ConfigMem.Inst_frame8_bit20.Q
+ _0358_ sg13g2_o21ai_1
X_0851_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit6.Q E2MID[3] E2END[3] E6END[3] _0079_
+ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit7.Q Inst_E_TT_IF_switch_matrix.N2BEG4 VPWR
+ VGND sg13g2_mux4_1
X_1196_ FrameStrobe[5] FrameStrobe_O[5] VPWR VGND sg13g2_buf_1
X_1265_ S2MID[6] S2BEGb[6] VPWR VGND sg13g2_buf_1
XFILLER_44_0 VPWR VGND sg13g2_fill_2
X_0765_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit23.Q E6END[5] _0069_ _0162_ _0070_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit21.Q
+ _0345_ VPWR VGND sg13g2_mux4_1
X_0903_ FrameData[1] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit1.Q VPWR
+ VGND sg13g2_dlhq_1
X_1050_ FrameData[20] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit20.Q VPWR
+ VGND sg13g2_dlhq_1
X_0834_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit29.Q UO_OUT_TT_PROJECT1 _0060_ UIO_OE_TT_PROJECT5
+ _0061_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit28.Q Inst_E_TT_IF_switch_matrix.WW4BEG1
+ VPWR VGND sg13g2_mux4_1
X_0696_ _0285_ VPWR _0286_ VGND UO_OUT_TT_PROJECT0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit19.Q
+ sg13g2_o21ai_1
XANTENNA_74 VPWR VGND S2MID[7] sg13g2_antennanp
XANTENNA_63 VPWR VGND N4END[5] sg13g2_antennanp
XANTENNA_52 VPWR VGND E6END[0] sg13g2_antennanp
X_1179_ FrameData[20] FrameData_O[20] VPWR VGND sg13g2_buf_1
XANTENNA_41 VPWR VGND N2MID[4] sg13g2_antennanp
XANTENNA_30 VPWR VGND E2MID[2] sg13g2_antennanp
X_1248_ Inst_E_TT_IF_switch_matrix.S1BEG1 S1BEG[1] VPWR VGND sg13g2_buf_1
X_1317_ Inst_E_TT_IF_switch_matrix.WW4BEG1 WW4BEG[1] VPWR VGND sg13g2_buf_1
X_0550_ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit12.Q N1END[2] N4END[2] S1END[2] S4END[2]
+ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit13.Q _0155_ VPWR VGND sg13g2_mux4_1
X_0481_ UIO_IN_TT_PROJECT3 _0094_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit19.Q _0092_
+ _0089_ VPWR VGND sg13g2_a22oi_1
X_1102_ FrameData[8] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit8.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_15_101 VPWR VGND sg13g2_fill_2
XFILLER_16_4 VPWR VGND sg13g2_fill_1
X_0748_ _0326_ _0329_ _0330_ VPWR VGND sg13g2_nor2_1
X_0817_ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit30.Q N4END[2] S4END[2] _0103_ _0069_
+ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit31.Q Inst_E_TT_IF_switch_matrix.W6BEG2 VPWR
+ VGND sg13g2_mux4_1
X_1033_ FrameData[3] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit3.Q VPWR
+ VGND sg13g2_dlhq_1
X_0679_ _0141_ _0088_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit22.Q _0270_ VPWR VGND
+ sg13g2_mux2_1
XFILLER_16_89 VPWR VGND sg13g2_fill_1
X_0464_ Inst_E_TT_IF_ConfigMem.Inst_frame0_bit16.Q N2MID[4] N2END[4] S2MID[4] S2END[4]
+ Inst_E_TT_IF_ConfigMem.Inst_frame0_bit17.Q _0079_ VPWR VGND sg13g2_mux4_1
X_0533_ UI_IN_TT_PROJECT5 _0140_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit1.Q _0138_
+ _0135_ VPWR VGND sg13g2_a22oi_1
X_0395_ VPWR _0014_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit12.Q VGND sg13g2_inv_1
XFILLER_7_185 VPWR VGND sg13g2_fill_1
X_1016_ FrameData[18] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit18.Q VPWR
+ VGND sg13g2_dlhq_1
X_0602_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame5_bit14.Q _0080_ _0201_ _0200_
+ sg13g2_a21oi_1
XFILLER_4_199 VPWR VGND sg13g2_fill_1
X_0447_ E1END[2] E2END[6] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit29.Q _0064_ VPWR VGND
+ sg13g2_mux2_1
X_0516_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit9.Q _0125_ _0126_ VPWR VGND sg13g2_nor2_1
X_1281_ Inst_E_TT_IF_switch_matrix.S4BEG2 S4BEG[14] VPWR VGND sg13g2_buf_1
X_0996_ FrameData[30] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit30.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_24_78 VPWR VGND sg13g2_fill_2
X_1195_ FrameStrobe[4] FrameStrobe_O[4] VPWR VGND sg13g2_buf_1
X_0850_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit9.Q E2MID[2] E6END[2] E2END[2] _0070_
+ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit8.Q Inst_E_TT_IF_switch_matrix.N2BEG5 VPWR
+ VGND sg13g2_mux4_1
X_0781_ _0357_ VPWR _0358_ VGND _0034_ _0060_ sg13g2_o21ai_1
XFILLER_36_198 VPWR VGND sg13g2_fill_2
X_1264_ S2MID[5] S2BEGb[5] VPWR VGND sg13g2_buf_1
X_0979_ FrameData[13] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit13.Q VPWR
+ VGND sg13g2_dlhq_1
X_0902_ FrameData[0] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit0.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_18_198 VPWR VGND sg13g2_fill_2
XFILLER_4_0 VPWR VGND sg13g2_fill_1
X_0833_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit31.Q UO_OUT_TT_PROJECT2 _0069_ UIO_OE_TT_PROJECT6
+ _0070_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit30.Q Inst_E_TT_IF_switch_matrix.WW4BEG2
+ VPWR VGND sg13g2_mux4_1
X_1178_ FrameData[19] FrameData_O[19] VPWR VGND sg13g2_buf_1
XANTENNA_64 VPWR VGND S2MID[5] sg13g2_antennanp
X_0764_ VGND VPWR _0342_ _0344_ Inst_E_TT_IF_switch_matrix.S4BEG2 _0340_ sg13g2_a21oi_1
XANTENNA_42 VPWR VGND N2MID[4] sg13g2_antennanp
XFILLER_37_0 VPWR VGND sg13g2_fill_2
XANTENNA_53 VPWR VGND E6END[0] sg13g2_antennanp
XFILLER_24_102 VPWR VGND sg13g2_decap_4
XANTENNA_31 VPWR VGND E2MID[2] sg13g2_antennanp
XANTENNA_20 VPWR VGND S2MID[0] sg13g2_antennanp
X_1247_ Inst_E_TT_IF_switch_matrix.S1BEG0 S1BEG[0] VPWR VGND sg13g2_buf_1
XANTENNA_75 VPWR VGND S2MID[7] sg13g2_antennanp
X_0695_ VGND VPWR _0026_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit19.Q _0285_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit20.Q
+ sg13g2_a21oi_1
X_1316_ Inst_E_TT_IF_switch_matrix.WW4BEG0 WW4BEG[0] VPWR VGND sg13g2_buf_1
X_0480_ _0094_ _0093_ _0011_ _0091_ _0087_ VPWR VGND sg13g2_a22oi_1
X_1101_ FrameData[7] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit7.Q VPWR
+ VGND sg13g2_dlhq_1
X_0747_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit28.Q VPWR _0329_ VGND Inst_E_TT_IF_ConfigMem.Inst_frame7_bit27.Q
+ _0328_ sg13g2_o21ai_1
X_0816_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit0.Q N4END[3] S4END[3] _0111_ _0078_
+ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit1.Q Inst_E_TT_IF_switch_matrix.W6BEG3 VPWR
+ VGND sg13g2_mux4_1
X_0678_ Inst_E_TT_IF_switch_matrix.W2BEG5 _0267_ _0269_ _0265_ _0260_ VPWR VGND sg13g2_a22oi_1
X_1032_ FrameData[2] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit2.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_32_89 VPWR VGND sg13g2_fill_1
X_0394_ VPWR _0013_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit15.Q VGND sg13g2_inv_1
X_0532_ _0140_ _0139_ _0016_ _0137_ _0134_ VPWR VGND sg13g2_a22oi_1
X_0601_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit15.Q VPWR _0200_ VGND Inst_E_TT_IF_ConfigMem.Inst_frame5_bit14.Q
+ _0088_ sg13g2_o21ai_1
X_0463_ Inst_E_TT_IF_ConfigMem.Inst_frame0_bit0.Q N1END[0] N4END[0] S1END[0] S4END[0]
+ Inst_E_TT_IF_ConfigMem.Inst_frame0_bit1.Q _0078_ VPWR VGND sg13g2_mux4_1
X_1015_ FrameData[17] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit17.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_8_91 VPWR VGND sg13g2_fill_1
X_0446_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit30.Q _0061_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit29.Q
+ _0063_ VPWR VGND sg13g2_nand3_1
X_0515_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit7.Q E2MID[7] E2END[7] EE4END[7] EE4END[15]
+ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit8.Q _0125_ VPWR VGND sg13g2_mux4_1
X_0995_ FrameData[29] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit29.Q VPWR
+ VGND sg13g2_dlhq_1
X_1280_ Inst_E_TT_IF_switch_matrix.S4BEG1 S4BEG[13] VPWR VGND sg13g2_buf_1
X_0429_ _0048_ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit5.Q E2END[5] VPWR VGND sg13g2_nand2b_1
X_0780_ VGND VPWR _0357_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit22.Q E6END[10] sg13g2_or2_1
X_1194_ FrameStrobe[3] FrameStrobe_O[3] VPWR VGND sg13g2_buf_1
X_1263_ S2MID[4] S2BEGb[4] VPWR VGND sg13g2_buf_1
XFILLER_51_103 VPWR VGND sg13g2_fill_2
XFILLER_42_136 VPWR VGND sg13g2_fill_2
XFILLER_27_199 VPWR VGND sg13g2_fill_1
XFILLER_10_37 VPWR VGND sg13g2_fill_2
X_0978_ FrameData[12] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit12.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_18_133 VPWR VGND sg13g2_decap_8
X_1246_ Inst_E_TT_IF_switch_matrix.N4BEG3 N4BEG[15] VPWR VGND sg13g2_buf_1
X_1177_ FrameData[18] FrameData_O[18] VPWR VGND sg13g2_buf_1
X_0763_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame7_bit24.Q _0343_ _0344_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit25.Q
+ sg13g2_a21oi_1
XANTENNA_10 VPWR VGND N4END[8] sg13g2_antennanp
XANTENNA_43 VPWR VGND N2MID[4] sg13g2_antennanp
XANTENNA_21 VPWR VGND S2MID[1] sg13g2_antennanp
X_0901_ FrameData[31] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit31.Q VPWR
+ VGND sg13g2_dlhq_1
XANTENNA_32 VPWR VGND E2MID[2] sg13g2_antennanp
X_1315_ Inst_E_TT_IF_switch_matrix.W6BEG11 W6BEG[11] VPWR VGND sg13g2_buf_1
XANTENNA_54 VPWR VGND E6END[0] sg13g2_antennanp
X_0832_ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit1.Q UO_OUT_TT_PROJECT3 _0078_ UIO_OE_TT_PROJECT7
+ _0079_ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit0.Q Inst_E_TT_IF_switch_matrix.WW4BEG3
+ VPWR VGND sg13g2_mux4_1
XANTENNA_65 VPWR VGND S2MID[5] sg13g2_antennanp
X_0694_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame6_bit20.Q _0281_ _0284_ _0027_
+ sg13g2_a21oi_1
XANTENNA_76 VPWR VGND S2MID[2] sg13g2_antennanp
X_1100_ FrameData[6] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit6.Q VPWR
+ VGND sg13g2_dlhq_1
X_0746_ _0327_ VPWR _0328_ VGND _0031_ _0051_ sg13g2_o21ai_1
X_0815_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit3.Q UIO_OUT_TT_PROJECT4 _0087_ _0120_
+ _0112_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit2.Q Inst_E_TT_IF_switch_matrix.W6BEG4
+ VPWR VGND sg13g2_mux4_1
X_1031_ FrameData[1] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit1.Q VPWR
+ VGND sg13g2_dlhq_1
X_1229_ N2MID[6] N2BEGb[6] VPWR VGND sg13g2_buf_1
X_0677_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame6_bit26.Q _0268_ _0269_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit27.Q
+ sg13g2_a21oi_1
X_0393_ VPWR _0012_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit18.Q VGND sg13g2_inv_1
X_0531_ E2END[5] EE4END[13] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit2.Q _0139_ VPWR
+ VGND sg13g2_mux2_1
X_0462_ UIO_IN_TT_PROJECT5 _0077_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit25.Q _0075_
+ _0072_ VPWR VGND sg13g2_a22oi_1
X_0600_ _0197_ _0199_ Inst_E_TT_IF_switch_matrix.W2BEGb5 VPWR VGND sg13g2_nor2_1
X_1014_ FrameData[16] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit16.Q VPWR
+ VGND sg13g2_dlhq_1
X_0729_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame6_bit11.Q _0315_ _0316_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit12.Q
+ sg13g2_a21oi_1
X_0445_ VPWR _0062_ _0061_ VGND sg13g2_inv_1
X_0514_ _0124_ _0123_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit7.Q VPWR VGND sg13g2_nand2b_1
XFILLER_12_0 VPWR VGND sg13g2_fill_2
XFILLER_38_34 VPWR VGND sg13g2_fill_1
X_0994_ FrameData[28] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit28.Q VPWR
+ VGND sg13g2_dlhq_1
X_0428_ _0047_ _0046_ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit6.Q _0039_ _0000_ VPWR
+ VGND sg13g2_a22oi_1
X_1331_ Inst_E_TT_IF_switch_matrix.WW4BEG15 WW4BEG[15] VPWR VGND sg13g2_buf_1
X_1193_ FrameStrobe[2] FrameStrobe_O[2] VPWR VGND sg13g2_buf_1
X_1262_ S2MID[3] S2BEGb[3] VPWR VGND sg13g2_buf_1
X_0977_ FrameData[11] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit11.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_42_115 VPWR VGND sg13g2_fill_1
X_1245_ Inst_E_TT_IF_switch_matrix.N4BEG2 N4BEG[14] VPWR VGND sg13g2_buf_1
X_1176_ FrameData[17] FrameData_O[17] VPWR VGND sg13g2_buf_1
X_0762_ EE4END[14] _0095_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit26.Q _0343_ VPWR VGND
+ sg13g2_mux2_1
X_0900_ FrameData[30] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit30.Q VPWR
+ VGND sg13g2_dlhq_1
X_1314_ Inst_E_TT_IF_switch_matrix.W6BEG10 W6BEG[10] VPWR VGND sg13g2_buf_1
X_0831_ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit3.Q UO_OUT_TT_PROJECT4 _0087_ UIO_OE_TT_PROJECT0
+ _0088_ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit2.Q Inst_E_TT_IF_switch_matrix.WW4BEG4
+ VPWR VGND sg13g2_mux4_1
X_0693_ _0283_ _0282_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit20.Q VPWR VGND sg13g2_nand2b_1
XANTENNA_66 VPWR VGND S2MID[5] sg13g2_antennanp
XANTENNA_11 VPWR VGND N4END[9] sg13g2_antennanp
XFILLER_46_89 VPWR VGND sg13g2_fill_2
XANTENNA_55 VPWR VGND E6END[0] sg13g2_antennanp
XANTENNA_33 VPWR VGND E2MID[2] sg13g2_antennanp
XANTENNA_44 VPWR VGND N2MID[4] sg13g2_antennanp
XANTENNA_22 VPWR VGND S2MID[1] sg13g2_antennanp
XANTENNA_77 VPWR VGND S2MID[2] sg13g2_antennanp
XFILLER_15_137 VPWR VGND sg13g2_fill_1
XFILLER_21_107 VPWR VGND sg13g2_fill_2
X_0814_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit5.Q UIO_OUT_TT_PROJECT5 _0095_ _0127_
+ _0104_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit4.Q Inst_E_TT_IF_switch_matrix.W6BEG5
+ VPWR VGND sg13g2_mux4_1
X_1030_ FrameData[0] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit0.Q VPWR
+ VGND sg13g2_dlhq_1
X_1228_ N2MID[5] N2BEGb[5] VPWR VGND sg13g2_buf_1
XFILLER_42_0 VPWR VGND sg13g2_fill_1
X_0745_ VGND VPWR _0327_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit29.Q E6END[7] sg13g2_or2_1
X_1159_ FrameData[0] FrameData_O[0] VPWR VGND sg13g2_buf_1
X_0676_ UIO_OUT_TT_PROJECT5 UIO_OE_TT_PROJECT2 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit25.Q
+ _0268_ VPWR VGND sg13g2_mux2_1
X_0530_ VPWR VGND E6END[5] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit1.Q _0137_ _0016_
+ _0138_ _0136_ sg13g2_a221oi_1
X_0392_ VPWR _0011_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit21.Q VGND sg13g2_inv_1
X_0461_ _0077_ _0076_ _0008_ _0074_ _0069_ VPWR VGND sg13g2_a22oi_1
X_0659_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit29.Q VPWR _0252_ VGND Inst_E_TT_IF_ConfigMem.Inst_frame6_bit28.Q
+ _0061_ sg13g2_o21ai_1
X_0728_ UIO_OUT_TT_PROJECT0 UIO_OE_TT_PROJECT7 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit10.Q
+ _0315_ VPWR VGND sg13g2_mux2_1
X_1013_ FrameData[15] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit15.Q VPWR
+ VGND sg13g2_dlhq_1
X_0444_ Inst_E_TT_IF_ConfigMem.Inst_frame0_bit20.Q N2MID[6] N2END[6] S2MID[6] S2END[6]
+ Inst_E_TT_IF_ConfigMem.Inst_frame0_bit21.Q _0061_ VPWR VGND sg13g2_mux4_1
X_0513_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame2_bit8.Q _0053_ _0123_ _0119_ sg13g2_a21oi_1
X_0993_ FrameData[27] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit27.Q VPWR
+ VGND sg13g2_dlhq_1
X_0427_ _0046_ S2END[2] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit5.Q VPWR VGND sg13g2_nand2b_1
XFILLER_39_198 VPWR VGND sg13g2_fill_2
X_1192_ FrameStrobe[1] FrameStrobe_O[1] VPWR VGND sg13g2_buf_1
X_1261_ S2MID[2] S2BEGb[2] VPWR VGND sg13g2_buf_1
X_0976_ FrameData[10] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit10.Q VPWR
+ VGND sg13g2_dlhq_1
X_1330_ Inst_E_TT_IF_switch_matrix.WW4BEG14 WW4BEG[14] VPWR VGND sg13g2_buf_1
XFILLER_50_193 VPWR VGND sg13g2_fill_1
XFILLER_27_135 VPWR VGND sg13g2_decap_4
X_1244_ Inst_E_TT_IF_switch_matrix.N4BEG1 N4BEG[13] VPWR VGND sg13g2_buf_1
X_0761_ _0341_ VPWR _0342_ VGND _0032_ _0127_ sg13g2_o21ai_1
XFILLER_25_80 VPWR VGND sg13g2_fill_2
X_1313_ Inst_E_TT_IF_switch_matrix.W6BEG9 W6BEG[9] VPWR VGND sg13g2_buf_1
X_0830_ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit5.Q UO_OUT_TT_PROJECT5 _0095_ UIO_OE_TT_PROJECT1
+ _0096_ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit4.Q Inst_E_TT_IF_switch_matrix.WW4BEG5
+ VPWR VGND sg13g2_mux4_1
X_0692_ _0148_ _0088_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit19.Q _0282_ VPWR VGND
+ sg13g2_mux2_1
X_1175_ FrameData[16] FrameData_O[16] VPWR VGND sg13g2_buf_1
XANTENNA_45 VPWR VGND N4END[13] sg13g2_antennanp
XANTENNA_56 VPWR VGND FrameStrobe[18] sg13g2_antennanp
XANTENNA_12 VPWR VGND S2MID[0] sg13g2_antennanp
XANTENNA_23 VPWR VGND S2MID[1] sg13g2_antennanp
XANTENNA_34 VPWR VGND E2MID[2] sg13g2_antennanp
XANTENNA_67 VPWR VGND S2MID[5] sg13g2_antennanp
X_0959_ FrameData[25] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit25.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_2_0 VPWR VGND sg13g2_fill_2
X_1227_ N2MID[4] N2BEGb[4] VPWR VGND sg13g2_buf_1
X_0744_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame7_bit29.Q _0053_ _0326_ _0325_
+ sg13g2_a21oi_1
X_1158_ clknet_1_0__leaf_UserCLK CLK_TT_PROJECT VPWR VGND sg13g2_buf_1
X_1089_ FrameData[27] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit27.Q VPWR
+ VGND sg13g2_dlhq_1
X_0813_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit7.Q UIO_OUT_TT_PROJECT6 _0103_ _0134_
+ _0096_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit6.Q Inst_E_TT_IF_switch_matrix.W6BEG6
+ VPWR VGND sg13g2_mux4_1
X_0675_ _0266_ VPWR _0267_ VGND UO_OUT_TT_PROJECT5 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit25.Q
+ sg13g2_o21ai_1
X_0460_ E2MID[5] EE4END[5] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit26.Q _0076_ VPWR
+ VGND sg13g2_mux2_1
X_0391_ VPWR _0010_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit24.Q VGND sg13g2_inv_1
X_0727_ _0313_ VPWR _0314_ VGND UO_OUT_TT_PROJECT0 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit10.Q
+ sg13g2_o21ai_1
X_1012_ FrameData[14] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit14.Q VPWR
+ VGND sg13g2_dlhq_1
X_0658_ VPWR _0251_ _0250_ VGND sg13g2_inv_1
X_0589_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit20.Q E2END[1] UIO_OUT_TT_PROJECT1 UIO_OUT_TT_PROJECT5
+ UIO_OUT_TT_PROJECT6 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit21.Q _0190_ VPWR VGND
+ sg13g2_mux4_1
X_0443_ Inst_E_TT_IF_ConfigMem.Inst_frame0_bit4.Q N1END[2] N4END[2] S1END[2] S4END[2]
+ Inst_E_TT_IF_ConfigMem.Inst_frame0_bit5.Q _0060_ VPWR VGND sg13g2_mux4_1
X_0512_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit9.Q _0121_ _0122_ VPWR VGND sg13g2_and2_1
XFILLER_1_129 VPWR VGND sg13g2_fill_2
X_0426_ _0043_ _0044_ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit4.Q _0045_ VPWR VGND sg13g2_nand3_1
X_0992_ FrameData[26] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit26.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_49_57 VPWR VGND sg13g2_fill_2
XFILLER_40_48 VPWR VGND sg13g2_fill_2
X_1191_ FrameStrobe[0] FrameStrobe_O[0] VPWR VGND sg13g2_buf_1
X_1260_ S2MID[1] S2BEGb[1] VPWR VGND sg13g2_buf_1
X_0975_ FrameData[9] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit9.Q VPWR
+ VGND sg13g2_dlhq_1
X_0409_ VPWR _0028_ UO_OUT_TT_PROJECT2 VGND sg13g2_inv_1
X_0760_ VGND VPWR _0004_ _0032_ _0341_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit24.Q
+ sg13g2_a21oi_1
XFILLER_18_169 VPWR VGND sg13g2_fill_2
XFILLER_18_147 VPWR VGND sg13g2_fill_1
X_0691_ _0079_ _0274_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit19.Q _0281_ VPWR VGND
+ sg13g2_mux2_1
X_1174_ FrameData[15] FrameData_O[15] VPWR VGND sg13g2_buf_1
XANTENNA_68 VPWR VGND S2MID[4] sg13g2_antennanp
XANTENNA_57 VPWR VGND FrameStrobe[19] sg13g2_antennanp
X_1243_ Inst_E_TT_IF_switch_matrix.N4BEG0 N4BEG[12] VPWR VGND sg13g2_buf_1
X_0889_ FrameData[19] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit19.Q VPWR
+ VGND sg13g2_dlhq_1
XANTENNA_13 VPWR VGND S2MID[0] sg13g2_antennanp
XANTENNA_46 VPWR VGND N4END[15] sg13g2_antennanp
XFILLER_24_106 VPWR VGND sg13g2_fill_2
X_1312_ Inst_E_TT_IF_switch_matrix.W6BEG8 W6BEG[8] VPWR VGND sg13g2_buf_1
XANTENNA_35 VPWR VGND E2MID[2] sg13g2_antennanp
XANTENNA_24 VPWR VGND S2MID[1] sg13g2_antennanp
X_0958_ FrameData[24] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit24.Q VPWR
+ VGND sg13g2_dlhq_1
X_1226_ N2MID[3] N2BEGb[3] VPWR VGND sg13g2_buf_1
X_1157_ FrameData[31] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit31.Q VPWR
+ VGND sg13g2_dlhq_1
X_0743_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit27.Q VPWR _0325_ VGND Inst_E_TT_IF_ConfigMem.Inst_frame7_bit29.Q
+ _0148_ sg13g2_o21ai_1
X_0674_ VGND VPWR _0023_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit25.Q _0266_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit26.Q
+ sg13g2_a21oi_1
X_0812_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit9.Q UIO_OUT_TT_PROJECT7 _0111_ _0141_
+ _0088_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit8.Q Inst_E_TT_IF_switch_matrix.W6BEG7
+ VPWR VGND sg13g2_mux4_1
X_1088_ FrameData[26] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit26.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_20_197 VPWR VGND sg13g2_fill_2
X_0390_ VPWR _0009_ S1END[0] VGND sg13g2_inv_1
X_1011_ FrameData[13] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit13.Q VPWR
+ VGND sg13g2_dlhq_1
X_1209_ FrameStrobe[18] FrameStrobe_O[18] VPWR VGND sg13g2_buf_1
X_0657_ VPWR VGND Inst_E_TT_IF_ConfigMem.Inst_frame0_bit26.Q _0248_ _0249_ _0007_
+ _0250_ Inst_E_TT_IF_ConfigMem.Inst_frame0_bit27.Q sg13g2_a221oi_1
X_0588_ _0185_ _0188_ _0189_ VPWR VGND sg13g2_nor2_1
X_0726_ VGND VPWR _0026_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit10.Q _0313_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit11.Q
+ sg13g2_a21oi_1
X_0511_ _0120_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit7.Q _0121_ VPWR VGND Inst_E_TT_IF_ConfigMem.Inst_frame2_bit8.Q
+ sg13g2_nand3b_1
X_0442_ UIO_IN_TT_PROJECT7 _0059_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit31.Q _0057_
+ _0054_ VPWR VGND sg13g2_a22oi_1
X_0709_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit14.Q VPWR _0297_ VGND Inst_E_TT_IF_ConfigMem.Inst_frame6_bit13.Q
+ _0061_ sg13g2_o21ai_1
X_0425_ _0044_ _0039_ E2END[4] S2END[3] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit6.Q
+ VPWR VGND sg13g2_a22oi_1
XFILLER_5_85 VPWR VGND sg13g2_fill_1
X_0991_ FrameData[25] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit25.Q VPWR
+ VGND sg13g2_dlhq_1
X_1190_ FrameData[31] FrameData_O[31] VPWR VGND sg13g2_buf_1
XFILLER_35_49 VPWR VGND sg13g2_fill_2
X_0974_ FrameData[8] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit8.Q VPWR
+ VGND sg13g2_dlhq_1
X_0408_ VPWR _0027_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit21.Q VGND sg13g2_inv_1
XFILLER_25_82 VPWR VGND sg13g2_fill_1
X_0690_ Inst_E_TT_IF_switch_matrix.W2BEG4 _0278_ _0280_ _0276_ _0271_ VPWR VGND sg13g2_a22oi_1
X_1173_ FrameData[14] FrameData_O[14] VPWR VGND sg13g2_buf_1
XANTENNA_25 VPWR VGND E2MID[2] sg13g2_antennanp
X_1242_ N4END[15] N4BEG[11] VPWR VGND sg13g2_buf_1
X_0888_ FrameData[18] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit18.Q VPWR
+ VGND sg13g2_dlhq_1
XANTENNA_58 VPWR VGND N2MID[5] sg13g2_antennanp
XANTENNA_47 VPWR VGND E6END[0] sg13g2_antennanp
XANTENNA_36 VPWR VGND E2MID[2] sg13g2_antennanp
XANTENNA_69 VPWR VGND S2MID[4] sg13g2_antennanp
XANTENNA_14 VPWR VGND S2MID[0] sg13g2_antennanp
X_0957_ FrameData[23] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit23.Q VPWR
+ VGND sg13g2_dlhq_1
X_1311_ Inst_E_TT_IF_switch_matrix.W6BEG7 W6BEG[7] VPWR VGND sg13g2_buf_1
XFILLER_23_140 VPWR VGND sg13g2_fill_1
X_0811_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit11.Q UIO_OUT_TT_PROJECT0 _0120_ _0148_
+ _0079_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit10.Q Inst_E_TT_IF_switch_matrix.W6BEG8
+ VPWR VGND sg13g2_mux4_1
X_0742_ _0324_ _0323_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit0.Q Inst_E_TT_IF_switch_matrix.W1BEG0
+ VPWR VGND sg13g2_mux2_1
X_0673_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame6_bit26.Q _0264_ _0265_ _0024_
+ sg13g2_a21oi_1
X_1225_ N2MID[2] N2BEGb[2] VPWR VGND sg13g2_buf_1
X_1156_ FrameData[30] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit30.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_32_17 VPWR VGND sg13g2_fill_2
X_1087_ FrameData[25] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit25.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_22_94 VPWR VGND sg13g2_decap_4
XFILLER_22_72 VPWR VGND sg13g2_fill_1
X_1010_ FrameData[12] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit12.Q VPWR
+ VGND sg13g2_dlhq_1
X_1208_ FrameStrobe[17] FrameStrobe_O[17] VPWR VGND sg13g2_buf_1
X_1139_ FrameData[13] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit13.Q VPWR
+ VGND sg13g2_dlhq_1
X_0656_ _0249_ E6END[1] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit27.Q VPWR VGND sg13g2_nand2b_1
X_0587_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit22.Q VPWR _0188_ VGND Inst_E_TT_IF_ConfigMem.Inst_frame5_bit21.Q
+ _0187_ sg13g2_o21ai_1
X_0725_ _0309_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit12.Q _0312_ VPWR VGND sg13g2_nor2b_1
X_0441_ _0059_ _0058_ _0003_ _0056_ _0051_ VPWR VGND sg13g2_a22oi_1
X_0510_ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit22.Q N1END[3] N4END[3] S1END[3] S4END[3]
+ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit23.Q _0120_ VPWR VGND sg13g2_mux4_1
X_0639_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit2.Q UIO_OE_TT_PROJECT0 _0234_ VPWR VGND
+ sg13g2_nor2b_1
X_0708_ Inst_E_TT_IF_switch_matrix.W2BEG2 _0294_ _0296_ _0292_ _0291_ VPWR VGND sg13g2_a22oi_1
X_0424_ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit5.Q VPWR _0043_ VGND Inst_E_TT_IF_ConfigMem.Inst_frame1_bit6.Q
+ S2MID[0] sg13g2_o21ai_1
X_0990_ FrameData[24] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit24.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_36_105 VPWR VGND sg13g2_fill_1
XFILLER_14_84 VPWR VGND sg13g2_fill_2
X_0973_ FrameData[7] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit7.Q VPWR
+ VGND sg13g2_dlhq_1
X_0407_ VPWR _0026_ UO_OUT_TT_PROJECT3 VGND sg13g2_inv_1
X_1241_ N4END[14] N4BEG[10] VPWR VGND sg13g2_buf_1
X_1172_ FrameData[13] FrameData_O[13] VPWR VGND sg13g2_buf_1
XANTENNA_59 VPWR VGND N2MID[5] sg13g2_antennanp
XANTENNA_37 VPWR VGND FrameStrobe[12] sg13g2_antennanp
XANTENNA_15 VPWR VGND S2MID[0] sg13g2_antennanp
XANTENNA_26 VPWR VGND E2MID[2] sg13g2_antennanp
XANTENNA_48 VPWR VGND E6END[0] sg13g2_antennanp
X_0956_ FrameData[22] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit22.Q VPWR
+ VGND sg13g2_dlhq_1
X_1310_ Inst_E_TT_IF_switch_matrix.W6BEG6 W6BEG[6] VPWR VGND sg13g2_buf_1
X_0887_ FrameData[17] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit17.Q VPWR
+ VGND sg13g2_dlhq_1
X_0810_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit13.Q UIO_OUT_TT_PROJECT1 _0127_ _0155_
+ _0070_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit12.Q Inst_E_TT_IF_switch_matrix.W6BEG9
+ VPWR VGND sg13g2_mux4_1
X_0741_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit30.Q N1END[0] S1END[0] UO_OUT_TT_PROJECT2
+ UO_OUT_TT_PROJECT7 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit31.Q _0324_ VPWR VGND sg13g2_mux4_1
X_0672_ _0070_ _0263_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit25.Q _0264_ VPWR VGND
+ sg13g2_mux2_1
XFILLER_14_185 VPWR VGND sg13g2_fill_1
X_1155_ FrameData[29] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit29.Q VPWR
+ VGND sg13g2_dlhq_1
X_1224_ N2MID[1] N2BEGb[1] VPWR VGND sg13g2_buf_1
X_1086_ FrameData[24] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit24.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_20_199 VPWR VGND sg13g2_fill_1
XFILLER_20_111 VPWR VGND sg13g2_decap_8
X_0939_ FrameData[5] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit5.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_0_0 VPWR VGND sg13g2_fill_2
XFILLER_11_100 VPWR VGND sg13g2_fill_1
X_1207_ FrameStrobe[16] FrameStrobe_O[16] VPWR VGND sg13g2_buf_1
X_0655_ N1END[1] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit26.Q Inst_E_TT_IF_ConfigMem.Inst_frame0_bit27.Q
+ _0248_ VPWR VGND sg13g2_nor3_1
X_0586_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame5_bit20.Q _0060_ _0187_ _0186_
+ sg13g2_a21oi_1
X_0724_ _0053_ _0030_ _0310_ _0311_ VPWR VGND sg13g2_a21o_1
X_1138_ FrameData[12] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit12.Q VPWR
+ VGND sg13g2_dlhq_1
X_1069_ FrameData[7] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit7.Q VPWR
+ VGND sg13g2_dlhq_1
X_0440_ E2MID[7] EE4END[7] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit0.Q _0058_ VPWR VGND
+ sg13g2_mux2_1
X_0569_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit19.Q _0021_ _0172_ VPWR VGND sg13g2_nor2_1
X_0707_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame6_bit17.Q _0295_ _0296_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit18.Q
+ sg13g2_a21oi_1
X_0638_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame5_bit2.Q _0053_ _0233_ _0232_ sg13g2_a21oi_1
XFILLER_44_71 VPWR VGND sg13g2_fill_1
XFILLER_0_198 VPWR VGND sg13g2_fill_2
X_0423_ _0041_ VPWR _0042_ VGND Inst_E_TT_IF_ConfigMem.Inst_frame1_bit6.Q _0040_ sg13g2_o21ai_1
X_0972_ FrameData[6] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit6.Q VPWR
+ VGND sg13g2_dlhq_1
X_0406_ VPWR _0025_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit24.Q VGND sg13g2_inv_1
X_1240_ N4END[13] N4BEG[9] VPWR VGND sg13g2_buf_1
X_1171_ FrameData[12] FrameData_O[12] VPWR VGND sg13g2_buf_1
XFILLER_25_73 VPWR VGND sg13g2_decap_8
XANTENNA_49 VPWR VGND E6END[0] sg13g2_antennanp
XANTENNA_38 VPWR VGND N2MID[2] sg13g2_antennanp
X_0886_ FrameData[16] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit16.Q VPWR
+ VGND sg13g2_dlhq_1
XANTENNA_16 VPWR VGND S2MID[0] sg13g2_antennanp
XFILLER_23_175 VPWR VGND sg13g2_fill_2
XANTENNA_27 VPWR VGND E2MID[2] sg13g2_antennanp
X_0955_ FrameData[21] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit21.Q VPWR
+ VGND sg13g2_dlhq_1
X_0740_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit30.Q UIO_OE_TT_PROJECT0 UIO_OE_TT_PROJECT2
+ UIO_OE_TT_PROJECT6 UIO_OE_TT_PROJECT7 Inst_E_TT_IF_ConfigMem.Inst_frame7_bit31.Q
+ _0323_ VPWR VGND sg13g2_mux4_1
XFILLER_11_42 VPWR VGND sg13g2_fill_1
X_0671_ VPWR VGND Inst_E_TT_IF_ConfigMem.Inst_frame0_bit28.Q _0262_ _0261_ _0005_
+ _0263_ Inst_E_TT_IF_ConfigMem.Inst_frame0_bit29.Q sg13g2_a221oi_1
X_1154_ FrameData[28] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit28.Q VPWR
+ VGND sg13g2_dlhq_1
X_1223_ N2MID[0] N2BEGb[0] VPWR VGND sg13g2_buf_1
X_0869_ FrameData[31] FrameStrobe[9] Inst_E_TT_IF_ConfigMem.Inst_frame9_bit31.Q VPWR
+ VGND sg13g2_dlhq_1
X_1085_ FrameData[23] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit23.Q VPWR
+ VGND sg13g2_dlhq_1
X_0938_ FrameData[4] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit4.Q VPWR
+ VGND sg13g2_dlhq_1
X_0585_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit20.Q UIO_OE_TT_PROJECT6 _0186_ VPWR
+ VGND sg13g2_nor2b_1
X_0654_ VGND VPWR _0245_ _0246_ _0247_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit29.Q
+ sg13g2_a21oi_1
X_0723_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit11.Q VPWR _0310_ VGND _0030_ _0242_
+ sg13g2_o21ai_1
X_1206_ FrameStrobe[15] FrameStrobe_O[15] VPWR VGND sg13g2_buf_1
X_1137_ FrameData[11] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit11.Q VPWR
+ VGND sg13g2_dlhq_1
X_1068_ FrameData[6] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit6.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_43_29 VPWR VGND sg13g2_fill_1
X_0499_ UIO_IN_TT_PROJECT1 _0110_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit13.Q _0108_
+ _0105_ VPWR VGND sg13g2_a22oi_1
X_0568_ E2MID[0] EE4END[0] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit19.Q _0171_ VPWR
+ VGND sg13g2_mux2_1
X_0637_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit3.Q VPWR _0232_ VGND Inst_E_TT_IF_ConfigMem.Inst_frame5_bit2.Q
+ _0112_ sg13g2_o21ai_1
X_0706_ UIO_OUT_TT_PROJECT2 UIO_OE_TT_PROJECT5 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit16.Q
+ _0295_ VPWR VGND sg13g2_mux2_1
X_0422_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame1_bit6.Q _0038_ _0041_ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit7.Q
+ sg13g2_a21oi_1
XFILLER_44_173 VPWR VGND sg13g2_fill_1
X_0971_ FrameData[5] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit5.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_50_198 VPWR VGND sg13g2_fill_2
XFILLER_50_187 VPWR VGND sg13g2_fill_2
X_0405_ VPWR _0024_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit27.Q VGND sg13g2_inv_1
XFILLER_41_198 VPWR VGND sg13g2_fill_2
X_1170_ FrameData[11] FrameData_O[11] VPWR VGND sg13g2_buf_1
XFILLER_2_23 VPWR VGND sg13g2_fill_2
XANTENNA_39 VPWR VGND N2MID[2] sg13g2_antennanp
XFILLER_32_110 VPWR VGND sg13g2_fill_2
X_0885_ FrameData[15] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit15.Q VPWR
+ VGND sg13g2_dlhq_1
XANTENNA_28 VPWR VGND E2MID[2] sg13g2_antennanp
X_1299_ Inst_E_TT_IF_switch_matrix.W2BEGb3 W2BEGb[3] VPWR VGND sg13g2_buf_1
XANTENNA_17 VPWR VGND S2MID[0] sg13g2_antennanp
X_0954_ FrameData[20] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit20.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_36_51 VPWR VGND sg13g2_fill_1
XFILLER_23_198 VPWR VGND sg13g2_fill_2
X_0670_ N1END[2] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit28.Q Inst_E_TT_IF_ConfigMem.Inst_frame0_bit29.Q
+ _0262_ VPWR VGND sg13g2_nor3_1
X_1222_ Inst_E_TT_IF_switch_matrix.N2BEG7 N2BEG[7] VPWR VGND sg13g2_buf_1
X_1153_ FrameData[27] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit27.Q VPWR
+ VGND sg13g2_dlhq_1
X_1084_ FrameData[22] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit22.Q VPWR
+ VGND sg13g2_dlhq_1
X_0868_ FrameData[30] FrameStrobe[9] Inst_E_TT_IF_ConfigMem.Inst_frame9_bit30.Q VPWR
+ VGND sg13g2_dlhq_1
X_0799_ _0373_ VPWR _0374_ VGND _0036_ _0078_ sg13g2_o21ai_1
X_0937_ FrameData[3] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit3.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_11_124 VPWR VGND sg13g2_fill_2
X_0653_ _0246_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit28.Q _0104_ VPWR VGND sg13g2_nand2_1
X_0722_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit11.Q _0307_ _0308_ _0309_ VPWR VGND
+ sg13g2_nor3_1
X_1136_ FrameData[10] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit10.Q VPWR
+ VGND sg13g2_dlhq_1
X_1067_ FrameData[5] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit5.Q VPWR
+ VGND sg13g2_dlhq_1
X_1205_ FrameStrobe[14] FrameStrobe_O[14] VPWR VGND sg13g2_buf_1
X_0584_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame5_bit20.Q _0062_ _0185_ _0184_
+ sg13g2_a21oi_1
X_0498_ _0110_ _0109_ _0013_ _0107_ _0103_ VPWR VGND sg13g2_a22oi_1
X_0567_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit20.Q _0112_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit19.Q
+ _0170_ VPWR VGND sg13g2_nand3_1
X_0636_ _0229_ _0231_ Inst_E_TT_IF_switch_matrix.W2BEGb1 VPWR VGND sg13g2_nor2_1
X_0705_ _0293_ VPWR _0294_ VGND UO_OUT_TT_PROJECT1 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit16.Q
+ sg13g2_o21ai_1
XFILLER_0_167 VPWR VGND sg13g2_fill_1
XFILLER_0_145 VPWR VGND sg13g2_fill_1
X_1119_ FrameData[25] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit25.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_47_193 VPWR VGND sg13g2_fill_2
X_0421_ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit4.Q N2MID[6] N2END[2] N2END[3] E2MID[0]
+ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit5.Q _0040_ VPWR VGND sg13g2_mux4_1
X_0619_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit9.Q VPWR _0216_ VGND Inst_E_TT_IF_ConfigMem.Inst_frame5_bit8.Q
+ _0096_ sg13g2_o21ai_1
XFILLER_39_95 VPWR VGND sg13g2_fill_1
X_0970_ FrameData[4] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit4.Q VPWR
+ VGND sg13g2_dlhq_1
X_0404_ VPWR _0023_ UO_OUT_TT_PROJECT6 VGND sg13g2_inv_1
XFILLER_25_20 VPWR VGND sg13g2_fill_1
XANTENNA_29 VPWR VGND E2MID[2] sg13g2_antennanp
XANTENNA_18 VPWR VGND S2MID[0] sg13g2_antennanp
X_0884_ FrameData[14] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit14.Q VPWR
+ VGND sg13g2_dlhq_1
X_0953_ FrameData[19] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit19.Q VPWR
+ VGND sg13g2_dlhq_1
X_1298_ Inst_E_TT_IF_switch_matrix.W2BEGb2 W2BEGb[2] VPWR VGND sg13g2_buf_1
X_1221_ Inst_E_TT_IF_switch_matrix.N2BEG6 N2BEG[6] VPWR VGND sg13g2_buf_1
X_1152_ FrameData[26] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit26.Q VPWR
+ VGND sg13g2_dlhq_1
X_1083_ FrameData[21] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit21.Q VPWR
+ VGND sg13g2_dlhq_1
X_0867_ FrameData[29] FrameStrobe[9] Inst_E_TT_IF_ConfigMem.Inst_frame9_bit29.Q VPWR
+ VGND sg13g2_dlhq_1
X_0798_ VGND VPWR _0373_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit16.Q E6END[8] sg13g2_or2_1
XFILLER_20_125 VPWR VGND sg13g2_fill_2
X_0936_ FrameData[2] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit2.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_22_98 VPWR VGND sg13g2_fill_1
X_1135_ FrameData[9] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit9.Q VPWR
+ VGND sg13g2_dlhq_1
X_1204_ FrameStrobe[13] FrameStrobe_O[13] VPWR VGND sg13g2_buf_1
X_1066_ FrameData[4] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit4.Q VPWR
+ VGND sg13g2_dlhq_1
X_0583_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit21.Q VPWR _0184_ VGND Inst_E_TT_IF_ConfigMem.Inst_frame5_bit20.Q
+ _0104_ sg13g2_o21ai_1
X_0919_ FrameData[17] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit17.Q VPWR
+ VGND sg13g2_dlhq_1
X_0652_ _0245_ _0127_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit28.Q VPWR VGND sg13g2_nand2b_1
X_0721_ _0030_ _0112_ _0308_ VPWR VGND sg13g2_nor2_1
XFILLER_33_20 VPWR VGND sg13g2_fill_1
XFILLER_31_0 VPWR VGND sg13g2_fill_2
X_0635_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit7.Q _0230_ _0231_ VPWR VGND sg13g2_nor2_1
X_0566_ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit8.Q N1END[0] N4END[0] S1END[0] S4END[0]
+ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit9.Q _0169_ VPWR VGND sg13g2_mux4_1
X_0704_ VGND VPWR _0028_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit16.Q _0293_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit17.Q
+ sg13g2_a21oi_1
X_0497_ E2END[1] EE4END[9] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit14.Q _0109_ VPWR
+ VGND sg13g2_mux2_1
X_1049_ FrameData[19] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit19.Q VPWR
+ VGND sg13g2_dlhq_1
X_1118_ FrameData[24] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit24.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_47_150 VPWR VGND sg13g2_fill_2
X_0420_ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit5.Q Inst_E_TT_IF_ConfigMem.Inst_frame1_bit6.Q
+ _0039_ VPWR VGND sg13g2_nor2_1
XFILLER_28_53 VPWR VGND sg13g2_fill_1
X_0549_ UI_IN_TT_PROJECT3 _0154_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit27.Q _0152_
+ _0149_ VPWR VGND sg13g2_a22oi_1
X_0618_ _0213_ _0215_ Inst_E_TT_IF_switch_matrix.W2BEGb3 VPWR VGND sg13g2_nor2_1
XFILLER_53_186 VPWR VGND sg13g2_fill_1
X_0403_ VPWR _0022_ UO_OUT_TT_PROJECT7 VGND sg13g2_inv_1
X_0883_ FrameData[13] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit13.Q VPWR
+ VGND sg13g2_dlhq_1
XANTENNA_19 VPWR VGND S2MID[0] sg13g2_antennanp
XFILLER_32_112 VPWR VGND sg13g2_fill_1
X_0952_ FrameData[18] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit18.Q VPWR
+ VGND sg13g2_dlhq_1
X_1297_ Inst_E_TT_IF_switch_matrix.W2BEGb1 W2BEGb[1] VPWR VGND sg13g2_buf_1
X_1220_ Inst_E_TT_IF_switch_matrix.N2BEG5 N2BEG[5] VPWR VGND sg13g2_buf_1
X_1151_ FrameData[25] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit25.Q VPWR
+ VGND sg13g2_dlhq_1
X_0866_ FrameData[28] FrameStrobe[9] Inst_E_TT_IF_ConfigMem.Inst_frame9_bit28.Q VPWR
+ VGND sg13g2_dlhq_1
X_1082_ FrameData[20] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit20.Q VPWR
+ VGND sg13g2_dlhq_1
X_0797_ _0112_ _0169_ _0036_ _0372_ VPWR VGND sg13g2_mux2_1
XFILLER_20_148 VPWR VGND sg13g2_fill_1
X_0935_ FrameData[1] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit1.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_47_96 VPWR VGND sg13g2_fill_2
X_1134_ FrameData[8] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit8.Q VPWR
+ VGND sg13g2_dlhq_1
X_1203_ FrameStrobe[12] FrameStrobe_O[12] VPWR VGND sg13g2_buf_1
X_1065_ FrameData[3] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit3.Q VPWR
+ VGND sg13g2_dlhq_1
X_0720_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit10.Q _0169_ _0307_ VPWR VGND sg13g2_nor2_1
X_0651_ _0244_ _0243_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit1.Q Inst_E_TT_IF_switch_matrix.W2BEG7
+ VPWR VGND sg13g2_mux2_1
X_0582_ _0181_ _0183_ Inst_E_TT_IF_switch_matrix.W2BEGb7 VPWR VGND sg13g2_nor2_1
X_0849_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit11.Q E2MID[1] E6END[1] E2END[1] _0061_
+ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit10.Q Inst_E_TT_IF_switch_matrix.N2BEG6 VPWR
+ VGND sg13g2_mux4_1
X_0918_ FrameData[16] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit16.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_3_100 VPWR VGND sg13g2_fill_2
X_0703_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame6_bit17.Q _0289_ _0292_ _0029_
+ sg13g2_a21oi_1
X_0565_ UI_IN_TT_PROJECT1 _0168_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit21.Q _0166_
+ _0163_ VPWR VGND sg13g2_a22oi_1
X_0496_ VPWR VGND E6END[9] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit13.Q _0107_ _0013_
+ _0108_ _0106_ sg13g2_a221oi_1
X_1048_ FrameData[18] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit18.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_24_0 VPWR VGND sg13g2_fill_1
X_0634_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit5.Q E2END[6] UIO_OUT_TT_PROJECT1 UIO_OUT_TT_PROJECT2
+ UIO_OUT_TT_PROJECT6 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit6.Q _0230_ VPWR VGND sg13g2_mux4_1
X_1117_ FrameData[23] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit23.Q VPWR
+ VGND sg13g2_dlhq_1
X_0548_ _0154_ _0153_ _0018_ _0151_ _0148_ VPWR VGND sg13g2_a22oi_1
X_0479_ E2END[3] EE4END[11] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit20.Q _0093_ VPWR
+ VGND sg13g2_mux2_1
X_0617_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit13.Q _0214_ _0215_ VPWR VGND sg13g2_nor2_1
XFILLER_44_198 VPWR VGND sg13g2_fill_2
XFILLER_35_110 VPWR VGND sg13g2_fill_1
X_0402_ VPWR _0021_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit20.Q VGND sg13g2_inv_1
X_0882_ FrameData[12] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit12.Q VPWR
+ VGND sg13g2_dlhq_1
X_0951_ FrameData[17] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit17.Q VPWR
+ VGND sg13g2_dlhq_1
X_1296_ Inst_E_TT_IF_switch_matrix.W2BEGb0 W2BEGb[0] VPWR VGND sg13g2_buf_1
X_0865_ FrameData[27] FrameStrobe[9] Inst_E_TT_IF_ConfigMem.Inst_frame9_bit27.Q VPWR
+ VGND sg13g2_dlhq_1
X_0796_ _0369_ _0371_ Inst_E_TT_IF_switch_matrix.N4BEG1 VPWR VGND sg13g2_nor2_1
X_1081_ FrameData[19] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit19.Q VPWR
+ VGND sg13g2_dlhq_1
X_0934_ FrameData[0] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit0.Q VPWR
+ VGND sg13g2_dlhq_1
X_1150_ FrameData[24] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit24.Q VPWR
+ VGND sg13g2_dlhq_1
X_1279_ Inst_E_TT_IF_switch_matrix.S4BEG0 S4BEG[12] VPWR VGND sg13g2_buf_1
X_1202_ FrameStrobe[11] FrameStrobe_O[11] VPWR VGND sg13g2_buf_1
X_1064_ FrameData[2] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit2.Q VPWR
+ VGND sg13g2_dlhq_1
X_1133_ FrameData[7] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit7.Q VPWR
+ VGND sg13g2_dlhq_1
X_0650_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit31.Q UO_OUT_TT_PROJECT4 UO_OUT_TT_PROJECT7
+ UIO_OUT_TT_PROJECT7 UIO_OE_TT_PROJECT0 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit0.Q
+ _0244_ VPWR VGND sg13g2_mux4_1
X_0581_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit25.Q _0182_ _0183_ VPWR VGND sg13g2_nor2_1
X_0779_ _0096_ _0155_ _0034_ _0356_ VPWR VGND sg13g2_mux2_1
X_0848_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit12.Q E2MID[0] E2END[0] E6END[0] _0052_
+ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit13.Q Inst_E_TT_IF_switch_matrix.N2BEG7 VPWR
+ VGND sg13g2_mux4_1
X_0917_ FrameData[15] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit15.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_17_67 VPWR VGND sg13g2_fill_1
X_0564_ _0168_ _0167_ _0020_ _0165_ _0162_ VPWR VGND sg13g2_a22oi_1
X_0495_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit14.Q _0013_ _0107_ VPWR VGND sg13g2_nor2_1
X_0633_ _0225_ _0228_ _0229_ VPWR VGND sg13g2_nor2_1
X_1116_ FrameData[22] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit22.Q VPWR
+ VGND sg13g2_dlhq_1
X_1047_ FrameData[17] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit17.Q VPWR
+ VGND sg13g2_dlhq_1
X_0702_ _0291_ _0290_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit17.Q VPWR VGND sg13g2_nand2b_1
X_0616_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit11.Q E2END[4] UIO_OUT_TT_PROJECT0 UIO_OUT_TT_PROJECT3
+ UIO_OUT_TT_PROJECT4 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit12.Q _0214_ VPWR VGND
+ sg13g2_mux4_1
XFILLER_53_199 VPWR VGND sg13g2_fill_1
X_0547_ E2END[3] EE4END[11] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit28.Q _0153_ VPWR
+ VGND sg13g2_mux2_1
X_0478_ VPWR VGND E6END[11] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit19.Q _0091_ _0011_
+ _0092_ _0090_ sg13g2_a221oi_1
XFILLER_44_155 VPWR VGND sg13g2_fill_1
X_0401_ VPWR _0020_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit23.Q VGND sg13g2_inv_1
XFILLER_26_144 VPWR VGND sg13g2_decap_4
XFILLER_6_91 VPWR VGND sg13g2_fill_2
X_0881_ FrameData[11] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit11.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_23_136 VPWR VGND sg13g2_decap_4
X_1295_ Inst_E_TT_IF_switch_matrix.W2BEG7 W2BEG[7] VPWR VGND sg13g2_buf_1
X_0950_ FrameData[16] FrameStrobe[6] Inst_E_TT_IF_ConfigMem.Inst_frame6_bit16.Q VPWR
+ VGND sg13g2_dlhq_1
X_0864_ FrameData[26] FrameStrobe[9] Inst_E_TT_IF_ConfigMem.Inst_frame9_bit26.Q VPWR
+ VGND sg13g2_dlhq_1
X_1080_ FrameData[18] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit18.Q VPWR
+ VGND sg13g2_dlhq_1
X_0795_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit18.Q _0370_ _0371_ VPWR VGND sg13g2_nor2_1
X_0933_ FrameData[31] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit31.Q VPWR
+ VGND sg13g2_dlhq_1
X_1278_ S4END[15] S4BEG[11] VPWR VGND sg13g2_buf_1
X_1201_ FrameStrobe[10] FrameStrobe_O[10] VPWR VGND sg13g2_buf_1
X_0580_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit23.Q E2END[0] UIO_OUT_TT_PROJECT0 UIO_OUT_TT_PROJECT4
+ UIO_OUT_TT_PROJECT7 Inst_E_TT_IF_ConfigMem.Inst_frame5_bit24.Q _0182_ VPWR VGND
+ sg13g2_mux4_1
X_0778_ _0353_ _0355_ Inst_E_TT_IF_switch_matrix.N4BEG3 VPWR VGND sg13g2_nor2_1
X_1063_ FrameData[1] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit1.Q VPWR
+ VGND sg13g2_dlhq_1
X_0847_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit26.Q E1END[0] E6END[8] _0078_ _0242_
+ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit27.Q Inst_E_TT_IF_switch_matrix.S1BEG0 VPWR
+ VGND sg13g2_mux4_1
X_1132_ FrameData[6] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit6.Q VPWR
+ VGND sg13g2_dlhq_1
X_0916_ FrameData[14] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit14.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_33_67 VPWR VGND sg13g2_fill_1
XFILLER_17_35 VPWR VGND sg13g2_fill_1
X_1115_ FrameData[21] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit21.Q VPWR
+ VGND sg13g2_dlhq_1
X_0563_ E2END[1] EE4END[9] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit22.Q _0167_ VPWR
+ VGND sg13g2_mux2_1
X_0494_ E2MID[1] EE4END[1] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit14.Q _0106_ VPWR
+ VGND sg13g2_mux2_1
X_0632_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit7.Q VPWR _0228_ VGND Inst_E_TT_IF_ConfigMem.Inst_frame5_bit6.Q
+ _0227_ sg13g2_o21ai_1
X_1046_ FrameData[16] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit16.Q VPWR
+ VGND sg13g2_dlhq_1
X_0701_ _0155_ _0096_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit16.Q _0290_ VPWR VGND
+ sg13g2_mux2_1
X_1029_ FrameData[31] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit31.Q VPWR
+ VGND sg13g2_dlhq_1
X_0546_ VPWR VGND E6END[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit27.Q _0151_ _0018_
+ _0152_ _0150_ sg13g2_a221oi_1
X_0477_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit20.Q _0011_ _0091_ VPWR VGND sg13g2_nor2_1
XFILLER_30_57 VPWR VGND sg13g2_fill_2
X_0615_ _0209_ _0212_ _0213_ VPWR VGND sg13g2_nor2_1
X_0400_ VPWR _0019_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit26.Q VGND sg13g2_inv_1
XFILLER_44_134 VPWR VGND sg13g2_fill_1
X_0529_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit2.Q _0016_ _0137_ VPWR VGND sg13g2_nor2_1
X_0880_ FrameData[10] FrameStrobe[8] Inst_E_TT_IF_ConfigMem.Inst_frame8_bit10.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_40_181 VPWR VGND sg13g2_fill_1
X_1294_ Inst_E_TT_IF_switch_matrix.W2BEG6 W2BEG[6] VPWR VGND sg13g2_buf_1
XFILLER_52_88 VPWR VGND sg13g2_fill_2
XFILLER_20_118 VPWR VGND sg13g2_decap_8
X_0932_ FrameData[30] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit30.Q VPWR
+ VGND sg13g2_dlhq_1
X_1277_ S4END[14] S4BEG[10] VPWR VGND sg13g2_buf_1
X_0863_ FrameData[25] FrameStrobe[9] Inst_E_TT_IF_ConfigMem.Inst_frame9_bit25.Q VPWR
+ VGND sg13g2_dlhq_1
X_0794_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit17.Q E1END[1] EE4END[1] _0134_ _0103_
+ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit19.Q _0370_ VPWR VGND sg13g2_mux4_1
X_1131_ FrameData[5] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit5.Q VPWR
+ VGND sg13g2_dlhq_1
X_1200_ FrameStrobe[9] FrameStrobe_O[9] VPWR VGND sg13g2_buf_1
X_0777_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit24.Q _0354_ _0355_ VPWR VGND sg13g2_nor2_1
X_0846_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit28.Q E1END[1] E6END[9] _0069_ _0250_
+ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit29.Q Inst_E_TT_IF_switch_matrix.S1BEG1 VPWR
+ VGND sg13g2_mux4_1
X_1062_ FrameData[0] FrameStrobe[2] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit0.Q VPWR
+ VGND sg13g2_dlhq_1
X_0915_ FrameData[13] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit13.Q VPWR
+ VGND sg13g2_dlhq_1
X_1329_ Inst_E_TT_IF_switch_matrix.WW4BEG13 WW4BEG[13] VPWR VGND sg13g2_buf_1
X_1114_ FrameData[20] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit20.Q VPWR
+ VGND sg13g2_dlhq_1
X_0562_ VPWR VGND E6END[1] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit21.Q _0165_ _0020_
+ _0166_ _0164_ sg13g2_a221oi_1
X_0493_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit15.Q _0104_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit14.Q
+ _0105_ VPWR VGND sg13g2_nand3_1
X_0631_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame5_bit5.Q _0103_ _0227_ _0226_ sg13g2_a21oi_1
X_0700_ _0070_ _0263_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit16.Q _0289_ VPWR VGND
+ sg13g2_mux2_1
X_1045_ FrameData[15] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit15.Q VPWR
+ VGND sg13g2_dlhq_1
X_0829_ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit7.Q UO_OUT_TT_PROJECT6 _0103_ UIO_OE_TT_PROJECT2
+ _0104_ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit6.Q Inst_E_TT_IF_switch_matrix.WW4BEG6
+ VPWR VGND sg13g2_mux4_1
X_1028_ FrameData[30] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit30.Q VPWR
+ VGND sg13g2_dlhq_1
X_0545_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit28.Q _0018_ _0151_ VPWR VGND sg13g2_nor2_1
X_0476_ E2MID[3] EE4END[3] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit20.Q _0090_ VPWR
+ VGND sg13g2_mux2_1
X_0614_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit13.Q VPWR _0212_ VGND Inst_E_TT_IF_ConfigMem.Inst_frame5_bit12.Q
+ _0211_ sg13g2_o21ai_1
XFILLER_29_110 VPWR VGND sg13g2_fill_1
X_0528_ E2MID[5] EE4END[5] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit2.Q _0136_ VPWR VGND
+ sg13g2_mux2_1
X_0459_ VPWR VGND EE4END[13] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit25.Q _0074_ _0008_
+ _0075_ _0073_ sg13g2_a221oi_1
XFILLER_40_160 VPWR VGND sg13g2_fill_1
X_1293_ Inst_E_TT_IF_switch_matrix.W2BEG5 W2BEG[5] VPWR VGND sg13g2_buf_1
XFILLER_52_45 VPWR VGND sg13g2_fill_1
XFILLER_14_138 VPWR VGND sg13g2_fill_1
X_1276_ S4END[13] S4BEG[9] VPWR VGND sg13g2_buf_1
X_0793_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame8_bit17.Q _0365_ _0369_ _0368_
+ sg13g2_a21oi_1
X_0862_ FrameData[24] FrameStrobe[9] Inst_E_TT_IF_ConfigMem.Inst_frame9_bit24.Q VPWR
+ VGND sg13g2_dlhq_1
X_0931_ FrameData[29] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit29.Q VPWR
+ VGND sg13g2_dlhq_1
X_1130_ FrameData[4] FrameStrobe[0] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit4.Q VPWR
+ VGND sg13g2_dlhq_1
X_1061_ FrameData[31] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit31.Q VPWR
+ VGND sg13g2_dlhq_1
X_0845_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit30.Q E1END[2] E6END[10] _0060_ _0263_
+ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit31.Q Inst_E_TT_IF_switch_matrix.S1BEG2 VPWR
+ VGND sg13g2_mux4_1
X_0914_ FrameData[12] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit12.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_52_0 VPWR VGND sg13g2_fill_2
X_0776_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit23.Q E1END[3] EE4END[3] _0120_ _0087_
+ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit25.Q _0354_ VPWR VGND sg13g2_mux4_1
X_1328_ Inst_E_TT_IF_switch_matrix.WW4BEG12 WW4BEG[12] VPWR VGND sg13g2_buf_1
X_1259_ S2MID[0] S2BEGb[0] VPWR VGND sg13g2_buf_1
X_0492_ Inst_E_TT_IF_ConfigMem.Inst_frame0_bit10.Q N2MID[1] N2END[1] S2MID[1] S2END[1]
+ Inst_E_TT_IF_ConfigMem.Inst_frame0_bit11.Q _0104_ VPWR VGND sg13g2_mux4_1
X_0561_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit22.Q _0020_ _0165_ VPWR VGND sg13g2_nor2_1
X_0630_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit5.Q UIO_OE_TT_PROJECT1 _0226_ VPWR VGND
+ sg13g2_nor2b_1
X_0759_ _0336_ _0339_ _0340_ VPWR VGND sg13g2_nor2_1
X_1113_ FrameData[19] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit19.Q VPWR
+ VGND sg13g2_dlhq_1
X_1044_ FrameData[14] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit14.Q VPWR
+ VGND sg13g2_dlhq_1
X_0828_ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit9.Q UO_OUT_TT_PROJECT7 _0111_ UIO_OE_TT_PROJECT3
+ _0112_ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit8.Q Inst_E_TT_IF_switch_matrix.WW4BEG7
+ VPWR VGND sg13g2_mux4_1
X_0544_ E2MID[3] EE4END[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit28.Q _0150_ VPWR
+ VGND sg13g2_mux2_1
X_0475_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit21.Q _0088_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit20.Q
+ _0089_ VPWR VGND sg13g2_nand3_1
X_1027_ FrameData[29] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit29.Q VPWR
+ VGND sg13g2_dlhq_1
X_0613_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame5_bit11.Q _0087_ _0211_ _0210_
+ sg13g2_a21oi_1
XFILLER_44_125 VPWR VGND sg13g2_fill_2
XFILLER_29_177 VPWR VGND sg13g2_fill_2
XFILLER_41_36 VPWR VGND sg13g2_fill_1
X_0527_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit3.Q _0070_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit2.Q
+ _0135_ VPWR VGND sg13g2_nand3_1
X_0458_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit26.Q _0008_ _0074_ VPWR VGND sg13g2_nor2_1
X_0389_ VPWR _0008_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit27.Q VGND sg13g2_inv_1
X_1292_ Inst_E_TT_IF_switch_matrix.W2BEG4 W2BEG[4] VPWR VGND sg13g2_buf_1
XFILLER_36_58 VPWR VGND sg13g2_fill_1
XFILLER_22_172 VPWR VGND sg13g2_fill_2
X_1275_ S4END[12] S4BEG[8] VPWR VGND sg13g2_buf_1
X_0792_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit18.Q VPWR _0368_ VGND Inst_E_TT_IF_ConfigMem.Inst_frame8_bit17.Q
+ _0367_ sg13g2_o21ai_1
X_0930_ FrameData[28] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit28.Q VPWR
+ VGND sg13g2_dlhq_1
X_0861_ FrameData[23] FrameStrobe[9] Inst_E_TT_IF_ConfigMem.Inst_frame9_bit23.Q VPWR
+ VGND sg13g2_dlhq_1
X_1060_ FrameData[30] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit30.Q VPWR
+ VGND sg13g2_dlhq_1
X_1189_ FrameData[30] FrameData_O[30] VPWR VGND sg13g2_buf_1
X_0775_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame8_bit23.Q _0349_ _0353_ _0352_
+ sg13g2_a21oi_1
X_0844_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit0.Q E1END[3] E6END[11] _0051_ _0274_
+ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit1.Q Inst_E_TT_IF_switch_matrix.S1BEG3 VPWR
+ VGND sg13g2_mux4_1
X_0913_ FrameData[11] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit11.Q VPWR
+ VGND sg13g2_dlhq_1
X_1258_ Inst_E_TT_IF_switch_matrix.S2BEG7 S2BEG[7] VPWR VGND sg13g2_buf_1
X_1327_ Inst_E_TT_IF_switch_matrix.WW4BEG11 WW4BEG[11] VPWR VGND sg13g2_buf_1
X_0758_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit25.Q VPWR _0339_ VGND Inst_E_TT_IF_ConfigMem.Inst_frame7_bit24.Q
+ _0338_ sg13g2_o21ai_1
X_0560_ E2MID[1] EE4END[1] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit22.Q _0164_ VPWR
+ VGND sg13g2_mux2_1
X_1112_ FrameData[18] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit18.Q VPWR
+ VGND sg13g2_dlhq_1
X_0491_ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit26.Q N1END[1] N4END[1] S1END[1] S4END[1]
+ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit27.Q _0103_ VPWR VGND sg13g2_mux4_1
X_1043_ FrameData[13] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit13.Q VPWR
+ VGND sg13g2_dlhq_1
X_0827_ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit11.Q UO_OUT_TT_PROJECT4 _0120_ UIO_OUT_TT_PROJECT0
+ _0052_ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit10.Q Inst_E_TT_IF_switch_matrix.WW4BEG8
+ VPWR VGND sg13g2_mux4_1
XFILLER_0_119 VPWR VGND sg13g2_fill_2
X_0689_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame6_bit23.Q _0279_ _0280_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit24.Q
+ sg13g2_a21oi_1
XFILLER_47_167 VPWR VGND sg13g2_fill_1
X_0474_ Inst_E_TT_IF_ConfigMem.Inst_frame0_bit15.Q N2MID[3] S2MID[3] N2END[3] S2END[3]
+ Inst_E_TT_IF_ConfigMem.Inst_frame0_bit14.Q _0088_ VPWR VGND sg13g2_mux4_1
X_0543_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit29.Q _0088_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit28.Q
+ _0149_ VPWR VGND sg13g2_nand3_1
X_0612_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit11.Q UIO_OE_TT_PROJECT3 _0210_ VPWR
+ VGND sg13g2_nor2b_1
X_1026_ FrameData[28] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit28.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_35_137 VPWR VGND sg13g2_fill_2
X_0388_ VPWR _0007_ S1END[1] VGND sg13g2_inv_1
X_0457_ E1END[1] E2END[5] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit26.Q _0073_ VPWR VGND
+ sg13g2_mux2_1
X_0526_ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit18.Q N1END[1] N4END[1] S1END[1] S4END[1]
+ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit19.Q _0134_ VPWR VGND sg13g2_mux4_1
XFILLER_26_126 VPWR VGND sg13g2_fill_1
X_1009_ FrameData[11] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit11.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_49_7 VPWR VGND sg13g2_fill_2
XFILLER_31_140 VPWR VGND sg13g2_fill_2
X_1291_ Inst_E_TT_IF_switch_matrix.W2BEG3 W2BEG[3] VPWR VGND sg13g2_buf_1
X_0509_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit8.Q E6END[7] _0119_ VPWR VGND sg13g2_nor2_1
X_0791_ _0366_ VPWR _0367_ VGND _0035_ _0069_ sg13g2_o21ai_1
X_0860_ FrameData[22] FrameStrobe[9] Inst_E_TT_IF_ConfigMem.Inst_frame9_bit22.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_26_70 VPWR VGND sg13g2_decap_8
XFILLER_3_52 VPWR VGND sg13g2_fill_1
XFILLER_9_100 VPWR VGND sg13g2_fill_1
XFILLER_9_199 VPWR VGND sg13g2_fill_1
X_1274_ S4END[11] S4BEG[7] VPWR VGND sg13g2_buf_1
X_0989_ FrameData[23] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit23.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_12_61 VPWR VGND sg13g2_fill_1
X_0774_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit24.Q VPWR _0352_ VGND Inst_E_TT_IF_ConfigMem.Inst_frame8_bit23.Q
+ _0351_ sg13g2_o21ai_1
X_1188_ FrameData[29] FrameData_O[29] VPWR VGND sg13g2_buf_1
X_0843_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit2.Q E2MID[7] E2END[7] E6END[8] _0112_
+ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit3.Q Inst_E_TT_IF_switch_matrix.S2BEG0 VPWR
+ VGND sg13g2_mux4_1
X_0912_ FrameData[10] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit10.Q VPWR
+ VGND sg13g2_dlhq_1
X_1326_ Inst_E_TT_IF_switch_matrix.WW4BEG10 WW4BEG[10] VPWR VGND sg13g2_buf_1
X_1257_ Inst_E_TT_IF_switch_matrix.S2BEG6 S2BEG[6] VPWR VGND sg13g2_buf_1
X_0490_ UIO_IN_TT_PROJECT2 _0102_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit16.Q _0100_
+ _0097_ VPWR VGND sg13g2_a22oi_1
X_1042_ FrameData[12] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit12.Q VPWR
+ VGND sg13g2_dlhq_1
X_1111_ FrameData[17] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit17.Q VPWR
+ VGND sg13g2_dlhq_1
X_0757_ _0337_ VPWR _0338_ VGND _0032_ _0060_ sg13g2_o21ai_1
XFILLER_44_48 VPWR VGND sg13g2_fill_2
X_0826_ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit13.Q UO_OUT_TT_PROJECT5 _0127_ UIO_OUT_TT_PROJECT1
+ _0061_ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit12.Q Inst_E_TT_IF_switch_matrix.WW4BEG9
+ VPWR VGND sg13g2_mux4_1
X_1309_ Inst_E_TT_IF_switch_matrix.W6BEG5 W6BEG[5] VPWR VGND sg13g2_buf_1
X_0688_ UIO_OUT_TT_PROJECT4 UIO_OE_TT_PROJECT3 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit22.Q
+ _0279_ VPWR VGND sg13g2_mux2_1
XFILLER_18_93 VPWR VGND sg13g2_fill_2
X_0542_ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit14.Q N1END[3] N4END[3] S1END[3] S4END[3]
+ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit15.Q _0148_ VPWR VGND sg13g2_mux4_1
X_0611_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame5_bit11.Q _0080_ _0209_ _0208_
+ sg13g2_a21oi_1
X_0473_ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit30.Q N1END[3] N4END[3] S1END[3] S4END[3]
+ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit31.Q _0087_ VPWR VGND sg13g2_mux4_1
X_0809_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit15.Q UIO_OUT_TT_PROJECT2 _0134_ _0162_
+ _0061_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit14.Q Inst_E_TT_IF_switch_matrix.W6BEG10
+ VPWR VGND sg13g2_mux4_1
X_1025_ FrameData[27] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit27.Q VPWR
+ VGND sg13g2_dlhq_1
X_0525_ UI_IN_TT_PROJECT6 _0133_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit4.Q _0131_
+ _0128_ VPWR VGND sg13g2_a22oi_1
XANTENNA_1 VPWR VGND FrameStrobe[10] sg13g2_antennanp
X_0387_ VPWR _0006_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit30.Q VGND sg13g2_inv_1
X_0456_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit27.Q _0070_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit26.Q
+ _0072_ VPWR VGND sg13g2_nand3_1
X_1008_ FrameData[10] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit10.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_31_93 VPWR VGND sg13g2_fill_1
X_1290_ Inst_E_TT_IF_switch_matrix.W2BEG2 W2BEG[2] VPWR VGND sg13g2_buf_1
X_0439_ VPWR VGND EE4END[15] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit31.Q _0056_ _0003_
+ _0057_ _0055_ sg13g2_a221oi_1
X_0508_ UIO_IN_TT_PROJECT0 _0118_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit10.Q _0116_
+ _0113_ VPWR VGND sg13g2_a22oi_1
X_0790_ VGND VPWR _0366_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit19.Q E6END[9] sg13g2_or2_1
X_1273_ S4END[10] S4BEG[6] VPWR VGND sg13g2_buf_1
X_0988_ FrameData[22] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit22.Q VPWR
+ VGND sg13g2_dlhq_1
X_0773_ _0350_ VPWR _0351_ VGND _0033_ _0051_ sg13g2_o21ai_1
X_0842_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit4.Q E2MID[6] E2END[6] E6END[9] _0104_
+ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit5.Q Inst_E_TT_IF_switch_matrix.S2BEG1 VPWR
+ VGND sg13g2_mux4_1
X_0911_ FrameData[9] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit9.Q VPWR
+ VGND sg13g2_dlhq_1
X_1325_ Inst_E_TT_IF_switch_matrix.WW4BEG9 WW4BEG[9] VPWR VGND sg13g2_buf_1
X_1256_ Inst_E_TT_IF_switch_matrix.S2BEG5 S2BEG[5] VPWR VGND sg13g2_buf_1
X_1187_ FrameData[28] FrameData_O[28] VPWR VGND sg13g2_buf_1
XFILLER_23_50 VPWR VGND sg13g2_fill_1
X_1041_ FrameData[11] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit11.Q VPWR
+ VGND sg13g2_dlhq_1
X_1110_ FrameData[16] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit16.Q VPWR
+ VGND sg13g2_dlhq_1
X_1239_ N4END[12] N4BEG[8] VPWR VGND sg13g2_buf_1
X_0756_ VGND VPWR _0337_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit26.Q E6END[6] sg13g2_or2_1
Xclkbuf_0_UserCLK UserCLK clknet_0_UserCLK VPWR VGND sg13g2_buf_8
XFILLER_28_17 VPWR VGND sg13g2_fill_1
X_1308_ Inst_E_TT_IF_switch_matrix.W6BEG4 W6BEG[4] VPWR VGND sg13g2_buf_1
X_0687_ _0277_ VPWR _0278_ VGND UO_OUT_TT_PROJECT4 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit22.Q
+ sg13g2_o21ai_1
X_0825_ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit15.Q UO_OUT_TT_PROJECT6 _0134_ UIO_OUT_TT_PROJECT2
+ _0070_ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit14.Q Inst_E_TT_IF_switch_matrix.WW4BEG10
+ VPWR VGND sg13g2_mux4_1
XFILLER_50_70 VPWR VGND sg13g2_fill_1
X_0541_ UI_IN_TT_PROJECT4 _0147_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit30.Q _0145_
+ _0142_ VPWR VGND sg13g2_a22oi_1
X_0472_ UIO_IN_TT_PROJECT4 _0086_ Inst_E_TT_IF_ConfigMem.Inst_frame2_bit22.Q _0084_
+ _0081_ VPWR VGND sg13g2_a22oi_1
X_0808_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit17.Q UIO_OUT_TT_PROJECT3 _0141_ _0169_
+ _0052_ Inst_E_TT_IF_ConfigMem.Inst_frame3_bit16.Q Inst_E_TT_IF_switch_matrix.W6BEG11
+ VPWR VGND sg13g2_mux4_1
X_1024_ FrameData[26] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit26.Q VPWR
+ VGND sg13g2_dlhq_1
X_0610_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit12.Q VPWR _0208_ VGND Inst_E_TT_IF_ConfigMem.Inst_frame5_bit11.Q
+ _0088_ sg13g2_o21ai_1
X_0739_ _0322_ _0321_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit3.Q Inst_E_TT_IF_switch_matrix.W1BEG1
+ VPWR VGND sg13g2_mux2_1
X_0524_ _0133_ _0132_ _0015_ _0130_ _0127_ VPWR VGND sg13g2_a22oi_1
XANTENNA_2 VPWR VGND FrameStrobe[11] sg13g2_antennanp
X_0455_ VPWR _0071_ _0070_ VGND sg13g2_inv_1
X_0386_ VPWR _0005_ S1END[2] VGND sg13g2_inv_1
X_1007_ FrameData[9] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit9.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_13_0 VPWR VGND sg13g2_fill_1
XFILLER_15_51 VPWR VGND sg13g2_fill_1
X_0438_ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit0.Q _0003_ _0056_ VPWR VGND sg13g2_nor2_1
X_0507_ _0118_ _0117_ _0014_ _0115_ _0111_ VPWR VGND sg13g2_a22oi_1
XFILLER_22_120 VPWR VGND sg13g2_fill_2
XFILLER_16_183 VPWR VGND sg13g2_fill_2
X_1272_ S4END[9] S4BEG[5] VPWR VGND sg13g2_buf_1
X_0987_ FrameData[21] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit21.Q VPWR
+ VGND sg13g2_dlhq_1
X_0772_ VGND VPWR _0350_ Inst_E_TT_IF_ConfigMem.Inst_frame8_bit25.Q E6END[11] sg13g2_or2_1
X_0910_ FrameData[8] FrameStrobe[7] Inst_E_TT_IF_ConfigMem.Inst_frame7_bit8.Q VPWR
+ VGND sg13g2_dlhq_1
X_0841_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit7.Q E2MID[5] E6END[10] E2END[5] _0096_
+ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit6.Q Inst_E_TT_IF_switch_matrix.S2BEG2 VPWR
+ VGND sg13g2_mux4_1
X_1186_ FrameData[27] FrameData_O[27] VPWR VGND sg13g2_buf_1
X_1255_ Inst_E_TT_IF_switch_matrix.S2BEG4 S2BEG[4] VPWR VGND sg13g2_buf_1
X_1324_ Inst_E_TT_IF_switch_matrix.WW4BEG8 WW4BEG[8] VPWR VGND sg13g2_buf_1
X_1040_ FrameData[10] FrameStrobe[3] Inst_E_TT_IF_ConfigMem.Inst_frame3_bit10.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_2_141 VPWR VGND sg13g2_fill_1
X_1238_ N4END[11] N4BEG[7] VPWR VGND sg13g2_buf_1
X_0755_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame7_bit26.Q _0062_ _0336_ _0335_
+ sg13g2_a21oi_1
X_1169_ FrameData[10] FrameData_O[10] VPWR VGND sg13g2_buf_1
X_0824_ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit17.Q UO_OUT_TT_PROJECT7 _0141_ UIO_OUT_TT_PROJECT3
+ _0079_ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit16.Q Inst_E_TT_IF_switch_matrix.WW4BEG11
+ VPWR VGND sg13g2_mux4_1
X_1307_ Inst_E_TT_IF_switch_matrix.W6BEG3 W6BEG[3] VPWR VGND sg13g2_buf_1
X_0686_ VGND VPWR _0022_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit22.Q _0277_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit23.Q
+ sg13g2_a21oi_1
XFILLER_34_50 VPWR VGND sg13g2_fill_1
X_0540_ _0147_ _0146_ _0017_ _0144_ _0141_ VPWR VGND sg13g2_a22oi_1
X_0471_ _0086_ _0085_ _0010_ _0083_ _0078_ VPWR VGND sg13g2_a22oi_1
X_1023_ FrameData[25] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit25.Q VPWR
+ VGND sg13g2_dlhq_1
X_0669_ _0261_ E6END[2] Inst_E_TT_IF_ConfigMem.Inst_frame0_bit29.Q VPWR VGND sg13g2_nand2b_1
XFILLER_29_159 VPWR VGND sg13g2_fill_1
X_0807_ _0379_ VPWR ENA_TT_PROJECT VGND Inst_E_TT_IF_ConfigMem.Inst_frame1_bit3.Q
+ _0380_ sg13g2_o21ai_1
X_0738_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit1.Q N1END[1] S1END[1] UO_OUT_TT_PROJECT3
+ UO_OUT_TT_PROJECT6 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit2.Q _0322_ VPWR VGND sg13g2_mux4_1
XANTENNA_3 VPWR VGND FrameStrobe[13] sg13g2_antennanp
X_0454_ Inst_E_TT_IF_ConfigMem.Inst_frame0_bit18.Q N2MID[5] N2END[5] S2MID[5] S2END[5]
+ Inst_E_TT_IF_ConfigMem.Inst_frame0_bit19.Q _0070_ VPWR VGND sg13g2_mux4_1
X_0385_ VPWR _0004_ E1END[2] VGND sg13g2_inv_1
X_0523_ E2END[6] EE4END[14] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit5.Q _0132_ VPWR
+ VGND sg13g2_mux2_1
X_1006_ FrameData[8] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit8.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_31_51 VPWR VGND sg13g2_fill_2
X_0437_ E1END[3] E2END[7] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit0.Q _0055_ VPWR VGND
+ sg13g2_mux2_1
XFILLER_31_198 VPWR VGND sg13g2_fill_2
X_0506_ E2END[0] EE4END[8] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit11.Q _0117_ VPWR
+ VGND sg13g2_mux2_1
XFILLER_26_84 VPWR VGND sg13g2_fill_1
X_1271_ S4END[8] S4BEG[4] VPWR VGND sg13g2_buf_1
XFILLER_47_39 VPWR VGND sg13g2_fill_1
X_0986_ FrameData[20] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit20.Q VPWR
+ VGND sg13g2_dlhq_1
X_0771_ _0088_ _0148_ _0033_ _0349_ VPWR VGND sg13g2_mux2_1
X_0840_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit9.Q E2MID[4] E6END[11] E2END[4] _0088_
+ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit8.Q Inst_E_TT_IF_switch_matrix.S2BEG3 VPWR
+ VGND sg13g2_mux4_1
X_1185_ FrameData[26] FrameData_O[26] VPWR VGND sg13g2_buf_1
X_1254_ Inst_E_TT_IF_switch_matrix.S2BEG3 S2BEG[3] VPWR VGND sg13g2_buf_1
X_0969_ FrameData[3] FrameStrobe[5] Inst_E_TT_IF_ConfigMem.Inst_frame5_bit3.Q VPWR
+ VGND sg13g2_dlhq_1
X_1323_ Inst_E_TT_IF_switch_matrix.WW4BEG7 WW4BEG[7] VPWR VGND sg13g2_buf_1
XFILLER_3_0 VPWR VGND sg13g2_fill_1
X_0754_ Inst_E_TT_IF_ConfigMem.Inst_frame7_bit24.Q VPWR _0335_ VGND Inst_E_TT_IF_ConfigMem.Inst_frame7_bit26.Q
+ _0155_ sg13g2_o21ai_1
XFILLER_36_0 VPWR VGND sg13g2_fill_1
X_1306_ Inst_E_TT_IF_switch_matrix.W6BEG2 W6BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_9_21 VPWR VGND sg13g2_fill_2
X_0685_ VGND VPWR Inst_E_TT_IF_ConfigMem.Inst_frame6_bit23.Q _0275_ _0276_ _0025_
+ sg13g2_a21oi_1
X_0823_ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit19.Q UO_OUT_TT_PROJECT0 _0148_ UIO_OUT_TT_PROJECT4
+ _0088_ Inst_E_TT_IF_ConfigMem.Inst_frame4_bit18.Q Inst_E_TT_IF_switch_matrix.WW4BEG12
+ VPWR VGND sg13g2_mux4_1
X_1237_ N4END[10] N4BEG[6] VPWR VGND sg13g2_buf_1
X_1099_ FrameData[5] FrameStrobe[1] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit5.Q VPWR
+ VGND sg13g2_dlhq_1
X_1168_ FrameData[9] FrameData_O[9] VPWR VGND sg13g2_buf_1
XFILLER_38_105 VPWR VGND sg13g2_fill_2
X_0470_ E2MID[4] EE4END[4] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit23.Q _0085_ VPWR
+ VGND sg13g2_mux2_1
X_1022_ FrameData[24] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit24.Q VPWR
+ VGND sg13g2_dlhq_1
X_0806_ _0380_ N2MID[6] Inst_E_TT_IF_ConfigMem.Inst_frame1_bit2.Q VPWR VGND sg13g2_nand2b_1
X_0737_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit1.Q UIO_OE_TT_PROJECT0 UIO_OE_TT_PROJECT1
+ UIO_OE_TT_PROJECT5 UIO_OE_TT_PROJECT6 Inst_E_TT_IF_ConfigMem.Inst_frame6_bit2.Q
+ _0321_ VPWR VGND sg13g2_mux4_1
X_0668_ _0260_ _0259_ Inst_E_TT_IF_ConfigMem.Inst_frame6_bit26.Q VPWR VGND sg13g2_nand2b_1
X_0599_ Inst_E_TT_IF_ConfigMem.Inst_frame5_bit19.Q _0198_ _0199_ VPWR VGND sg13g2_nor2_1
X_0522_ VPWR VGND E6END[6] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit4.Q _0130_ _0015_
+ _0131_ _0129_ sg13g2_a221oi_1
XANTENNA_4 VPWR VGND FrameStrobe[17] sg13g2_antennanp
X_0453_ Inst_E_TT_IF_ConfigMem.Inst_frame0_bit2.Q N1END[1] N4END[1] S1END[1] S4END[1]
+ Inst_E_TT_IF_ConfigMem.Inst_frame0_bit3.Q _0069_ VPWR VGND sg13g2_mux4_1
X_0384_ VPWR _0003_ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit1.Q VGND sg13g2_inv_1
XFILLER_26_119 VPWR VGND sg13g2_decap_8
X_1005_ FrameData[7] FrameStrobe[4] Inst_E_TT_IF_ConfigMem.Inst_frame4_bit7.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_31_74 VPWR VGND sg13g2_fill_1
X_0436_ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit1.Q _0052_ Inst_E_TT_IF_ConfigMem.Inst_frame1_bit0.Q
+ _0054_ VPWR VGND sg13g2_nand3_1
XFILLER_31_122 VPWR VGND sg13g2_fill_1
X_0505_ VPWR VGND E6END[8] Inst_E_TT_IF_ConfigMem.Inst_frame2_bit10.Q _0115_ _0014_
+ _0116_ _0114_ sg13g2_a221oi_1
XFILLER_16_163 VPWR VGND sg13g2_fill_2
XFILLER_16_185 VPWR VGND sg13g2_fill_1
.ends

