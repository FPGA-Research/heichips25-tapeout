VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO E_TT_IF
  CLASS BLOCK ;
  FOREIGN E_TT_IF ;
  ORIGIN 0.000 0.000 ;
  SIZE 107.520 BY 215.040 ;
  PIN CLK_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 116.980 107.520 117.380 ;
    END
  END CLK_TT_PROJECT
  PIN E1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.292200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 80.860 0.400 81.260 ;
    END
  END E1END[0]
  PIN E1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.292200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 82.540 0.400 82.940 ;
    END
  END E1END[1]
  PIN E1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.107600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 84.220 0.400 84.620 ;
    END
  END E1END[2]
  PIN E1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.320800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 85.900 0.400 86.300 ;
    END
  END E1END[3]
  PIN E2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.092000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 101.020 0.400 101.420 ;
    END
  END E2END[0]
  PIN E2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.305200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 102.700 0.400 103.100 ;
    END
  END E2END[1]
  PIN E2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.305200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 104.380 0.400 104.780 ;
    END
  END E2END[2]
  PIN E2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.333800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 106.060 0.400 106.460 ;
    END
  END E2END[3]
  PIN E2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.333800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 107.740 0.400 108.140 ;
    END
  END E2END[4]
  PIN E2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.272700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 109.420 0.400 109.820 ;
    END
  END E2END[5]
  PIN E2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.092000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 111.100 0.400 111.500 ;
    END
  END E2END[6]
  PIN E2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.079000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 112.780 0.400 113.180 ;
    END
  END E2END[7]
  PIN E2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.092000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 87.580 0.400 87.980 ;
    END
  END E2MID[0]
  PIN E2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.878800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 89.260 0.400 89.660 ;
    END
  END E2MID[1]
  PIN E2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 8.179600 ;
    ANTENNADIFFAREA 24.184799 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 90.940 0.400 91.340 ;
    END
  END E2MID[2]
  PIN E2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.092000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 92.620 0.400 93.020 ;
    END
  END E2MID[3]
  PIN E2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.878800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 94.300 0.400 94.700 ;
    END
  END E2MID[4]
  PIN E2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.878800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 95.980 0.400 96.380 ;
    END
  END E2MID[5]
  PIN E2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.371000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 97.660 0.400 98.060 ;
    END
  END E2MID[6]
  PIN E2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.865800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 99.340 0.400 99.740 ;
    END
  END E2MID[7]
  PIN E6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.172400 ;
    ANTENNADIFFAREA 18.138599 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 141.340 0.400 141.740 ;
    END
  END E6END[0]
  PIN E6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.848900 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 158.140 0.400 158.540 ;
    END
  END E6END[10]
  PIN E6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.848900 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 159.820 0.400 160.220 ;
    END
  END E6END[11]
  PIN E6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.696800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 143.020 0.400 143.420 ;
    END
  END E6END[1]
  PIN E6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.696800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 144.700 0.400 145.100 ;
    END
  END E6END[2]
  PIN E6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.696800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 146.380 0.400 146.780 ;
    END
  END E6END[3]
  PIN E6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.881400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 148.060 0.400 148.460 ;
    END
  END E6END[4]
  PIN E6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.881400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 149.740 0.400 150.140 ;
    END
  END E6END[5]
  PIN E6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.848900 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 151.420 0.400 151.820 ;
    END
  END E6END[6]
  PIN E6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.848900 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 153.100 0.400 153.500 ;
    END
  END E6END[7]
  PIN E6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.848900 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 154.780 0.400 155.180 ;
    END
  END E6END[8]
  PIN E6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.848900 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 156.460 0.400 156.860 ;
    END
  END E6END[9]
  PIN EE4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.665600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 114.460 0.400 114.860 ;
    END
  END EE4END[0]
  PIN EE4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.452400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 131.260 0.400 131.660 ;
    END
  END EE4END[10]
  PIN EE4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.452400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 132.940 0.400 133.340 ;
    END
  END EE4END[11]
  PIN EE4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.681200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 134.620 0.400 135.020 ;
    END
  END EE4END[12]
  PIN EE4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.681200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 136.300 0.400 136.700 ;
    END
  END EE4END[13]
  PIN EE4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.694200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 137.980 0.400 138.380 ;
    END
  END EE4END[14]
  PIN EE4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.681200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 139.660 0.400 140.060 ;
    END
  END EE4END[15]
  PIN EE4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.665600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 116.140 0.400 116.540 ;
    END
  END EE4END[1]
  PIN EE4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.678600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 117.820 0.400 118.220 ;
    END
  END EE4END[2]
  PIN EE4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.665600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 119.500 0.400 119.900 ;
    END
  END EE4END[3]
  PIN EE4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.452400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 121.180 0.400 121.580 ;
    END
  END EE4END[4]
  PIN EE4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.452400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 122.860 0.400 123.260 ;
    END
  END EE4END[5]
  PIN EE4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.452400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 124.540 0.400 124.940 ;
    END
  END EE4END[6]
  PIN EE4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.439400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 126.220 0.400 126.620 ;
    END
  END EE4END[7]
  PIN EE4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.452400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 127.900 0.400 128.300 ;
    END
  END EE4END[8]
  PIN EE4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.452400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 129.580 0.400 129.980 ;
    END
  END EE4END[9]
  PIN ENA_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 114.460 107.520 114.860 ;
    END
  END ENA_TT_PROJECT
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 161.500 0.400 161.900 ;
    END
  END FrameData[0]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 178.300 0.400 178.700 ;
    END
  END FrameData[10]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 179.980 0.400 180.380 ;
    END
  END FrameData[11]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 181.660 0.400 182.060 ;
    END
  END FrameData[12]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 183.340 0.400 183.740 ;
    END
  END FrameData[13]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 185.020 0.400 185.420 ;
    END
  END FrameData[14]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 186.700 0.400 187.100 ;
    END
  END FrameData[15]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 188.380 0.400 188.780 ;
    END
  END FrameData[16]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 190.060 0.400 190.460 ;
    END
  END FrameData[17]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 191.740 0.400 192.140 ;
    END
  END FrameData[18]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 193.420 0.400 193.820 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 163.180 0.400 163.580 ;
    END
  END FrameData[1]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 195.100 0.400 195.500 ;
    END
  END FrameData[20]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 196.780 0.400 197.180 ;
    END
  END FrameData[21]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.987700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 198.460 0.400 198.860 ;
    END
  END FrameData[22]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.987700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 200.140 0.400 200.540 ;
    END
  END FrameData[23]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.987700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 201.820 0.400 202.220 ;
    END
  END FrameData[24]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.987700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 203.500 0.400 203.900 ;
    END
  END FrameData[25]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.987700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 205.180 0.400 205.580 ;
    END
  END FrameData[26]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.987700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 206.860 0.400 207.260 ;
    END
  END FrameData[27]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.987700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 208.540 0.400 208.940 ;
    END
  END FrameData[28]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.987700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 210.220 0.400 210.620 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 164.860 0.400 165.260 ;
    END
  END FrameData[2]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.987700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 211.900 0.400 212.300 ;
    END
  END FrameData[30]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.987700 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 213.580 0.400 213.980 ;
    END
  END FrameData[31]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 166.540 0.400 166.940 ;
    END
  END FrameData[3]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 168.220 0.400 168.620 ;
    END
  END FrameData[4]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 169.900 0.400 170.300 ;
    END
  END FrameData[5]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 171.580 0.400 171.980 ;
    END
  END FrameData[6]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 173.260 0.400 173.660 ;
    END
  END FrameData[7]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 174.940 0.400 175.340 ;
    END
  END FrameData[8]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.807000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 176.620 0.400 177.020 ;
    END
  END FrameData[9]
  PIN FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 122.020 107.520 122.420 ;
    END
  END FrameData_O[0]
  PIN FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 147.220 107.520 147.620 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 149.740 107.520 150.140 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 152.260 107.520 152.660 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 154.780 107.520 155.180 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 157.300 107.520 157.700 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 159.820 107.520 160.220 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 162.340 107.520 162.740 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 164.860 107.520 165.260 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 167.380 107.520 167.780 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 169.900 107.520 170.300 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 124.540 107.520 124.940 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 172.420 107.520 172.820 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 174.940 107.520 175.340 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 177.460 107.520 177.860 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 179.980 107.520 180.380 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 182.500 107.520 182.900 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 185.020 107.520 185.420 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 187.540 107.520 187.940 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 190.060 107.520 190.460 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 192.580 107.520 192.980 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 195.100 107.520 195.500 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 127.060 107.520 127.460 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 197.620 107.520 198.020 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 200.140 107.520 200.540 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 129.580 107.520 129.980 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 132.100 107.520 132.500 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 134.620 107.520 135.020 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 137.140 107.520 137.540 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 139.660 107.520 140.060 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 142.180 107.520 142.580 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 144.700 107.520 145.100 ;
    END
  END FrameData_O[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.753500 ;
    PORT
      LAYER Metal2 ;
        RECT 79.000 0.000 79.400 0.400 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.789100 ;
    ANTENNADIFFAREA 2.015400 ;
    PORT
      LAYER Metal2 ;
        RECT 88.600 0.000 89.000 0.400 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.789100 ;
    ANTENNADIFFAREA 2.015400 ;
    PORT
      LAYER Metal2 ;
        RECT 89.560 0.000 89.960 0.400 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.789100 ;
    ANTENNADIFFAREA 2.015400 ;
    PORT
      LAYER Metal2 ;
        RECT 90.520 0.000 90.920 0.400 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.789100 ;
    ANTENNADIFFAREA 2.015400 ;
    PORT
      LAYER Metal2 ;
        RECT 91.480 0.000 91.880 0.400 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 92.440 0.000 92.840 0.400 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 93.400 0.000 93.800 0.400 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 94.360 0.000 94.760 0.400 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.789100 ;
    ANTENNADIFFAREA 2.015400 ;
    PORT
      LAYER Metal2 ;
        RECT 95.320 0.000 95.720 0.400 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.789100 ;
    ANTENNADIFFAREA 2.015400 ;
    PORT
      LAYER Metal2 ;
        RECT 96.280 0.000 96.680 0.400 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.789100 ;
    ANTENNADIFFAREA 2.015400 ;
    PORT
      LAYER Metal2 ;
        RECT 97.240 0.000 97.640 0.400 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.753500 ;
    PORT
      LAYER Metal2 ;
        RECT 79.960 0.000 80.360 0.400 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.753500 ;
    PORT
      LAYER Metal2 ;
        RECT 80.920 0.000 81.320 0.400 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.753500 ;
    PORT
      LAYER Metal2 ;
        RECT 81.880 0.000 82.280 0.400 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.753500 ;
    PORT
      LAYER Metal2 ;
        RECT 82.840 0.000 83.240 0.400 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.753500 ;
    PORT
      LAYER Metal2 ;
        RECT 83.800 0.000 84.200 0.400 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.753500 ;
    PORT
      LAYER Metal2 ;
        RECT 84.760 0.000 85.160 0.400 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.753500 ;
    PORT
      LAYER Metal2 ;
        RECT 85.720 0.000 86.120 0.400 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.753500 ;
    PORT
      LAYER Metal2 ;
        RECT 86.680 0.000 87.080 0.400 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.234700 ;
    PORT
      LAYER Metal2 ;
        RECT 87.640 0.000 88.040 0.400 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 79.000 214.640 79.400 215.040 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 88.600 214.640 89.000 215.040 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 89.560 214.640 89.960 215.040 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 90.520 214.640 90.920 215.040 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 91.480 214.640 91.880 215.040 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 92.440 214.640 92.840 215.040 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 93.400 214.640 93.800 215.040 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 94.360 214.640 94.760 215.040 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 95.320 214.640 95.720 215.040 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 96.280 214.640 96.680 215.040 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 97.240 214.640 97.640 215.040 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 79.960 214.640 80.360 215.040 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 80.920 214.640 81.320 215.040 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 81.880 214.640 82.280 215.040 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 82.840 214.640 83.240 215.040 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 83.800 214.640 84.200 215.040 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 84.760 214.640 85.160 215.040 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 85.720 214.640 86.120 215.040 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 86.680 214.640 87.080 215.040 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 87.640 214.640 88.040 215.040 ;
    END
  END FrameStrobe_O[9]
  PIN N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 8.920 214.640 9.320 215.040 ;
    END
  END N1BEG[0]
  PIN N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 9.880 214.640 10.280 215.040 ;
    END
  END N1BEG[1]
  PIN N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 10.840 214.640 11.240 215.040 ;
    END
  END N1BEG[2]
  PIN N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 11.800 214.640 12.200 215.040 ;
    END
  END N1BEG[3]
  PIN N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.311700 ;
    PORT
      LAYER Metal2 ;
        RECT 8.920 0.000 9.320 0.400 ;
    END
  END N1END[0]
  PIN N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.311700 ;
    PORT
      LAYER Metal2 ;
        RECT 9.880 0.000 10.280 0.400 ;
    END
  END N1END[1]
  PIN N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.311700 ;
    PORT
      LAYER Metal2 ;
        RECT 10.840 0.000 11.240 0.400 ;
    END
  END N1END[2]
  PIN N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.311700 ;
    PORT
      LAYER Metal2 ;
        RECT 11.800 0.000 12.200 0.400 ;
    END
  END N1END[3]
  PIN N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 12.760 214.640 13.160 215.040 ;
    END
  END N2BEG[0]
  PIN N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 13.720 214.640 14.120 215.040 ;
    END
  END N2BEG[1]
  PIN N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 14.680 214.640 15.080 215.040 ;
    END
  END N2BEG[2]
  PIN N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 15.640 214.640 16.040 215.040 ;
    END
  END N2BEG[3]
  PIN N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 16.600 214.640 17.000 215.040 ;
    END
  END N2BEG[4]
  PIN N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 17.560 214.640 17.960 215.040 ;
    END
  END N2BEG[5]
  PIN N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 18.520 214.640 18.920 215.040 ;
    END
  END N2BEG[6]
  PIN N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 19.480 214.640 19.880 215.040 ;
    END
  END N2BEG[7]
  PIN N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 20.440 214.640 20.840 215.040 ;
    END
  END N2BEGb[0]
  PIN N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 21.400 214.640 21.800 215.040 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 22.360 214.640 22.760 215.040 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 23.320 214.640 23.720 215.040 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 24.280 214.640 24.680 215.040 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 25.240 214.640 25.640 215.040 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 26.200 214.640 26.600 215.040 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 27.160 214.640 27.560 215.040 ;
    END
  END N2BEGb[7]
  PIN N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.821600 ;
    ANTENNADIFFAREA 2.015400 ;
    PORT
      LAYER Metal2 ;
        RECT 20.440 0.000 20.840 0.400 ;
    END
  END N2END[0]
  PIN N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 21.400 0.000 21.800 0.400 ;
    END
  END N2END[1]
  PIN N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal2 ;
        RECT 22.360 0.000 22.760 0.400 ;
    END
  END N2END[2]
  PIN N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal2 ;
        RECT 23.320 0.000 23.720 0.400 ;
    END
  END N2END[3]
  PIN N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 24.280 0.000 24.680 0.400 ;
    END
  END N2END[4]
  PIN N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 25.240 0.000 25.640 0.400 ;
    END
  END N2END[5]
  PIN N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 26.200 0.000 26.600 0.400 ;
    END
  END N2END[6]
  PIN N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 27.160 0.000 27.560 0.400 ;
    END
  END N2END[7]
  PIN N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.393900 ;
    PORT
      LAYER Metal2 ;
        RECT 12.760 0.000 13.160 0.400 ;
    END
  END N2MID[0]
  PIN N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.393900 ;
    PORT
      LAYER Metal2 ;
        RECT 13.720 0.000 14.120 0.400 ;
    END
  END N2MID[1]
  PIN N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.219100 ;
    ANTENNADIFFAREA 6.046200 ;
    PORT
      LAYER Metal2 ;
        RECT 14.680 0.000 15.080 0.400 ;
    END
  END N2MID[2]
  PIN N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.393900 ;
    PORT
      LAYER Metal2 ;
        RECT 15.640 0.000 16.040 0.400 ;
    END
  END N2MID[3]
  PIN N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.827500 ;
    ANTENNADIFFAREA 8.061600 ;
    PORT
      LAYER Metal2 ;
        RECT 16.600 0.000 17.000 0.400 ;
    END
  END N2MID[4]
  PIN N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.219100 ;
    ANTENNADIFFAREA 6.046200 ;
    PORT
      LAYER Metal2 ;
        RECT 17.560 0.000 17.960 0.400 ;
    END
  END N2MID[5]
  PIN N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.848900 ;
    PORT
      LAYER Metal2 ;
        RECT 18.520 0.000 18.920 0.400 ;
    END
  END N2MID[6]
  PIN N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.393900 ;
    PORT
      LAYER Metal2 ;
        RECT 19.480 0.000 19.880 0.400 ;
    END
  END N2MID[7]
  PIN N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 28.120 214.640 28.520 215.040 ;
    END
  END N4BEG[0]
  PIN N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 37.720 214.640 38.120 215.040 ;
    END
  END N4BEG[10]
  PIN N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 38.680 214.640 39.080 215.040 ;
    END
  END N4BEG[11]
  PIN N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 39.640 214.640 40.040 215.040 ;
    END
  END N4BEG[12]
  PIN N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 40.600 214.640 41.000 215.040 ;
    END
  END N4BEG[13]
  PIN N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 41.560 214.640 41.960 215.040 ;
    END
  END N4BEG[14]
  PIN N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 42.520 214.640 42.920 215.040 ;
    END
  END N4BEG[15]
  PIN N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 29.080 214.640 29.480 215.040 ;
    END
  END N4BEG[1]
  PIN N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 30.040 214.640 30.440 215.040 ;
    END
  END N4BEG[2]
  PIN N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 31.000 214.640 31.400 215.040 ;
    END
  END N4BEG[3]
  PIN N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 31.960 214.640 32.360 215.040 ;
    END
  END N4BEG[4]
  PIN N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 32.920 214.640 33.320 215.040 ;
    END
  END N4BEG[5]
  PIN N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 33.880 214.640 34.280 215.040 ;
    END
  END N4BEG[6]
  PIN N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 34.840 214.640 35.240 215.040 ;
    END
  END N4BEG[7]
  PIN N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 35.800 214.640 36.200 215.040 ;
    END
  END N4BEG[8]
  PIN N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 36.760 214.640 37.160 215.040 ;
    END
  END N4BEG[9]
  PIN N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal2 ;
        RECT 28.120 0.000 28.520 0.400 ;
    END
  END N4END[0]
  PIN N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.789100 ;
    ANTENNADIFFAREA 2.015400 ;
    PORT
      LAYER Metal2 ;
        RECT 37.720 0.000 38.120 0.400 ;
    END
  END N4END[10]
  PIN N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.789100 ;
    ANTENNADIFFAREA 2.015400 ;
    PORT
      LAYER Metal2 ;
        RECT 38.680 0.000 39.080 0.400 ;
    END
  END N4END[11]
  PIN N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.789100 ;
    ANTENNADIFFAREA 2.015400 ;
    PORT
      LAYER Metal2 ;
        RECT 39.640 0.000 40.040 0.400 ;
    END
  END N4END[12]
  PIN N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.789100 ;
    ANTENNADIFFAREA 2.015400 ;
    PORT
      LAYER Metal2 ;
        RECT 40.600 0.000 41.000 0.400 ;
    END
  END N4END[13]
  PIN N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 41.560 0.000 41.960 0.400 ;
    END
  END N4END[14]
  PIN N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.789100 ;
    ANTENNADIFFAREA 2.015400 ;
    PORT
      LAYER Metal2 ;
        RECT 42.520 0.000 42.920 0.400 ;
    END
  END N4END[15]
  PIN N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal2 ;
        RECT 29.080 0.000 29.480 0.400 ;
    END
  END N4END[1]
  PIN N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal2 ;
        RECT 30.040 0.000 30.440 0.400 ;
    END
  END N4END[2]
  PIN N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal2 ;
        RECT 31.000 0.000 31.400 0.400 ;
    END
  END N4END[3]
  PIN N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.789100 ;
    ANTENNADIFFAREA 2.015400 ;
    PORT
      LAYER Metal2 ;
        RECT 31.960 0.000 32.360 0.400 ;
    END
  END N4END[4]
  PIN N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.789100 ;
    ANTENNADIFFAREA 2.015400 ;
    PORT
      LAYER Metal2 ;
        RECT 32.920 0.000 33.320 0.400 ;
    END
  END N4END[5]
  PIN N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 33.880 0.000 34.280 0.400 ;
    END
  END N4END[6]
  PIN N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.789100 ;
    ANTENNADIFFAREA 2.015400 ;
    PORT
      LAYER Metal2 ;
        RECT 34.840 0.000 35.240 0.400 ;
    END
  END N4END[7]
  PIN N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.789100 ;
    ANTENNADIFFAREA 2.015400 ;
    PORT
      LAYER Metal2 ;
        RECT 35.800 0.000 36.200 0.400 ;
    END
  END N4END[8]
  PIN N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.789100 ;
    ANTENNADIFFAREA 2.015400 ;
    PORT
      LAYER Metal2 ;
        RECT 36.760 0.000 37.160 0.400 ;
    END
  END N4END[9]
  PIN RST_N_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 119.500 107.520 119.900 ;
    END
  END RST_N_TT_PROJECT
  PIN S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 43.480 0.000 43.880 0.400 ;
    END
  END S1BEG[0]
  PIN S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 44.440 0.000 44.840 0.400 ;
    END
  END S1BEG[1]
  PIN S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 45.400 0.000 45.800 0.400 ;
    END
  END S1BEG[2]
  PIN S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 46.360 0.000 46.760 0.400 ;
    END
  END S1BEG[3]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.307800 ;
    PORT
      LAYER Metal2 ;
        RECT 43.480 214.640 43.880 215.040 ;
    END
  END S1END[0]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.307800 ;
    PORT
      LAYER Metal2 ;
        RECT 44.440 214.640 44.840 215.040 ;
    END
  END S1END[1]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.307800 ;
    PORT
      LAYER Metal2 ;
        RECT 45.400 214.640 45.800 215.040 ;
    END
  END S1END[2]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.307800 ;
    PORT
      LAYER Metal2 ;
        RECT 46.360 214.640 46.760 215.040 ;
    END
  END S1END[3]
  PIN S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 47.320 0.000 47.720 0.400 ;
    END
  END S2BEG[0]
  PIN S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 48.280 0.000 48.680 0.400 ;
    END
  END S2BEG[1]
  PIN S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 49.240 0.000 49.640 0.400 ;
    END
  END S2BEG[2]
  PIN S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 50.200 0.000 50.600 0.400 ;
    END
  END S2BEG[3]
  PIN S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 51.160 0.000 51.560 0.400 ;
    END
  END S2BEG[4]
  PIN S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 52.120 0.000 52.520 0.400 ;
    END
  END S2BEG[5]
  PIN S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 53.080 0.000 53.480 0.400 ;
    END
  END S2BEG[6]
  PIN S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 54.040 0.000 54.440 0.400 ;
    END
  END S2BEG[7]
  PIN S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 55.000 0.000 55.400 0.400 ;
    END
  END S2BEGb[0]
  PIN S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 55.960 0.000 56.360 0.400 ;
    END
  END S2BEGb[1]
  PIN S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 56.920 0.000 57.320 0.400 ;
    END
  END S2BEGb[2]
  PIN S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 57.880 0.000 58.280 0.400 ;
    END
  END S2BEGb[3]
  PIN S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 58.840 0.000 59.240 0.400 ;
    END
  END S2BEGb[4]
  PIN S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 59.800 0.000 60.200 0.400 ;
    END
  END S2BEGb[5]
  PIN S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 60.760 0.000 61.160 0.400 ;
    END
  END S2BEGb[6]
  PIN S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 61.720 0.000 62.120 0.400 ;
    END
  END S2BEGb[7]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 55.000 214.640 55.400 215.040 ;
    END
  END S2END[0]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 55.960 214.640 56.360 215.040 ;
    END
  END S2END[1]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.455000 ;
    PORT
      LAYER Metal2 ;
        RECT 56.920 214.640 57.320 215.040 ;
    END
  END S2END[2]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.455000 ;
    PORT
      LAYER Metal2 ;
        RECT 57.880 214.640 58.280 215.040 ;
    END
  END S2END[3]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 58.840 214.640 59.240 215.040 ;
    END
  END S2END[4]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 59.800 214.640 60.200 215.040 ;
    END
  END S2END[5]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 60.760 214.640 61.160 215.040 ;
    END
  END S2END[6]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 61.720 214.640 62.120 215.040 ;
    END
  END S2END[7]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.148500 ;
    ANTENNADIFFAREA 18.138599 ;
    PORT
      LAYER Metal2 ;
        RECT 47.320 214.640 47.720 215.040 ;
    END
  END S2MID[0]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.827500 ;
    ANTENNADIFFAREA 8.061600 ;
    PORT
      LAYER Metal2 ;
        RECT 48.280 214.640 48.680 215.040 ;
    END
  END S2MID[1]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.610700 ;
    ANTENNADIFFAREA 4.030800 ;
    PORT
      LAYER Metal2 ;
        RECT 49.240 214.640 49.640 215.040 ;
    END
  END S2MID[2]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.393900 ;
    PORT
      LAYER Metal2 ;
        RECT 50.200 214.640 50.600 215.040 ;
    END
  END S2MID[3]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.610700 ;
    ANTENNADIFFAREA 4.030800 ;
    PORT
      LAYER Metal2 ;
        RECT 51.160 214.640 51.560 215.040 ;
    END
  END S2MID[4]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.827500 ;
    ANTENNADIFFAREA 8.061600 ;
    PORT
      LAYER Metal2 ;
        RECT 52.120 214.640 52.520 215.040 ;
    END
  END S2MID[5]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.827500 ;
    ANTENNADIFFAREA 8.061600 ;
    PORT
      LAYER Metal2 ;
        RECT 53.080 214.640 53.480 215.040 ;
    END
  END S2MID[6]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.610700 ;
    ANTENNADIFFAREA 4.030800 ;
    PORT
      LAYER Metal2 ;
        RECT 54.040 214.640 54.440 215.040 ;
    END
  END S2MID[7]
  PIN S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 62.680 0.000 63.080 0.400 ;
    END
  END S4BEG[0]
  PIN S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 72.280 0.000 72.680 0.400 ;
    END
  END S4BEG[10]
  PIN S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 73.240 0.000 73.640 0.400 ;
    END
  END S4BEG[11]
  PIN S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 74.200 0.000 74.600 0.400 ;
    END
  END S4BEG[12]
  PIN S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 75.160 0.000 75.560 0.400 ;
    END
  END S4BEG[13]
  PIN S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 76.120 0.000 76.520 0.400 ;
    END
  END S4BEG[14]
  PIN S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 77.080 0.000 77.480 0.400 ;
    END
  END S4BEG[15]
  PIN S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 63.640 0.000 64.040 0.400 ;
    END
  END S4BEG[1]
  PIN S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 64.600 0.000 65.000 0.400 ;
    END
  END S4BEG[2]
  PIN S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 65.560 0.000 65.960 0.400 ;
    END
  END S4BEG[3]
  PIN S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 66.520 0.000 66.920 0.400 ;
    END
  END S4BEG[4]
  PIN S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 67.480 0.000 67.880 0.400 ;
    END
  END S4BEG[5]
  PIN S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 68.440 0.000 68.840 0.400 ;
    END
  END S4BEG[6]
  PIN S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 69.400 0.000 69.800 0.400 ;
    END
  END S4BEG[7]
  PIN S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 70.360 0.000 70.760 0.400 ;
    END
  END S4BEG[8]
  PIN S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 71.320 0.000 71.720 0.400 ;
    END
  END S4BEG[9]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal2 ;
        RECT 62.680 214.640 63.080 215.040 ;
    END
  END S4END[0]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 72.280 214.640 72.680 215.040 ;
    END
  END S4END[10]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 73.240 214.640 73.640 215.040 ;
    END
  END S4END[11]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 74.200 214.640 74.600 215.040 ;
    END
  END S4END[12]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 75.160 214.640 75.560 215.040 ;
    END
  END S4END[13]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 76.120 214.640 76.520 215.040 ;
    END
  END S4END[14]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 77.080 214.640 77.480 215.040 ;
    END
  END S4END[15]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal2 ;
        RECT 63.640 214.640 64.040 215.040 ;
    END
  END S4END[1]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal2 ;
        RECT 64.600 214.640 65.000 215.040 ;
    END
  END S4END[2]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal2 ;
        RECT 65.560 214.640 65.960 215.040 ;
    END
  END S4END[3]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 66.520 214.640 66.920 215.040 ;
    END
  END S4END[4]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 67.480 214.640 67.880 215.040 ;
    END
  END S4END[5]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 68.440 214.640 68.840 215.040 ;
    END
  END S4END[6]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 69.400 214.640 69.800 215.040 ;
    END
  END S4END[7]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 70.360 214.640 70.760 215.040 ;
    END
  END S4END[8]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 71.320 214.640 71.720 215.040 ;
    END
  END S4END[9]
  PIN UIO_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.958400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 94.300 107.520 94.700 ;
    END
  END UIO_IN_TT_PROJECT0
  PIN UIO_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.958400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 96.820 107.520 97.220 ;
    END
  END UIO_IN_TT_PROJECT1
  PIN UIO_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.958400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 99.340 107.520 99.740 ;
    END
  END UIO_IN_TT_PROJECT2
  PIN UIO_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.958400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 101.860 107.520 102.260 ;
    END
  END UIO_IN_TT_PROJECT3
  PIN UIO_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.958400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 104.380 107.520 104.780 ;
    END
  END UIO_IN_TT_PROJECT4
  PIN UIO_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.958400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 106.900 107.520 107.300 ;
    END
  END UIO_IN_TT_PROJECT5
  PIN UIO_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.958400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 109.420 107.520 109.820 ;
    END
  END UIO_IN_TT_PROJECT6
  PIN UIO_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.958400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 111.940 107.520 112.340 ;
    END
  END UIO_IN_TT_PROJECT7
  PIN UIO_OE_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.033500 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 53.980 107.520 54.380 ;
    END
  END UIO_OE_TT_PROJECT0
  PIN UIO_OE_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.046500 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 56.500 107.520 56.900 ;
    END
  END UIO_OE_TT_PROJECT1
  PIN UIO_OE_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.046500 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 59.020 107.520 59.420 ;
    END
  END UIO_OE_TT_PROJECT2
  PIN UIO_OE_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.046500 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 61.540 107.520 61.940 ;
    END
  END UIO_OE_TT_PROJECT3
  PIN UIO_OE_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.046500 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 64.060 107.520 64.460 ;
    END
  END UIO_OE_TT_PROJECT4
  PIN UIO_OE_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.046500 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 66.580 107.520 66.980 ;
    END
  END UIO_OE_TT_PROJECT5
  PIN UIO_OE_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.046500 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 69.100 107.520 69.500 ;
    END
  END UIO_OE_TT_PROJECT6
  PIN UIO_OE_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.046500 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 71.620 107.520 72.020 ;
    END
  END UIO_OE_TT_PROJECT7
  PIN UIO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.292200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 33.820 107.520 34.220 ;
    END
  END UIO_OUT_TT_PROJECT0
  PIN UIO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.292200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 36.340 107.520 36.740 ;
    END
  END UIO_OUT_TT_PROJECT1
  PIN UIO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.292200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 38.860 107.520 39.260 ;
    END
  END UIO_OUT_TT_PROJECT2
  PIN UIO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.292200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 41.380 107.520 41.780 ;
    END
  END UIO_OUT_TT_PROJECT3
  PIN UIO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.292200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 43.900 107.520 44.300 ;
    END
  END UIO_OUT_TT_PROJECT4
  PIN UIO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.292200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 46.420 107.520 46.820 ;
    END
  END UIO_OUT_TT_PROJECT5
  PIN UIO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.292200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 48.940 107.520 49.340 ;
    END
  END UIO_OUT_TT_PROJECT6
  PIN UIO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 51.460 107.520 51.860 ;
    END
  END UIO_OUT_TT_PROJECT7
  PIN UI_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.958400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 74.140 107.520 74.540 ;
    END
  END UI_IN_TT_PROJECT0
  PIN UI_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.958400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 76.660 107.520 77.060 ;
    END
  END UI_IN_TT_PROJECT1
  PIN UI_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.958400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 79.180 107.520 79.580 ;
    END
  END UI_IN_TT_PROJECT2
  PIN UI_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.958400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 81.700 107.520 82.100 ;
    END
  END UI_IN_TT_PROJECT3
  PIN UI_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.958400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 84.220 107.520 84.620 ;
    END
  END UI_IN_TT_PROJECT4
  PIN UI_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.958400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 86.740 107.520 87.140 ;
    END
  END UI_IN_TT_PROJECT5
  PIN UI_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.958400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 89.260 107.520 89.660 ;
    END
  END UI_IN_TT_PROJECT6
  PIN UI_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.662000 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 91.780 107.520 92.180 ;
    END
  END UI_IN_TT_PROJECT7
  PIN UO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.197600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 13.660 107.520 14.060 ;
    END
  END UO_OUT_TT_PROJECT0
  PIN UO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.197600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 16.180 107.520 16.580 ;
    END
  END UO_OUT_TT_PROJECT1
  PIN UO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.881400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 18.700 107.520 19.100 ;
    END
  END UO_OUT_TT_PROJECT2
  PIN UO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.881400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 21.220 107.520 21.620 ;
    END
  END UO_OUT_TT_PROJECT3
  PIN UO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.131800 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 23.740 107.520 24.140 ;
    END
  END UO_OUT_TT_PROJECT4
  PIN UO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.197600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 26.260 107.520 26.660 ;
    END
  END UO_OUT_TT_PROJECT5
  PIN UO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.881400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 28.780 107.520 29.180 ;
    END
  END UO_OUT_TT_PROJECT6
  PIN UO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.094600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 31.300 107.520 31.700 ;
    END
  END UO_OUT_TT_PROJECT7
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.725400 ;
    PORT
      LAYER Metal2 ;
        RECT 78.040 0.000 78.440 0.400 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 78.040 214.640 78.440 215.040 ;
    END
  END UserCLKo
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER TopMetal1 ;
        RECT 24.460 0.000 26.660 215.040 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 100.060 0.000 102.260 215.040 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER TopMetal1 ;
        RECT 18.260 0.000 20.460 215.040 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 93.860 0.000 96.060 215.040 ;
    END
  END VPWR
  PIN W1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 0.220 0.400 0.620 ;
    END
  END W1BEG[0]
  PIN W1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1.900 0.400 2.300 ;
    END
  END W1BEG[1]
  PIN W1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 3.580 0.400 3.980 ;
    END
  END W1BEG[2]
  PIN W1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 5.260 0.400 5.660 ;
    END
  END W1BEG[3]
  PIN W2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 6.940 0.400 7.340 ;
    END
  END W2BEG[0]
  PIN W2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 8.620 0.400 9.020 ;
    END
  END W2BEG[1]
  PIN W2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 10.300 0.400 10.700 ;
    END
  END W2BEG[2]
  PIN W2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 11.980 0.400 12.380 ;
    END
  END W2BEG[3]
  PIN W2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 13.660 0.400 14.060 ;
    END
  END W2BEG[4]
  PIN W2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 15.340 0.400 15.740 ;
    END
  END W2BEG[5]
  PIN W2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 17.020 0.400 17.420 ;
    END
  END W2BEG[6]
  PIN W2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 18.700 0.400 19.100 ;
    END
  END W2BEG[7]
  PIN W2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 20.380 0.400 20.780 ;
    END
  END W2BEGb[0]
  PIN W2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 22.060 0.400 22.460 ;
    END
  END W2BEGb[1]
  PIN W2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 23.740 0.400 24.140 ;
    END
  END W2BEGb[2]
  PIN W2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 25.420 0.400 25.820 ;
    END
  END W2BEGb[3]
  PIN W2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 27.100 0.400 27.500 ;
    END
  END W2BEGb[4]
  PIN W2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 28.780 0.400 29.180 ;
    END
  END W2BEGb[5]
  PIN W2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 30.460 0.400 30.860 ;
    END
  END W2BEGb[6]
  PIN W2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 32.140 0.400 32.540 ;
    END
  END W2BEGb[7]
  PIN W6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 60.700 0.400 61.100 ;
    END
  END W6BEG[0]
  PIN W6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 77.500 0.400 77.900 ;
    END
  END W6BEG[10]
  PIN W6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 79.180 0.400 79.580 ;
    END
  END W6BEG[11]
  PIN W6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 62.380 0.400 62.780 ;
    END
  END W6BEG[1]
  PIN W6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 64.060 0.400 64.460 ;
    END
  END W6BEG[2]
  PIN W6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 65.740 0.400 66.140 ;
    END
  END W6BEG[3]
  PIN W6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 67.420 0.400 67.820 ;
    END
  END W6BEG[4]
  PIN W6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 69.100 0.400 69.500 ;
    END
  END W6BEG[5]
  PIN W6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 70.780 0.400 71.180 ;
    END
  END W6BEG[6]
  PIN W6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 72.460 0.400 72.860 ;
    END
  END W6BEG[7]
  PIN W6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 74.140 0.400 74.540 ;
    END
  END W6BEG[8]
  PIN W6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 75.820 0.400 76.220 ;
    END
  END W6BEG[9]
  PIN WW4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 33.820 0.400 34.220 ;
    END
  END WW4BEG[0]
  PIN WW4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 50.620 0.400 51.020 ;
    END
  END WW4BEG[10]
  PIN WW4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 52.300 0.400 52.700 ;
    END
  END WW4BEG[11]
  PIN WW4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 53.980 0.400 54.380 ;
    END
  END WW4BEG[12]
  PIN WW4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 55.660 0.400 56.060 ;
    END
  END WW4BEG[13]
  PIN WW4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 57.340 0.400 57.740 ;
    END
  END WW4BEG[14]
  PIN WW4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 59.020 0.400 59.420 ;
    END
  END WW4BEG[15]
  PIN WW4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 35.500 0.400 35.900 ;
    END
  END WW4BEG[1]
  PIN WW4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 37.180 0.400 37.580 ;
    END
  END WW4BEG[2]
  PIN WW4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 38.860 0.400 39.260 ;
    END
  END WW4BEG[3]
  PIN WW4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 40.540 0.400 40.940 ;
    END
  END WW4BEG[4]
  PIN WW4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 42.220 0.400 42.620 ;
    END
  END WW4BEG[5]
  PIN WW4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 43.900 0.400 44.300 ;
    END
  END WW4BEG[6]
  PIN WW4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 45.580 0.400 45.980 ;
    END
  END WW4BEG[7]
  PIN WW4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 47.260 0.400 47.660 ;
    END
  END WW4BEG[8]
  PIN WW4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 48.940 0.400 49.340 ;
    END
  END WW4BEG[9]
  OBS
      LAYER GatPoly ;
        RECT 5.760 3.630 101.760 208.050 ;
      LAYER Metal1 ;
        RECT 5.760 3.560 102.260 208.120 ;
      LAYER Metal2 ;
        RECT 0.375 214.430 8.710 214.640 ;
        RECT 9.530 214.430 9.670 214.640 ;
        RECT 10.490 214.430 10.630 214.640 ;
        RECT 11.450 214.430 11.590 214.640 ;
        RECT 12.410 214.430 12.550 214.640 ;
        RECT 13.370 214.430 13.510 214.640 ;
        RECT 14.330 214.430 14.470 214.640 ;
        RECT 15.290 214.430 15.430 214.640 ;
        RECT 16.250 214.430 16.390 214.640 ;
        RECT 17.210 214.430 17.350 214.640 ;
        RECT 18.170 214.430 18.310 214.640 ;
        RECT 19.130 214.430 19.270 214.640 ;
        RECT 20.090 214.430 20.230 214.640 ;
        RECT 21.050 214.430 21.190 214.640 ;
        RECT 22.010 214.430 22.150 214.640 ;
        RECT 22.970 214.430 23.110 214.640 ;
        RECT 23.930 214.430 24.070 214.640 ;
        RECT 24.890 214.430 25.030 214.640 ;
        RECT 25.850 214.430 25.990 214.640 ;
        RECT 26.810 214.430 26.950 214.640 ;
        RECT 27.770 214.430 27.910 214.640 ;
        RECT 28.730 214.430 28.870 214.640 ;
        RECT 29.690 214.430 29.830 214.640 ;
        RECT 30.650 214.430 30.790 214.640 ;
        RECT 31.610 214.430 31.750 214.640 ;
        RECT 32.570 214.430 32.710 214.640 ;
        RECT 33.530 214.430 33.670 214.640 ;
        RECT 34.490 214.430 34.630 214.640 ;
        RECT 35.450 214.430 35.590 214.640 ;
        RECT 36.410 214.430 36.550 214.640 ;
        RECT 37.370 214.430 37.510 214.640 ;
        RECT 38.330 214.430 38.470 214.640 ;
        RECT 39.290 214.430 39.430 214.640 ;
        RECT 40.250 214.430 40.390 214.640 ;
        RECT 41.210 214.430 41.350 214.640 ;
        RECT 42.170 214.430 42.310 214.640 ;
        RECT 43.130 214.430 43.270 214.640 ;
        RECT 44.090 214.430 44.230 214.640 ;
        RECT 45.050 214.430 45.190 214.640 ;
        RECT 46.010 214.430 46.150 214.640 ;
        RECT 46.970 214.430 47.110 214.640 ;
        RECT 47.930 214.430 48.070 214.640 ;
        RECT 48.890 214.430 49.030 214.640 ;
        RECT 49.850 214.430 49.990 214.640 ;
        RECT 50.810 214.430 50.950 214.640 ;
        RECT 51.770 214.430 51.910 214.640 ;
        RECT 52.730 214.430 52.870 214.640 ;
        RECT 53.690 214.430 53.830 214.640 ;
        RECT 54.650 214.430 54.790 214.640 ;
        RECT 55.610 214.430 55.750 214.640 ;
        RECT 56.570 214.430 56.710 214.640 ;
        RECT 57.530 214.430 57.670 214.640 ;
        RECT 58.490 214.430 58.630 214.640 ;
        RECT 59.450 214.430 59.590 214.640 ;
        RECT 60.410 214.430 60.550 214.640 ;
        RECT 61.370 214.430 61.510 214.640 ;
        RECT 62.330 214.430 62.470 214.640 ;
        RECT 63.290 214.430 63.430 214.640 ;
        RECT 64.250 214.430 64.390 214.640 ;
        RECT 65.210 214.430 65.350 214.640 ;
        RECT 66.170 214.430 66.310 214.640 ;
        RECT 67.130 214.430 67.270 214.640 ;
        RECT 68.090 214.430 68.230 214.640 ;
        RECT 69.050 214.430 69.190 214.640 ;
        RECT 70.010 214.430 70.150 214.640 ;
        RECT 70.970 214.430 71.110 214.640 ;
        RECT 71.930 214.430 72.070 214.640 ;
        RECT 72.890 214.430 73.030 214.640 ;
        RECT 73.850 214.430 73.990 214.640 ;
        RECT 74.810 214.430 74.950 214.640 ;
        RECT 75.770 214.430 75.910 214.640 ;
        RECT 76.730 214.430 76.870 214.640 ;
        RECT 77.690 214.430 77.830 214.640 ;
        RECT 78.650 214.430 78.790 214.640 ;
        RECT 79.610 214.430 79.750 214.640 ;
        RECT 80.570 214.430 80.710 214.640 ;
        RECT 81.530 214.430 81.670 214.640 ;
        RECT 82.490 214.430 82.630 214.640 ;
        RECT 83.450 214.430 83.590 214.640 ;
        RECT 84.410 214.430 84.550 214.640 ;
        RECT 85.370 214.430 85.510 214.640 ;
        RECT 86.330 214.430 86.470 214.640 ;
        RECT 87.290 214.430 87.430 214.640 ;
        RECT 88.250 214.430 88.390 214.640 ;
        RECT 89.210 214.430 89.350 214.640 ;
        RECT 90.170 214.430 90.310 214.640 ;
        RECT 91.130 214.430 91.270 214.640 ;
        RECT 92.090 214.430 92.230 214.640 ;
        RECT 93.050 214.430 93.190 214.640 ;
        RECT 94.010 214.430 94.150 214.640 ;
        RECT 94.970 214.430 95.110 214.640 ;
        RECT 95.930 214.430 96.070 214.640 ;
        RECT 96.890 214.430 97.030 214.640 ;
        RECT 97.850 214.430 107.145 214.640 ;
        RECT 0.375 0.610 107.145 214.430 ;
        RECT 0.375 0.400 8.710 0.610 ;
        RECT 9.530 0.400 9.670 0.610 ;
        RECT 10.490 0.400 10.630 0.610 ;
        RECT 11.450 0.400 11.590 0.610 ;
        RECT 12.410 0.400 12.550 0.610 ;
        RECT 13.370 0.400 13.510 0.610 ;
        RECT 14.330 0.400 14.470 0.610 ;
        RECT 15.290 0.400 15.430 0.610 ;
        RECT 16.250 0.400 16.390 0.610 ;
        RECT 17.210 0.400 17.350 0.610 ;
        RECT 18.170 0.400 18.310 0.610 ;
        RECT 19.130 0.400 19.270 0.610 ;
        RECT 20.090 0.400 20.230 0.610 ;
        RECT 21.050 0.400 21.190 0.610 ;
        RECT 22.010 0.400 22.150 0.610 ;
        RECT 22.970 0.400 23.110 0.610 ;
        RECT 23.930 0.400 24.070 0.610 ;
        RECT 24.890 0.400 25.030 0.610 ;
        RECT 25.850 0.400 25.990 0.610 ;
        RECT 26.810 0.400 26.950 0.610 ;
        RECT 27.770 0.400 27.910 0.610 ;
        RECT 28.730 0.400 28.870 0.610 ;
        RECT 29.690 0.400 29.830 0.610 ;
        RECT 30.650 0.400 30.790 0.610 ;
        RECT 31.610 0.400 31.750 0.610 ;
        RECT 32.570 0.400 32.710 0.610 ;
        RECT 33.530 0.400 33.670 0.610 ;
        RECT 34.490 0.400 34.630 0.610 ;
        RECT 35.450 0.400 35.590 0.610 ;
        RECT 36.410 0.400 36.550 0.610 ;
        RECT 37.370 0.400 37.510 0.610 ;
        RECT 38.330 0.400 38.470 0.610 ;
        RECT 39.290 0.400 39.430 0.610 ;
        RECT 40.250 0.400 40.390 0.610 ;
        RECT 41.210 0.400 41.350 0.610 ;
        RECT 42.170 0.400 42.310 0.610 ;
        RECT 43.130 0.400 43.270 0.610 ;
        RECT 44.090 0.400 44.230 0.610 ;
        RECT 45.050 0.400 45.190 0.610 ;
        RECT 46.010 0.400 46.150 0.610 ;
        RECT 46.970 0.400 47.110 0.610 ;
        RECT 47.930 0.400 48.070 0.610 ;
        RECT 48.890 0.400 49.030 0.610 ;
        RECT 49.850 0.400 49.990 0.610 ;
        RECT 50.810 0.400 50.950 0.610 ;
        RECT 51.770 0.400 51.910 0.610 ;
        RECT 52.730 0.400 52.870 0.610 ;
        RECT 53.690 0.400 53.830 0.610 ;
        RECT 54.650 0.400 54.790 0.610 ;
        RECT 55.610 0.400 55.750 0.610 ;
        RECT 56.570 0.400 56.710 0.610 ;
        RECT 57.530 0.400 57.670 0.610 ;
        RECT 58.490 0.400 58.630 0.610 ;
        RECT 59.450 0.400 59.590 0.610 ;
        RECT 60.410 0.400 60.550 0.610 ;
        RECT 61.370 0.400 61.510 0.610 ;
        RECT 62.330 0.400 62.470 0.610 ;
        RECT 63.290 0.400 63.430 0.610 ;
        RECT 64.250 0.400 64.390 0.610 ;
        RECT 65.210 0.400 65.350 0.610 ;
        RECT 66.170 0.400 66.310 0.610 ;
        RECT 67.130 0.400 67.270 0.610 ;
        RECT 68.090 0.400 68.230 0.610 ;
        RECT 69.050 0.400 69.190 0.610 ;
        RECT 70.010 0.400 70.150 0.610 ;
        RECT 70.970 0.400 71.110 0.610 ;
        RECT 71.930 0.400 72.070 0.610 ;
        RECT 72.890 0.400 73.030 0.610 ;
        RECT 73.850 0.400 73.990 0.610 ;
        RECT 74.810 0.400 74.950 0.610 ;
        RECT 75.770 0.400 75.910 0.610 ;
        RECT 76.730 0.400 76.870 0.610 ;
        RECT 77.690 0.400 77.830 0.610 ;
        RECT 78.650 0.400 78.790 0.610 ;
        RECT 79.610 0.400 79.750 0.610 ;
        RECT 80.570 0.400 80.710 0.610 ;
        RECT 81.530 0.400 81.670 0.610 ;
        RECT 82.490 0.400 82.630 0.610 ;
        RECT 83.450 0.400 83.590 0.610 ;
        RECT 84.410 0.400 84.550 0.610 ;
        RECT 85.370 0.400 85.510 0.610 ;
        RECT 86.330 0.400 86.470 0.610 ;
        RECT 87.290 0.400 87.430 0.610 ;
        RECT 88.250 0.400 88.390 0.610 ;
        RECT 89.210 0.400 89.350 0.610 ;
        RECT 90.170 0.400 90.310 0.610 ;
        RECT 91.130 0.400 91.270 0.610 ;
        RECT 92.090 0.400 92.230 0.610 ;
        RECT 93.050 0.400 93.190 0.610 ;
        RECT 94.010 0.400 94.150 0.610 ;
        RECT 94.970 0.400 95.110 0.610 ;
        RECT 95.930 0.400 96.070 0.610 ;
        RECT 96.890 0.400 97.030 0.610 ;
        RECT 97.850 0.400 107.145 0.610 ;
      LAYER Metal3 ;
        RECT 0.335 214.190 107.420 214.720 ;
        RECT 0.610 213.370 107.420 214.190 ;
        RECT 0.335 212.510 107.420 213.370 ;
        RECT 0.610 211.690 107.420 212.510 ;
        RECT 0.335 210.830 107.420 211.690 ;
        RECT 0.610 210.010 107.420 210.830 ;
        RECT 0.335 209.150 107.420 210.010 ;
        RECT 0.610 208.330 107.420 209.150 ;
        RECT 0.335 207.470 107.420 208.330 ;
        RECT 0.610 206.650 107.420 207.470 ;
        RECT 0.335 205.790 107.420 206.650 ;
        RECT 0.610 204.970 107.420 205.790 ;
        RECT 0.335 204.110 107.420 204.970 ;
        RECT 0.610 203.290 107.420 204.110 ;
        RECT 0.335 202.430 107.420 203.290 ;
        RECT 0.610 201.610 107.420 202.430 ;
        RECT 0.335 200.750 107.420 201.610 ;
        RECT 0.610 199.930 106.910 200.750 ;
        RECT 0.335 199.070 107.420 199.930 ;
        RECT 0.610 198.250 107.420 199.070 ;
        RECT 0.335 198.230 107.420 198.250 ;
        RECT 0.335 197.410 106.910 198.230 ;
        RECT 0.335 197.390 107.420 197.410 ;
        RECT 0.610 196.570 107.420 197.390 ;
        RECT 0.335 195.710 107.420 196.570 ;
        RECT 0.610 194.890 106.910 195.710 ;
        RECT 0.335 194.030 107.420 194.890 ;
        RECT 0.610 193.210 107.420 194.030 ;
        RECT 0.335 193.190 107.420 193.210 ;
        RECT 0.335 192.370 106.910 193.190 ;
        RECT 0.335 192.350 107.420 192.370 ;
        RECT 0.610 191.530 107.420 192.350 ;
        RECT 0.335 190.670 107.420 191.530 ;
        RECT 0.610 189.850 106.910 190.670 ;
        RECT 0.335 188.990 107.420 189.850 ;
        RECT 0.610 188.170 107.420 188.990 ;
        RECT 0.335 188.150 107.420 188.170 ;
        RECT 0.335 187.330 106.910 188.150 ;
        RECT 0.335 187.310 107.420 187.330 ;
        RECT 0.610 186.490 107.420 187.310 ;
        RECT 0.335 185.630 107.420 186.490 ;
        RECT 0.610 184.810 106.910 185.630 ;
        RECT 0.335 183.950 107.420 184.810 ;
        RECT 0.610 183.130 107.420 183.950 ;
        RECT 0.335 183.110 107.420 183.130 ;
        RECT 0.335 182.290 106.910 183.110 ;
        RECT 0.335 182.270 107.420 182.290 ;
        RECT 0.610 181.450 107.420 182.270 ;
        RECT 0.335 180.590 107.420 181.450 ;
        RECT 0.610 179.770 106.910 180.590 ;
        RECT 0.335 178.910 107.420 179.770 ;
        RECT 0.610 178.090 107.420 178.910 ;
        RECT 0.335 178.070 107.420 178.090 ;
        RECT 0.335 177.250 106.910 178.070 ;
        RECT 0.335 177.230 107.420 177.250 ;
        RECT 0.610 176.410 107.420 177.230 ;
        RECT 0.335 175.550 107.420 176.410 ;
        RECT 0.610 174.730 106.910 175.550 ;
        RECT 0.335 173.870 107.420 174.730 ;
        RECT 0.610 173.050 107.420 173.870 ;
        RECT 0.335 173.030 107.420 173.050 ;
        RECT 0.335 172.210 106.910 173.030 ;
        RECT 0.335 172.190 107.420 172.210 ;
        RECT 0.610 171.370 107.420 172.190 ;
        RECT 0.335 170.510 107.420 171.370 ;
        RECT 0.610 169.690 106.910 170.510 ;
        RECT 0.335 168.830 107.420 169.690 ;
        RECT 0.610 168.010 107.420 168.830 ;
        RECT 0.335 167.990 107.420 168.010 ;
        RECT 0.335 167.170 106.910 167.990 ;
        RECT 0.335 167.150 107.420 167.170 ;
        RECT 0.610 166.330 107.420 167.150 ;
        RECT 0.335 165.470 107.420 166.330 ;
        RECT 0.610 164.650 106.910 165.470 ;
        RECT 0.335 163.790 107.420 164.650 ;
        RECT 0.610 162.970 107.420 163.790 ;
        RECT 0.335 162.950 107.420 162.970 ;
        RECT 0.335 162.130 106.910 162.950 ;
        RECT 0.335 162.110 107.420 162.130 ;
        RECT 0.610 161.290 107.420 162.110 ;
        RECT 0.335 160.430 107.420 161.290 ;
        RECT 0.610 159.610 106.910 160.430 ;
        RECT 0.335 158.750 107.420 159.610 ;
        RECT 0.610 157.930 107.420 158.750 ;
        RECT 0.335 157.910 107.420 157.930 ;
        RECT 0.335 157.090 106.910 157.910 ;
        RECT 0.335 157.070 107.420 157.090 ;
        RECT 0.610 156.250 107.420 157.070 ;
        RECT 0.335 155.390 107.420 156.250 ;
        RECT 0.610 154.570 106.910 155.390 ;
        RECT 0.335 153.710 107.420 154.570 ;
        RECT 0.610 152.890 107.420 153.710 ;
        RECT 0.335 152.870 107.420 152.890 ;
        RECT 0.335 152.050 106.910 152.870 ;
        RECT 0.335 152.030 107.420 152.050 ;
        RECT 0.610 151.210 107.420 152.030 ;
        RECT 0.335 150.350 107.420 151.210 ;
        RECT 0.610 149.530 106.910 150.350 ;
        RECT 0.335 148.670 107.420 149.530 ;
        RECT 0.610 147.850 107.420 148.670 ;
        RECT 0.335 147.830 107.420 147.850 ;
        RECT 0.335 147.010 106.910 147.830 ;
        RECT 0.335 146.990 107.420 147.010 ;
        RECT 0.610 146.170 107.420 146.990 ;
        RECT 0.335 145.310 107.420 146.170 ;
        RECT 0.610 144.490 106.910 145.310 ;
        RECT 0.335 143.630 107.420 144.490 ;
        RECT 0.610 142.810 107.420 143.630 ;
        RECT 0.335 142.790 107.420 142.810 ;
        RECT 0.335 141.970 106.910 142.790 ;
        RECT 0.335 141.950 107.420 141.970 ;
        RECT 0.610 141.130 107.420 141.950 ;
        RECT 0.335 140.270 107.420 141.130 ;
        RECT 0.610 139.450 106.910 140.270 ;
        RECT 0.335 138.590 107.420 139.450 ;
        RECT 0.610 137.770 107.420 138.590 ;
        RECT 0.335 137.750 107.420 137.770 ;
        RECT 0.335 136.930 106.910 137.750 ;
        RECT 0.335 136.910 107.420 136.930 ;
        RECT 0.610 136.090 107.420 136.910 ;
        RECT 0.335 135.230 107.420 136.090 ;
        RECT 0.610 134.410 106.910 135.230 ;
        RECT 0.335 133.550 107.420 134.410 ;
        RECT 0.610 132.730 107.420 133.550 ;
        RECT 0.335 132.710 107.420 132.730 ;
        RECT 0.335 131.890 106.910 132.710 ;
        RECT 0.335 131.870 107.420 131.890 ;
        RECT 0.610 131.050 107.420 131.870 ;
        RECT 0.335 130.190 107.420 131.050 ;
        RECT 0.610 129.370 106.910 130.190 ;
        RECT 0.335 128.510 107.420 129.370 ;
        RECT 0.610 127.690 107.420 128.510 ;
        RECT 0.335 127.670 107.420 127.690 ;
        RECT 0.335 126.850 106.910 127.670 ;
        RECT 0.335 126.830 107.420 126.850 ;
        RECT 0.610 126.010 107.420 126.830 ;
        RECT 0.335 125.150 107.420 126.010 ;
        RECT 0.610 124.330 106.910 125.150 ;
        RECT 0.335 123.470 107.420 124.330 ;
        RECT 0.610 122.650 107.420 123.470 ;
        RECT 0.335 122.630 107.420 122.650 ;
        RECT 0.335 121.810 106.910 122.630 ;
        RECT 0.335 121.790 107.420 121.810 ;
        RECT 0.610 120.970 107.420 121.790 ;
        RECT 0.335 120.110 107.420 120.970 ;
        RECT 0.610 119.290 106.910 120.110 ;
        RECT 0.335 118.430 107.420 119.290 ;
        RECT 0.610 117.610 107.420 118.430 ;
        RECT 0.335 117.590 107.420 117.610 ;
        RECT 0.335 116.770 106.910 117.590 ;
        RECT 0.335 116.750 107.420 116.770 ;
        RECT 0.610 115.930 107.420 116.750 ;
        RECT 0.335 115.070 107.420 115.930 ;
        RECT 0.610 114.250 106.910 115.070 ;
        RECT 0.335 113.390 107.420 114.250 ;
        RECT 0.610 112.570 107.420 113.390 ;
        RECT 0.335 112.550 107.420 112.570 ;
        RECT 0.335 111.730 106.910 112.550 ;
        RECT 0.335 111.710 107.420 111.730 ;
        RECT 0.610 110.890 107.420 111.710 ;
        RECT 0.335 110.030 107.420 110.890 ;
        RECT 0.610 109.210 106.910 110.030 ;
        RECT 0.335 108.350 107.420 109.210 ;
        RECT 0.610 107.530 107.420 108.350 ;
        RECT 0.335 107.510 107.420 107.530 ;
        RECT 0.335 106.690 106.910 107.510 ;
        RECT 0.335 106.670 107.420 106.690 ;
        RECT 0.610 105.850 107.420 106.670 ;
        RECT 0.335 104.990 107.420 105.850 ;
        RECT 0.610 104.170 106.910 104.990 ;
        RECT 0.335 103.310 107.420 104.170 ;
        RECT 0.610 102.490 107.420 103.310 ;
        RECT 0.335 102.470 107.420 102.490 ;
        RECT 0.335 101.650 106.910 102.470 ;
        RECT 0.335 101.630 107.420 101.650 ;
        RECT 0.610 100.810 107.420 101.630 ;
        RECT 0.335 99.950 107.420 100.810 ;
        RECT 0.610 99.130 106.910 99.950 ;
        RECT 0.335 98.270 107.420 99.130 ;
        RECT 0.610 97.450 107.420 98.270 ;
        RECT 0.335 97.430 107.420 97.450 ;
        RECT 0.335 96.610 106.910 97.430 ;
        RECT 0.335 96.590 107.420 96.610 ;
        RECT 0.610 95.770 107.420 96.590 ;
        RECT 0.335 94.910 107.420 95.770 ;
        RECT 0.610 94.090 106.910 94.910 ;
        RECT 0.335 93.230 107.420 94.090 ;
        RECT 0.610 92.410 107.420 93.230 ;
        RECT 0.335 92.390 107.420 92.410 ;
        RECT 0.335 91.570 106.910 92.390 ;
        RECT 0.335 91.550 107.420 91.570 ;
        RECT 0.610 90.730 107.420 91.550 ;
        RECT 0.335 89.870 107.420 90.730 ;
        RECT 0.610 89.050 106.910 89.870 ;
        RECT 0.335 88.190 107.420 89.050 ;
        RECT 0.610 87.370 107.420 88.190 ;
        RECT 0.335 87.350 107.420 87.370 ;
        RECT 0.335 86.530 106.910 87.350 ;
        RECT 0.335 86.510 107.420 86.530 ;
        RECT 0.610 85.690 107.420 86.510 ;
        RECT 0.335 84.830 107.420 85.690 ;
        RECT 0.610 84.010 106.910 84.830 ;
        RECT 0.335 83.150 107.420 84.010 ;
        RECT 0.610 82.330 107.420 83.150 ;
        RECT 0.335 82.310 107.420 82.330 ;
        RECT 0.335 81.490 106.910 82.310 ;
        RECT 0.335 81.470 107.420 81.490 ;
        RECT 0.610 80.650 107.420 81.470 ;
        RECT 0.335 79.790 107.420 80.650 ;
        RECT 0.610 78.970 106.910 79.790 ;
        RECT 0.335 78.110 107.420 78.970 ;
        RECT 0.610 77.290 107.420 78.110 ;
        RECT 0.335 77.270 107.420 77.290 ;
        RECT 0.335 76.450 106.910 77.270 ;
        RECT 0.335 76.430 107.420 76.450 ;
        RECT 0.610 75.610 107.420 76.430 ;
        RECT 0.335 74.750 107.420 75.610 ;
        RECT 0.610 73.930 106.910 74.750 ;
        RECT 0.335 73.070 107.420 73.930 ;
        RECT 0.610 72.250 107.420 73.070 ;
        RECT 0.335 72.230 107.420 72.250 ;
        RECT 0.335 71.410 106.910 72.230 ;
        RECT 0.335 71.390 107.420 71.410 ;
        RECT 0.610 70.570 107.420 71.390 ;
        RECT 0.335 69.710 107.420 70.570 ;
        RECT 0.610 68.890 106.910 69.710 ;
        RECT 0.335 68.030 107.420 68.890 ;
        RECT 0.610 67.210 107.420 68.030 ;
        RECT 0.335 67.190 107.420 67.210 ;
        RECT 0.335 66.370 106.910 67.190 ;
        RECT 0.335 66.350 107.420 66.370 ;
        RECT 0.610 65.530 107.420 66.350 ;
        RECT 0.335 64.670 107.420 65.530 ;
        RECT 0.610 63.850 106.910 64.670 ;
        RECT 0.335 62.990 107.420 63.850 ;
        RECT 0.610 62.170 107.420 62.990 ;
        RECT 0.335 62.150 107.420 62.170 ;
        RECT 0.335 61.330 106.910 62.150 ;
        RECT 0.335 61.310 107.420 61.330 ;
        RECT 0.610 60.490 107.420 61.310 ;
        RECT 0.335 59.630 107.420 60.490 ;
        RECT 0.610 58.810 106.910 59.630 ;
        RECT 0.335 57.950 107.420 58.810 ;
        RECT 0.610 57.130 107.420 57.950 ;
        RECT 0.335 57.110 107.420 57.130 ;
        RECT 0.335 56.290 106.910 57.110 ;
        RECT 0.335 56.270 107.420 56.290 ;
        RECT 0.610 55.450 107.420 56.270 ;
        RECT 0.335 54.590 107.420 55.450 ;
        RECT 0.610 53.770 106.910 54.590 ;
        RECT 0.335 52.910 107.420 53.770 ;
        RECT 0.610 52.090 107.420 52.910 ;
        RECT 0.335 52.070 107.420 52.090 ;
        RECT 0.335 51.250 106.910 52.070 ;
        RECT 0.335 51.230 107.420 51.250 ;
        RECT 0.610 50.410 107.420 51.230 ;
        RECT 0.335 49.550 107.420 50.410 ;
        RECT 0.610 48.730 106.910 49.550 ;
        RECT 0.335 47.870 107.420 48.730 ;
        RECT 0.610 47.050 107.420 47.870 ;
        RECT 0.335 47.030 107.420 47.050 ;
        RECT 0.335 46.210 106.910 47.030 ;
        RECT 0.335 46.190 107.420 46.210 ;
        RECT 0.610 45.370 107.420 46.190 ;
        RECT 0.335 44.510 107.420 45.370 ;
        RECT 0.610 43.690 106.910 44.510 ;
        RECT 0.335 42.830 107.420 43.690 ;
        RECT 0.610 42.010 107.420 42.830 ;
        RECT 0.335 41.990 107.420 42.010 ;
        RECT 0.335 41.170 106.910 41.990 ;
        RECT 0.335 41.150 107.420 41.170 ;
        RECT 0.610 40.330 107.420 41.150 ;
        RECT 0.335 39.470 107.420 40.330 ;
        RECT 0.610 38.650 106.910 39.470 ;
        RECT 0.335 37.790 107.420 38.650 ;
        RECT 0.610 36.970 107.420 37.790 ;
        RECT 0.335 36.950 107.420 36.970 ;
        RECT 0.335 36.130 106.910 36.950 ;
        RECT 0.335 36.110 107.420 36.130 ;
        RECT 0.610 35.290 107.420 36.110 ;
        RECT 0.335 34.430 107.420 35.290 ;
        RECT 0.610 33.610 106.910 34.430 ;
        RECT 0.335 32.750 107.420 33.610 ;
        RECT 0.610 31.930 107.420 32.750 ;
        RECT 0.335 31.910 107.420 31.930 ;
        RECT 0.335 31.090 106.910 31.910 ;
        RECT 0.335 31.070 107.420 31.090 ;
        RECT 0.610 30.250 107.420 31.070 ;
        RECT 0.335 29.390 107.420 30.250 ;
        RECT 0.610 28.570 106.910 29.390 ;
        RECT 0.335 27.710 107.420 28.570 ;
        RECT 0.610 26.890 107.420 27.710 ;
        RECT 0.335 26.870 107.420 26.890 ;
        RECT 0.335 26.050 106.910 26.870 ;
        RECT 0.335 26.030 107.420 26.050 ;
        RECT 0.610 25.210 107.420 26.030 ;
        RECT 0.335 24.350 107.420 25.210 ;
        RECT 0.610 23.530 106.910 24.350 ;
        RECT 0.335 22.670 107.420 23.530 ;
        RECT 0.610 21.850 107.420 22.670 ;
        RECT 0.335 21.830 107.420 21.850 ;
        RECT 0.335 21.010 106.910 21.830 ;
        RECT 0.335 20.990 107.420 21.010 ;
        RECT 0.610 20.170 107.420 20.990 ;
        RECT 0.335 19.310 107.420 20.170 ;
        RECT 0.610 18.490 106.910 19.310 ;
        RECT 0.335 17.630 107.420 18.490 ;
        RECT 0.610 16.810 107.420 17.630 ;
        RECT 0.335 16.790 107.420 16.810 ;
        RECT 0.335 15.970 106.910 16.790 ;
        RECT 0.335 15.950 107.420 15.970 ;
        RECT 0.610 15.130 107.420 15.950 ;
        RECT 0.335 14.270 107.420 15.130 ;
        RECT 0.610 13.450 106.910 14.270 ;
        RECT 0.335 12.590 107.420 13.450 ;
        RECT 0.610 11.770 107.420 12.590 ;
        RECT 0.335 10.910 107.420 11.770 ;
        RECT 0.610 10.090 107.420 10.910 ;
        RECT 0.335 9.230 107.420 10.090 ;
        RECT 0.610 8.410 107.420 9.230 ;
        RECT 0.335 7.550 107.420 8.410 ;
        RECT 0.610 6.730 107.420 7.550 ;
        RECT 0.335 5.870 107.420 6.730 ;
        RECT 0.610 5.050 107.420 5.870 ;
        RECT 0.335 4.190 107.420 5.050 ;
        RECT 0.610 3.370 107.420 4.190 ;
        RECT 0.335 2.510 107.420 3.370 ;
        RECT 0.610 1.690 107.420 2.510 ;
        RECT 0.335 0.830 107.420 1.690 ;
        RECT 0.610 0.315 107.420 0.830 ;
      LAYER Metal4 ;
        RECT 0.375 0.265 107.140 214.345 ;
      LAYER Metal5 ;
        RECT 0.335 0.320 106.705 208.210 ;
      LAYER TopMetal1 ;
        RECT 0.820 0.020 16.620 205.780 ;
        RECT 22.100 0.020 22.820 205.780 ;
        RECT 28.300 0.020 86.820 205.780 ;
  END
END E_TT_IF
END LIBRARY

