magic
tech ihp-sg13g2
magscale 1 2
timestamp 1753877276
<< metal1 >>
rect 1152 9848 41856 9872
rect 1152 9808 4928 9848
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 5296 9808 20048 9848
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20416 9808 35168 9848
rect 35208 9808 35250 9848
rect 35290 9808 35332 9848
rect 35372 9808 35414 9848
rect 35454 9808 35496 9848
rect 35536 9808 41856 9848
rect 1152 9784 41856 9808
rect 6411 9680 6453 9689
rect 6411 9640 6412 9680
rect 6452 9640 6453 9680
rect 6411 9631 6453 9640
rect 7651 9680 7709 9681
rect 7651 9640 7660 9680
rect 7700 9640 7709 9680
rect 7651 9639 7709 9640
rect 8995 9680 9053 9681
rect 8995 9640 9004 9680
rect 9044 9640 9053 9680
rect 8995 9639 9053 9640
rect 9387 9680 9429 9689
rect 9387 9640 9388 9680
rect 9428 9640 9429 9680
rect 9387 9631 9429 9640
rect 9771 9680 9813 9689
rect 9771 9640 9772 9680
rect 9812 9640 9813 9680
rect 9771 9631 9813 9640
rect 10155 9680 10197 9689
rect 10155 9640 10156 9680
rect 10196 9640 10197 9680
rect 10155 9631 10197 9640
rect 12651 9680 12693 9689
rect 12651 9640 12652 9680
rect 12692 9640 12693 9680
rect 12651 9631 12693 9640
rect 13035 9680 13077 9689
rect 13035 9640 13036 9680
rect 13076 9640 13077 9680
rect 13035 9631 13077 9640
rect 14763 9680 14805 9689
rect 14763 9640 14764 9680
rect 14804 9640 14805 9680
rect 14763 9631 14805 9640
rect 18795 9680 18837 9689
rect 18795 9640 18796 9680
rect 18836 9640 18837 9680
rect 18795 9631 18837 9640
rect 25035 9680 25077 9689
rect 25035 9640 25036 9680
rect 25076 9640 25077 9680
rect 25035 9631 25077 9640
rect 27051 9680 27093 9689
rect 27051 9640 27052 9680
rect 27092 9640 27093 9680
rect 27051 9631 27093 9640
rect 3243 9596 3285 9605
rect 3243 9556 3244 9596
rect 3284 9556 3285 9596
rect 3243 9547 3285 9556
rect 22923 9596 22965 9605
rect 22923 9556 22924 9596
rect 22964 9556 22965 9596
rect 22923 9547 22965 9556
rect 1603 9512 1661 9513
rect 1603 9472 1612 9512
rect 1652 9472 1661 9512
rect 1603 9471 1661 9472
rect 2851 9512 2909 9513
rect 2851 9472 2860 9512
rect 2900 9472 2909 9512
rect 2851 9471 2909 9472
rect 3427 9512 3485 9513
rect 3427 9472 3436 9512
rect 3476 9472 3485 9512
rect 3427 9471 3485 9472
rect 4675 9512 4733 9513
rect 4675 9472 4684 9512
rect 4724 9472 4733 9512
rect 4675 9471 4733 9472
rect 4875 9512 4917 9521
rect 4875 9472 4876 9512
rect 4916 9472 4917 9512
rect 4875 9463 4917 9472
rect 4971 9512 5013 9521
rect 4971 9472 4972 9512
rect 5012 9472 5013 9512
rect 4971 9463 5013 9472
rect 5067 9512 5109 9521
rect 5067 9472 5068 9512
rect 5108 9472 5109 9512
rect 5067 9463 5109 9472
rect 5163 9512 5205 9521
rect 5163 9472 5164 9512
rect 5204 9472 5205 9512
rect 5163 9463 5205 9472
rect 6219 9512 6261 9521
rect 6219 9472 6220 9512
rect 6260 9472 6261 9512
rect 6219 9463 6261 9472
rect 6595 9512 6653 9513
rect 6595 9472 6604 9512
rect 6644 9472 6653 9512
rect 6595 9471 6653 9472
rect 6691 9512 6749 9513
rect 6691 9472 6700 9512
rect 6740 9472 6749 9512
rect 6691 9471 6749 9472
rect 6891 9512 6933 9521
rect 6891 9472 6892 9512
rect 6932 9472 6933 9512
rect 6891 9463 6933 9472
rect 6987 9512 7029 9521
rect 6987 9472 6988 9512
rect 7028 9472 7029 9512
rect 6987 9463 7029 9472
rect 7080 9512 7138 9513
rect 7080 9472 7089 9512
rect 7129 9472 7138 9512
rect 7080 9471 7138 9472
rect 7371 9512 7413 9521
rect 7371 9472 7372 9512
rect 7412 9472 7413 9512
rect 7371 9463 7413 9472
rect 7467 9512 7509 9521
rect 7467 9472 7468 9512
rect 7508 9472 7509 9512
rect 7467 9463 7509 9472
rect 8139 9512 8181 9521
rect 8139 9472 8140 9512
rect 8180 9472 8181 9512
rect 8139 9463 8181 9472
rect 8235 9512 8277 9521
rect 8235 9472 8236 9512
rect 8276 9472 8277 9512
rect 8235 9463 8277 9472
rect 8331 9512 8373 9521
rect 8331 9472 8332 9512
rect 8372 9472 8373 9512
rect 8331 9463 8373 9472
rect 8427 9512 8469 9521
rect 8427 9472 8428 9512
rect 8468 9472 8469 9512
rect 8427 9463 8469 9472
rect 8715 9512 8757 9521
rect 8715 9472 8716 9512
rect 8756 9472 8757 9512
rect 8715 9463 8757 9472
rect 8811 9512 8853 9521
rect 8811 9472 8812 9512
rect 8852 9472 8853 9512
rect 8811 9463 8853 9472
rect 15139 9512 15197 9513
rect 15139 9472 15148 9512
rect 15188 9472 15197 9512
rect 15139 9471 15197 9472
rect 16387 9512 16445 9513
rect 16387 9472 16396 9512
rect 16436 9472 16445 9512
rect 16387 9471 16445 9472
rect 16771 9512 16829 9513
rect 16771 9472 16780 9512
rect 16820 9472 16829 9512
rect 16771 9471 16829 9472
rect 18019 9512 18077 9513
rect 18019 9472 18028 9512
rect 18068 9472 18077 9512
rect 18019 9471 18077 9472
rect 19459 9512 19517 9513
rect 19459 9472 19468 9512
rect 19508 9472 19517 9512
rect 19459 9471 19517 9472
rect 20707 9512 20765 9513
rect 20707 9472 20716 9512
rect 20756 9472 20765 9512
rect 20707 9471 20765 9472
rect 21195 9512 21237 9521
rect 21195 9472 21196 9512
rect 21236 9472 21237 9512
rect 21195 9463 21237 9472
rect 21291 9512 21333 9521
rect 21291 9472 21292 9512
rect 21332 9472 21333 9512
rect 21291 9463 21333 9472
rect 21675 9512 21717 9521
rect 21675 9472 21676 9512
rect 21716 9472 21717 9512
rect 21675 9463 21717 9472
rect 22243 9512 22301 9513
rect 22243 9472 22252 9512
rect 22292 9472 22301 9512
rect 23299 9512 23357 9513
rect 22243 9471 22301 9472
rect 22731 9498 22773 9507
rect 22731 9458 22732 9498
rect 22772 9458 22773 9498
rect 23299 9472 23308 9512
rect 23348 9472 23357 9512
rect 23299 9471 23357 9472
rect 24547 9512 24605 9513
rect 24547 9472 24556 9512
rect 24596 9472 24605 9512
rect 24547 9471 24605 9472
rect 25411 9512 25469 9513
rect 25411 9472 25420 9512
rect 25460 9472 25469 9512
rect 25411 9471 25469 9472
rect 26659 9512 26717 9513
rect 26659 9472 26668 9512
rect 26708 9472 26717 9512
rect 26659 9471 26717 9472
rect 29347 9512 29405 9513
rect 29347 9472 29356 9512
rect 29396 9472 29405 9512
rect 29347 9471 29405 9472
rect 30595 9512 30653 9513
rect 30595 9472 30604 9512
rect 30644 9472 30653 9512
rect 30595 9471 30653 9472
rect 31171 9512 31229 9513
rect 31171 9472 31180 9512
rect 31220 9472 31229 9512
rect 31171 9471 31229 9472
rect 32419 9512 32477 9513
rect 32419 9472 32428 9512
rect 32468 9472 32477 9512
rect 32419 9471 32477 9472
rect 32803 9512 32861 9513
rect 32803 9472 32812 9512
rect 32852 9472 32861 9512
rect 32803 9471 32861 9472
rect 34051 9512 34109 9513
rect 34051 9472 34060 9512
rect 34100 9472 34109 9512
rect 34051 9471 34109 9472
rect 34435 9512 34493 9513
rect 34435 9472 34444 9512
rect 34484 9472 34493 9512
rect 34435 9471 34493 9472
rect 35683 9512 35741 9513
rect 35683 9472 35692 9512
rect 35732 9472 35741 9512
rect 35683 9471 35741 9472
rect 36067 9512 36125 9513
rect 36067 9472 36076 9512
rect 36116 9472 36125 9512
rect 36067 9471 36125 9472
rect 37315 9512 37373 9513
rect 37315 9472 37324 9512
rect 37364 9472 37373 9512
rect 37315 9471 37373 9472
rect 37891 9512 37949 9513
rect 37891 9472 37900 9512
rect 37940 9472 37949 9512
rect 37891 9471 37949 9472
rect 39139 9512 39197 9513
rect 39139 9472 39148 9512
rect 39188 9472 39197 9512
rect 39139 9471 39197 9472
rect 39331 9512 39389 9513
rect 39331 9472 39340 9512
rect 39380 9472 39389 9512
rect 39331 9471 39389 9472
rect 40579 9512 40637 9513
rect 40579 9472 40588 9512
rect 40628 9472 40637 9512
rect 40579 9471 40637 9472
rect 22731 9449 22773 9458
rect 9571 9428 9629 9429
rect 9571 9388 9580 9428
rect 9620 9388 9629 9428
rect 9571 9387 9629 9388
rect 9955 9428 10013 9429
rect 9955 9388 9964 9428
rect 10004 9388 10013 9428
rect 9955 9387 10013 9388
rect 10339 9428 10397 9429
rect 10339 9388 10348 9428
rect 10388 9388 10397 9428
rect 10339 9387 10397 9388
rect 12835 9428 12893 9429
rect 12835 9388 12844 9428
rect 12884 9388 12893 9428
rect 12835 9387 12893 9388
rect 13219 9428 13277 9429
rect 13219 9388 13228 9428
rect 13268 9388 13277 9428
rect 13219 9387 13277 9388
rect 14947 9428 15005 9429
rect 14947 9388 14956 9428
rect 14996 9388 15005 9428
rect 14947 9387 15005 9388
rect 18595 9428 18653 9429
rect 18595 9388 18604 9428
rect 18644 9388 18653 9428
rect 18595 9387 18653 9388
rect 21771 9428 21813 9437
rect 21771 9388 21772 9428
rect 21812 9388 21813 9428
rect 21771 9379 21813 9388
rect 25219 9428 25277 9429
rect 25219 9388 25228 9428
rect 25268 9388 25277 9428
rect 25219 9387 25277 9388
rect 27235 9428 27293 9429
rect 27235 9388 27244 9428
rect 27284 9388 27293 9428
rect 27235 9387 27293 9388
rect 40963 9428 41021 9429
rect 40963 9388 40972 9428
rect 41012 9388 41021 9428
rect 40963 9387 41021 9388
rect 6219 9344 6261 9353
rect 6219 9304 6220 9344
rect 6260 9304 6261 9344
rect 6219 9295 6261 9304
rect 26859 9344 26901 9353
rect 26859 9304 26860 9344
rect 26900 9304 26901 9344
rect 26859 9295 26901 9304
rect 41355 9344 41397 9353
rect 41355 9304 41356 9344
rect 41396 9304 41397 9344
rect 41355 9295 41397 9304
rect 3051 9260 3093 9269
rect 3051 9220 3052 9260
rect 3092 9220 3093 9260
rect 3051 9211 3093 9220
rect 6603 9260 6645 9269
rect 6603 9220 6604 9260
rect 6644 9220 6645 9260
rect 6603 9211 6645 9220
rect 16587 9260 16629 9269
rect 16587 9220 16588 9260
rect 16628 9220 16629 9260
rect 16587 9211 16629 9220
rect 18219 9260 18261 9269
rect 18219 9220 18220 9260
rect 18260 9220 18261 9260
rect 18219 9211 18261 9220
rect 20907 9260 20949 9269
rect 20907 9220 20908 9260
rect 20948 9220 20949 9260
rect 20907 9211 20949 9220
rect 23115 9260 23157 9269
rect 23115 9220 23116 9260
rect 23156 9220 23157 9260
rect 23115 9211 23157 9220
rect 30795 9260 30837 9269
rect 30795 9220 30796 9260
rect 30836 9220 30837 9260
rect 30795 9211 30837 9220
rect 30987 9260 31029 9269
rect 30987 9220 30988 9260
rect 31028 9220 31029 9260
rect 30987 9211 31029 9220
rect 32619 9260 32661 9269
rect 32619 9220 32620 9260
rect 32660 9220 32661 9260
rect 32619 9211 32661 9220
rect 34251 9260 34293 9269
rect 34251 9220 34252 9260
rect 34292 9220 34293 9260
rect 34251 9211 34293 9220
rect 37515 9260 37557 9269
rect 37515 9220 37516 9260
rect 37556 9220 37557 9260
rect 37515 9211 37557 9220
rect 37707 9260 37749 9269
rect 37707 9220 37708 9260
rect 37748 9220 37749 9260
rect 37707 9211 37749 9220
rect 40779 9260 40821 9269
rect 40779 9220 40780 9260
rect 40820 9220 40821 9260
rect 40779 9211 40821 9220
rect 41163 9260 41205 9269
rect 41163 9220 41164 9260
rect 41204 9220 41205 9260
rect 41163 9211 41205 9220
rect 1152 9092 41856 9116
rect 1152 9052 3688 9092
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 4056 9052 18808 9092
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 19176 9052 33928 9092
rect 33968 9052 34010 9092
rect 34050 9052 34092 9092
rect 34132 9052 34174 9092
rect 34214 9052 34256 9092
rect 34296 9052 41856 9092
rect 1152 9028 41856 9052
rect 9475 8924 9533 8925
rect 9475 8884 9484 8924
rect 9524 8884 9533 8924
rect 9475 8883 9533 8884
rect 9867 8840 9909 8849
rect 9867 8800 9868 8840
rect 9908 8800 9909 8840
rect 9867 8791 9909 8800
rect 10635 8840 10677 8849
rect 10635 8800 10636 8840
rect 10676 8800 10677 8840
rect 10635 8791 10677 8800
rect 10827 8840 10869 8849
rect 10827 8800 10828 8840
rect 10868 8800 10869 8840
rect 10827 8791 10869 8800
rect 11211 8840 11253 8849
rect 11211 8800 11212 8840
rect 11252 8800 11253 8840
rect 11211 8791 11253 8800
rect 11787 8840 11829 8849
rect 11787 8800 11788 8840
rect 11828 8800 11829 8840
rect 11787 8791 11829 8800
rect 12171 8840 12213 8849
rect 12171 8800 12172 8840
rect 12212 8800 12213 8840
rect 12171 8791 12213 8800
rect 30027 8840 30069 8849
rect 30027 8800 30028 8840
rect 30068 8800 30069 8840
rect 30027 8791 30069 8800
rect 9667 8756 9725 8757
rect 9667 8716 9676 8756
rect 9716 8716 9725 8756
rect 9667 8715 9725 8716
rect 10051 8756 10109 8757
rect 10051 8716 10060 8756
rect 10100 8716 10109 8756
rect 10051 8715 10109 8716
rect 10435 8756 10493 8757
rect 10435 8716 10444 8756
rect 10484 8716 10493 8756
rect 10435 8715 10493 8716
rect 11011 8756 11069 8757
rect 11011 8716 11020 8756
rect 11060 8716 11069 8756
rect 11011 8715 11069 8716
rect 11395 8756 11453 8757
rect 11395 8716 11404 8756
rect 11444 8716 11453 8756
rect 11395 8715 11453 8716
rect 11587 8756 11645 8757
rect 11587 8716 11596 8756
rect 11636 8716 11645 8756
rect 11587 8715 11645 8716
rect 11971 8756 12029 8757
rect 11971 8716 11980 8756
rect 12020 8716 12029 8756
rect 11971 8715 12029 8716
rect 15243 8756 15285 8765
rect 15243 8716 15244 8756
rect 15284 8716 15285 8756
rect 15243 8707 15285 8716
rect 18891 8756 18933 8765
rect 18891 8716 18892 8756
rect 18932 8716 18933 8756
rect 18891 8707 18933 8716
rect 24363 8756 24405 8765
rect 24363 8716 24364 8756
rect 24404 8716 24405 8756
rect 24363 8707 24405 8716
rect 26475 8756 26517 8765
rect 26475 8716 26476 8756
rect 26516 8716 26517 8756
rect 26475 8707 26517 8716
rect 29443 8756 29501 8757
rect 29443 8716 29452 8756
rect 29492 8716 29501 8756
rect 29443 8715 29501 8716
rect 29827 8756 29885 8757
rect 29827 8716 29836 8756
rect 29876 8716 29885 8756
rect 29827 8715 29885 8716
rect 31467 8756 31509 8765
rect 31467 8716 31468 8756
rect 31508 8716 31509 8756
rect 31467 8707 31509 8716
rect 32515 8756 32573 8757
rect 32515 8716 32524 8756
rect 32564 8716 32573 8756
rect 32515 8715 32573 8716
rect 32899 8756 32957 8757
rect 32899 8716 32908 8756
rect 32948 8716 32957 8756
rect 32899 8715 32957 8716
rect 35395 8756 35453 8757
rect 35395 8716 35404 8756
rect 35444 8716 35453 8756
rect 35395 8715 35453 8716
rect 41347 8756 41405 8757
rect 41347 8716 41356 8756
rect 41396 8716 41405 8756
rect 41347 8715 41405 8716
rect 1899 8672 1941 8681
rect 1899 8632 1900 8672
rect 1940 8632 1941 8672
rect 1899 8623 1941 8632
rect 1995 8672 2037 8681
rect 1995 8632 1996 8672
rect 2036 8632 2037 8672
rect 1995 8623 2037 8632
rect 2091 8672 2133 8681
rect 2091 8632 2092 8672
rect 2132 8632 2133 8672
rect 2091 8623 2133 8632
rect 2475 8672 2517 8681
rect 2475 8632 2476 8672
rect 2516 8632 2517 8672
rect 2475 8623 2517 8632
rect 2571 8672 2613 8681
rect 2571 8632 2572 8672
rect 2612 8632 2613 8672
rect 2571 8623 2613 8632
rect 2859 8672 2901 8681
rect 2859 8632 2860 8672
rect 2900 8632 2901 8672
rect 2859 8623 2901 8632
rect 2955 8672 2997 8681
rect 2955 8632 2956 8672
rect 2996 8632 2997 8672
rect 2955 8623 2997 8632
rect 3339 8672 3381 8681
rect 3339 8632 3340 8672
rect 3380 8632 3381 8672
rect 3339 8623 3381 8632
rect 3435 8672 3477 8681
rect 4395 8677 4437 8686
rect 3435 8632 3436 8672
rect 3476 8632 3477 8672
rect 3435 8623 3477 8632
rect 3907 8672 3965 8673
rect 3907 8632 3916 8672
rect 3956 8632 3965 8672
rect 3907 8631 3965 8632
rect 4395 8637 4396 8677
rect 4436 8637 4437 8677
rect 4395 8628 4437 8637
rect 4771 8672 4829 8673
rect 4771 8632 4780 8672
rect 4820 8632 4829 8672
rect 4771 8631 4829 8632
rect 6019 8672 6077 8673
rect 6019 8632 6028 8672
rect 6068 8632 6077 8672
rect 6019 8631 6077 8632
rect 6795 8672 6837 8681
rect 6795 8632 6796 8672
rect 6836 8632 6837 8672
rect 6795 8623 6837 8632
rect 6891 8672 6933 8681
rect 6891 8632 6892 8672
rect 6932 8632 6933 8672
rect 6891 8623 6933 8632
rect 7275 8672 7317 8681
rect 7275 8632 7276 8672
rect 7316 8632 7317 8672
rect 7275 8623 7317 8632
rect 7371 8672 7413 8681
rect 8331 8677 8373 8686
rect 14139 8681 14181 8690
rect 17931 8686 17973 8695
rect 23307 8686 23349 8695
rect 7371 8632 7372 8672
rect 7412 8632 7413 8672
rect 7371 8623 7413 8632
rect 7843 8672 7901 8673
rect 7843 8632 7852 8672
rect 7892 8632 7901 8672
rect 7843 8631 7901 8632
rect 8331 8637 8332 8677
rect 8372 8637 8373 8677
rect 8331 8628 8373 8637
rect 8803 8672 8861 8673
rect 8803 8632 8812 8672
rect 8852 8632 8861 8672
rect 8803 8631 8861 8632
rect 9099 8672 9141 8681
rect 9099 8632 9100 8672
rect 9140 8632 9141 8672
rect 9099 8623 9141 8632
rect 12355 8672 12413 8673
rect 12355 8632 12364 8672
rect 12404 8632 12413 8672
rect 12355 8631 12413 8632
rect 13603 8672 13661 8673
rect 13603 8632 13612 8672
rect 13652 8632 13661 8672
rect 14139 8641 14140 8681
rect 14180 8641 14181 8681
rect 14139 8632 14181 8641
rect 14659 8672 14717 8673
rect 14659 8632 14668 8672
rect 14708 8632 14717 8672
rect 13603 8631 13661 8632
rect 14659 8631 14717 8632
rect 15147 8672 15189 8681
rect 15147 8632 15148 8672
rect 15188 8632 15189 8672
rect 15147 8623 15189 8632
rect 15627 8672 15669 8681
rect 15627 8632 15628 8672
rect 15668 8632 15669 8672
rect 15627 8623 15669 8632
rect 15723 8672 15765 8681
rect 15723 8632 15724 8672
rect 15764 8632 15765 8672
rect 15723 8623 15765 8632
rect 16395 8672 16437 8681
rect 16395 8632 16396 8672
rect 16436 8632 16437 8672
rect 16395 8623 16437 8632
rect 16491 8672 16533 8681
rect 16491 8632 16492 8672
rect 16532 8632 16533 8672
rect 16491 8623 16533 8632
rect 16875 8672 16917 8681
rect 16875 8632 16876 8672
rect 16916 8632 16917 8672
rect 16875 8623 16917 8632
rect 16971 8672 17013 8681
rect 16971 8632 16972 8672
rect 17012 8632 17013 8672
rect 16971 8623 17013 8632
rect 17443 8672 17501 8673
rect 17443 8632 17452 8672
rect 17492 8632 17501 8672
rect 17931 8646 17932 8686
rect 17972 8646 17973 8686
rect 17931 8637 17973 8646
rect 18411 8672 18453 8681
rect 17443 8631 17501 8632
rect 18411 8632 18412 8672
rect 18452 8632 18453 8672
rect 18411 8623 18453 8632
rect 18507 8672 18549 8681
rect 18507 8632 18508 8672
rect 18548 8632 18549 8672
rect 18507 8623 18549 8632
rect 18987 8672 19029 8681
rect 19947 8677 19989 8686
rect 18987 8632 18988 8672
rect 19028 8632 19029 8672
rect 18987 8623 19029 8632
rect 19459 8672 19517 8673
rect 19459 8632 19468 8672
rect 19508 8632 19517 8672
rect 19459 8631 19517 8632
rect 19947 8637 19948 8677
rect 19988 8637 19989 8677
rect 19947 8628 19989 8637
rect 21771 8672 21813 8681
rect 21771 8632 21772 8672
rect 21812 8632 21813 8672
rect 21771 8623 21813 8632
rect 21867 8672 21909 8681
rect 21867 8632 21868 8672
rect 21908 8632 21909 8672
rect 21867 8623 21909 8632
rect 22251 8672 22293 8681
rect 22251 8632 22252 8672
rect 22292 8632 22293 8672
rect 22251 8623 22293 8632
rect 22347 8672 22389 8681
rect 22347 8632 22348 8672
rect 22388 8632 22389 8672
rect 22347 8623 22389 8632
rect 22819 8672 22877 8673
rect 22819 8632 22828 8672
rect 22868 8632 22877 8672
rect 23307 8646 23308 8686
rect 23348 8646 23349 8686
rect 25467 8681 25509 8690
rect 27483 8681 27525 8690
rect 23307 8637 23349 8646
rect 23883 8672 23925 8681
rect 22819 8631 22877 8632
rect 23883 8632 23884 8672
rect 23924 8632 23925 8672
rect 23883 8623 23925 8632
rect 23979 8672 24021 8681
rect 23979 8632 23980 8672
rect 24020 8632 24021 8672
rect 23979 8623 24021 8632
rect 24459 8672 24501 8681
rect 24459 8632 24460 8672
rect 24500 8632 24501 8672
rect 24459 8623 24501 8632
rect 24931 8672 24989 8673
rect 24931 8632 24940 8672
rect 24980 8632 24989 8672
rect 25467 8641 25468 8681
rect 25508 8641 25509 8681
rect 25467 8632 25509 8641
rect 25899 8672 25941 8681
rect 25899 8632 25900 8672
rect 25940 8632 25941 8672
rect 24931 8631 24989 8632
rect 25899 8623 25941 8632
rect 25995 8672 26037 8681
rect 25995 8632 25996 8672
rect 26036 8632 26037 8672
rect 25995 8623 26037 8632
rect 26379 8672 26421 8681
rect 26379 8632 26380 8672
rect 26420 8632 26421 8672
rect 26379 8623 26421 8632
rect 26947 8672 27005 8673
rect 26947 8632 26956 8672
rect 26996 8632 27005 8672
rect 27483 8641 27484 8681
rect 27524 8641 27525 8681
rect 30507 8686 30549 8695
rect 27483 8632 27525 8641
rect 28003 8672 28061 8673
rect 28003 8632 28012 8672
rect 28052 8632 28061 8672
rect 26947 8631 27005 8632
rect 28003 8631 28061 8632
rect 29251 8672 29309 8673
rect 29251 8632 29260 8672
rect 29300 8632 29309 8672
rect 30507 8646 30508 8686
rect 30548 8646 30549 8686
rect 34827 8686 34869 8695
rect 30507 8637 30549 8646
rect 30979 8672 31037 8673
rect 29251 8631 29309 8632
rect 30979 8632 30988 8672
rect 31028 8632 31037 8672
rect 30979 8631 31037 8632
rect 31563 8672 31605 8681
rect 31563 8632 31564 8672
rect 31604 8632 31605 8672
rect 32043 8672 32085 8681
rect 31563 8623 31605 8632
rect 31947 8652 31989 8661
rect 31947 8612 31948 8652
rect 31988 8612 31989 8652
rect 32043 8632 32044 8672
rect 32084 8632 32085 8672
rect 32043 8623 32085 8632
rect 33291 8672 33333 8681
rect 33291 8632 33292 8672
rect 33332 8632 33333 8672
rect 33291 8623 33333 8632
rect 33387 8672 33429 8681
rect 33387 8632 33388 8672
rect 33428 8632 33429 8672
rect 33387 8623 33429 8632
rect 33771 8672 33813 8681
rect 33771 8632 33772 8672
rect 33812 8632 33813 8672
rect 33771 8623 33813 8632
rect 33867 8672 33909 8681
rect 33867 8632 33868 8672
rect 33908 8632 33909 8672
rect 33867 8623 33909 8632
rect 34339 8672 34397 8673
rect 34339 8632 34348 8672
rect 34388 8632 34397 8672
rect 34827 8646 34828 8686
rect 34868 8646 34869 8686
rect 37371 8681 37413 8690
rect 39339 8686 39381 8695
rect 34827 8637 34869 8646
rect 35787 8672 35829 8681
rect 34339 8631 34397 8632
rect 35787 8632 35788 8672
rect 35828 8632 35829 8672
rect 35787 8623 35829 8632
rect 35883 8672 35925 8681
rect 35883 8632 35884 8672
rect 35924 8632 35925 8672
rect 35883 8623 35925 8632
rect 36267 8672 36309 8681
rect 36267 8632 36268 8672
rect 36308 8632 36309 8672
rect 36267 8623 36309 8632
rect 36363 8672 36405 8681
rect 36363 8632 36364 8672
rect 36404 8632 36405 8672
rect 36363 8623 36405 8632
rect 36835 8672 36893 8673
rect 36835 8632 36844 8672
rect 36884 8632 36893 8672
rect 37371 8641 37372 8681
rect 37412 8641 37413 8681
rect 37371 8632 37413 8641
rect 37803 8672 37845 8681
rect 37803 8632 37804 8672
rect 37844 8632 37845 8672
rect 36835 8631 36893 8632
rect 37803 8623 37845 8632
rect 37899 8672 37941 8681
rect 37899 8632 37900 8672
rect 37940 8632 37941 8672
rect 37899 8623 37941 8632
rect 38283 8672 38325 8681
rect 38283 8632 38284 8672
rect 38324 8632 38325 8672
rect 38283 8623 38325 8632
rect 38379 8672 38421 8681
rect 38379 8632 38380 8672
rect 38420 8632 38421 8672
rect 38379 8623 38421 8632
rect 38851 8672 38909 8673
rect 38851 8632 38860 8672
rect 38900 8632 38909 8672
rect 39339 8646 39340 8686
rect 39380 8646 39381 8686
rect 39339 8637 39381 8646
rect 39907 8672 39965 8673
rect 38851 8631 38909 8632
rect 39907 8632 39916 8672
rect 39956 8632 39965 8672
rect 39907 8631 39965 8632
rect 41155 8672 41213 8673
rect 41155 8632 41164 8672
rect 41204 8632 41213 8672
rect 41155 8631 41213 8632
rect 31947 8603 31989 8612
rect 8523 8588 8565 8597
rect 8523 8548 8524 8588
rect 8564 8548 8565 8588
rect 8523 8539 8565 8548
rect 9195 8588 9237 8597
rect 9195 8548 9196 8588
rect 9236 8548 9237 8588
rect 9195 8539 9237 8548
rect 18123 8588 18165 8597
rect 18123 8548 18124 8588
rect 18164 8548 18165 8588
rect 18123 8539 18165 8548
rect 20139 8588 20181 8597
rect 20139 8548 20140 8588
rect 20180 8548 20181 8588
rect 20139 8539 20181 8548
rect 25611 8588 25653 8597
rect 25611 8548 25612 8588
rect 25652 8548 25653 8588
rect 25611 8539 25653 8548
rect 27627 8588 27669 8597
rect 27627 8548 27628 8588
rect 27668 8548 27669 8588
rect 27627 8539 27669 8548
rect 30315 8588 30357 8597
rect 30315 8548 30316 8588
rect 30356 8548 30357 8588
rect 30315 8539 30357 8548
rect 1795 8504 1853 8505
rect 1795 8464 1804 8504
rect 1844 8464 1853 8504
rect 1795 8463 1853 8464
rect 2275 8504 2333 8505
rect 2275 8464 2284 8504
rect 2324 8464 2333 8504
rect 2275 8463 2333 8464
rect 4587 8504 4629 8513
rect 4587 8464 4588 8504
rect 4628 8464 4629 8504
rect 4587 8455 4629 8464
rect 6219 8504 6261 8513
rect 6219 8464 6220 8504
rect 6260 8464 6261 8504
rect 6219 8455 6261 8464
rect 10251 8504 10293 8513
rect 10251 8464 10252 8504
rect 10292 8464 10293 8504
rect 10251 8455 10293 8464
rect 13803 8504 13845 8513
rect 13803 8464 13804 8504
rect 13844 8464 13845 8504
rect 13803 8455 13845 8464
rect 13995 8504 14037 8513
rect 13995 8464 13996 8504
rect 14036 8464 14037 8504
rect 13995 8455 14037 8464
rect 20323 8504 20381 8505
rect 20323 8464 20332 8504
rect 20372 8464 20381 8504
rect 20323 8463 20381 8464
rect 23499 8504 23541 8513
rect 23499 8464 23500 8504
rect 23540 8464 23541 8504
rect 23499 8455 23541 8464
rect 27819 8504 27861 8513
rect 27819 8464 27820 8504
rect 27860 8464 27861 8504
rect 27819 8455 27861 8464
rect 29643 8504 29685 8513
rect 29643 8464 29644 8504
rect 29684 8464 29685 8504
rect 29643 8455 29685 8464
rect 32331 8504 32373 8513
rect 32331 8464 32332 8504
rect 32372 8464 32373 8504
rect 32331 8455 32373 8464
rect 32715 8504 32757 8513
rect 32715 8464 32716 8504
rect 32756 8464 32757 8504
rect 32715 8455 32757 8464
rect 35019 8504 35061 8513
rect 35019 8464 35020 8504
rect 35060 8464 35061 8504
rect 35019 8455 35061 8464
rect 35211 8504 35253 8513
rect 35211 8464 35212 8504
rect 35252 8464 35253 8504
rect 35211 8455 35253 8464
rect 37515 8504 37557 8513
rect 37515 8464 37516 8504
rect 37556 8464 37557 8504
rect 37515 8455 37557 8464
rect 39531 8504 39573 8513
rect 39531 8464 39532 8504
rect 39572 8464 39573 8504
rect 39531 8455 39573 8464
rect 39723 8504 39765 8513
rect 39723 8464 39724 8504
rect 39764 8464 39765 8504
rect 39723 8455 39765 8464
rect 41547 8504 41589 8513
rect 41547 8464 41548 8504
rect 41588 8464 41589 8504
rect 41547 8455 41589 8464
rect 1152 8336 41856 8360
rect 1152 8296 4928 8336
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 5296 8296 20048 8336
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20416 8296 35168 8336
rect 35208 8296 35250 8336
rect 35290 8296 35332 8336
rect 35372 8296 35414 8336
rect 35454 8296 35496 8336
rect 35536 8296 41856 8336
rect 1152 8272 41856 8296
rect 4099 8210 4157 8211
rect 3339 8168 3381 8177
rect 4099 8170 4108 8210
rect 4148 8170 4157 8210
rect 4099 8169 4157 8170
rect 3339 8128 3340 8168
rect 3380 8128 3381 8168
rect 3339 8119 3381 8128
rect 8427 8168 8469 8177
rect 8427 8128 8428 8168
rect 8468 8128 8469 8168
rect 8427 8119 8469 8128
rect 11115 8168 11157 8177
rect 11115 8128 11116 8168
rect 11156 8128 11157 8168
rect 11115 8119 11157 8128
rect 13995 8168 14037 8177
rect 13995 8128 13996 8168
rect 14036 8128 14037 8168
rect 13995 8119 14037 8128
rect 17739 8168 17781 8177
rect 17739 8128 17740 8168
rect 17780 8128 17781 8168
rect 17739 8119 17781 8128
rect 19371 8168 19413 8177
rect 19371 8128 19372 8168
rect 19412 8128 19413 8168
rect 19371 8119 19413 8128
rect 21003 8168 21045 8177
rect 21003 8128 21004 8168
rect 21044 8128 21045 8168
rect 21003 8119 21045 8128
rect 23211 8168 23253 8177
rect 23211 8128 23212 8168
rect 23252 8128 23253 8168
rect 23211 8119 23253 8128
rect 25515 8168 25557 8177
rect 25515 8128 25516 8168
rect 25556 8128 25557 8168
rect 25515 8119 25557 8128
rect 25707 8168 25749 8177
rect 25707 8128 25708 8168
rect 25748 8128 25749 8168
rect 25707 8119 25749 8128
rect 26283 8168 26325 8177
rect 26283 8128 26284 8168
rect 26324 8128 26325 8168
rect 26283 8119 26325 8128
rect 30411 8168 30453 8177
rect 30411 8128 30412 8168
rect 30452 8128 30453 8168
rect 30411 8119 30453 8128
rect 30795 8168 30837 8177
rect 30795 8128 30796 8168
rect 30836 8128 30837 8168
rect 30795 8119 30837 8128
rect 33195 8168 33237 8177
rect 33195 8128 33196 8168
rect 33236 8128 33237 8168
rect 33195 8119 33237 8128
rect 35691 8168 35733 8177
rect 35691 8128 35692 8168
rect 35732 8128 35733 8168
rect 35691 8119 35733 8128
rect 37899 8168 37941 8177
rect 37899 8128 37900 8168
rect 37940 8128 37941 8168
rect 37899 8119 37941 8128
rect 40683 8168 40725 8177
rect 40683 8128 40684 8168
rect 40724 8128 40725 8168
rect 40683 8119 40725 8128
rect 10923 8084 10965 8093
rect 10923 8044 10924 8084
rect 10964 8044 10965 8084
rect 10923 8035 10965 8044
rect 23019 8084 23061 8093
rect 23019 8044 23020 8084
rect 23060 8044 23061 8084
rect 23019 8035 23061 8044
rect 28587 8084 28629 8093
rect 28587 8044 28588 8084
rect 28628 8044 28629 8084
rect 28587 8035 28629 8044
rect 1891 8000 1949 8001
rect 1891 7960 1900 8000
rect 1940 7960 1949 8000
rect 1891 7959 1949 7960
rect 3139 8000 3197 8001
rect 3139 7960 3148 8000
rect 3188 7960 3197 8000
rect 3139 7959 3197 7960
rect 3819 8000 3861 8009
rect 3819 7960 3820 8000
rect 3860 7960 3861 8000
rect 3819 7951 3861 7960
rect 3915 8001 3957 8010
rect 32515 8009 32573 8010
rect 3915 7961 3916 8001
rect 3956 7961 3957 8001
rect 3915 7952 3957 7961
rect 4299 8000 4341 8009
rect 4299 7960 4300 8000
rect 4340 7960 4341 8000
rect 4299 7951 4341 7960
rect 4395 8000 4437 8009
rect 4395 7960 4396 8000
rect 4436 7960 4437 8000
rect 4395 7951 4437 7960
rect 4491 8000 4533 8009
rect 4491 7960 4492 8000
rect 4532 7960 4533 8000
rect 4491 7951 4533 7960
rect 4587 8000 4629 8009
rect 4587 7960 4588 8000
rect 4628 7960 4629 8000
rect 4587 7951 4629 7960
rect 4771 8000 4829 8001
rect 4771 7960 4780 8000
rect 4820 7960 4829 8000
rect 4771 7959 4829 7960
rect 6019 8000 6077 8001
rect 6019 7960 6028 8000
rect 6068 7960 6077 8000
rect 6019 7959 6077 7960
rect 6699 8000 6741 8009
rect 6699 7960 6700 8000
rect 6740 7960 6741 8000
rect 6699 7951 6741 7960
rect 6795 8000 6837 8009
rect 6795 7960 6796 8000
rect 6836 7960 6837 8000
rect 6795 7951 6837 7960
rect 7747 8000 7805 8001
rect 7747 7960 7756 8000
rect 7796 7960 7805 8000
rect 8619 8000 8661 8009
rect 7747 7959 7805 7960
rect 8235 7986 8277 7995
rect 8235 7946 8236 7986
rect 8276 7946 8277 7986
rect 8619 7960 8620 8000
rect 8660 7960 8661 8000
rect 8619 7951 8661 7960
rect 8715 8000 8757 8009
rect 8715 7960 8716 8000
rect 8756 7960 8757 8000
rect 8715 7951 8757 7960
rect 8811 8000 8853 8009
rect 8811 7960 8812 8000
rect 8852 7960 8853 8000
rect 8811 7951 8853 7960
rect 8907 8000 8949 8009
rect 8907 7960 8908 8000
rect 8948 7960 8949 8000
rect 8907 7951 8949 7960
rect 9099 8000 9141 8009
rect 9099 7960 9100 8000
rect 9140 7960 9141 8000
rect 9099 7951 9141 7960
rect 9283 8000 9341 8001
rect 9283 7960 9292 8000
rect 9332 7960 9341 8000
rect 9283 7959 9341 7960
rect 9475 8000 9533 8001
rect 9475 7960 9484 8000
rect 9524 7960 9533 8000
rect 9475 7959 9533 7960
rect 10723 8000 10781 8001
rect 10723 7960 10732 8000
rect 10772 7960 10781 8000
rect 11779 8000 11837 8001
rect 10723 7959 10781 7960
rect 11259 7990 11301 7999
rect 8235 7937 8277 7946
rect 11259 7950 11260 7990
rect 11300 7950 11301 7990
rect 11779 7960 11788 8000
rect 11828 7960 11837 8000
rect 11779 7959 11837 7960
rect 12267 8000 12309 8009
rect 12267 7960 12268 8000
rect 12308 7960 12309 8000
rect 12267 7951 12309 7960
rect 12747 8000 12789 8009
rect 12747 7960 12748 8000
rect 12788 7960 12789 8000
rect 12747 7951 12789 7960
rect 12843 8000 12885 8009
rect 12843 7960 12844 8000
rect 12884 7960 12885 8000
rect 12843 7951 12885 7960
rect 14179 8000 14237 8001
rect 14179 7960 14188 8000
rect 14228 7960 14237 8000
rect 14179 7959 14237 7960
rect 15427 8000 15485 8001
rect 15427 7960 15436 8000
rect 15476 7960 15485 8000
rect 15427 7959 15485 7960
rect 16291 8000 16349 8001
rect 16291 7960 16300 8000
rect 16340 7960 16349 8000
rect 16291 7959 16349 7960
rect 17539 8000 17597 8001
rect 17539 7960 17548 8000
rect 17588 7960 17597 8000
rect 17539 7959 17597 7960
rect 17923 8000 17981 8001
rect 17923 7960 17932 8000
rect 17972 7960 17981 8000
rect 17923 7959 17981 7960
rect 19171 8000 19229 8001
rect 19171 7960 19180 8000
rect 19220 7960 19229 8000
rect 19171 7959 19229 7960
rect 19555 8000 19613 8001
rect 19555 7960 19564 8000
rect 19604 7960 19613 8000
rect 19555 7959 19613 7960
rect 20803 8000 20861 8001
rect 20803 7960 20812 8000
rect 20852 7960 20861 8000
rect 20803 7959 20861 7960
rect 21291 8000 21333 8009
rect 21291 7960 21292 8000
rect 21332 7960 21333 8000
rect 21291 7951 21333 7960
rect 21387 8000 21429 8009
rect 21387 7960 21388 8000
rect 21428 7960 21429 8000
rect 21387 7951 21429 7960
rect 21771 8000 21813 8009
rect 21771 7960 21772 8000
rect 21812 7960 21813 8000
rect 21771 7951 21813 7960
rect 21867 8000 21909 8009
rect 21867 7960 21868 8000
rect 21908 7960 21909 8000
rect 21867 7951 21909 7960
rect 22339 8000 22397 8001
rect 22339 7960 22348 8000
rect 22388 7960 22397 8000
rect 24067 8000 24125 8001
rect 22339 7959 22397 7960
rect 22827 7986 22869 7995
rect 11259 7941 11301 7950
rect 22827 7946 22828 7986
rect 22868 7946 22869 7986
rect 24067 7960 24076 8000
rect 24116 7960 24125 8000
rect 24067 7959 24125 7960
rect 25315 8000 25373 8001
rect 25315 7960 25324 8000
rect 25364 7960 25373 8000
rect 25315 7959 25373 7960
rect 26859 8000 26901 8009
rect 26859 7960 26860 8000
rect 26900 7960 26901 8000
rect 26859 7951 26901 7960
rect 26955 8000 26997 8009
rect 26955 7960 26956 8000
rect 26996 7960 26997 8000
rect 26955 7951 26997 7960
rect 27435 8000 27477 8009
rect 27435 7960 27436 8000
rect 27476 7960 27477 8000
rect 27435 7951 27477 7960
rect 27907 8000 27965 8001
rect 27907 7960 27916 8000
rect 27956 7960 27965 8000
rect 27907 7959 27965 7960
rect 28395 7995 28437 8004
rect 28395 7955 28396 7995
rect 28436 7955 28437 7995
rect 28771 8000 28829 8001
rect 28771 7960 28780 8000
rect 28820 7960 28829 8000
rect 28771 7959 28829 7960
rect 30019 8000 30077 8001
rect 30019 7960 30028 8000
rect 30068 7960 30077 8000
rect 30019 7959 30077 7960
rect 31467 8000 31509 8009
rect 31467 7960 31468 8000
rect 31508 7960 31509 8000
rect 28395 7946 28437 7955
rect 31467 7951 31509 7960
rect 31563 8000 31605 8009
rect 31563 7960 31564 8000
rect 31604 7960 31605 8000
rect 31563 7951 31605 7960
rect 31947 8000 31989 8009
rect 31947 7960 31948 8000
rect 31988 7960 31989 8000
rect 31947 7951 31989 7960
rect 32043 8000 32085 8009
rect 32043 7960 32044 8000
rect 32084 7960 32085 8000
rect 32515 7969 32524 8009
rect 32564 7969 32573 8009
rect 34051 8000 34109 8001
rect 32515 7968 32573 7969
rect 33051 7990 33093 7999
rect 32043 7951 32085 7960
rect 33051 7950 33052 7990
rect 33092 7950 33093 7990
rect 34051 7960 34060 8000
rect 34100 7960 34109 8000
rect 34051 7959 34109 7960
rect 35299 8000 35357 8001
rect 35299 7960 35308 8000
rect 35348 7960 35357 8000
rect 35299 7959 35357 7960
rect 35875 8000 35933 8001
rect 35875 7960 35884 8000
rect 35924 7960 35933 8000
rect 35875 7959 35933 7960
rect 37123 8000 37181 8001
rect 37123 7960 37132 8000
rect 37172 7960 37181 8000
rect 37123 7959 37181 7960
rect 38955 8000 38997 8009
rect 38955 7960 38956 8000
rect 38996 7960 38997 8000
rect 38955 7951 38997 7960
rect 39051 8000 39093 8009
rect 39051 7960 39052 8000
rect 39092 7960 39093 8000
rect 39051 7951 39093 7960
rect 39435 8000 39477 8009
rect 39435 7960 39436 8000
rect 39476 7960 39477 8000
rect 39435 7951 39477 7960
rect 39531 8000 39573 8009
rect 39531 7960 39532 8000
rect 39572 7960 39573 8000
rect 39531 7951 39573 7960
rect 40003 8000 40061 8001
rect 40003 7960 40012 8000
rect 40052 7960 40061 8000
rect 40003 7959 40061 7960
rect 40491 7986 40533 7995
rect 22827 7937 22869 7946
rect 33051 7941 33093 7950
rect 40491 7946 40492 7986
rect 40532 7946 40533 7986
rect 40491 7937 40533 7946
rect 7179 7916 7221 7925
rect 7179 7876 7180 7916
rect 7220 7876 7221 7916
rect 7179 7867 7221 7876
rect 7275 7916 7317 7925
rect 7275 7876 7276 7916
rect 7316 7876 7317 7916
rect 7275 7867 7317 7876
rect 12363 7916 12405 7925
rect 12363 7876 12364 7916
rect 12404 7876 12405 7916
rect 12363 7867 12405 7876
rect 23395 7916 23453 7917
rect 23395 7876 23404 7916
rect 23444 7876 23453 7916
rect 23395 7875 23453 7876
rect 25891 7916 25949 7917
rect 25891 7876 25900 7916
rect 25940 7876 25949 7916
rect 27339 7916 27381 7925
rect 25891 7875 25949 7876
rect 26083 7905 26141 7906
rect 26083 7865 26092 7905
rect 26132 7865 26141 7905
rect 27339 7876 27340 7916
rect 27380 7876 27381 7916
rect 27339 7867 27381 7876
rect 30595 7916 30653 7917
rect 30595 7876 30604 7916
rect 30644 7876 30653 7916
rect 30595 7875 30653 7876
rect 30979 7916 31037 7917
rect 30979 7876 30988 7916
rect 31028 7876 31037 7916
rect 30979 7875 31037 7876
rect 33859 7916 33917 7917
rect 33859 7876 33868 7916
rect 33908 7876 33917 7916
rect 33859 7875 33917 7876
rect 37507 7916 37565 7917
rect 37507 7876 37516 7916
rect 37556 7876 37565 7916
rect 37507 7875 37565 7876
rect 37699 7916 37757 7917
rect 37699 7876 37708 7916
rect 37748 7876 37757 7916
rect 37699 7875 37757 7876
rect 38275 7916 38333 7917
rect 38275 7876 38284 7916
rect 38324 7876 38333 7916
rect 38275 7875 38333 7876
rect 38659 7916 38717 7917
rect 38659 7876 38668 7916
rect 38708 7876 38717 7916
rect 38659 7875 38717 7876
rect 40867 7916 40925 7917
rect 40867 7876 40876 7916
rect 40916 7876 40925 7916
rect 40867 7875 40925 7876
rect 41251 7916 41309 7917
rect 41251 7876 41260 7916
rect 41300 7876 41309 7916
rect 41251 7875 41309 7876
rect 26083 7864 26141 7865
rect 33675 7832 33717 7841
rect 33675 7792 33676 7832
rect 33716 7792 33717 7832
rect 33675 7783 33717 7792
rect 41451 7832 41493 7841
rect 41451 7792 41452 7832
rect 41492 7792 41493 7832
rect 41451 7783 41493 7792
rect 6219 7748 6261 7757
rect 6219 7708 6220 7748
rect 6260 7708 6261 7748
rect 6219 7699 6261 7708
rect 9195 7748 9237 7757
rect 9195 7708 9196 7748
rect 9236 7708 9237 7748
rect 9195 7699 9237 7708
rect 30219 7748 30261 7757
rect 30219 7708 30220 7748
rect 30260 7708 30261 7748
rect 30219 7699 30261 7708
rect 35499 7748 35541 7757
rect 35499 7708 35500 7748
rect 35540 7708 35541 7748
rect 35499 7699 35541 7708
rect 37323 7748 37365 7757
rect 37323 7708 37324 7748
rect 37364 7708 37365 7748
rect 37323 7699 37365 7708
rect 38091 7748 38133 7757
rect 38091 7708 38092 7748
rect 38132 7708 38133 7748
rect 38091 7699 38133 7708
rect 38475 7748 38517 7757
rect 38475 7708 38476 7748
rect 38516 7708 38517 7748
rect 38475 7699 38517 7708
rect 41067 7748 41109 7757
rect 41067 7708 41068 7748
rect 41108 7708 41109 7748
rect 41067 7699 41109 7708
rect 1152 7580 41856 7604
rect 1152 7540 3688 7580
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 4056 7540 18808 7580
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 19176 7540 33928 7580
rect 33968 7540 34010 7580
rect 34050 7540 34092 7580
rect 34132 7540 34174 7580
rect 34214 7540 34256 7580
rect 34296 7540 41856 7580
rect 1152 7516 41856 7540
rect 6027 7412 6069 7421
rect 6027 7372 6028 7412
rect 6068 7372 6069 7412
rect 6027 7363 6069 7372
rect 6979 7412 7037 7413
rect 6979 7372 6988 7412
rect 7028 7372 7037 7412
rect 6979 7371 7037 7372
rect 7371 7412 7413 7421
rect 7371 7372 7372 7412
rect 7412 7372 7413 7412
rect 7371 7363 7413 7372
rect 7851 7412 7893 7421
rect 7851 7372 7852 7412
rect 7892 7372 7893 7412
rect 7851 7363 7893 7372
rect 10443 7412 10485 7421
rect 10443 7372 10444 7412
rect 10484 7372 10485 7412
rect 10443 7363 10485 7372
rect 10827 7412 10869 7421
rect 10827 7372 10828 7412
rect 10868 7372 10869 7412
rect 10827 7363 10869 7372
rect 11019 7412 11061 7421
rect 11019 7372 11020 7412
rect 11060 7372 11061 7412
rect 11019 7363 11061 7372
rect 12651 7412 12693 7421
rect 12651 7372 12652 7412
rect 12692 7372 12693 7412
rect 12651 7363 12693 7372
rect 15723 7412 15765 7421
rect 15723 7372 15724 7412
rect 15764 7372 15765 7412
rect 15723 7363 15765 7372
rect 22443 7412 22485 7421
rect 22443 7372 22444 7412
rect 22484 7372 22485 7412
rect 22443 7363 22485 7372
rect 24075 7412 24117 7421
rect 24075 7372 24076 7412
rect 24116 7372 24117 7412
rect 24075 7363 24117 7372
rect 26187 7412 26229 7421
rect 26187 7372 26188 7412
rect 26228 7372 26229 7412
rect 26187 7363 26229 7372
rect 31851 7412 31893 7421
rect 31851 7372 31852 7412
rect 31892 7372 31893 7412
rect 31851 7363 31893 7372
rect 33483 7412 33525 7421
rect 33483 7372 33484 7412
rect 33524 7372 33525 7412
rect 33483 7363 33525 7372
rect 35403 7412 35445 7421
rect 35403 7372 35404 7412
rect 35444 7372 35445 7412
rect 35403 7363 35445 7372
rect 41259 7412 41301 7421
rect 41259 7372 41260 7412
rect 41300 7372 41301 7412
rect 41259 7363 41301 7372
rect 10243 7244 10301 7245
rect 10243 7204 10252 7244
rect 10292 7204 10301 7244
rect 10243 7203 10301 7204
rect 10627 7244 10685 7245
rect 10627 7204 10636 7244
rect 10676 7204 10685 7244
rect 10627 7203 10685 7204
rect 12835 7244 12893 7245
rect 12835 7204 12844 7244
rect 12884 7204 12893 7244
rect 12835 7203 12893 7204
rect 13803 7244 13845 7253
rect 13803 7204 13804 7244
rect 13844 7204 13845 7244
rect 13803 7195 13845 7204
rect 15523 7244 15581 7245
rect 15523 7204 15532 7244
rect 15572 7204 15581 7244
rect 15523 7203 15581 7204
rect 18603 7244 18645 7253
rect 18603 7204 18604 7244
rect 18644 7204 18645 7244
rect 18603 7195 18645 7204
rect 28299 7244 28341 7253
rect 28299 7204 28300 7244
rect 28340 7204 28341 7244
rect 28299 7195 28341 7204
rect 28395 7244 28437 7253
rect 28395 7204 28396 7244
rect 28436 7204 28437 7244
rect 28395 7195 28437 7204
rect 29827 7244 29885 7245
rect 29827 7204 29836 7244
rect 29876 7204 29885 7244
rect 29827 7203 29885 7204
rect 35587 7244 35645 7245
rect 35587 7204 35596 7244
rect 35636 7204 35645 7244
rect 35587 7203 35645 7204
rect 35779 7244 35837 7245
rect 35779 7204 35788 7244
rect 35828 7204 35837 7244
rect 35779 7203 35837 7204
rect 36355 7244 36413 7245
rect 36355 7204 36364 7244
rect 36404 7204 36413 7244
rect 36355 7203 36413 7204
rect 41443 7244 41501 7245
rect 41443 7204 41452 7244
rect 41492 7204 41501 7244
rect 41443 7203 41501 7204
rect 1323 7160 1365 7169
rect 1323 7120 1324 7160
rect 1364 7120 1365 7160
rect 1323 7111 1365 7120
rect 1515 7160 1557 7169
rect 1515 7120 1516 7160
rect 1556 7120 1557 7160
rect 1515 7111 1557 7120
rect 1699 7160 1757 7161
rect 1699 7120 1708 7160
rect 1748 7120 1757 7160
rect 1699 7119 1757 7120
rect 2947 7160 3005 7161
rect 2947 7120 2956 7160
rect 2996 7120 3005 7160
rect 2947 7119 3005 7120
rect 3435 7160 3477 7169
rect 3435 7120 3436 7160
rect 3476 7120 3477 7160
rect 3435 7111 3477 7120
rect 3531 7160 3573 7169
rect 3531 7120 3532 7160
rect 3572 7120 3573 7160
rect 3531 7111 3573 7120
rect 3627 7160 3669 7169
rect 3627 7120 3628 7160
rect 3668 7120 3669 7160
rect 3627 7111 3669 7120
rect 4107 7160 4149 7169
rect 4107 7120 4108 7160
rect 4148 7120 4149 7160
rect 4107 7111 4149 7120
rect 4203 7160 4245 7169
rect 4203 7120 4204 7160
rect 4244 7120 4245 7160
rect 4203 7111 4245 7120
rect 4579 7160 4637 7161
rect 4579 7120 4588 7160
rect 4628 7120 4637 7160
rect 4579 7119 4637 7120
rect 5827 7160 5885 7161
rect 5827 7120 5836 7160
rect 5876 7120 5885 7160
rect 5827 7119 5885 7120
rect 6307 7160 6365 7161
rect 6307 7120 6316 7160
rect 6356 7120 6365 7160
rect 6307 7119 6365 7120
rect 6603 7160 6645 7169
rect 6603 7120 6604 7160
rect 6644 7120 6645 7160
rect 6603 7111 6645 7120
rect 6699 7160 6741 7169
rect 6699 7120 6700 7160
rect 6740 7120 6741 7160
rect 6699 7111 6741 7120
rect 7371 7160 7413 7169
rect 7371 7120 7372 7160
rect 7412 7120 7413 7160
rect 7371 7111 7413 7120
rect 7563 7160 7605 7169
rect 7563 7120 7564 7160
rect 7604 7120 7605 7160
rect 7563 7111 7605 7120
rect 7651 7160 7709 7161
rect 7651 7120 7660 7160
rect 7700 7120 7709 7160
rect 7651 7119 7709 7120
rect 8035 7160 8093 7161
rect 8035 7120 8044 7160
rect 8084 7120 8093 7160
rect 8035 7119 8093 7120
rect 9283 7160 9341 7161
rect 9283 7120 9292 7160
rect 9332 7120 9341 7160
rect 9283 7119 9341 7120
rect 9483 7160 9525 7169
rect 9483 7120 9484 7160
rect 9524 7120 9525 7160
rect 9483 7111 9525 7120
rect 9675 7160 9717 7169
rect 9675 7120 9676 7160
rect 9716 7120 9717 7160
rect 9675 7111 9717 7120
rect 9763 7160 9821 7161
rect 9763 7120 9772 7160
rect 9812 7120 9821 7160
rect 9763 7119 9821 7120
rect 10051 7160 10109 7161
rect 10051 7120 10060 7160
rect 10100 7120 10109 7160
rect 10051 7119 10109 7120
rect 11203 7160 11261 7161
rect 11203 7120 11212 7160
rect 11252 7120 11261 7160
rect 11203 7119 11261 7120
rect 12451 7160 12509 7161
rect 12451 7120 12460 7160
rect 12500 7120 12509 7160
rect 12451 7119 12509 7120
rect 13323 7160 13365 7169
rect 13323 7120 13324 7160
rect 13364 7120 13365 7160
rect 13323 7111 13365 7120
rect 13419 7160 13461 7169
rect 13419 7120 13420 7160
rect 13460 7120 13461 7160
rect 13419 7111 13461 7120
rect 13899 7160 13941 7169
rect 14859 7165 14901 7174
rect 13899 7120 13900 7160
rect 13940 7120 13941 7160
rect 13899 7111 13941 7120
rect 14371 7160 14429 7161
rect 14371 7120 14380 7160
rect 14420 7120 14429 7160
rect 14371 7119 14429 7120
rect 14859 7125 14860 7165
rect 14900 7125 14901 7165
rect 14859 7116 14901 7125
rect 15907 7160 15965 7161
rect 15907 7120 15916 7160
rect 15956 7120 15965 7160
rect 15907 7119 15965 7120
rect 17155 7160 17213 7161
rect 17155 7120 17164 7160
rect 17204 7120 17213 7160
rect 17155 7119 17213 7120
rect 18123 7160 18165 7169
rect 18123 7120 18124 7160
rect 18164 7120 18165 7160
rect 18123 7111 18165 7120
rect 18219 7160 18261 7169
rect 18219 7120 18220 7160
rect 18260 7120 18261 7160
rect 18219 7111 18261 7120
rect 18699 7160 18741 7169
rect 19659 7165 19701 7174
rect 18699 7120 18700 7160
rect 18740 7120 18741 7160
rect 18699 7111 18741 7120
rect 19171 7160 19229 7161
rect 19171 7120 19180 7160
rect 19220 7120 19229 7160
rect 19171 7119 19229 7120
rect 19659 7125 19660 7165
rect 19700 7125 19701 7165
rect 19659 7116 19701 7125
rect 20995 7160 21053 7161
rect 20995 7120 21004 7160
rect 21044 7120 21053 7160
rect 20995 7119 21053 7120
rect 22243 7160 22301 7161
rect 22243 7120 22252 7160
rect 22292 7120 22301 7160
rect 22243 7119 22301 7120
rect 22627 7160 22685 7161
rect 22627 7120 22636 7160
rect 22676 7120 22685 7160
rect 22627 7119 22685 7120
rect 23875 7160 23933 7161
rect 23875 7120 23884 7160
rect 23924 7120 23933 7160
rect 23875 7119 23933 7120
rect 24739 7160 24797 7161
rect 24739 7120 24748 7160
rect 24788 7120 24797 7160
rect 24739 7119 24797 7120
rect 25987 7160 26045 7161
rect 25987 7120 25996 7160
rect 26036 7120 26045 7160
rect 25987 7119 26045 7120
rect 27819 7160 27861 7169
rect 27819 7120 27820 7160
rect 27860 7120 27861 7160
rect 27819 7111 27861 7120
rect 27915 7160 27957 7169
rect 29355 7165 29397 7174
rect 27915 7120 27916 7160
rect 27956 7120 27957 7160
rect 27915 7111 27957 7120
rect 28867 7160 28925 7161
rect 28867 7120 28876 7160
rect 28916 7120 28925 7160
rect 28867 7119 28925 7120
rect 29355 7125 29356 7165
rect 29396 7125 29397 7165
rect 29355 7116 29397 7125
rect 30211 7160 30269 7161
rect 30211 7120 30220 7160
rect 30260 7120 30269 7160
rect 30211 7119 30269 7120
rect 31459 7160 31517 7161
rect 31459 7120 31468 7160
rect 31508 7120 31517 7160
rect 31459 7119 31517 7120
rect 32035 7160 32093 7161
rect 32035 7120 32044 7160
rect 32084 7120 32093 7160
rect 32035 7119 32093 7120
rect 33283 7160 33341 7161
rect 33283 7120 33292 7160
rect 33332 7120 33341 7160
rect 33283 7119 33341 7120
rect 33667 7160 33725 7161
rect 33667 7120 33676 7160
rect 33716 7120 33725 7160
rect 33667 7119 33725 7120
rect 34915 7160 34973 7161
rect 34915 7120 34924 7160
rect 34964 7120 34973 7160
rect 34915 7119 34973 7120
rect 36547 7160 36605 7161
rect 36547 7120 36556 7160
rect 36596 7120 36605 7160
rect 36547 7119 36605 7120
rect 37795 7160 37853 7161
rect 37795 7120 37804 7160
rect 37844 7120 37853 7160
rect 37795 7119 37853 7120
rect 38371 7160 38429 7161
rect 38371 7120 38380 7160
rect 38420 7120 38429 7160
rect 38371 7119 38429 7120
rect 39619 7160 39677 7161
rect 39619 7120 39628 7160
rect 39668 7120 39677 7160
rect 39619 7119 39677 7120
rect 39811 7160 39869 7161
rect 39811 7120 39820 7160
rect 39860 7120 39869 7160
rect 39811 7119 39869 7120
rect 41059 7160 41117 7161
rect 41059 7120 41068 7160
rect 41108 7120 41117 7160
rect 41059 7119 41117 7120
rect 3147 7076 3189 7085
rect 3147 7036 3148 7076
rect 3188 7036 3189 7076
rect 3147 7027 3189 7036
rect 15051 7076 15093 7085
rect 15051 7036 15052 7076
rect 15092 7036 15093 7076
rect 15051 7027 15093 7036
rect 19851 7076 19893 7085
rect 19851 7036 19852 7076
rect 19892 7036 19893 7076
rect 19851 7027 19893 7036
rect 1419 6992 1461 7001
rect 1419 6952 1420 6992
rect 1460 6952 1461 6992
rect 1419 6943 1461 6952
rect 3715 6992 3773 6993
rect 3715 6952 3724 6992
rect 3764 6952 3773 6992
rect 3715 6951 3773 6952
rect 3907 6992 3965 6993
rect 3907 6952 3916 6992
rect 3956 6952 3965 6992
rect 3907 6951 3965 6952
rect 9571 6992 9629 6993
rect 9571 6952 9580 6992
rect 9620 6952 9629 6992
rect 9571 6951 9629 6952
rect 9963 6992 10005 7001
rect 9963 6952 9964 6992
rect 10004 6952 10005 6992
rect 9963 6943 10005 6952
rect 17355 6992 17397 7001
rect 17355 6952 17356 6992
rect 17396 6952 17397 6992
rect 17355 6943 17397 6952
rect 29547 6992 29589 7001
rect 29547 6952 29548 6992
rect 29588 6952 29589 6992
rect 29547 6943 29589 6952
rect 30027 6992 30069 7001
rect 30027 6952 30028 6992
rect 30068 6952 30069 6992
rect 30027 6943 30069 6952
rect 31659 6992 31701 7001
rect 31659 6952 31660 6992
rect 31700 6952 31701 6992
rect 31659 6943 31701 6952
rect 35979 6992 36021 7001
rect 35979 6952 35980 6992
rect 36020 6952 36021 6992
rect 35979 6943 36021 6952
rect 36171 6992 36213 7001
rect 36171 6952 36172 6992
rect 36212 6952 36213 6992
rect 36171 6943 36213 6952
rect 37995 6992 38037 7001
rect 37995 6952 37996 6992
rect 38036 6952 38037 6992
rect 37995 6943 38037 6952
rect 38187 6992 38229 7001
rect 38187 6952 38188 6992
rect 38228 6952 38229 6992
rect 38187 6943 38229 6952
rect 41643 6992 41685 7001
rect 41643 6952 41644 6992
rect 41684 6952 41685 6992
rect 41643 6943 41685 6952
rect 1152 6824 41856 6848
rect 1152 6784 4928 6824
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 5296 6784 20048 6824
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20416 6784 35168 6824
rect 35208 6784 35250 6824
rect 35290 6784 35332 6824
rect 35372 6784 35414 6824
rect 35454 6784 35496 6824
rect 35536 6784 41856 6824
rect 1152 6760 41856 6784
rect 4683 6656 4725 6665
rect 4683 6616 4684 6656
rect 4724 6616 4725 6656
rect 4683 6607 4725 6616
rect 5155 6656 5213 6657
rect 5155 6616 5164 6656
rect 5204 6616 5213 6656
rect 5155 6615 5213 6616
rect 5923 6656 5981 6657
rect 5923 6616 5932 6656
rect 5972 6616 5981 6656
rect 5923 6615 5981 6616
rect 8419 6656 8477 6657
rect 8419 6616 8428 6656
rect 8468 6616 8477 6656
rect 8419 6615 8477 6616
rect 10251 6656 10293 6665
rect 10251 6616 10252 6656
rect 10292 6616 10293 6656
rect 10251 6607 10293 6616
rect 12459 6656 12501 6665
rect 12459 6616 12460 6656
rect 12500 6616 12501 6656
rect 12459 6607 12501 6616
rect 14091 6656 14133 6665
rect 14091 6616 14092 6656
rect 14132 6616 14133 6656
rect 14091 6607 14133 6616
rect 17739 6656 17781 6665
rect 17739 6616 17740 6656
rect 17780 6616 17781 6656
rect 17739 6607 17781 6616
rect 25707 6656 25749 6665
rect 25707 6616 25708 6656
rect 25748 6616 25749 6656
rect 25707 6607 25749 6616
rect 31563 6656 31605 6665
rect 31563 6616 31564 6656
rect 31604 6616 31605 6656
rect 31563 6607 31605 6616
rect 31947 6656 31989 6665
rect 31947 6616 31948 6656
rect 31988 6616 31989 6656
rect 31947 6607 31989 6616
rect 32523 6656 32565 6665
rect 32523 6616 32524 6656
rect 32564 6616 32565 6656
rect 32523 6607 32565 6616
rect 34731 6656 34773 6665
rect 34731 6616 34732 6656
rect 34772 6616 34773 6656
rect 34731 6607 34773 6616
rect 36843 6656 36885 6665
rect 36843 6616 36844 6656
rect 36884 6616 36885 6656
rect 36843 6607 36885 6616
rect 37419 6656 37461 6665
rect 37419 6616 37420 6656
rect 37460 6616 37461 6656
rect 37419 6607 37461 6616
rect 39435 6656 39477 6665
rect 39435 6616 39436 6656
rect 39476 6616 39477 6656
rect 39435 6607 39477 6616
rect 41067 6656 41109 6665
rect 41067 6616 41068 6656
rect 41108 6616 41109 6656
rect 41067 6607 41109 6616
rect 6507 6572 6549 6581
rect 6507 6532 6508 6572
rect 6548 6532 6549 6572
rect 6507 6523 6549 6532
rect 15723 6572 15765 6581
rect 15723 6532 15724 6572
rect 15764 6532 15765 6572
rect 15723 6523 15765 6532
rect 20619 6572 20661 6581
rect 20619 6532 20620 6572
rect 20660 6532 20661 6572
rect 20619 6523 20661 6532
rect 23691 6572 23733 6581
rect 23691 6532 23692 6572
rect 23732 6532 23733 6572
rect 23691 6523 23733 6532
rect 27531 6572 27573 6581
rect 27531 6532 27532 6572
rect 27572 6532 27573 6572
rect 27531 6523 27573 6532
rect 29547 6572 29589 6581
rect 29547 6532 29548 6572
rect 29588 6532 29589 6572
rect 29547 6523 29589 6532
rect 1219 6488 1277 6489
rect 1219 6448 1228 6488
rect 1268 6448 1277 6488
rect 1219 6447 1277 6448
rect 2467 6488 2525 6489
rect 2467 6448 2476 6488
rect 2516 6448 2525 6488
rect 2467 6447 2525 6448
rect 2955 6488 2997 6497
rect 2955 6448 2956 6488
rect 2996 6448 2997 6488
rect 2955 6439 2997 6448
rect 3051 6488 3093 6497
rect 3051 6448 3052 6488
rect 3092 6448 3093 6488
rect 3051 6439 3093 6448
rect 3435 6488 3477 6497
rect 3435 6448 3436 6488
rect 3476 6448 3477 6488
rect 3435 6439 3477 6448
rect 4003 6488 4061 6489
rect 4003 6448 4012 6488
rect 4052 6448 4061 6488
rect 4003 6447 4061 6448
rect 4491 6483 4533 6492
rect 4491 6443 4492 6483
rect 4532 6443 4533 6483
rect 4491 6434 4533 6443
rect 4875 6488 4917 6497
rect 4875 6448 4876 6488
rect 4916 6448 4917 6488
rect 4875 6439 4917 6448
rect 4971 6488 5013 6497
rect 4971 6448 4972 6488
rect 5012 6448 5013 6488
rect 4971 6439 5013 6448
rect 5067 6488 5109 6497
rect 5067 6448 5068 6488
rect 5108 6448 5109 6488
rect 5067 6439 5109 6448
rect 5355 6488 5397 6497
rect 5355 6448 5356 6488
rect 5396 6448 5397 6488
rect 5355 6439 5397 6448
rect 5539 6488 5597 6489
rect 5539 6448 5548 6488
rect 5588 6448 5597 6488
rect 5539 6447 5597 6448
rect 5731 6488 5789 6489
rect 5731 6448 5740 6488
rect 5780 6448 5789 6488
rect 5731 6447 5789 6448
rect 5835 6488 5877 6497
rect 5835 6448 5836 6488
rect 5876 6448 5877 6488
rect 5835 6439 5877 6448
rect 6027 6488 6069 6497
rect 6027 6448 6028 6488
rect 6068 6448 6069 6488
rect 6027 6439 6069 6448
rect 6219 6488 6261 6497
rect 6219 6448 6220 6488
rect 6260 6448 6261 6488
rect 6219 6439 6261 6448
rect 6315 6488 6357 6497
rect 6315 6448 6316 6488
rect 6356 6448 6357 6488
rect 6315 6439 6357 6448
rect 6411 6488 6453 6497
rect 6411 6448 6412 6488
rect 6452 6448 6453 6488
rect 6411 6439 6453 6448
rect 6699 6488 6741 6497
rect 6699 6448 6700 6488
rect 6740 6448 6741 6488
rect 6699 6439 6741 6448
rect 6891 6488 6933 6497
rect 6891 6448 6892 6488
rect 6932 6448 6933 6488
rect 6891 6439 6933 6448
rect 6987 6488 7029 6497
rect 6987 6448 6988 6488
rect 7028 6448 7029 6488
rect 6987 6439 7029 6448
rect 7267 6488 7325 6489
rect 7267 6448 7276 6488
rect 7316 6448 7325 6488
rect 7267 6447 7325 6448
rect 7563 6488 7605 6497
rect 7563 6448 7564 6488
rect 7604 6448 7605 6488
rect 7563 6439 7605 6448
rect 7659 6488 7701 6497
rect 7659 6448 7660 6488
rect 7700 6448 7701 6488
rect 7659 6439 7701 6448
rect 8139 6488 8181 6497
rect 8139 6448 8140 6488
rect 8180 6448 8181 6488
rect 8139 6439 8181 6448
rect 8235 6488 8277 6497
rect 8235 6448 8236 6488
rect 8276 6448 8277 6488
rect 8235 6439 8277 6448
rect 8331 6488 8373 6497
rect 8331 6448 8332 6488
rect 8372 6448 8373 6488
rect 8331 6439 8373 6448
rect 8803 6488 8861 6489
rect 8803 6448 8812 6488
rect 8852 6448 8861 6488
rect 8803 6447 8861 6448
rect 10051 6488 10109 6489
rect 10051 6448 10060 6488
rect 10100 6448 10109 6488
rect 10051 6447 10109 6448
rect 10443 6488 10485 6497
rect 10443 6448 10444 6488
rect 10484 6448 10485 6488
rect 10443 6439 10485 6448
rect 10635 6488 10677 6497
rect 10635 6448 10636 6488
rect 10676 6448 10677 6488
rect 10635 6439 10677 6448
rect 10723 6488 10781 6489
rect 10723 6448 10732 6488
rect 10772 6448 10781 6488
rect 10723 6447 10781 6448
rect 11011 6488 11069 6489
rect 11011 6448 11020 6488
rect 11060 6448 11069 6488
rect 11011 6447 11069 6448
rect 12259 6488 12317 6489
rect 12259 6448 12268 6488
rect 12308 6448 12317 6488
rect 12259 6447 12317 6448
rect 12643 6488 12701 6489
rect 12643 6448 12652 6488
rect 12692 6448 12701 6488
rect 12643 6447 12701 6448
rect 13891 6488 13949 6489
rect 13891 6448 13900 6488
rect 13940 6448 13949 6488
rect 13891 6447 13949 6448
rect 14275 6488 14333 6489
rect 14275 6448 14284 6488
rect 14324 6448 14333 6488
rect 14275 6447 14333 6448
rect 15523 6488 15581 6489
rect 15523 6448 15532 6488
rect 15572 6448 15581 6488
rect 15523 6447 15581 6448
rect 16011 6488 16053 6497
rect 16011 6448 16012 6488
rect 16052 6448 16053 6488
rect 16011 6439 16053 6448
rect 16107 6488 16149 6497
rect 16107 6448 16108 6488
rect 16148 6448 16149 6488
rect 16107 6439 16149 6448
rect 16491 6488 16533 6497
rect 16491 6448 16492 6488
rect 16532 6448 16533 6488
rect 16491 6439 16533 6448
rect 17059 6488 17117 6489
rect 17059 6448 17068 6488
rect 17108 6448 17117 6488
rect 17059 6447 17117 6448
rect 17547 6483 17589 6492
rect 17547 6443 17548 6483
rect 17588 6443 17589 6483
rect 17547 6434 17589 6443
rect 18891 6488 18933 6497
rect 18891 6448 18892 6488
rect 18932 6448 18933 6488
rect 18891 6439 18933 6448
rect 18987 6488 19029 6497
rect 18987 6448 18988 6488
rect 19028 6448 19029 6488
rect 18987 6439 19029 6448
rect 19371 6488 19413 6497
rect 19371 6448 19372 6488
rect 19412 6448 19413 6488
rect 19371 6439 19413 6448
rect 19467 6488 19509 6497
rect 19467 6448 19468 6488
rect 19508 6448 19509 6488
rect 19467 6439 19509 6448
rect 19939 6488 19997 6489
rect 19939 6448 19948 6488
rect 19988 6448 19997 6488
rect 22243 6488 22301 6489
rect 19939 6447 19997 6448
rect 20427 6474 20469 6483
rect 20427 6434 20428 6474
rect 20468 6434 20469 6474
rect 22243 6448 22252 6488
rect 22292 6448 22301 6488
rect 22243 6447 22301 6448
rect 23491 6488 23549 6489
rect 23491 6448 23500 6488
rect 23540 6448 23549 6488
rect 23491 6447 23549 6448
rect 23979 6488 24021 6497
rect 23979 6448 23980 6488
rect 24020 6448 24021 6488
rect 23979 6439 24021 6448
rect 24075 6488 24117 6497
rect 24075 6448 24076 6488
rect 24116 6448 24117 6488
rect 24075 6439 24117 6448
rect 24459 6488 24501 6497
rect 24459 6448 24460 6488
rect 24500 6448 24501 6488
rect 24459 6439 24501 6448
rect 25027 6488 25085 6489
rect 25027 6448 25036 6488
rect 25076 6448 25085 6488
rect 26083 6488 26141 6489
rect 25027 6447 25085 6448
rect 25563 6478 25605 6487
rect 20427 6425 20469 6434
rect 25563 6438 25564 6478
rect 25604 6438 25605 6478
rect 26083 6448 26092 6488
rect 26132 6448 26141 6488
rect 26083 6447 26141 6448
rect 27331 6488 27389 6489
rect 27331 6448 27340 6488
rect 27380 6448 27389 6488
rect 27331 6447 27389 6448
rect 27819 6488 27861 6497
rect 27819 6448 27820 6488
rect 27860 6448 27861 6488
rect 27819 6439 27861 6448
rect 27915 6488 27957 6497
rect 27915 6448 27916 6488
rect 27956 6448 27957 6488
rect 27915 6439 27957 6448
rect 28395 6488 28437 6497
rect 28395 6448 28396 6488
rect 28436 6448 28437 6488
rect 28395 6439 28437 6448
rect 28867 6488 28925 6489
rect 28867 6448 28876 6488
rect 28916 6448 28925 6488
rect 29835 6488 29877 6497
rect 28867 6447 28925 6448
rect 29355 6474 29397 6483
rect 25563 6429 25605 6438
rect 29355 6434 29356 6474
rect 29396 6434 29397 6474
rect 29835 6448 29836 6488
rect 29876 6448 29877 6488
rect 29835 6439 29877 6448
rect 29931 6488 29973 6497
rect 29931 6448 29932 6488
rect 29972 6448 29973 6488
rect 29931 6439 29973 6448
rect 30411 6488 30453 6497
rect 30411 6448 30412 6488
rect 30452 6448 30453 6488
rect 30411 6439 30453 6448
rect 30883 6488 30941 6489
rect 30883 6448 30892 6488
rect 30932 6448 30941 6488
rect 33003 6488 33045 6497
rect 30883 6447 30941 6448
rect 31419 6478 31461 6487
rect 29355 6425 29397 6434
rect 31419 6438 31420 6478
rect 31460 6438 31461 6478
rect 33003 6448 33004 6488
rect 33044 6448 33045 6488
rect 33003 6439 33045 6448
rect 33099 6488 33141 6497
rect 33099 6448 33100 6488
rect 33140 6448 33141 6488
rect 33099 6439 33141 6448
rect 33579 6488 33621 6497
rect 33579 6448 33580 6488
rect 33620 6448 33621 6488
rect 33579 6439 33621 6448
rect 34051 6488 34109 6489
rect 34051 6448 34060 6488
rect 34100 6448 34109 6488
rect 35115 6488 35157 6497
rect 34051 6447 34109 6448
rect 34587 6446 34629 6455
rect 31419 6429 31461 6438
rect 3531 6404 3573 6413
rect 3531 6364 3532 6404
rect 3572 6364 3573 6404
rect 3531 6355 3573 6364
rect 16587 6404 16629 6413
rect 16587 6364 16588 6404
rect 16628 6364 16629 6404
rect 16587 6355 16629 6364
rect 24555 6404 24597 6413
rect 24555 6364 24556 6404
rect 24596 6364 24597 6404
rect 24555 6355 24597 6364
rect 28299 6404 28341 6413
rect 28299 6364 28300 6404
rect 28340 6364 28341 6404
rect 28299 6355 28341 6364
rect 30315 6404 30357 6413
rect 30315 6364 30316 6404
rect 30356 6364 30357 6404
rect 30315 6355 30357 6364
rect 31747 6404 31805 6405
rect 31747 6364 31756 6404
rect 31796 6364 31805 6404
rect 31747 6363 31805 6364
rect 32131 6404 32189 6405
rect 32131 6364 32140 6404
rect 32180 6364 32189 6404
rect 32131 6363 32189 6364
rect 32707 6404 32765 6405
rect 32707 6364 32716 6404
rect 32756 6364 32765 6404
rect 32707 6363 32765 6364
rect 33483 6404 33525 6413
rect 33483 6364 33484 6404
rect 33524 6364 33525 6404
rect 34587 6406 34588 6446
rect 34628 6406 34629 6446
rect 35115 6448 35116 6488
rect 35156 6448 35157 6488
rect 35115 6439 35157 6448
rect 35211 6488 35253 6497
rect 35211 6448 35212 6488
rect 35252 6448 35253 6488
rect 35211 6439 35253 6448
rect 35595 6488 35637 6497
rect 35595 6448 35596 6488
rect 35636 6448 35637 6488
rect 36163 6488 36221 6489
rect 35595 6439 35637 6448
rect 35691 6446 35733 6455
rect 36163 6448 36172 6488
rect 36212 6448 36221 6488
rect 37707 6488 37749 6497
rect 36163 6447 36221 6448
rect 36651 6474 36693 6483
rect 34587 6397 34629 6406
rect 35691 6406 35692 6446
rect 35732 6406 35733 6446
rect 36651 6434 36652 6474
rect 36692 6434 36693 6474
rect 37707 6448 37708 6488
rect 37748 6448 37749 6488
rect 37707 6439 37749 6448
rect 37803 6488 37845 6497
rect 37803 6448 37804 6488
rect 37844 6448 37845 6488
rect 37803 6439 37845 6448
rect 38187 6488 38229 6497
rect 38187 6448 38188 6488
rect 38228 6448 38229 6488
rect 38187 6439 38229 6448
rect 38283 6488 38325 6497
rect 38283 6448 38284 6488
rect 38324 6448 38325 6488
rect 38283 6439 38325 6448
rect 38755 6488 38813 6489
rect 38755 6448 38764 6488
rect 38804 6448 38813 6488
rect 38755 6447 38813 6448
rect 39243 6483 39285 6492
rect 39243 6443 39244 6483
rect 39284 6443 39285 6483
rect 39243 6434 39285 6443
rect 36651 6425 36693 6434
rect 35691 6397 35733 6406
rect 37219 6404 37277 6405
rect 33483 6355 33525 6364
rect 37219 6364 37228 6404
rect 37268 6364 37277 6404
rect 37219 6363 37277 6364
rect 39811 6404 39869 6405
rect 39811 6364 39820 6404
rect 39860 6364 39869 6404
rect 39811 6363 39869 6364
rect 40387 6404 40445 6405
rect 40387 6364 40396 6404
rect 40436 6364 40445 6404
rect 40387 6363 40445 6364
rect 40867 6404 40925 6405
rect 40867 6364 40876 6404
rect 40916 6364 40925 6404
rect 40867 6363 40925 6364
rect 41251 6404 41309 6405
rect 41251 6364 41260 6404
rect 41300 6364 41309 6404
rect 41251 6363 41309 6364
rect 2667 6320 2709 6329
rect 2667 6280 2668 6320
rect 2708 6280 2709 6320
rect 2667 6271 2709 6280
rect 5451 6320 5493 6329
rect 5451 6280 5452 6320
rect 5492 6280 5493 6320
rect 5451 6271 5493 6280
rect 40011 6320 40053 6329
rect 40011 6280 40012 6320
rect 40052 6280 40053 6320
rect 40011 6271 40053 6280
rect 40203 6320 40245 6329
rect 40203 6280 40204 6320
rect 40244 6280 40245 6320
rect 40203 6271 40245 6280
rect 41451 6320 41493 6329
rect 41451 6280 41452 6320
rect 41492 6280 41493 6320
rect 41451 6271 41493 6280
rect 7939 6236 7997 6237
rect 7939 6196 7948 6236
rect 7988 6196 7997 6236
rect 7939 6195 7997 6196
rect 10443 6236 10485 6245
rect 10443 6196 10444 6236
rect 10484 6196 10485 6236
rect 10443 6187 10485 6196
rect 32331 6236 32373 6245
rect 32331 6196 32332 6236
rect 32372 6196 32373 6236
rect 32331 6187 32373 6196
rect 1152 6068 41856 6092
rect 1152 6028 3688 6068
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 4056 6028 18808 6068
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 19176 6028 33928 6068
rect 33968 6028 34010 6068
rect 34050 6028 34092 6068
rect 34132 6028 34174 6068
rect 34214 6028 34256 6068
rect 34296 6028 41856 6068
rect 1152 6004 41856 6028
rect 2763 5900 2805 5909
rect 2763 5860 2764 5900
rect 2804 5860 2805 5900
rect 2763 5851 2805 5860
rect 9763 5900 9821 5901
rect 9763 5860 9772 5900
rect 9812 5860 9821 5900
rect 9763 5859 9821 5860
rect 10539 5900 10581 5909
rect 10539 5860 10540 5900
rect 10580 5860 10581 5900
rect 10539 5851 10581 5860
rect 11499 5900 11541 5909
rect 11499 5860 11500 5900
rect 11540 5860 11541 5900
rect 11499 5851 11541 5860
rect 11883 5900 11925 5909
rect 11883 5860 11884 5900
rect 11924 5860 11925 5900
rect 11883 5851 11925 5860
rect 12267 5900 12309 5909
rect 12267 5860 12268 5900
rect 12308 5860 12309 5900
rect 12267 5851 12309 5860
rect 13227 5900 13269 5909
rect 13227 5860 13228 5900
rect 13268 5860 13269 5900
rect 13227 5851 13269 5860
rect 13803 5900 13845 5909
rect 13803 5860 13804 5900
rect 13844 5860 13845 5900
rect 13803 5851 13845 5860
rect 17931 5900 17973 5909
rect 17931 5860 17932 5900
rect 17972 5860 17973 5900
rect 17931 5851 17973 5860
rect 19563 5900 19605 5909
rect 19563 5860 19564 5900
rect 19604 5860 19605 5900
rect 19563 5851 19605 5860
rect 21195 5900 21237 5909
rect 21195 5860 21196 5900
rect 21236 5860 21237 5900
rect 21195 5851 21237 5860
rect 22827 5900 22869 5909
rect 22827 5860 22828 5900
rect 22868 5860 22869 5900
rect 22827 5851 22869 5860
rect 25803 5900 25845 5909
rect 25803 5860 25804 5900
rect 25844 5860 25845 5900
rect 25803 5851 25845 5860
rect 27531 5900 27573 5909
rect 27531 5860 27532 5900
rect 27572 5860 27573 5900
rect 27531 5851 27573 5860
rect 27723 5900 27765 5909
rect 27723 5860 27724 5900
rect 27764 5860 27765 5900
rect 27723 5851 27765 5860
rect 29355 5900 29397 5909
rect 29355 5860 29356 5900
rect 29396 5860 29397 5900
rect 29355 5851 29397 5860
rect 31659 5900 31701 5909
rect 31659 5860 31660 5900
rect 31700 5860 31701 5900
rect 31659 5851 31701 5860
rect 34923 5900 34965 5909
rect 34923 5860 34924 5900
rect 34964 5860 34965 5900
rect 34923 5851 34965 5860
rect 37035 5900 37077 5909
rect 37035 5860 37036 5900
rect 37076 5860 37077 5900
rect 37035 5851 37077 5860
rect 38187 5900 38229 5909
rect 38187 5860 38188 5900
rect 38228 5860 38229 5900
rect 38187 5851 38229 5860
rect 38571 5900 38613 5909
rect 38571 5860 38572 5900
rect 38612 5860 38613 5900
rect 38571 5851 38613 5860
rect 41067 5900 41109 5909
rect 41067 5860 41068 5900
rect 41108 5860 41109 5900
rect 41067 5851 41109 5860
rect 11211 5816 11253 5825
rect 11211 5776 11212 5816
rect 11252 5776 11253 5816
rect 11211 5767 11253 5776
rect 41451 5816 41493 5825
rect 41451 5776 41452 5816
rect 41492 5776 41493 5816
rect 41451 5767 41493 5776
rect 11683 5732 11741 5733
rect 11683 5692 11692 5732
rect 11732 5692 11741 5732
rect 11683 5691 11741 5692
rect 12067 5732 12125 5733
rect 12067 5692 12076 5732
rect 12116 5692 12125 5732
rect 12067 5691 12125 5692
rect 12451 5732 12509 5733
rect 12451 5692 12460 5732
rect 12500 5692 12509 5732
rect 12451 5691 12509 5692
rect 13411 5732 13469 5733
rect 13411 5692 13420 5732
rect 13460 5692 13469 5732
rect 13411 5691 13469 5692
rect 13603 5732 13661 5733
rect 13603 5692 13612 5732
rect 13652 5692 13661 5732
rect 13603 5691 13661 5692
rect 16291 5732 16349 5733
rect 16291 5692 16300 5732
rect 16340 5692 16349 5732
rect 16291 5691 16349 5692
rect 31075 5732 31133 5733
rect 31075 5692 31084 5732
rect 31124 5692 31133 5732
rect 31075 5691 31133 5692
rect 31459 5732 31517 5733
rect 31459 5692 31468 5732
rect 31508 5692 31517 5732
rect 31459 5691 31517 5692
rect 35203 5732 35261 5733
rect 35203 5692 35212 5732
rect 35252 5692 35261 5732
rect 35203 5691 35261 5692
rect 37411 5732 37469 5733
rect 37411 5692 37420 5732
rect 37460 5692 37469 5732
rect 37411 5691 37469 5692
rect 37603 5732 37661 5733
rect 37603 5692 37612 5732
rect 37652 5692 37661 5732
rect 37603 5691 37661 5692
rect 37987 5732 38045 5733
rect 37987 5692 37996 5732
rect 38036 5692 38045 5732
rect 37987 5691 38045 5692
rect 38371 5732 38429 5733
rect 38371 5692 38380 5732
rect 38420 5692 38429 5732
rect 38371 5691 38429 5692
rect 39339 5732 39381 5741
rect 39339 5692 39340 5732
rect 39380 5692 39381 5732
rect 39339 5683 39381 5692
rect 39435 5732 39477 5741
rect 39435 5692 39436 5732
rect 39476 5692 39477 5732
rect 39435 5683 39477 5692
rect 40867 5732 40925 5733
rect 40867 5692 40876 5732
rect 40916 5692 40925 5732
rect 40867 5691 40925 5692
rect 41251 5732 41309 5733
rect 41251 5692 41260 5732
rect 41300 5692 41309 5732
rect 41251 5691 41309 5692
rect 9997 5663 10039 5672
rect 1315 5648 1373 5649
rect 1315 5608 1324 5648
rect 1364 5608 1373 5648
rect 1315 5607 1373 5608
rect 2563 5648 2621 5649
rect 2563 5608 2572 5648
rect 2612 5608 2621 5648
rect 3339 5648 3381 5657
rect 2563 5607 2621 5608
rect 3243 5627 3285 5636
rect 3243 5587 3244 5627
rect 3284 5587 3285 5627
rect 3339 5608 3340 5648
rect 3380 5608 3381 5648
rect 3339 5599 3381 5608
rect 3435 5648 3477 5657
rect 3435 5608 3436 5648
rect 3476 5608 3477 5648
rect 3435 5599 3477 5608
rect 3723 5648 3765 5657
rect 3723 5608 3724 5648
rect 3764 5608 3765 5648
rect 3723 5599 3765 5608
rect 3819 5648 3861 5657
rect 3819 5608 3820 5648
rect 3860 5608 3861 5648
rect 3819 5599 3861 5608
rect 3915 5648 3957 5657
rect 3915 5608 3916 5648
rect 3956 5608 3957 5648
rect 3915 5599 3957 5608
rect 4011 5648 4053 5657
rect 4011 5608 4012 5648
rect 4052 5608 4053 5648
rect 4011 5599 4053 5608
rect 4203 5648 4245 5657
rect 4203 5608 4204 5648
rect 4244 5608 4245 5648
rect 4203 5599 4245 5608
rect 4299 5648 4341 5657
rect 4299 5608 4300 5648
rect 4340 5608 4341 5648
rect 4299 5599 4341 5608
rect 4683 5648 4725 5657
rect 4683 5608 4684 5648
rect 4724 5608 4725 5648
rect 4683 5599 4725 5608
rect 4779 5648 4821 5657
rect 4779 5608 4780 5648
rect 4820 5608 4821 5648
rect 4779 5599 4821 5608
rect 4875 5648 4917 5657
rect 4875 5608 4876 5648
rect 4916 5608 4917 5648
rect 4875 5599 4917 5608
rect 5155 5648 5213 5649
rect 5155 5608 5164 5648
rect 5204 5608 5213 5648
rect 5155 5607 5213 5608
rect 6403 5648 6461 5649
rect 6403 5608 6412 5648
rect 6452 5608 6461 5648
rect 6403 5607 6461 5608
rect 6787 5648 6845 5649
rect 6787 5608 6796 5648
rect 6836 5608 6845 5648
rect 6787 5607 6845 5608
rect 8035 5648 8093 5649
rect 8035 5608 8044 5648
rect 8084 5608 8093 5648
rect 8035 5607 8093 5608
rect 8523 5648 8565 5657
rect 8523 5608 8524 5648
rect 8564 5608 8565 5648
rect 8523 5599 8565 5608
rect 8619 5648 8661 5657
rect 8619 5608 8620 5648
rect 8660 5608 8661 5648
rect 8619 5599 8661 5608
rect 9091 5648 9149 5649
rect 9091 5608 9100 5648
rect 9140 5608 9149 5648
rect 9091 5607 9149 5608
rect 9387 5648 9429 5657
rect 9387 5608 9388 5648
rect 9428 5608 9429 5648
rect 9997 5623 9998 5663
rect 10038 5623 10039 5663
rect 9997 5614 10039 5623
rect 10155 5648 10197 5657
rect 9387 5599 9429 5608
rect 10155 5608 10156 5648
rect 10196 5608 10197 5648
rect 10155 5599 10197 5608
rect 10251 5648 10293 5657
rect 10251 5608 10252 5648
rect 10292 5608 10293 5648
rect 10251 5599 10293 5608
rect 10435 5648 10493 5649
rect 10435 5608 10444 5648
rect 10484 5608 10493 5648
rect 10435 5607 10493 5608
rect 10531 5648 10589 5649
rect 10531 5608 10540 5648
rect 10580 5608 10589 5648
rect 10531 5607 10589 5608
rect 10819 5648 10877 5649
rect 10819 5608 10828 5648
rect 10868 5608 10877 5648
rect 10819 5607 10877 5608
rect 10923 5648 10965 5657
rect 10923 5608 10924 5648
rect 10964 5608 10965 5648
rect 10923 5599 10965 5608
rect 13987 5648 14045 5649
rect 13987 5608 13996 5648
rect 14036 5608 14045 5648
rect 13987 5607 14045 5608
rect 15235 5648 15293 5649
rect 15235 5608 15244 5648
rect 15284 5608 15293 5648
rect 15235 5607 15293 5608
rect 16483 5648 16541 5649
rect 16483 5608 16492 5648
rect 16532 5608 16541 5648
rect 16483 5607 16541 5608
rect 17731 5648 17789 5649
rect 17731 5608 17740 5648
rect 17780 5608 17789 5648
rect 17731 5607 17789 5608
rect 18115 5648 18173 5649
rect 18115 5608 18124 5648
rect 18164 5608 18173 5648
rect 18115 5607 18173 5608
rect 19363 5648 19421 5649
rect 19363 5608 19372 5648
rect 19412 5608 19421 5648
rect 19363 5607 19421 5608
rect 19747 5648 19805 5649
rect 19747 5608 19756 5648
rect 19796 5608 19805 5648
rect 19747 5607 19805 5608
rect 20995 5648 21053 5649
rect 20995 5608 21004 5648
rect 21044 5608 21053 5648
rect 20995 5607 21053 5608
rect 21379 5648 21437 5649
rect 21379 5608 21388 5648
rect 21428 5608 21437 5648
rect 21379 5607 21437 5608
rect 22627 5648 22685 5649
rect 22627 5608 22636 5648
rect 22676 5608 22685 5648
rect 22627 5607 22685 5608
rect 24355 5648 24413 5649
rect 24355 5608 24364 5648
rect 24404 5608 24413 5648
rect 24355 5607 24413 5608
rect 25603 5648 25661 5649
rect 25603 5608 25612 5648
rect 25652 5608 25661 5648
rect 25603 5607 25661 5608
rect 26083 5648 26141 5649
rect 26083 5608 26092 5648
rect 26132 5608 26141 5648
rect 26083 5607 26141 5608
rect 27331 5648 27389 5649
rect 27331 5608 27340 5648
rect 27380 5608 27389 5648
rect 27331 5607 27389 5608
rect 27907 5648 27965 5649
rect 27907 5608 27916 5648
rect 27956 5608 27965 5648
rect 27907 5607 27965 5608
rect 29155 5648 29213 5649
rect 29155 5608 29164 5648
rect 29204 5608 29213 5648
rect 29155 5607 29213 5608
rect 29539 5648 29597 5649
rect 29539 5608 29548 5648
rect 29588 5608 29597 5648
rect 29539 5607 29597 5608
rect 30787 5648 30845 5649
rect 30787 5608 30796 5648
rect 30836 5608 30845 5648
rect 30787 5607 30845 5608
rect 31843 5648 31901 5649
rect 31843 5608 31852 5648
rect 31892 5608 31901 5648
rect 31843 5607 31901 5608
rect 33091 5648 33149 5649
rect 33091 5608 33100 5648
rect 33140 5608 33149 5648
rect 33091 5607 33149 5608
rect 33475 5648 33533 5649
rect 33475 5608 33484 5648
rect 33524 5608 33533 5648
rect 33475 5607 33533 5608
rect 34723 5648 34781 5649
rect 34723 5608 34732 5648
rect 34772 5608 34781 5648
rect 34723 5607 34781 5608
rect 35587 5648 35645 5649
rect 35587 5608 35596 5648
rect 35636 5608 35645 5648
rect 35587 5607 35645 5608
rect 36835 5648 36893 5649
rect 36835 5608 36844 5648
rect 36884 5608 36893 5648
rect 36835 5607 36893 5608
rect 38859 5648 38901 5657
rect 38859 5608 38860 5648
rect 38900 5608 38901 5648
rect 38859 5599 38901 5608
rect 38955 5648 38997 5657
rect 40395 5653 40437 5662
rect 38955 5608 38956 5648
rect 38996 5608 38997 5648
rect 38955 5599 38997 5608
rect 39907 5648 39965 5649
rect 39907 5608 39916 5648
rect 39956 5608 39965 5648
rect 39907 5607 39965 5608
rect 40395 5613 40396 5653
rect 40436 5613 40437 5653
rect 40395 5604 40437 5613
rect 3243 5578 3285 5587
rect 8235 5564 8277 5573
rect 8235 5524 8236 5564
rect 8276 5524 8277 5564
rect 8235 5515 8277 5524
rect 9483 5564 9525 5573
rect 9483 5524 9484 5564
rect 9524 5524 9525 5564
rect 9483 5515 9525 5524
rect 40587 5564 40629 5573
rect 40587 5524 40588 5564
rect 40628 5524 40629 5564
rect 40587 5515 40629 5524
rect 3523 5480 3581 5481
rect 3523 5440 3532 5480
rect 3572 5440 3581 5480
rect 3523 5439 3581 5440
rect 4483 5480 4541 5481
rect 4483 5440 4492 5480
rect 4532 5440 4541 5480
rect 4483 5439 4541 5440
rect 4963 5480 5021 5481
rect 4963 5440 4972 5480
rect 5012 5440 5021 5480
rect 4963 5439 5021 5440
rect 6603 5480 6645 5489
rect 6603 5440 6604 5480
rect 6644 5440 6645 5480
rect 6603 5431 6645 5440
rect 8803 5480 8861 5481
rect 8803 5440 8812 5480
rect 8852 5440 8861 5480
rect 8803 5439 8861 5440
rect 15435 5480 15477 5489
rect 15435 5440 15436 5480
rect 15476 5440 15477 5480
rect 15435 5431 15477 5440
rect 16107 5480 16149 5489
rect 16107 5440 16108 5480
rect 16148 5440 16149 5480
rect 16107 5431 16149 5440
rect 31275 5480 31317 5489
rect 31275 5440 31276 5480
rect 31316 5440 31317 5480
rect 31275 5431 31317 5440
rect 33291 5480 33333 5489
rect 33291 5440 33292 5480
rect 33332 5440 33333 5480
rect 33291 5431 33333 5440
rect 35403 5480 35445 5489
rect 35403 5440 35404 5480
rect 35444 5440 35445 5480
rect 35403 5431 35445 5440
rect 37227 5480 37269 5489
rect 37227 5440 37228 5480
rect 37268 5440 37269 5480
rect 37227 5431 37269 5440
rect 37803 5480 37845 5489
rect 37803 5440 37804 5480
rect 37844 5440 37845 5480
rect 37803 5431 37845 5440
rect 10731 5422 10773 5431
rect 10731 5382 10732 5422
rect 10772 5382 10773 5422
rect 10731 5373 10773 5382
rect 1152 5312 41856 5336
rect 1152 5272 4928 5312
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 5296 5272 20048 5312
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20416 5272 35168 5312
rect 35208 5272 35250 5312
rect 35290 5272 35332 5312
rect 35372 5272 35414 5312
rect 35454 5272 35496 5312
rect 35536 5272 41856 5312
rect 1152 5248 41856 5272
rect 4683 5144 4725 5153
rect 4683 5104 4684 5144
rect 4724 5104 4725 5144
rect 4683 5095 4725 5104
rect 10435 5144 10493 5145
rect 10435 5104 10444 5144
rect 10484 5104 10493 5144
rect 10435 5103 10493 5104
rect 20619 5144 20661 5153
rect 20619 5104 20620 5144
rect 20660 5104 20661 5144
rect 20619 5095 20661 5104
rect 37227 5144 37269 5153
rect 37227 5104 37228 5144
rect 37268 5104 37269 5144
rect 37227 5095 37269 5104
rect 40971 5144 41013 5153
rect 40971 5104 40972 5144
rect 41012 5104 41013 5144
rect 40971 5095 41013 5104
rect 2667 5060 2709 5069
rect 2667 5020 2668 5060
rect 2708 5020 2709 5060
rect 2667 5011 2709 5020
rect 9003 5060 9045 5069
rect 9003 5020 9004 5060
rect 9044 5020 9045 5060
rect 9003 5011 9045 5020
rect 12075 5060 12117 5069
rect 12075 5020 12076 5060
rect 12116 5020 12117 5060
rect 12075 5011 12117 5020
rect 14091 5060 14133 5069
rect 14091 5020 14092 5060
rect 14132 5020 14133 5060
rect 14091 5011 14133 5020
rect 16491 5060 16533 5069
rect 16491 5020 16492 5060
rect 16532 5020 16533 5060
rect 16491 5011 16533 5020
rect 16779 5060 16821 5069
rect 16779 5020 16780 5060
rect 16820 5020 16821 5060
rect 16779 5011 16821 5020
rect 25515 5060 25557 5069
rect 25515 5020 25516 5060
rect 25556 5020 25557 5060
rect 25515 5011 25557 5020
rect 30891 5060 30933 5069
rect 30891 5020 30892 5060
rect 30932 5020 30933 5060
rect 30891 5011 30933 5020
rect 37419 5060 37461 5069
rect 37419 5020 37420 5060
rect 37460 5020 37461 5060
rect 37419 5011 37461 5020
rect 1219 4976 1277 4977
rect 1219 4936 1228 4976
rect 1268 4936 1277 4976
rect 1219 4935 1277 4936
rect 2467 4976 2525 4977
rect 2467 4936 2476 4976
rect 2516 4936 2525 4976
rect 2467 4935 2525 4936
rect 2955 4976 2997 4985
rect 2955 4936 2956 4976
rect 2996 4936 2997 4976
rect 2955 4927 2997 4936
rect 3051 4976 3093 4985
rect 3051 4936 3052 4976
rect 3092 4936 3093 4976
rect 3051 4927 3093 4936
rect 4003 4976 4061 4977
rect 4003 4936 4012 4976
rect 4052 4936 4061 4976
rect 4003 4935 4061 4936
rect 4491 4971 4533 4980
rect 4491 4931 4492 4971
rect 4532 4931 4533 4971
rect 5155 4976 5213 4977
rect 5155 4936 5164 4976
rect 5204 4936 5213 4976
rect 5155 4935 5213 4936
rect 6403 4976 6461 4977
rect 6403 4936 6412 4976
rect 6452 4936 6461 4976
rect 6403 4935 6461 4936
rect 6795 4976 6837 4985
rect 6795 4936 6796 4976
rect 6836 4936 6837 4976
rect 4491 4922 4533 4931
rect 6795 4927 6837 4936
rect 6987 4976 7029 4985
rect 6987 4936 6988 4976
rect 7028 4936 7029 4976
rect 6987 4927 7029 4936
rect 7275 4976 7317 4985
rect 7275 4936 7276 4976
rect 7316 4936 7317 4976
rect 7275 4927 7317 4936
rect 7371 4976 7413 4985
rect 7371 4936 7372 4976
rect 7412 4936 7413 4976
rect 7371 4927 7413 4936
rect 8323 4976 8381 4977
rect 8323 4936 8332 4976
rect 8372 4936 8381 4976
rect 8323 4935 8381 4936
rect 8811 4971 8853 4980
rect 8811 4931 8812 4971
rect 8852 4931 8853 4971
rect 9283 4976 9341 4977
rect 9283 4936 9292 4976
rect 9332 4936 9341 4976
rect 9283 4935 9341 4936
rect 9579 4976 9621 4985
rect 9579 4936 9580 4976
rect 9620 4936 9621 4976
rect 8811 4922 8853 4931
rect 9579 4927 9621 4936
rect 9675 4976 9717 4985
rect 9675 4936 9676 4976
rect 9716 4936 9717 4976
rect 9675 4927 9717 4936
rect 10155 4976 10197 4985
rect 10155 4936 10156 4976
rect 10196 4936 10197 4976
rect 10155 4927 10197 4936
rect 10251 4976 10293 4985
rect 10251 4936 10252 4976
rect 10292 4936 10293 4976
rect 10251 4927 10293 4936
rect 10627 4976 10685 4977
rect 10627 4936 10636 4976
rect 10676 4936 10685 4976
rect 10627 4935 10685 4936
rect 11875 4976 11933 4977
rect 11875 4936 11884 4976
rect 11924 4936 11933 4976
rect 11875 4935 11933 4936
rect 12363 4976 12405 4985
rect 12363 4936 12364 4976
rect 12404 4936 12405 4976
rect 12363 4927 12405 4936
rect 12459 4976 12501 4985
rect 12459 4936 12460 4976
rect 12500 4936 12501 4976
rect 12459 4927 12501 4936
rect 13411 4976 13469 4977
rect 13411 4936 13420 4976
rect 13460 4936 13469 4976
rect 14763 4976 14805 4985
rect 13411 4935 13469 4936
rect 13899 4962 13941 4971
rect 13899 4922 13900 4962
rect 13940 4922 13941 4962
rect 14763 4936 14764 4976
rect 14804 4936 14805 4976
rect 14763 4927 14805 4936
rect 14859 4976 14901 4985
rect 14859 4936 14860 4976
rect 14900 4936 14901 4976
rect 14859 4927 14901 4936
rect 15339 4976 15381 4985
rect 15339 4936 15340 4976
rect 15380 4936 15381 4976
rect 15339 4927 15381 4936
rect 15811 4976 15869 4977
rect 15811 4936 15820 4976
rect 15860 4936 15869 4976
rect 17443 4976 17501 4977
rect 15811 4935 15869 4936
rect 16299 4962 16341 4971
rect 13899 4913 13941 4922
rect 16299 4922 16300 4962
rect 16340 4922 16341 4962
rect 16299 4913 16341 4922
rect 16971 4962 17013 4971
rect 16971 4922 16972 4962
rect 17012 4922 17013 4962
rect 17443 4936 17452 4976
rect 17492 4936 17501 4976
rect 17443 4935 17501 4936
rect 17931 4976 17973 4985
rect 17931 4936 17932 4976
rect 17972 4936 17973 4976
rect 17931 4927 17973 4936
rect 18411 4976 18453 4985
rect 18411 4936 18412 4976
rect 18452 4936 18453 4976
rect 18411 4927 18453 4936
rect 18507 4976 18549 4985
rect 18507 4936 18508 4976
rect 18548 4936 18549 4976
rect 18507 4927 18549 4936
rect 19171 4976 19229 4977
rect 19171 4936 19180 4976
rect 19220 4936 19229 4976
rect 19171 4935 19229 4936
rect 20419 4976 20477 4977
rect 20419 4936 20428 4976
rect 20468 4936 20477 4976
rect 20419 4935 20477 4936
rect 21667 4976 21725 4977
rect 21667 4936 21676 4976
rect 21716 4936 21725 4976
rect 21667 4935 21725 4936
rect 22915 4976 22973 4977
rect 22915 4936 22924 4976
rect 22964 4936 22973 4976
rect 22915 4935 22973 4936
rect 23787 4976 23829 4985
rect 23787 4936 23788 4976
rect 23828 4936 23829 4976
rect 23787 4927 23829 4936
rect 23883 4976 23925 4985
rect 23883 4936 23884 4976
rect 23924 4936 23925 4976
rect 23883 4927 23925 4936
rect 24267 4976 24309 4985
rect 24267 4936 24268 4976
rect 24308 4936 24309 4976
rect 24267 4927 24309 4936
rect 24363 4976 24405 4985
rect 24363 4936 24364 4976
rect 24404 4936 24405 4976
rect 24363 4927 24405 4936
rect 24835 4976 24893 4977
rect 24835 4936 24844 4976
rect 24884 4936 24893 4976
rect 25891 4976 25949 4977
rect 24835 4935 24893 4936
rect 25371 4934 25413 4943
rect 25891 4936 25900 4976
rect 25940 4936 25949 4976
rect 25891 4935 25949 4936
rect 27139 4976 27197 4977
rect 27139 4936 27148 4976
rect 27188 4936 27197 4976
rect 27139 4935 27197 4936
rect 27907 4976 27965 4977
rect 27907 4936 27916 4976
rect 27956 4936 27965 4976
rect 27907 4935 27965 4936
rect 28867 4976 28925 4977
rect 28867 4936 28876 4976
rect 28916 4936 28925 4976
rect 28867 4935 28925 4936
rect 29163 4976 29205 4985
rect 29163 4936 29164 4976
rect 29204 4936 29205 4976
rect 16971 4913 17013 4922
rect 3435 4892 3477 4901
rect 3435 4852 3436 4892
rect 3476 4852 3477 4892
rect 3435 4843 3477 4852
rect 3531 4892 3573 4901
rect 3531 4852 3532 4892
rect 3572 4852 3573 4892
rect 3531 4843 3573 4852
rect 7755 4892 7797 4901
rect 7755 4852 7756 4892
rect 7796 4852 7797 4892
rect 7755 4843 7797 4852
rect 7851 4892 7893 4901
rect 7851 4852 7852 4892
rect 7892 4852 7893 4892
rect 7851 4843 7893 4852
rect 12843 4892 12885 4901
rect 12843 4852 12844 4892
rect 12884 4852 12885 4892
rect 12843 4843 12885 4852
rect 12939 4892 12981 4901
rect 12939 4852 12940 4892
rect 12980 4852 12981 4892
rect 12939 4843 12981 4852
rect 15243 4892 15285 4901
rect 15243 4852 15244 4892
rect 15284 4852 15285 4892
rect 15243 4843 15285 4852
rect 18027 4892 18069 4901
rect 25371 4894 25372 4934
rect 25412 4894 25413 4934
rect 29163 4927 29205 4936
rect 29259 4976 29301 4985
rect 29259 4936 29260 4976
rect 29300 4936 29301 4976
rect 29259 4927 29301 4936
rect 29739 4976 29781 4985
rect 29739 4936 29740 4976
rect 29780 4936 29781 4976
rect 29739 4927 29781 4936
rect 30211 4976 30269 4977
rect 30211 4936 30220 4976
rect 30260 4936 30269 4976
rect 31267 4976 31325 4977
rect 30211 4935 30269 4936
rect 30699 4962 30741 4971
rect 30699 4922 30700 4962
rect 30740 4922 30741 4962
rect 31267 4936 31276 4976
rect 31316 4936 31325 4976
rect 31267 4935 31325 4936
rect 32515 4976 32573 4977
rect 32515 4936 32524 4976
rect 32564 4936 32573 4976
rect 32515 4935 32573 4936
rect 33283 4976 33341 4977
rect 33283 4936 33292 4976
rect 33332 4936 33341 4976
rect 33283 4935 33341 4936
rect 34531 4976 34589 4977
rect 34531 4936 34540 4976
rect 34580 4936 34589 4976
rect 34531 4935 34589 4936
rect 35499 4976 35541 4985
rect 35499 4936 35500 4976
rect 35540 4936 35541 4976
rect 35499 4927 35541 4936
rect 35595 4976 35637 4985
rect 35595 4936 35596 4976
rect 35636 4936 35637 4976
rect 35595 4927 35637 4936
rect 36547 4976 36605 4977
rect 36547 4936 36556 4976
rect 36596 4936 36605 4976
rect 37603 4976 37661 4977
rect 36547 4935 36605 4936
rect 37083 4966 37125 4975
rect 30699 4913 30741 4922
rect 37083 4926 37084 4966
rect 37124 4926 37125 4966
rect 37603 4936 37612 4976
rect 37652 4936 37661 4976
rect 37603 4935 37661 4936
rect 38851 4976 38909 4977
rect 38851 4936 38860 4976
rect 38900 4936 38909 4976
rect 38851 4935 38909 4936
rect 40771 4976 40829 4977
rect 40771 4936 40780 4976
rect 40820 4936 40829 4976
rect 40771 4935 40829 4936
rect 37083 4917 37125 4926
rect 39523 4934 39581 4935
rect 18027 4852 18028 4892
rect 18068 4852 18069 4892
rect 18027 4843 18069 4852
rect 18787 4892 18845 4893
rect 18787 4852 18796 4892
rect 18836 4852 18845 4892
rect 18787 4851 18845 4852
rect 23491 4892 23549 4893
rect 23491 4852 23500 4892
rect 23540 4852 23549 4892
rect 25371 4885 25413 4894
rect 27427 4892 27485 4893
rect 23491 4851 23549 4852
rect 27427 4852 27436 4892
rect 27476 4852 27485 4892
rect 27427 4851 27485 4852
rect 29643 4892 29685 4901
rect 29643 4852 29644 4892
rect 29684 4852 29685 4892
rect 29643 4843 29685 4852
rect 33091 4892 33149 4893
rect 33091 4852 33100 4892
rect 33140 4852 33149 4892
rect 33091 4851 33149 4852
rect 35107 4892 35165 4893
rect 35107 4852 35116 4892
rect 35156 4852 35165 4892
rect 35107 4851 35165 4852
rect 35979 4892 36021 4901
rect 35979 4852 35980 4892
rect 36020 4852 36021 4892
rect 35979 4843 36021 4852
rect 36075 4892 36117 4901
rect 39523 4894 39532 4934
rect 39572 4894 39581 4934
rect 39523 4893 39581 4894
rect 36075 4852 36076 4892
rect 36116 4852 36117 4892
rect 36075 4843 36117 4852
rect 39139 4892 39197 4893
rect 39139 4852 39148 4892
rect 39188 4852 39197 4892
rect 39139 4851 39197 4852
rect 41155 4892 41213 4893
rect 41155 4852 41164 4892
rect 41204 4852 41213 4892
rect 41155 4851 41213 4852
rect 41731 4892 41789 4893
rect 41731 4852 41740 4892
rect 41780 4852 41789 4892
rect 41731 4851 41789 4852
rect 9955 4808 10013 4809
rect 9955 4768 9964 4808
rect 10004 4768 10013 4808
rect 9955 4767 10013 4768
rect 18987 4808 19029 4817
rect 18987 4768 18988 4808
rect 19028 4768 19029 4808
rect 18987 4759 19029 4768
rect 23307 4808 23349 4817
rect 23307 4768 23308 4808
rect 23348 4768 23349 4808
rect 23307 4759 23349 4768
rect 25707 4808 25749 4817
rect 25707 4768 25708 4808
rect 25748 4768 25749 4808
rect 25707 4759 25749 4768
rect 34923 4808 34965 4817
rect 34923 4768 34924 4808
rect 34964 4768 34965 4808
rect 34923 4759 34965 4768
rect 39339 4808 39381 4817
rect 39339 4768 39340 4808
rect 39380 4768 39381 4808
rect 39339 4759 39381 4768
rect 41355 4808 41397 4817
rect 41355 4768 41356 4808
rect 41396 4768 41397 4808
rect 41355 4759 41397 4768
rect 6603 4724 6645 4733
rect 6603 4684 6604 4724
rect 6644 4684 6645 4724
rect 6603 4675 6645 4684
rect 6795 4724 6837 4733
rect 6795 4684 6796 4724
rect 6836 4684 6837 4724
rect 6795 4675 6837 4684
rect 23115 4724 23157 4733
rect 23115 4684 23116 4724
rect 23156 4684 23157 4724
rect 23115 4675 23157 4684
rect 27627 4724 27669 4733
rect 27627 4684 27628 4724
rect 27668 4684 27669 4724
rect 27627 4675 27669 4684
rect 32715 4724 32757 4733
rect 32715 4684 32716 4724
rect 32756 4684 32757 4724
rect 32715 4675 32757 4684
rect 32907 4724 32949 4733
rect 32907 4684 32908 4724
rect 32948 4684 32949 4724
rect 32907 4675 32949 4684
rect 34731 4724 34773 4733
rect 34731 4684 34732 4724
rect 34772 4684 34773 4724
rect 34731 4675 34773 4684
rect 41547 4724 41589 4733
rect 41547 4684 41548 4724
rect 41588 4684 41589 4724
rect 41547 4675 41589 4684
rect 1152 4556 41856 4580
rect 1152 4516 3688 4556
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 4056 4516 18808 4556
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 19176 4516 33928 4556
rect 33968 4516 34010 4556
rect 34050 4516 34092 4556
rect 34132 4516 34174 4556
rect 34214 4516 34256 4556
rect 34296 4516 41856 4556
rect 1152 4492 41856 4516
rect 2763 4388 2805 4397
rect 2763 4348 2764 4388
rect 2804 4348 2805 4388
rect 2763 4339 2805 4348
rect 4875 4388 4917 4397
rect 4875 4348 4876 4388
rect 4916 4348 4917 4388
rect 4875 4339 4917 4348
rect 5259 4388 5301 4397
rect 5259 4348 5260 4388
rect 5300 4348 5301 4388
rect 5259 4339 5301 4348
rect 6883 4388 6941 4389
rect 6883 4348 6892 4388
rect 6932 4348 6941 4388
rect 6883 4347 6941 4348
rect 7843 4388 7901 4389
rect 7843 4348 7852 4388
rect 7892 4348 7901 4388
rect 7843 4347 7901 4348
rect 8803 4388 8861 4389
rect 8803 4348 8812 4388
rect 8852 4348 8861 4388
rect 8803 4347 8861 4348
rect 8995 4388 9053 4389
rect 8995 4348 9004 4388
rect 9044 4348 9053 4388
rect 8995 4347 9053 4348
rect 13611 4388 13653 4397
rect 13611 4348 13612 4388
rect 13652 4348 13653 4388
rect 13611 4339 13653 4348
rect 16491 4388 16533 4397
rect 16491 4348 16492 4388
rect 16532 4348 16533 4388
rect 16491 4339 16533 4348
rect 17067 4388 17109 4397
rect 17067 4348 17068 4388
rect 17108 4348 17109 4388
rect 17067 4339 17109 4348
rect 18891 4388 18933 4397
rect 18891 4348 18892 4388
rect 18932 4348 18933 4388
rect 18891 4339 18933 4348
rect 28587 4388 28629 4397
rect 28587 4348 28588 4388
rect 28628 4348 28629 4388
rect 28587 4339 28629 4348
rect 30411 4388 30453 4397
rect 30411 4348 30412 4388
rect 30452 4348 30453 4388
rect 30411 4339 30453 4348
rect 41547 4388 41589 4397
rect 41547 4348 41548 4388
rect 41588 4348 41589 4388
rect 41547 4339 41589 4348
rect 14667 4220 14709 4229
rect 14667 4180 14668 4220
rect 14708 4180 14709 4220
rect 14667 4171 14709 4180
rect 14763 4220 14805 4229
rect 14763 4180 14764 4220
rect 14804 4180 14805 4220
rect 14763 4171 14805 4180
rect 16291 4220 16349 4221
rect 16291 4180 16300 4220
rect 16340 4180 16349 4220
rect 16291 4179 16349 4180
rect 17251 4220 17309 4221
rect 17251 4180 17260 4220
rect 17300 4180 17309 4220
rect 17251 4179 17309 4180
rect 20235 4220 20277 4229
rect 20235 4180 20236 4220
rect 20276 4180 20277 4220
rect 20235 4171 20277 4180
rect 20331 4220 20373 4229
rect 20331 4180 20332 4220
rect 20372 4180 20373 4220
rect 20331 4171 20373 4180
rect 21867 4220 21909 4229
rect 21867 4180 21868 4220
rect 21908 4180 21909 4220
rect 21867 4171 21909 4180
rect 21963 4220 22005 4229
rect 21963 4180 21964 4220
rect 22004 4180 22005 4220
rect 25131 4220 25173 4229
rect 21963 4171 22005 4180
rect 22971 4178 23013 4187
rect 15723 4150 15765 4159
rect 1315 4136 1373 4137
rect 1315 4096 1324 4136
rect 1364 4096 1373 4136
rect 1315 4095 1373 4096
rect 2563 4136 2621 4137
rect 2563 4096 2572 4136
rect 2612 4096 2621 4136
rect 2563 4095 2621 4096
rect 2955 4136 2997 4145
rect 2955 4096 2956 4136
rect 2996 4096 2997 4136
rect 2955 4087 2997 4096
rect 3051 4136 3093 4145
rect 3051 4096 3052 4136
rect 3092 4096 3093 4136
rect 3051 4087 3093 4096
rect 3147 4136 3189 4145
rect 3147 4096 3148 4136
rect 3188 4096 3189 4136
rect 3147 4087 3189 4096
rect 3427 4136 3485 4137
rect 3427 4096 3436 4136
rect 3476 4096 3485 4136
rect 3427 4095 3485 4096
rect 4675 4136 4733 4137
rect 4675 4096 4684 4136
rect 4724 4096 4733 4136
rect 4675 4095 4733 4096
rect 5059 4136 5117 4137
rect 5059 4096 5068 4136
rect 5108 4096 5117 4136
rect 5059 4095 5117 4096
rect 5259 4136 5301 4145
rect 5259 4096 5260 4136
rect 5300 4096 5301 4136
rect 5259 4087 5301 4096
rect 5347 4136 5405 4137
rect 5347 4096 5356 4136
rect 5396 4096 5405 4136
rect 5347 4095 5405 4096
rect 5539 4136 5597 4137
rect 5539 4096 5548 4136
rect 5588 4096 5597 4136
rect 5539 4095 5597 4096
rect 5643 4136 5685 4145
rect 5643 4096 5644 4136
rect 5684 4096 5685 4136
rect 5643 4087 5685 4096
rect 5835 4136 5877 4145
rect 5835 4096 5836 4136
rect 5876 4096 5877 4136
rect 5835 4087 5877 4096
rect 6211 4136 6269 4137
rect 6211 4096 6220 4136
rect 6260 4096 6269 4136
rect 6211 4095 6269 4096
rect 6507 4136 6549 4145
rect 6507 4096 6508 4136
rect 6548 4096 6549 4136
rect 6507 4087 6549 4096
rect 6603 4136 6645 4145
rect 6603 4096 6604 4136
rect 6644 4096 6645 4136
rect 6603 4087 6645 4096
rect 7171 4136 7229 4137
rect 7171 4096 7180 4136
rect 7220 4096 7229 4136
rect 7171 4095 7229 4096
rect 7467 4136 7509 4145
rect 7467 4096 7468 4136
rect 7508 4096 7509 4136
rect 7467 4087 7509 4096
rect 7563 4136 7605 4145
rect 7563 4096 7564 4136
rect 7604 4096 7605 4136
rect 7563 4087 7605 4096
rect 8131 4136 8189 4137
rect 8131 4096 8140 4136
rect 8180 4096 8189 4136
rect 8131 4095 8189 4096
rect 8427 4136 8469 4145
rect 8427 4096 8428 4136
rect 8468 4096 8469 4136
rect 8427 4087 8469 4096
rect 8523 4136 8565 4145
rect 8523 4096 8524 4136
rect 8564 4096 8565 4136
rect 8523 4087 8565 4096
rect 9387 4136 9429 4145
rect 9387 4096 9388 4136
rect 9428 4096 9429 4136
rect 9387 4087 9429 4096
rect 9667 4136 9725 4137
rect 9667 4096 9676 4136
rect 9716 4096 9725 4136
rect 9667 4095 9725 4096
rect 10059 4136 10101 4145
rect 10059 4096 10060 4136
rect 10100 4096 10101 4136
rect 10059 4087 10101 4096
rect 10347 4136 10389 4145
rect 10347 4096 10348 4136
rect 10388 4096 10389 4136
rect 10347 4087 10389 4096
rect 10531 4136 10589 4137
rect 10531 4096 10540 4136
rect 10580 4096 10589 4136
rect 10531 4095 10589 4096
rect 11779 4136 11837 4137
rect 11779 4096 11788 4136
rect 11828 4096 11837 4136
rect 11779 4095 11837 4096
rect 12163 4136 12221 4137
rect 12163 4096 12172 4136
rect 12212 4096 12221 4136
rect 12163 4095 12221 4096
rect 13411 4136 13469 4137
rect 13411 4096 13420 4136
rect 13460 4096 13469 4136
rect 13411 4095 13469 4096
rect 14187 4136 14229 4145
rect 14187 4096 14188 4136
rect 14228 4096 14229 4136
rect 14187 4087 14229 4096
rect 14283 4136 14325 4145
rect 14283 4096 14284 4136
rect 14324 4096 14325 4136
rect 14283 4087 14325 4096
rect 15235 4136 15293 4137
rect 15235 4096 15244 4136
rect 15284 4096 15293 4136
rect 15723 4110 15724 4150
rect 15764 4110 15765 4150
rect 19275 4141 19317 4150
rect 15723 4101 15765 4110
rect 17443 4136 17501 4137
rect 15235 4095 15293 4096
rect 17443 4096 17452 4136
rect 17492 4096 17501 4136
rect 17443 4095 17501 4096
rect 18691 4136 18749 4137
rect 18691 4096 18700 4136
rect 18740 4096 18749 4136
rect 18691 4095 18749 4096
rect 19275 4101 19276 4141
rect 19316 4101 19317 4141
rect 19275 4092 19317 4101
rect 19747 4136 19805 4137
rect 19747 4096 19756 4136
rect 19796 4096 19805 4136
rect 19747 4095 19805 4096
rect 20715 4136 20757 4145
rect 20715 4096 20716 4136
rect 20756 4096 20757 4136
rect 20715 4087 20757 4096
rect 20811 4136 20853 4145
rect 20811 4096 20812 4136
rect 20852 4096 20853 4136
rect 20811 4087 20853 4096
rect 21387 4136 21429 4145
rect 21387 4096 21388 4136
rect 21428 4096 21429 4136
rect 21387 4087 21429 4096
rect 21483 4136 21525 4145
rect 22971 4138 22972 4178
rect 23012 4138 23013 4178
rect 25131 4180 25132 4220
rect 25172 4180 25173 4220
rect 25131 4171 25173 4180
rect 27147 4220 27189 4229
rect 27147 4180 27148 4220
rect 27188 4180 27189 4220
rect 27147 4171 27189 4180
rect 27243 4220 27285 4229
rect 27243 4180 27244 4220
rect 27284 4180 27285 4220
rect 27243 4171 27285 4180
rect 30211 4220 30269 4221
rect 30211 4180 30220 4220
rect 30260 4180 30269 4220
rect 30211 4179 30269 4180
rect 31275 4220 31317 4229
rect 31275 4180 31276 4220
rect 31316 4180 31317 4220
rect 31275 4171 31317 4180
rect 33291 4220 33333 4229
rect 33291 4180 33292 4220
rect 33332 4180 33333 4220
rect 36459 4220 36501 4229
rect 33291 4171 33333 4180
rect 34299 4178 34341 4187
rect 21483 4096 21484 4136
rect 21524 4096 21525 4136
rect 21483 4087 21525 4096
rect 22435 4136 22493 4137
rect 22435 4096 22444 4136
rect 22484 4096 22493 4136
rect 22971 4129 23013 4138
rect 24555 4136 24597 4145
rect 22435 4095 22493 4096
rect 24555 4096 24556 4136
rect 24596 4096 24597 4136
rect 24555 4087 24597 4096
rect 24651 4136 24693 4145
rect 24651 4096 24652 4136
rect 24692 4096 24693 4136
rect 24651 4087 24693 4096
rect 25035 4136 25077 4145
rect 26091 4141 26133 4150
rect 25035 4096 25036 4136
rect 25076 4096 25077 4136
rect 25035 4087 25077 4096
rect 25603 4136 25661 4137
rect 25603 4096 25612 4136
rect 25652 4096 25661 4136
rect 25603 4095 25661 4096
rect 26091 4101 26092 4141
rect 26132 4101 26133 4141
rect 26091 4092 26133 4101
rect 26667 4136 26709 4145
rect 26667 4096 26668 4136
rect 26708 4096 26709 4136
rect 26667 4087 26709 4096
rect 26763 4136 26805 4145
rect 28203 4141 28245 4150
rect 26763 4096 26764 4136
rect 26804 4096 26805 4136
rect 26763 4087 26805 4096
rect 27715 4136 27773 4137
rect 27715 4096 27724 4136
rect 27764 4096 27773 4136
rect 27715 4095 27773 4096
rect 28203 4101 28204 4141
rect 28244 4101 28245 4141
rect 28203 4092 28245 4101
rect 28771 4136 28829 4137
rect 28771 4096 28780 4136
rect 28820 4096 28829 4136
rect 28771 4095 28829 4096
rect 30019 4136 30077 4137
rect 30019 4096 30028 4136
rect 30068 4096 30077 4136
rect 30019 4095 30077 4096
rect 30699 4136 30741 4145
rect 30699 4096 30700 4136
rect 30740 4096 30741 4136
rect 30699 4087 30741 4096
rect 30795 4136 30837 4145
rect 30795 4096 30796 4136
rect 30836 4096 30837 4136
rect 30795 4087 30837 4096
rect 31179 4136 31221 4145
rect 32235 4141 32277 4150
rect 31179 4096 31180 4136
rect 31220 4096 31221 4136
rect 31179 4087 31221 4096
rect 31747 4136 31805 4137
rect 31747 4096 31756 4136
rect 31796 4096 31805 4136
rect 31747 4095 31805 4096
rect 32235 4101 32236 4141
rect 32276 4101 32277 4141
rect 32235 4092 32277 4101
rect 32715 4136 32757 4145
rect 32715 4096 32716 4136
rect 32756 4096 32757 4136
rect 32715 4087 32757 4096
rect 32811 4136 32853 4145
rect 32811 4096 32812 4136
rect 32852 4096 32853 4136
rect 32811 4087 32853 4096
rect 33195 4136 33237 4145
rect 34299 4138 34300 4178
rect 34340 4138 34341 4178
rect 36459 4180 36460 4220
rect 36500 4180 36501 4220
rect 36459 4171 36501 4180
rect 36555 4220 36597 4229
rect 36555 4180 36556 4220
rect 36596 4180 36597 4220
rect 36555 4171 36597 4180
rect 38083 4220 38141 4221
rect 38083 4180 38092 4220
rect 38132 4180 38141 4220
rect 38083 4179 38141 4180
rect 38275 4220 38333 4221
rect 38275 4180 38284 4220
rect 38324 4180 38333 4220
rect 38275 4179 38333 4180
rect 39531 4220 39573 4229
rect 39531 4180 39532 4220
rect 39572 4180 39573 4220
rect 39531 4171 39573 4180
rect 39627 4220 39669 4229
rect 39627 4180 39628 4220
rect 39668 4180 39669 4220
rect 39627 4171 39669 4180
rect 40963 4220 41021 4221
rect 40963 4180 40972 4220
rect 41012 4180 41021 4220
rect 40963 4179 41021 4180
rect 41347 4220 41405 4221
rect 41347 4180 41356 4220
rect 41396 4180 41405 4220
rect 41347 4179 41405 4180
rect 37563 4145 37605 4154
rect 33195 4096 33196 4136
rect 33236 4096 33237 4136
rect 33195 4087 33237 4096
rect 33763 4136 33821 4137
rect 33763 4096 33772 4136
rect 33812 4096 33821 4136
rect 34299 4129 34341 4138
rect 35587 4136 35645 4137
rect 33763 4095 33821 4096
rect 35587 4096 35596 4136
rect 35636 4096 35645 4136
rect 35587 4095 35645 4096
rect 35979 4136 36021 4145
rect 35979 4096 35980 4136
rect 36020 4096 36021 4136
rect 35979 4087 36021 4096
rect 36075 4136 36117 4145
rect 36075 4096 36076 4136
rect 36116 4096 36117 4136
rect 36075 4087 36117 4096
rect 37027 4136 37085 4137
rect 37027 4096 37036 4136
rect 37076 4096 37085 4136
rect 37563 4105 37564 4145
rect 37604 4105 37605 4145
rect 37563 4096 37605 4105
rect 39051 4136 39093 4145
rect 39051 4096 39052 4136
rect 39092 4096 39093 4136
rect 37027 4095 37085 4096
rect 39051 4087 39093 4096
rect 39147 4136 39189 4145
rect 40587 4141 40629 4150
rect 39147 4096 39148 4136
rect 39188 4096 39189 4136
rect 39147 4087 39189 4096
rect 40099 4136 40157 4137
rect 40099 4096 40108 4136
rect 40148 4096 40157 4136
rect 40099 4095 40157 4096
rect 40587 4101 40588 4141
rect 40628 4101 40629 4141
rect 40587 4092 40629 4101
rect 9291 4052 9333 4061
rect 9291 4012 9292 4052
rect 9332 4012 9333 4052
rect 9291 4003 9333 4012
rect 19083 4052 19125 4061
rect 19083 4012 19084 4052
rect 19124 4012 19125 4052
rect 19083 4003 19125 4012
rect 23115 4052 23157 4061
rect 23115 4012 23116 4052
rect 23156 4012 23157 4052
rect 23115 4003 23157 4012
rect 32427 4052 32469 4061
rect 32427 4012 32428 4052
rect 32468 4012 32469 4052
rect 32427 4003 32469 4012
rect 34443 4052 34485 4061
rect 34443 4012 34444 4052
rect 34484 4012 34485 4052
rect 34443 4003 34485 4012
rect 40779 4052 40821 4061
rect 40779 4012 40780 4052
rect 40820 4012 40821 4052
rect 40779 4003 40821 4012
rect 3235 3968 3293 3969
rect 3235 3928 3244 3968
rect 3284 3928 3293 3968
rect 3235 3927 3293 3928
rect 5731 3968 5789 3969
rect 5731 3928 5740 3968
rect 5780 3928 5789 3968
rect 5731 3927 5789 3928
rect 10251 3968 10293 3977
rect 10251 3928 10252 3968
rect 10292 3928 10293 3968
rect 10251 3919 10293 3928
rect 11979 3968 12021 3977
rect 11979 3928 11980 3968
rect 12020 3928 12021 3968
rect 11979 3919 12021 3928
rect 15915 3968 15957 3977
rect 15915 3928 15916 3968
rect 15956 3928 15957 3968
rect 15915 3919 15957 3928
rect 26283 3968 26325 3977
rect 26283 3928 26284 3968
rect 26324 3928 26325 3968
rect 26283 3919 26325 3928
rect 28395 3968 28437 3977
rect 28395 3928 28396 3968
rect 28436 3928 28437 3968
rect 28395 3919 28437 3928
rect 35115 3968 35157 3977
rect 35115 3928 35116 3968
rect 35156 3928 35157 3968
rect 35115 3919 35157 3928
rect 37707 3968 37749 3977
rect 37707 3928 37708 3968
rect 37748 3928 37749 3968
rect 37707 3919 37749 3928
rect 37899 3968 37941 3977
rect 37899 3928 37900 3968
rect 37940 3928 37941 3968
rect 37899 3919 37941 3928
rect 38475 3968 38517 3977
rect 38475 3928 38476 3968
rect 38516 3928 38517 3968
rect 38475 3919 38517 3928
rect 41163 3968 41205 3977
rect 41163 3928 41164 3968
rect 41204 3928 41205 3968
rect 41163 3919 41205 3928
rect 1152 3800 41856 3824
rect 1152 3760 4928 3800
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 5296 3760 20048 3800
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20416 3760 35168 3800
rect 35208 3760 35250 3800
rect 35290 3760 35332 3800
rect 35372 3760 35414 3800
rect 35454 3760 35496 3800
rect 35536 3760 41856 3800
rect 1152 3736 41856 3760
rect 2763 3632 2805 3641
rect 2763 3592 2764 3632
rect 2804 3592 2805 3632
rect 2763 3583 2805 3592
rect 5251 3632 5309 3633
rect 5251 3592 5260 3632
rect 5300 3592 5309 3632
rect 5251 3591 5309 3592
rect 8331 3632 8373 3641
rect 8331 3592 8332 3632
rect 8372 3592 8373 3632
rect 8331 3583 8373 3592
rect 8907 3632 8949 3641
rect 8907 3592 8908 3632
rect 8948 3592 8949 3632
rect 8907 3583 8949 3592
rect 12355 3632 12413 3633
rect 12355 3592 12364 3632
rect 12404 3592 12413 3632
rect 12355 3591 12413 3592
rect 13995 3632 14037 3641
rect 13995 3592 13996 3632
rect 14036 3592 14037 3632
rect 13995 3583 14037 3592
rect 14187 3632 14229 3641
rect 14187 3592 14188 3632
rect 14228 3592 14229 3632
rect 14187 3583 14229 3592
rect 16203 3632 16245 3641
rect 16203 3592 16204 3632
rect 16244 3592 16245 3632
rect 16203 3583 16245 3592
rect 16395 3632 16437 3641
rect 16395 3592 16396 3632
rect 16436 3592 16437 3632
rect 16395 3583 16437 3592
rect 16779 3632 16821 3641
rect 16779 3592 16780 3632
rect 16820 3592 16821 3632
rect 16779 3583 16821 3592
rect 19851 3632 19893 3641
rect 19851 3592 19852 3632
rect 19892 3592 19893 3632
rect 19851 3583 19893 3592
rect 21483 3632 21525 3641
rect 21483 3592 21484 3632
rect 21524 3592 21525 3632
rect 21483 3583 21525 3592
rect 21675 3632 21717 3641
rect 21675 3592 21676 3632
rect 21716 3592 21717 3632
rect 21675 3583 21717 3592
rect 23979 3632 24021 3641
rect 23979 3592 23980 3632
rect 24020 3592 24021 3632
rect 23979 3583 24021 3592
rect 26955 3632 26997 3641
rect 26955 3592 26956 3632
rect 26996 3592 26997 3632
rect 26955 3583 26997 3592
rect 28587 3632 28629 3641
rect 28587 3592 28588 3632
rect 28628 3592 28629 3632
rect 28587 3583 28629 3592
rect 28779 3632 28821 3641
rect 28779 3592 28780 3632
rect 28820 3592 28821 3632
rect 28779 3583 28821 3592
rect 30411 3632 30453 3641
rect 30411 3592 30412 3632
rect 30452 3592 30453 3632
rect 30411 3583 30453 3592
rect 32043 3632 32085 3641
rect 32043 3592 32044 3632
rect 32084 3592 32085 3632
rect 32043 3583 32085 3592
rect 33675 3632 33717 3641
rect 33675 3592 33676 3632
rect 33716 3592 33717 3632
rect 33675 3583 33717 3592
rect 35691 3632 35733 3641
rect 35691 3592 35692 3632
rect 35732 3592 35733 3632
rect 35691 3583 35733 3592
rect 37611 3632 37653 3641
rect 37611 3592 37612 3632
rect 37652 3592 37653 3632
rect 37611 3583 37653 3592
rect 39723 3632 39765 3641
rect 39723 3592 39724 3632
rect 39764 3592 39765 3632
rect 39723 3583 39765 3592
rect 39915 3632 39957 3641
rect 39915 3592 39916 3632
rect 39956 3592 39957 3632
rect 39915 3583 39957 3592
rect 4395 3548 4437 3557
rect 4395 3508 4396 3548
rect 4436 3508 4437 3548
rect 4395 3499 4437 3508
rect 4683 3548 4725 3557
rect 4683 3508 4684 3548
rect 4724 3508 4725 3548
rect 4683 3499 4725 3508
rect 7371 3548 7413 3557
rect 7371 3508 7372 3548
rect 7412 3508 7413 3548
rect 7371 3499 7413 3508
rect 10923 3548 10965 3557
rect 10923 3508 10924 3548
rect 10964 3508 10965 3548
rect 10923 3499 10965 3508
rect 10242 3473 10300 3474
rect 1315 3464 1373 3465
rect 1315 3424 1324 3464
rect 1364 3424 1373 3464
rect 1315 3423 1373 3424
rect 2563 3464 2621 3465
rect 2563 3424 2572 3464
rect 2612 3424 2621 3464
rect 2563 3423 2621 3424
rect 2947 3464 3005 3465
rect 2947 3424 2956 3464
rect 2996 3424 3005 3464
rect 2947 3423 3005 3424
rect 4195 3464 4253 3465
rect 4195 3424 4204 3464
rect 4244 3424 4253 3464
rect 4195 3423 4253 3424
rect 4579 3464 4637 3465
rect 4579 3424 4588 3464
rect 4628 3424 4637 3464
rect 4579 3423 4637 3424
rect 4779 3464 4821 3473
rect 4779 3424 4780 3464
rect 4820 3424 4821 3464
rect 4779 3415 4821 3424
rect 4971 3464 5013 3473
rect 4971 3424 4972 3464
rect 5012 3424 5013 3464
rect 4971 3415 5013 3424
rect 5067 3464 5109 3473
rect 5067 3424 5068 3464
rect 5108 3424 5109 3464
rect 5067 3415 5109 3424
rect 5547 3464 5589 3473
rect 5547 3424 5548 3464
rect 5588 3424 5589 3464
rect 5547 3415 5589 3424
rect 5931 3464 5973 3473
rect 5931 3424 5932 3464
rect 5972 3424 5973 3464
rect 5931 3415 5973 3424
rect 6123 3464 6165 3473
rect 6123 3424 6124 3464
rect 6164 3424 6165 3464
rect 6123 3415 6165 3424
rect 6211 3464 6269 3465
rect 6211 3424 6220 3464
rect 6260 3424 6269 3464
rect 6211 3423 6269 3424
rect 6411 3464 6453 3473
rect 6411 3424 6412 3464
rect 6452 3424 6453 3464
rect 6411 3415 6453 3424
rect 6699 3464 6741 3473
rect 6699 3424 6700 3464
rect 6740 3424 6741 3464
rect 6699 3415 6741 3424
rect 6979 3464 7037 3465
rect 6979 3424 6988 3464
rect 7028 3424 7037 3464
rect 6979 3423 7037 3424
rect 7275 3464 7317 3473
rect 7275 3424 7276 3464
rect 7316 3424 7317 3464
rect 7275 3415 7317 3424
rect 7851 3464 7893 3473
rect 7851 3424 7852 3464
rect 7892 3424 7893 3464
rect 7851 3415 7893 3424
rect 7947 3464 7989 3473
rect 7947 3424 7948 3464
rect 7988 3424 7989 3464
rect 7947 3415 7989 3424
rect 8043 3464 8085 3473
rect 8043 3424 8044 3464
rect 8084 3424 8085 3464
rect 8043 3415 8085 3424
rect 8139 3464 8181 3473
rect 8139 3424 8140 3464
rect 8180 3424 8181 3464
rect 8139 3415 8181 3424
rect 8323 3464 8381 3465
rect 8323 3424 8332 3464
rect 8372 3424 8381 3464
rect 8323 3423 8381 3424
rect 8523 3464 8565 3473
rect 8523 3424 8524 3464
rect 8564 3424 8565 3464
rect 8523 3415 8565 3424
rect 8611 3464 8669 3465
rect 8611 3424 8620 3464
rect 8660 3424 8669 3464
rect 8611 3423 8669 3424
rect 8803 3464 8861 3465
rect 8803 3424 8812 3464
rect 8852 3424 8861 3464
rect 8803 3423 8861 3424
rect 9195 3464 9237 3473
rect 9195 3424 9196 3464
rect 9236 3424 9237 3464
rect 9195 3415 9237 3424
rect 9291 3464 9333 3473
rect 9291 3424 9292 3464
rect 9332 3424 9333 3464
rect 10242 3433 10251 3473
rect 10291 3433 10300 3473
rect 11203 3464 11261 3465
rect 10242 3432 10300 3433
rect 10731 3450 10773 3459
rect 9291 3415 9333 3424
rect 10731 3410 10732 3450
rect 10772 3410 10773 3450
rect 11203 3424 11212 3464
rect 11252 3424 11261 3464
rect 11203 3423 11261 3424
rect 11499 3464 11541 3473
rect 11499 3424 11500 3464
rect 11540 3424 11541 3464
rect 11499 3415 11541 3424
rect 11595 3464 11637 3473
rect 11595 3424 11596 3464
rect 11636 3424 11637 3464
rect 11595 3415 11637 3424
rect 12075 3464 12117 3473
rect 12075 3424 12076 3464
rect 12116 3424 12117 3464
rect 12075 3415 12117 3424
rect 12171 3464 12213 3473
rect 12171 3424 12172 3464
rect 12212 3424 12213 3464
rect 12171 3415 12213 3424
rect 12547 3464 12605 3465
rect 12547 3424 12556 3464
rect 12596 3424 12605 3464
rect 12547 3423 12605 3424
rect 14755 3464 14813 3465
rect 14755 3424 14764 3464
rect 14804 3424 14813 3464
rect 14755 3423 14813 3424
rect 16003 3464 16061 3465
rect 16003 3424 16012 3464
rect 16052 3424 16061 3464
rect 16003 3423 16061 3424
rect 16963 3464 17021 3465
rect 16963 3424 16972 3464
rect 17012 3424 17021 3464
rect 16963 3423 17021 3424
rect 18211 3464 18269 3465
rect 18211 3424 18220 3464
rect 18260 3424 18269 3464
rect 18211 3423 18269 3424
rect 18403 3464 18461 3465
rect 18403 3424 18412 3464
rect 18452 3424 18461 3464
rect 18403 3423 18461 3424
rect 19651 3464 19709 3465
rect 19651 3424 19660 3464
rect 19700 3424 19709 3464
rect 19651 3423 19709 3424
rect 20035 3464 20093 3465
rect 20035 3424 20044 3464
rect 20084 3424 20093 3464
rect 20035 3423 20093 3424
rect 21283 3464 21341 3465
rect 21283 3424 21292 3464
rect 21332 3424 21341 3464
rect 21283 3423 21341 3424
rect 22531 3464 22589 3465
rect 22531 3424 22540 3464
rect 22580 3424 22589 3464
rect 22531 3423 22589 3424
rect 23779 3464 23837 3465
rect 23779 3424 23788 3464
rect 23828 3424 23837 3464
rect 23779 3423 23837 3424
rect 25507 3464 25565 3465
rect 25507 3424 25516 3464
rect 25556 3424 25565 3464
rect 25507 3423 25565 3424
rect 26755 3464 26813 3465
rect 26755 3424 26764 3464
rect 26804 3424 26813 3464
rect 26755 3423 26813 3424
rect 27139 3464 27197 3465
rect 27139 3424 27148 3464
rect 27188 3424 27197 3464
rect 27139 3423 27197 3424
rect 28387 3464 28445 3465
rect 28387 3424 28396 3464
rect 28436 3424 28445 3464
rect 28387 3423 28445 3424
rect 28963 3464 29021 3465
rect 28963 3424 28972 3464
rect 29012 3424 29021 3464
rect 28963 3423 29021 3424
rect 30211 3464 30269 3465
rect 30211 3424 30220 3464
rect 30260 3424 30269 3464
rect 30211 3423 30269 3424
rect 30595 3464 30653 3465
rect 30595 3424 30604 3464
rect 30644 3424 30653 3464
rect 30595 3423 30653 3424
rect 31843 3464 31901 3465
rect 31843 3424 31852 3464
rect 31892 3424 31901 3464
rect 31843 3423 31901 3424
rect 32227 3464 32285 3465
rect 32227 3424 32236 3464
rect 32276 3424 32285 3464
rect 32227 3423 32285 3424
rect 33475 3464 33533 3465
rect 33475 3424 33484 3464
rect 33524 3424 33533 3464
rect 33475 3423 33533 3424
rect 34243 3464 34301 3465
rect 34243 3424 34252 3464
rect 34292 3424 34301 3464
rect 34243 3423 34301 3424
rect 35491 3464 35549 3465
rect 35491 3424 35500 3464
rect 35540 3424 35549 3464
rect 35491 3423 35549 3424
rect 36163 3464 36221 3465
rect 36163 3424 36172 3464
rect 36212 3424 36221 3464
rect 36163 3423 36221 3424
rect 37411 3464 37469 3465
rect 37411 3424 37420 3464
rect 37460 3424 37469 3464
rect 37411 3423 37469 3424
rect 38275 3464 38333 3465
rect 38275 3424 38284 3464
rect 38324 3424 38333 3464
rect 38275 3423 38333 3424
rect 39523 3464 39581 3465
rect 39523 3424 39532 3464
rect 39572 3424 39581 3464
rect 39523 3423 39581 3424
rect 40099 3464 40157 3465
rect 40099 3424 40108 3464
rect 40148 3424 40157 3464
rect 40099 3423 40157 3424
rect 41347 3464 41405 3465
rect 41347 3424 41356 3464
rect 41396 3424 41405 3464
rect 41347 3423 41405 3424
rect 13795 3422 13853 3423
rect 10731 3401 10773 3410
rect 9675 3380 9717 3389
rect 9675 3340 9676 3380
rect 9716 3340 9717 3380
rect 9675 3331 9717 3340
rect 9771 3380 9813 3389
rect 13795 3382 13804 3422
rect 13844 3382 13853 3422
rect 13795 3381 13853 3382
rect 9771 3340 9772 3380
rect 9812 3340 9813 3380
rect 9771 3331 9813 3340
rect 14371 3380 14429 3381
rect 14371 3340 14380 3380
rect 14420 3340 14429 3380
rect 14371 3339 14429 3340
rect 16579 3380 16637 3381
rect 16579 3340 16588 3380
rect 16628 3340 16637 3380
rect 16579 3339 16637 3340
rect 21859 3380 21917 3381
rect 21859 3340 21868 3380
rect 21908 3340 21917 3380
rect 21859 3339 21917 3340
rect 24355 3380 24413 3381
rect 24355 3340 24364 3380
rect 24404 3340 24413 3380
rect 24355 3339 24413 3340
rect 24739 3380 24797 3381
rect 24739 3340 24748 3380
rect 24788 3340 24797 3380
rect 24739 3339 24797 3340
rect 25123 3380 25181 3381
rect 25123 3340 25132 3380
rect 25172 3340 25181 3380
rect 25123 3339 25181 3340
rect 33859 3380 33917 3381
rect 33859 3340 33868 3380
rect 33908 3340 33917 3380
rect 33859 3339 33917 3340
rect 38083 3380 38141 3381
rect 38083 3340 38092 3380
rect 38132 3340 38141 3380
rect 38083 3339 38141 3340
rect 5547 3296 5589 3305
rect 5547 3256 5548 3296
rect 5588 3256 5589 3296
rect 5547 3247 5589 3256
rect 11875 3296 11933 3297
rect 11875 3256 11884 3296
rect 11924 3256 11933 3296
rect 11875 3255 11933 3256
rect 24939 3296 24981 3305
rect 24939 3256 24940 3296
rect 24980 3256 24981 3296
rect 24939 3247 24981 3256
rect 25323 3296 25365 3305
rect 25323 3256 25324 3296
rect 25364 3256 25365 3296
rect 25323 3247 25365 3256
rect 41547 3296 41589 3305
rect 41547 3256 41548 3296
rect 41588 3256 41589 3296
rect 41547 3247 41589 3256
rect 2763 3212 2805 3221
rect 2763 3172 2764 3212
rect 2804 3172 2805 3212
rect 2763 3163 2805 3172
rect 5739 3212 5781 3221
rect 5739 3172 5740 3212
rect 5780 3172 5781 3212
rect 5739 3163 5781 3172
rect 5931 3212 5973 3221
rect 5931 3172 5932 3212
rect 5972 3172 5973 3212
rect 5931 3163 5973 3172
rect 6699 3212 6741 3221
rect 6699 3172 6700 3212
rect 6740 3172 6741 3212
rect 6699 3163 6741 3172
rect 7651 3212 7709 3213
rect 7651 3172 7660 3212
rect 7700 3172 7709 3212
rect 7651 3171 7709 3172
rect 24555 3212 24597 3221
rect 24555 3172 24556 3212
rect 24596 3172 24597 3212
rect 24555 3163 24597 3172
rect 37899 3212 37941 3221
rect 37899 3172 37900 3212
rect 37940 3172 37941 3212
rect 37899 3163 37941 3172
rect 1152 3044 41856 3068
rect 1152 3004 3688 3044
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 4056 3004 18808 3044
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 19176 3004 33928 3044
rect 33968 3004 34010 3044
rect 34050 3004 34092 3044
rect 34132 3004 34174 3044
rect 34214 3004 34256 3044
rect 34296 3004 41856 3044
rect 1152 2980 41856 3004
rect 2955 2876 2997 2885
rect 2955 2836 2956 2876
rect 2996 2836 2997 2876
rect 2955 2827 2997 2836
rect 6219 2876 6261 2885
rect 6219 2836 6220 2876
rect 6260 2836 6261 2876
rect 6219 2827 6261 2836
rect 9963 2876 10005 2885
rect 9963 2836 9964 2876
rect 10004 2836 10005 2876
rect 9963 2827 10005 2836
rect 13899 2876 13941 2885
rect 13899 2836 13900 2876
rect 13940 2836 13941 2876
rect 13899 2827 13941 2836
rect 16299 2876 16341 2885
rect 16299 2836 16300 2876
rect 16340 2836 16341 2876
rect 16299 2827 16341 2836
rect 26667 2876 26709 2885
rect 26667 2836 26668 2876
rect 26708 2836 26709 2876
rect 26667 2827 26709 2836
rect 29547 2876 29589 2885
rect 29547 2836 29548 2876
rect 29588 2836 29589 2876
rect 29547 2827 29589 2836
rect 30027 2876 30069 2885
rect 30027 2836 30028 2876
rect 30068 2836 30069 2876
rect 30027 2827 30069 2836
rect 31659 2876 31701 2885
rect 31659 2836 31660 2876
rect 31700 2836 31701 2876
rect 31659 2827 31701 2836
rect 32043 2876 32085 2885
rect 32043 2836 32044 2876
rect 32084 2836 32085 2876
rect 32043 2827 32085 2836
rect 36363 2876 36405 2885
rect 36363 2836 36364 2876
rect 36404 2836 36405 2876
rect 36363 2827 36405 2836
rect 36939 2876 36981 2885
rect 36939 2836 36940 2876
rect 36980 2836 36981 2876
rect 36939 2827 36981 2836
rect 37603 2876 37661 2877
rect 37603 2836 37612 2876
rect 37652 2836 37661 2876
rect 37603 2835 37661 2836
rect 6019 2792 6077 2793
rect 6019 2752 6028 2792
rect 6068 2752 6077 2792
rect 6019 2751 6077 2752
rect 41643 2792 41685 2801
rect 41643 2752 41644 2792
rect 41684 2752 41685 2792
rect 41643 2743 41685 2752
rect 4299 2708 4341 2717
rect 4299 2668 4300 2708
rect 4340 2668 4341 2708
rect 4299 2659 4341 2668
rect 4395 2708 4437 2717
rect 4395 2668 4396 2708
rect 4436 2668 4437 2708
rect 7083 2708 7125 2717
rect 4395 2659 4437 2668
rect 5643 2666 5685 2675
rect 3339 2629 3381 2638
rect 1507 2624 1565 2625
rect 1507 2584 1516 2624
rect 1556 2584 1565 2624
rect 1507 2583 1565 2584
rect 2755 2624 2813 2625
rect 2755 2584 2764 2624
rect 2804 2584 2813 2624
rect 2755 2583 2813 2584
rect 3339 2589 3340 2629
rect 3380 2589 3381 2629
rect 3339 2580 3381 2589
rect 3811 2624 3869 2625
rect 3811 2584 3820 2624
rect 3860 2584 3869 2624
rect 3811 2583 3869 2584
rect 4779 2624 4821 2633
rect 4779 2584 4780 2624
rect 4820 2584 4821 2624
rect 4779 2575 4821 2584
rect 4875 2624 4917 2633
rect 5643 2626 5644 2666
rect 5684 2626 5685 2666
rect 7083 2668 7084 2708
rect 7124 2668 7125 2708
rect 7083 2659 7125 2668
rect 7179 2708 7221 2717
rect 7179 2668 7180 2708
rect 7220 2668 7221 2708
rect 7179 2659 7221 2668
rect 10827 2708 10869 2717
rect 10827 2668 10828 2708
rect 10868 2668 10869 2708
rect 10827 2659 10869 2668
rect 14667 2708 14709 2717
rect 14667 2668 14668 2708
rect 14708 2668 14709 2708
rect 14667 2659 14709 2668
rect 14763 2708 14805 2717
rect 14763 2668 14764 2708
rect 14804 2668 14805 2708
rect 14763 2659 14805 2668
rect 16099 2708 16157 2709
rect 16099 2668 16108 2708
rect 16148 2668 16157 2708
rect 16099 2667 16157 2668
rect 17067 2708 17109 2717
rect 17067 2668 17068 2708
rect 17108 2668 17109 2708
rect 17067 2659 17109 2668
rect 17163 2708 17205 2717
rect 17163 2668 17164 2708
rect 17204 2668 17205 2708
rect 17163 2659 17205 2668
rect 19179 2708 19221 2717
rect 19179 2668 19180 2708
rect 19220 2668 19221 2708
rect 19179 2659 19221 2668
rect 21195 2708 21237 2717
rect 21195 2668 21196 2708
rect 21236 2668 21237 2708
rect 21195 2659 21237 2668
rect 21291 2708 21333 2717
rect 21291 2668 21292 2708
rect 21332 2668 21333 2708
rect 21291 2659 21333 2668
rect 23787 2708 23829 2717
rect 23787 2668 23788 2708
rect 23828 2668 23829 2708
rect 23787 2659 23829 2668
rect 23883 2708 23925 2717
rect 23883 2668 23884 2708
rect 23924 2668 23925 2708
rect 23883 2659 23925 2668
rect 27043 2708 27101 2709
rect 27043 2668 27052 2708
rect 27092 2668 27101 2708
rect 27043 2667 27101 2668
rect 28011 2708 28053 2717
rect 28011 2668 28012 2708
rect 28052 2668 28053 2708
rect 28011 2659 28053 2668
rect 28107 2708 28149 2717
rect 28107 2668 28108 2708
rect 28148 2668 28149 2708
rect 28107 2659 28149 2668
rect 29731 2708 29789 2709
rect 29731 2668 29740 2708
rect 29780 2668 29789 2708
rect 29731 2667 29789 2668
rect 31843 2708 31901 2709
rect 31843 2668 31852 2708
rect 31892 2668 31901 2708
rect 31843 2667 31901 2668
rect 32227 2708 32285 2709
rect 32227 2668 32236 2708
rect 32276 2668 32285 2708
rect 32227 2667 32285 2668
rect 33291 2708 33333 2717
rect 33291 2668 33292 2708
rect 33332 2668 33333 2708
rect 33291 2659 33333 2668
rect 33387 2708 33429 2717
rect 33387 2668 33388 2708
rect 33428 2668 33429 2708
rect 33387 2659 33429 2668
rect 36547 2708 36605 2709
rect 36547 2668 36556 2708
rect 36596 2668 36605 2708
rect 36547 2667 36605 2668
rect 37123 2708 37181 2709
rect 37123 2668 37132 2708
rect 37172 2668 37181 2708
rect 37123 2667 37181 2668
rect 4875 2584 4876 2624
rect 4916 2584 4917 2624
rect 4875 2575 4917 2584
rect 5347 2624 5405 2625
rect 5347 2584 5356 2624
rect 5396 2584 5405 2624
rect 5643 2617 5685 2626
rect 5739 2624 5781 2633
rect 5347 2583 5405 2584
rect 5739 2584 5740 2624
rect 5780 2584 5781 2624
rect 5739 2575 5781 2584
rect 6307 2624 6365 2625
rect 6307 2584 6316 2624
rect 6356 2584 6365 2624
rect 6307 2583 6365 2584
rect 6603 2624 6645 2633
rect 6603 2584 6604 2624
rect 6644 2584 6645 2624
rect 6603 2575 6645 2584
rect 6699 2624 6741 2633
rect 8139 2629 8181 2638
rect 6699 2584 6700 2624
rect 6740 2584 6741 2624
rect 6699 2575 6741 2584
rect 7651 2624 7709 2625
rect 7651 2584 7660 2624
rect 7700 2584 7709 2624
rect 7651 2583 7709 2584
rect 8139 2589 8140 2629
rect 8180 2589 8181 2629
rect 8139 2580 8181 2589
rect 8515 2624 8573 2625
rect 8515 2584 8524 2624
rect 8564 2584 8573 2624
rect 8515 2583 8573 2584
rect 9763 2624 9821 2625
rect 9763 2584 9772 2624
rect 9812 2584 9821 2624
rect 9763 2583 9821 2584
rect 10251 2624 10293 2633
rect 10251 2584 10252 2624
rect 10292 2584 10293 2624
rect 10251 2575 10293 2584
rect 10347 2624 10389 2633
rect 10347 2584 10348 2624
rect 10388 2584 10389 2624
rect 10347 2575 10389 2584
rect 10731 2624 10773 2633
rect 11787 2629 11829 2638
rect 10731 2584 10732 2624
rect 10772 2584 10773 2624
rect 10731 2575 10773 2584
rect 11299 2624 11357 2625
rect 11299 2584 11308 2624
rect 11348 2584 11357 2624
rect 11299 2583 11357 2584
rect 11787 2589 11788 2629
rect 11828 2589 11829 2629
rect 11787 2580 11829 2589
rect 12259 2624 12317 2625
rect 12259 2584 12268 2624
rect 12308 2584 12317 2624
rect 12259 2583 12317 2584
rect 12451 2624 12509 2625
rect 12451 2584 12460 2624
rect 12500 2584 12509 2624
rect 12451 2583 12509 2584
rect 13699 2624 13757 2625
rect 13699 2584 13708 2624
rect 13748 2584 13757 2624
rect 13699 2583 13757 2584
rect 14187 2624 14229 2633
rect 14187 2584 14188 2624
rect 14228 2584 14229 2624
rect 14187 2575 14229 2584
rect 14283 2624 14325 2633
rect 15723 2629 15765 2638
rect 14283 2584 14284 2624
rect 14324 2584 14325 2624
rect 14283 2575 14325 2584
rect 15235 2624 15293 2625
rect 15235 2584 15244 2624
rect 15284 2584 15293 2624
rect 15235 2583 15293 2584
rect 15723 2589 15724 2629
rect 15764 2589 15765 2629
rect 15723 2580 15765 2589
rect 16587 2624 16629 2633
rect 16587 2584 16588 2624
rect 16628 2584 16629 2624
rect 16587 2575 16629 2584
rect 16683 2624 16725 2633
rect 18123 2629 18165 2638
rect 20283 2633 20325 2642
rect 22299 2633 22341 2642
rect 16683 2584 16684 2624
rect 16724 2584 16725 2624
rect 16683 2575 16725 2584
rect 17635 2624 17693 2625
rect 17635 2584 17644 2624
rect 17684 2584 17693 2624
rect 17635 2583 17693 2584
rect 18123 2589 18124 2629
rect 18164 2589 18165 2629
rect 18123 2580 18165 2589
rect 18699 2624 18741 2633
rect 18699 2584 18700 2624
rect 18740 2584 18741 2624
rect 18699 2575 18741 2584
rect 18795 2624 18837 2633
rect 18795 2584 18796 2624
rect 18836 2584 18837 2624
rect 18795 2575 18837 2584
rect 19275 2624 19317 2633
rect 19275 2584 19276 2624
rect 19316 2584 19317 2624
rect 19275 2575 19317 2584
rect 19747 2624 19805 2625
rect 19747 2584 19756 2624
rect 19796 2584 19805 2624
rect 20283 2593 20284 2633
rect 20324 2593 20325 2633
rect 20283 2584 20325 2593
rect 20715 2624 20757 2633
rect 20715 2584 20716 2624
rect 20756 2584 20757 2624
rect 19747 2583 19805 2584
rect 20715 2575 20757 2584
rect 20811 2624 20853 2633
rect 20811 2584 20812 2624
rect 20852 2584 20853 2624
rect 20811 2575 20853 2584
rect 21763 2624 21821 2625
rect 21763 2584 21772 2624
rect 21812 2584 21821 2624
rect 22299 2593 22300 2633
rect 22340 2593 22341 2633
rect 22299 2584 22341 2593
rect 23307 2624 23349 2633
rect 23307 2584 23308 2624
rect 23348 2584 23349 2624
rect 21763 2583 21821 2584
rect 23307 2575 23349 2584
rect 23403 2624 23445 2633
rect 24843 2629 24885 2638
rect 29115 2633 29157 2642
rect 34395 2633 34437 2642
rect 23403 2584 23404 2624
rect 23444 2584 23445 2624
rect 23403 2575 23445 2584
rect 24355 2624 24413 2625
rect 24355 2584 24364 2624
rect 24404 2584 24413 2624
rect 24355 2583 24413 2584
rect 24843 2589 24844 2629
rect 24884 2589 24885 2629
rect 24843 2580 24885 2589
rect 25219 2624 25277 2625
rect 25219 2584 25228 2624
rect 25268 2584 25277 2624
rect 25219 2583 25277 2584
rect 26467 2624 26525 2625
rect 26467 2584 26476 2624
rect 26516 2584 26525 2624
rect 26467 2583 26525 2584
rect 27531 2624 27573 2633
rect 27531 2584 27532 2624
rect 27572 2584 27573 2624
rect 27531 2575 27573 2584
rect 27627 2624 27669 2633
rect 27627 2584 27628 2624
rect 27668 2584 27669 2624
rect 27627 2575 27669 2584
rect 28579 2624 28637 2625
rect 28579 2584 28588 2624
rect 28628 2584 28637 2624
rect 29115 2593 29116 2633
rect 29156 2593 29157 2633
rect 29115 2584 29157 2593
rect 30211 2624 30269 2625
rect 30211 2584 30220 2624
rect 30260 2584 30269 2624
rect 28579 2583 28637 2584
rect 30211 2583 30269 2584
rect 31459 2624 31517 2625
rect 31459 2584 31468 2624
rect 31508 2584 31517 2624
rect 31459 2583 31517 2584
rect 32811 2624 32853 2633
rect 32811 2584 32812 2624
rect 32852 2584 32853 2624
rect 32811 2575 32853 2584
rect 32907 2624 32949 2633
rect 32907 2584 32908 2624
rect 32948 2584 32949 2624
rect 32907 2575 32949 2584
rect 33859 2624 33917 2625
rect 33859 2584 33868 2624
rect 33908 2584 33917 2624
rect 34395 2593 34396 2633
rect 34436 2593 34437 2633
rect 34395 2584 34437 2593
rect 34915 2624 34973 2625
rect 34915 2584 34924 2624
rect 34964 2584 34973 2624
rect 33859 2583 33917 2584
rect 34915 2583 34973 2584
rect 36163 2624 36221 2625
rect 36163 2584 36172 2624
rect 36212 2584 36221 2624
rect 36163 2583 36221 2584
rect 38755 2624 38813 2625
rect 38755 2584 38764 2624
rect 38804 2584 38813 2624
rect 38755 2583 38813 2584
rect 39619 2624 39677 2625
rect 39619 2584 39628 2624
rect 39668 2584 39677 2624
rect 39619 2583 39677 2584
rect 40011 2624 40053 2633
rect 40011 2584 40012 2624
rect 40052 2584 40053 2624
rect 40011 2575 40053 2584
rect 40195 2624 40253 2625
rect 40195 2584 40204 2624
rect 40244 2584 40253 2624
rect 40195 2583 40253 2584
rect 41443 2624 41501 2625
rect 41443 2584 41452 2624
rect 41492 2584 41501 2624
rect 41443 2583 41501 2584
rect 3147 2540 3189 2549
rect 3147 2500 3148 2540
rect 3188 2500 3189 2540
rect 3147 2491 3189 2500
rect 15915 2540 15957 2549
rect 15915 2500 15916 2540
rect 15956 2500 15957 2540
rect 15915 2491 15957 2500
rect 18315 2540 18357 2549
rect 18315 2500 18316 2540
rect 18356 2500 18357 2540
rect 18315 2491 18357 2500
rect 25035 2540 25077 2549
rect 25035 2500 25036 2540
rect 25076 2500 25077 2540
rect 25035 2491 25077 2500
rect 29259 2540 29301 2549
rect 29259 2500 29260 2540
rect 29300 2500 29301 2540
rect 29259 2491 29301 2500
rect 8331 2456 8373 2465
rect 8331 2416 8332 2456
rect 8372 2416 8373 2456
rect 8331 2407 8373 2416
rect 11979 2456 12021 2465
rect 11979 2416 11980 2456
rect 12020 2416 12021 2456
rect 11979 2407 12021 2416
rect 12171 2456 12213 2465
rect 12171 2416 12172 2456
rect 12212 2416 12213 2456
rect 22443 2456 22485 2465
rect 12171 2407 12213 2416
rect 20427 2414 20469 2423
rect 20427 2374 20428 2414
rect 20468 2374 20469 2414
rect 22443 2416 22444 2456
rect 22484 2416 22485 2456
rect 22443 2407 22485 2416
rect 27243 2456 27285 2465
rect 27243 2416 27244 2456
rect 27284 2416 27285 2456
rect 27243 2407 27285 2416
rect 34539 2456 34581 2465
rect 34539 2416 34540 2456
rect 34580 2416 34581 2456
rect 34539 2407 34581 2416
rect 36747 2456 36789 2465
rect 36747 2416 36748 2456
rect 36788 2416 36789 2456
rect 36747 2407 36789 2416
rect 20427 2365 20469 2374
rect 1152 2288 41856 2312
rect 1152 2248 4928 2288
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 5296 2248 20048 2288
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20416 2248 35168 2288
rect 35208 2248 35250 2288
rect 35290 2248 35332 2288
rect 35372 2248 35414 2288
rect 35454 2248 35496 2288
rect 35536 2248 41856 2288
rect 1152 2224 41856 2248
rect 2955 2120 2997 2129
rect 2955 2080 2956 2120
rect 2996 2080 2997 2120
rect 2955 2071 2997 2080
rect 3523 2120 3581 2121
rect 3523 2080 3532 2120
rect 3572 2080 3581 2120
rect 3523 2079 3581 2080
rect 5923 2120 5981 2121
rect 5923 2080 5932 2120
rect 5972 2080 5981 2120
rect 5923 2079 5981 2080
rect 10923 2120 10965 2129
rect 10923 2080 10924 2120
rect 10964 2080 10965 2120
rect 10923 2071 10965 2080
rect 14091 2120 14133 2129
rect 14091 2080 14092 2120
rect 14132 2080 14133 2120
rect 14091 2071 14133 2080
rect 16011 2120 16053 2129
rect 16011 2080 16012 2120
rect 16052 2080 16053 2120
rect 16011 2071 16053 2080
rect 17643 2120 17685 2129
rect 17643 2080 17644 2120
rect 17684 2080 17685 2120
rect 17643 2071 17685 2080
rect 19275 2120 19317 2129
rect 19275 2080 19276 2120
rect 19316 2080 19317 2120
rect 19275 2071 19317 2080
rect 21003 2120 21045 2129
rect 21003 2080 21004 2120
rect 21044 2080 21045 2120
rect 21003 2071 21045 2080
rect 22635 2120 22677 2129
rect 22635 2080 22636 2120
rect 22676 2080 22677 2120
rect 22635 2071 22677 2080
rect 24267 2120 24309 2129
rect 24267 2080 24268 2120
rect 24308 2080 24309 2120
rect 24267 2071 24309 2080
rect 26283 2120 26325 2129
rect 26283 2080 26284 2120
rect 26324 2080 26325 2120
rect 26283 2071 26325 2080
rect 30123 2120 30165 2129
rect 30123 2080 30124 2120
rect 30164 2080 30165 2120
rect 30123 2071 30165 2080
rect 33195 2120 33237 2129
rect 33195 2080 33196 2120
rect 33236 2080 33237 2120
rect 33195 2071 33237 2080
rect 36067 2120 36125 2121
rect 36067 2080 36076 2120
rect 36116 2080 36125 2120
rect 36067 2079 36125 2080
rect 38947 2120 39005 2121
rect 38947 2080 38956 2120
rect 38996 2080 39005 2120
rect 38947 2079 39005 2080
rect 41259 2120 41301 2129
rect 41259 2080 41260 2120
rect 41300 2080 41301 2120
rect 41259 2071 41301 2080
rect 3243 2036 3285 2045
rect 3243 1996 3244 2036
rect 3284 1996 3285 2036
rect 3243 1987 3285 1996
rect 8523 2036 8565 2045
rect 8523 1996 8524 2036
rect 8564 1996 8565 2036
rect 8523 1987 8565 1996
rect 11883 2036 11925 2045
rect 11883 1996 11884 2036
rect 11924 1996 11925 2036
rect 11883 1987 11925 1996
rect 26475 2036 26517 2045
rect 26475 1996 26476 2036
rect 26516 1996 26517 2036
rect 26475 1987 26517 1996
rect 29931 2036 29973 2045
rect 29931 1996 29932 2036
rect 29972 1996 29973 2036
rect 29931 1987 29973 1996
rect 33675 2036 33717 2045
rect 33675 1996 33676 2036
rect 33716 1996 33717 2036
rect 33675 1987 33717 1996
rect 36555 2036 36597 2045
rect 36555 1996 36556 2036
rect 36596 1996 36597 2036
rect 36555 1987 36597 1996
rect 1507 1952 1565 1953
rect 1507 1912 1516 1952
rect 1556 1912 1565 1952
rect 1507 1911 1565 1912
rect 2755 1952 2813 1953
rect 2755 1912 2764 1952
rect 2804 1912 2813 1952
rect 2755 1911 2813 1912
rect 3139 1952 3197 1953
rect 3139 1912 3148 1952
rect 3188 1912 3197 1952
rect 3139 1911 3197 1912
rect 3339 1952 3381 1961
rect 3339 1912 3340 1952
rect 3380 1912 3381 1952
rect 3339 1903 3381 1912
rect 3627 1952 3669 1961
rect 3627 1912 3628 1952
rect 3668 1912 3669 1952
rect 3627 1903 3669 1912
rect 3723 1952 3765 1961
rect 3723 1912 3724 1952
rect 3764 1912 3765 1952
rect 3723 1903 3765 1912
rect 3819 1952 3861 1961
rect 3819 1912 3820 1952
rect 3860 1912 3861 1952
rect 3819 1903 3861 1912
rect 4195 1952 4253 1953
rect 4195 1912 4204 1952
rect 4244 1912 4253 1952
rect 4195 1911 4253 1912
rect 5443 1952 5501 1953
rect 5443 1912 5452 1952
rect 5492 1912 5501 1952
rect 5443 1911 5501 1912
rect 5731 1952 5789 1953
rect 5731 1912 5740 1952
rect 5780 1912 5789 1952
rect 5731 1911 5789 1912
rect 5827 1952 5885 1953
rect 5827 1912 5836 1952
rect 5876 1912 5885 1952
rect 5827 1911 5885 1912
rect 6027 1952 6069 1961
rect 6027 1912 6028 1952
rect 6068 1912 6069 1952
rect 6027 1903 6069 1912
rect 6123 1952 6165 1961
rect 6123 1912 6124 1952
rect 6164 1912 6165 1952
rect 6123 1903 6165 1912
rect 6280 1945 6322 1954
rect 6280 1905 6281 1945
rect 6321 1905 6322 1945
rect 6280 1896 6322 1905
rect 6795 1952 6837 1961
rect 6795 1912 6796 1952
rect 6836 1912 6837 1952
rect 6795 1903 6837 1912
rect 6891 1952 6933 1961
rect 6891 1912 6892 1952
rect 6932 1912 6933 1952
rect 6891 1903 6933 1912
rect 7275 1952 7317 1961
rect 7275 1912 7276 1952
rect 7316 1912 7317 1952
rect 7275 1903 7317 1912
rect 7371 1952 7413 1961
rect 7371 1912 7372 1952
rect 7412 1912 7413 1952
rect 7371 1903 7413 1912
rect 7843 1952 7901 1953
rect 7843 1912 7852 1952
rect 7892 1912 7901 1952
rect 9195 1952 9237 1961
rect 7843 1911 7901 1912
rect 8331 1942 8373 1951
rect 8331 1902 8332 1942
rect 8372 1902 8373 1942
rect 9195 1912 9196 1952
rect 9236 1912 9237 1952
rect 9195 1903 9237 1912
rect 9291 1952 9333 1961
rect 9291 1912 9292 1952
rect 9332 1912 9333 1952
rect 9291 1903 9333 1912
rect 9675 1952 9717 1961
rect 9675 1912 9676 1952
rect 9716 1912 9717 1952
rect 9675 1903 9717 1912
rect 9771 1952 9813 1961
rect 9771 1912 9772 1952
rect 9812 1912 9813 1952
rect 9771 1903 9813 1912
rect 10243 1952 10301 1953
rect 10243 1912 10252 1952
rect 10292 1912 10301 1952
rect 11115 1952 11157 1961
rect 10243 1911 10301 1912
rect 10731 1938 10773 1947
rect 8331 1893 8373 1902
rect 10731 1898 10732 1938
rect 10772 1898 10773 1938
rect 11115 1912 11116 1952
rect 11156 1912 11157 1952
rect 11115 1903 11157 1912
rect 11211 1952 11253 1961
rect 11211 1912 11212 1952
rect 11252 1912 11253 1952
rect 11211 1903 11253 1912
rect 11307 1952 11349 1961
rect 11307 1912 11308 1952
rect 11348 1912 11349 1952
rect 11307 1903 11349 1912
rect 11403 1952 11445 1961
rect 11403 1912 11404 1952
rect 11444 1912 11445 1952
rect 11403 1903 11445 1912
rect 11979 1952 12021 1961
rect 11979 1912 11980 1952
rect 12020 1912 12021 1952
rect 11979 1903 12021 1912
rect 12259 1952 12317 1953
rect 12259 1912 12268 1952
rect 12308 1912 12317 1952
rect 12259 1911 12317 1912
rect 12643 1952 12701 1953
rect 12643 1912 12652 1952
rect 12692 1912 12701 1952
rect 12643 1911 12701 1912
rect 13891 1952 13949 1953
rect 13891 1912 13900 1952
rect 13940 1912 13949 1952
rect 13891 1911 13949 1912
rect 14563 1952 14621 1953
rect 14563 1912 14572 1952
rect 14612 1912 14621 1952
rect 14563 1911 14621 1912
rect 15811 1952 15869 1953
rect 15811 1912 15820 1952
rect 15860 1912 15869 1952
rect 15811 1911 15869 1912
rect 16195 1952 16253 1953
rect 16195 1912 16204 1952
rect 16244 1912 16253 1952
rect 16195 1911 16253 1912
rect 17443 1952 17501 1953
rect 17443 1912 17452 1952
rect 17492 1912 17501 1952
rect 17443 1911 17501 1912
rect 17827 1952 17885 1953
rect 17827 1912 17836 1952
rect 17876 1912 17885 1952
rect 17827 1911 17885 1912
rect 19075 1952 19133 1953
rect 19075 1912 19084 1952
rect 19124 1912 19133 1952
rect 19075 1911 19133 1912
rect 19555 1952 19613 1953
rect 19555 1912 19564 1952
rect 19604 1912 19613 1952
rect 19555 1911 19613 1912
rect 20803 1952 20861 1953
rect 20803 1912 20812 1952
rect 20852 1912 20861 1952
rect 20803 1911 20861 1912
rect 21187 1952 21245 1953
rect 21187 1912 21196 1952
rect 21236 1912 21245 1952
rect 21187 1911 21245 1912
rect 22435 1952 22493 1953
rect 22435 1912 22444 1952
rect 22484 1912 22493 1952
rect 22435 1911 22493 1912
rect 22819 1952 22877 1953
rect 22819 1912 22828 1952
rect 22868 1912 22877 1952
rect 22819 1911 22877 1912
rect 24067 1952 24125 1953
rect 24067 1912 24076 1952
rect 24116 1912 24125 1952
rect 24067 1911 24125 1912
rect 24555 1952 24597 1961
rect 24555 1912 24556 1952
rect 24596 1912 24597 1952
rect 24555 1903 24597 1912
rect 24651 1952 24693 1961
rect 24651 1912 24652 1952
rect 24692 1912 24693 1952
rect 24651 1903 24693 1912
rect 25035 1952 25077 1961
rect 25035 1912 25036 1952
rect 25076 1912 25077 1952
rect 25035 1903 25077 1912
rect 25131 1952 25173 1961
rect 25131 1912 25132 1952
rect 25172 1912 25173 1952
rect 25131 1903 25173 1912
rect 25603 1952 25661 1953
rect 25603 1912 25612 1952
rect 25652 1912 25661 1952
rect 25603 1911 25661 1912
rect 26091 1947 26133 1956
rect 26091 1907 26092 1947
rect 26132 1907 26133 1947
rect 26659 1952 26717 1953
rect 26659 1912 26668 1952
rect 26708 1912 26717 1952
rect 26659 1911 26717 1912
rect 27907 1952 27965 1953
rect 27907 1912 27916 1952
rect 27956 1912 27965 1952
rect 27907 1911 27965 1912
rect 28203 1952 28245 1961
rect 28203 1912 28204 1952
rect 28244 1912 28245 1952
rect 26091 1898 26133 1907
rect 28203 1903 28245 1912
rect 28299 1952 28341 1961
rect 28299 1912 28300 1952
rect 28340 1912 28341 1952
rect 28299 1903 28341 1912
rect 28683 1952 28725 1961
rect 28683 1912 28684 1952
rect 28724 1912 28725 1952
rect 28683 1903 28725 1912
rect 28779 1952 28821 1961
rect 28779 1912 28780 1952
rect 28820 1912 28821 1952
rect 28779 1903 28821 1912
rect 29251 1952 29309 1953
rect 29251 1912 29260 1952
rect 29300 1912 29309 1952
rect 30307 1952 30365 1953
rect 29251 1911 29309 1912
rect 29739 1938 29781 1947
rect 29739 1898 29740 1938
rect 29780 1898 29781 1938
rect 30307 1912 30316 1952
rect 30356 1912 30365 1952
rect 30307 1911 30365 1912
rect 31555 1952 31613 1953
rect 31555 1912 31564 1952
rect 31604 1912 31613 1952
rect 31555 1911 31613 1912
rect 31747 1952 31805 1953
rect 31747 1912 31756 1952
rect 31796 1912 31805 1952
rect 31747 1911 31805 1912
rect 32995 1952 33053 1953
rect 32995 1912 33004 1952
rect 33044 1912 33053 1952
rect 32995 1911 33053 1912
rect 34051 1952 34109 1953
rect 34051 1912 34060 1952
rect 34100 1912 34109 1952
rect 34051 1911 34109 1912
rect 34915 1952 34973 1953
rect 34915 1912 34924 1952
rect 34964 1912 34973 1952
rect 34915 1911 34973 1912
rect 36931 1952 36989 1953
rect 36931 1912 36940 1952
rect 36980 1912 36989 1952
rect 36931 1911 36989 1912
rect 37795 1952 37853 1953
rect 37795 1912 37804 1952
rect 37844 1912 37853 1952
rect 37795 1911 37853 1912
rect 39235 1952 39293 1953
rect 39235 1912 39244 1952
rect 39284 1912 39293 1952
rect 39235 1911 39293 1912
rect 40771 1952 40829 1953
rect 40771 1912 40780 1952
rect 40820 1912 40829 1952
rect 40771 1911 40829 1912
rect 10731 1889 10773 1898
rect 29739 1889 29781 1898
rect 4011 1700 4053 1709
rect 4011 1660 4012 1700
rect 4052 1660 4053 1700
rect 4011 1651 4053 1660
rect 11587 1700 11645 1701
rect 11587 1660 11596 1700
rect 11636 1660 11645 1700
rect 11587 1659 11645 1660
rect 39531 1700 39573 1709
rect 39531 1660 39532 1700
rect 39572 1660 39573 1700
rect 39531 1651 39573 1660
rect 1152 1532 41856 1556
rect 1152 1492 3688 1532
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 4056 1492 18808 1532
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 19176 1492 33928 1532
rect 33968 1492 34010 1532
rect 34050 1492 34092 1532
rect 34132 1492 34174 1532
rect 34214 1492 34256 1532
rect 34296 1492 41856 1532
rect 1152 1468 41856 1492
rect 3339 1364 3381 1373
rect 3339 1324 3340 1364
rect 3380 1324 3381 1364
rect 3339 1315 3381 1324
rect 11211 1364 11253 1373
rect 11211 1324 11212 1364
rect 11252 1324 11253 1364
rect 11211 1315 11253 1324
rect 20907 1364 20949 1373
rect 20907 1324 20908 1364
rect 20948 1324 20949 1364
rect 20907 1315 20949 1324
rect 24459 1364 24501 1373
rect 24459 1324 24460 1364
rect 24500 1324 24501 1364
rect 24459 1315 24501 1324
rect 27915 1364 27957 1373
rect 27915 1324 27916 1364
rect 27956 1324 27957 1364
rect 27915 1315 27957 1324
rect 29547 1364 29589 1373
rect 29547 1324 29548 1364
rect 29588 1324 29589 1364
rect 29547 1315 29589 1324
rect 31563 1364 31605 1373
rect 31563 1324 31564 1364
rect 31604 1324 31605 1364
rect 31563 1315 31605 1324
rect 41547 1364 41589 1373
rect 41547 1324 41548 1364
rect 41588 1324 41589 1364
rect 41547 1315 41589 1324
rect 5259 1280 5301 1289
rect 5259 1240 5260 1280
rect 5300 1240 5301 1280
rect 5259 1231 5301 1240
rect 7171 1280 7229 1281
rect 7171 1240 7180 1280
rect 7220 1240 7229 1280
rect 7171 1239 7229 1240
rect 9579 1280 9621 1289
rect 9579 1240 9580 1280
rect 9620 1240 9621 1280
rect 9579 1231 9621 1240
rect 11691 1280 11733 1289
rect 11691 1240 11692 1280
rect 11732 1240 11733 1280
rect 11691 1231 11733 1240
rect 13611 1280 13653 1289
rect 13611 1240 13612 1280
rect 13652 1240 13653 1280
rect 13611 1231 13653 1240
rect 15435 1280 15477 1289
rect 15435 1240 15436 1280
rect 15476 1240 15477 1280
rect 15435 1231 15477 1240
rect 17355 1280 17397 1289
rect 17355 1240 17356 1280
rect 17396 1240 17397 1280
rect 17355 1231 17397 1240
rect 19083 1280 19125 1289
rect 19083 1240 19084 1280
rect 19124 1240 19125 1280
rect 19083 1231 19125 1240
rect 22539 1280 22581 1289
rect 22539 1240 22540 1280
rect 22580 1240 22581 1280
rect 22539 1231 22581 1240
rect 24651 1280 24693 1289
rect 24651 1240 24652 1280
rect 24692 1240 24693 1280
rect 24651 1231 24693 1240
rect 27723 1280 27765 1289
rect 27723 1240 27724 1280
rect 27764 1240 27765 1280
rect 27723 1231 27765 1240
rect 32427 1280 32469 1289
rect 32427 1240 32428 1280
rect 32468 1240 32469 1280
rect 32427 1231 32469 1240
rect 32811 1280 32853 1289
rect 32811 1240 32812 1280
rect 32852 1240 32853 1280
rect 32811 1231 32853 1240
rect 34827 1280 34869 1289
rect 34827 1240 34828 1280
rect 34868 1240 34869 1280
rect 34827 1231 34869 1240
rect 36267 1280 36309 1289
rect 36267 1240 36268 1280
rect 36308 1240 36309 1280
rect 36267 1231 36309 1240
rect 36835 1280 36893 1281
rect 36835 1240 36844 1280
rect 36884 1240 36893 1280
rect 36835 1239 36893 1240
rect 40203 1280 40245 1289
rect 40203 1240 40204 1280
rect 40244 1240 40245 1280
rect 40203 1231 40245 1240
rect 40587 1280 40629 1289
rect 40587 1240 40588 1280
rect 40628 1240 40629 1280
rect 40587 1231 40629 1240
rect 13795 1196 13853 1197
rect 13795 1156 13804 1196
rect 13844 1156 13853 1196
rect 13795 1155 13853 1156
rect 32611 1196 32669 1197
rect 32611 1156 32620 1196
rect 32660 1156 32669 1196
rect 32611 1155 32669 1156
rect 32995 1196 33053 1197
rect 32995 1156 33004 1196
rect 33044 1156 33053 1196
rect 32995 1155 33053 1156
rect 35203 1196 35261 1197
rect 35203 1156 35212 1196
rect 35252 1156 35261 1196
rect 35203 1155 35261 1156
rect 39619 1196 39677 1197
rect 39619 1156 39628 1196
rect 39668 1156 39677 1196
rect 39619 1155 39677 1156
rect 40003 1196 40061 1197
rect 40003 1156 40012 1196
rect 40052 1156 40061 1196
rect 40003 1155 40061 1156
rect 41155 1196 41213 1197
rect 41155 1156 41164 1196
rect 41204 1156 41213 1196
rect 41155 1155 41213 1156
rect 41347 1196 41405 1197
rect 41347 1156 41356 1196
rect 41396 1156 41405 1196
rect 41347 1155 41405 1156
rect 1515 1112 1557 1121
rect 1515 1072 1516 1112
rect 1556 1072 1557 1112
rect 1515 1063 1557 1072
rect 1611 1112 1653 1121
rect 1611 1072 1612 1112
rect 1652 1072 1653 1112
rect 1611 1063 1653 1072
rect 1707 1112 1749 1121
rect 1707 1072 1708 1112
rect 1748 1072 1749 1112
rect 1707 1063 1749 1072
rect 1891 1112 1949 1113
rect 1891 1072 1900 1112
rect 1940 1072 1949 1112
rect 1891 1071 1949 1072
rect 3139 1112 3197 1113
rect 3139 1072 3148 1112
rect 3188 1072 3197 1112
rect 3139 1071 3197 1072
rect 3811 1112 3869 1113
rect 3811 1072 3820 1112
rect 3860 1072 3869 1112
rect 3811 1071 3869 1072
rect 5059 1112 5117 1113
rect 5059 1072 5068 1112
rect 5108 1072 5117 1112
rect 5059 1071 5117 1072
rect 5739 1112 5781 1121
rect 5739 1072 5740 1112
rect 5780 1072 5781 1112
rect 5739 1063 5781 1072
rect 5835 1112 5877 1121
rect 5835 1072 5836 1112
rect 5876 1072 5877 1112
rect 5835 1063 5877 1072
rect 6219 1112 6261 1121
rect 6219 1072 6220 1112
rect 6260 1072 6261 1112
rect 6219 1063 6261 1072
rect 6315 1112 6357 1121
rect 6315 1072 6316 1112
rect 6356 1072 6357 1112
rect 6315 1063 6357 1072
rect 6411 1112 6453 1121
rect 6411 1072 6412 1112
rect 6452 1072 6453 1112
rect 6411 1063 6453 1072
rect 6699 1112 6741 1121
rect 6699 1072 6700 1112
rect 6740 1072 6741 1112
rect 6699 1063 6741 1072
rect 6795 1112 6837 1121
rect 6795 1072 6796 1112
rect 6836 1072 6837 1112
rect 6795 1063 6837 1072
rect 6891 1112 6933 1121
rect 6891 1072 6892 1112
rect 6932 1072 6933 1112
rect 6891 1063 6933 1072
rect 6987 1112 7029 1121
rect 6987 1072 6988 1112
rect 7028 1072 7029 1112
rect 6987 1063 7029 1072
rect 7467 1112 7509 1121
rect 7467 1072 7468 1112
rect 7508 1072 7509 1112
rect 7467 1063 7509 1072
rect 7563 1112 7605 1121
rect 7563 1072 7564 1112
rect 7604 1072 7605 1112
rect 7563 1063 7605 1072
rect 7843 1112 7901 1113
rect 7843 1072 7852 1112
rect 7892 1072 7901 1112
rect 7843 1071 7901 1072
rect 8131 1112 8189 1113
rect 8131 1072 8140 1112
rect 8180 1072 8189 1112
rect 8131 1071 8189 1072
rect 9379 1112 9437 1113
rect 9379 1072 9388 1112
rect 9428 1072 9437 1112
rect 9379 1071 9437 1072
rect 9763 1112 9821 1113
rect 9763 1072 9772 1112
rect 9812 1072 9821 1112
rect 9763 1071 9821 1072
rect 11011 1112 11069 1113
rect 11011 1072 11020 1112
rect 11060 1072 11069 1112
rect 11011 1071 11069 1072
rect 11395 1112 11453 1113
rect 11395 1072 11404 1112
rect 11444 1072 11453 1112
rect 11395 1071 11453 1072
rect 11499 1112 11541 1121
rect 11499 1072 11500 1112
rect 11540 1072 11541 1112
rect 11499 1063 11541 1072
rect 11691 1112 11733 1121
rect 11691 1072 11692 1112
rect 11732 1072 11733 1112
rect 11691 1063 11733 1072
rect 11883 1112 11925 1121
rect 11883 1072 11884 1112
rect 11924 1072 11925 1112
rect 11883 1063 11925 1072
rect 11979 1112 12021 1121
rect 11979 1072 11980 1112
rect 12020 1072 12021 1112
rect 11979 1063 12021 1072
rect 12075 1112 12117 1121
rect 12075 1072 12076 1112
rect 12116 1072 12117 1112
rect 12075 1063 12117 1072
rect 12363 1112 12405 1121
rect 12363 1072 12364 1112
rect 12404 1072 12405 1112
rect 12363 1063 12405 1072
rect 12459 1112 12501 1121
rect 12459 1072 12460 1112
rect 12500 1072 12501 1112
rect 12459 1063 12501 1072
rect 12555 1112 12597 1121
rect 12555 1072 12556 1112
rect 12596 1072 12597 1112
rect 12555 1063 12597 1072
rect 12651 1112 12693 1121
rect 12651 1072 12652 1112
rect 12692 1072 12693 1112
rect 12651 1063 12693 1072
rect 12843 1112 12885 1121
rect 12843 1072 12844 1112
rect 12884 1072 12885 1112
rect 12843 1063 12885 1072
rect 12939 1112 12981 1121
rect 12939 1072 12940 1112
rect 12980 1072 12981 1112
rect 12939 1063 12981 1072
rect 13035 1112 13077 1121
rect 13035 1072 13036 1112
rect 13076 1072 13077 1112
rect 13035 1063 13077 1072
rect 13131 1112 13173 1121
rect 13131 1072 13132 1112
rect 13172 1072 13173 1112
rect 13131 1063 13173 1072
rect 13987 1112 14045 1113
rect 13987 1072 13996 1112
rect 14036 1072 14045 1112
rect 13987 1071 14045 1072
rect 15235 1112 15293 1113
rect 15235 1072 15244 1112
rect 15284 1072 15293 1112
rect 15235 1071 15293 1072
rect 15907 1112 15965 1113
rect 15907 1072 15916 1112
rect 15956 1072 15965 1112
rect 15907 1071 15965 1072
rect 17155 1112 17213 1113
rect 17155 1072 17164 1112
rect 17204 1072 17213 1112
rect 17155 1071 17213 1072
rect 17635 1112 17693 1113
rect 17635 1072 17644 1112
rect 17684 1072 17693 1112
rect 17635 1071 17693 1072
rect 18883 1112 18941 1113
rect 18883 1072 18892 1112
rect 18932 1072 18941 1112
rect 18883 1071 18941 1072
rect 19459 1112 19517 1113
rect 19459 1072 19468 1112
rect 19508 1072 19517 1112
rect 19459 1071 19517 1072
rect 20707 1112 20765 1113
rect 20707 1072 20716 1112
rect 20756 1072 20765 1112
rect 20707 1071 20765 1072
rect 21091 1112 21149 1113
rect 21091 1072 21100 1112
rect 21140 1072 21149 1112
rect 21091 1071 21149 1072
rect 22339 1112 22397 1113
rect 22339 1072 22348 1112
rect 22388 1072 22397 1112
rect 22339 1071 22397 1072
rect 23011 1112 23069 1113
rect 23011 1072 23020 1112
rect 23060 1072 23069 1112
rect 23011 1071 23069 1072
rect 24259 1112 24317 1113
rect 24259 1072 24268 1112
rect 24308 1072 24317 1112
rect 24259 1071 24317 1072
rect 24835 1112 24893 1113
rect 24835 1072 24844 1112
rect 24884 1072 24893 1112
rect 24835 1071 24893 1072
rect 26083 1112 26141 1113
rect 26083 1072 26092 1112
rect 26132 1072 26141 1112
rect 26083 1071 26141 1072
rect 26275 1112 26333 1113
rect 26275 1072 26284 1112
rect 26324 1072 26333 1112
rect 26275 1071 26333 1072
rect 27523 1112 27581 1113
rect 27523 1072 27532 1112
rect 27572 1072 27581 1112
rect 27523 1071 27581 1072
rect 28099 1112 28157 1113
rect 28099 1072 28108 1112
rect 28148 1072 28157 1112
rect 28099 1071 28157 1072
rect 29347 1112 29405 1113
rect 29347 1072 29356 1112
rect 29396 1072 29405 1112
rect 29347 1071 29405 1072
rect 29731 1112 29789 1113
rect 29731 1072 29740 1112
rect 29780 1072 29789 1112
rect 29731 1071 29789 1072
rect 30979 1112 31037 1113
rect 30979 1072 30988 1112
rect 31028 1072 31037 1112
rect 30979 1071 31037 1072
rect 31267 1112 31325 1113
rect 31267 1072 31276 1112
rect 31316 1072 31325 1112
rect 31267 1071 31325 1072
rect 33379 1112 33437 1113
rect 33379 1072 33388 1112
rect 33428 1072 33437 1112
rect 33379 1071 33437 1072
rect 34627 1112 34685 1113
rect 34627 1072 34636 1112
rect 34676 1072 34685 1112
rect 34627 1071 34685 1072
rect 35587 1112 35645 1113
rect 35587 1072 35596 1112
rect 35636 1072 35645 1112
rect 35587 1071 35645 1072
rect 36547 1112 36605 1113
rect 36547 1072 36556 1112
rect 36596 1072 36605 1112
rect 36547 1071 36605 1072
rect 37987 1112 38045 1113
rect 37987 1072 37996 1112
rect 38036 1072 38045 1112
rect 37987 1071 38045 1072
rect 38851 1112 38909 1113
rect 38851 1072 38860 1112
rect 38900 1072 38909 1112
rect 38851 1071 38909 1072
rect 39243 1112 39285 1121
rect 39243 1072 39244 1112
rect 39284 1072 39285 1112
rect 39243 1063 39285 1072
rect 1411 944 1469 945
rect 1411 904 1420 944
rect 1460 904 1469 944
rect 1411 903 1469 904
rect 6019 944 6077 945
rect 6019 904 6028 944
rect 6068 904 6077 944
rect 6019 903 6077 904
rect 6499 944 6557 945
rect 6499 904 6508 944
rect 6548 904 6557 944
rect 6499 903 6557 904
rect 12163 944 12221 945
rect 12163 904 12172 944
rect 12212 904 12221 944
rect 12163 903 12221 904
rect 35019 944 35061 953
rect 35019 904 35020 944
rect 35060 904 35061 944
rect 35019 895 35061 904
rect 39435 944 39477 953
rect 39435 904 39436 944
rect 39476 904 39477 944
rect 39435 895 39477 904
rect 39819 944 39861 953
rect 39819 904 39820 944
rect 39860 904 39861 944
rect 39819 895 39861 904
rect 40971 944 41013 953
rect 40971 904 40972 944
rect 41012 904 41013 944
rect 40971 895 41013 904
rect 1152 776 41856 800
rect 1152 736 4928 776
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 5296 736 20048 776
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20416 736 35168 776
rect 35208 736 35250 776
rect 35290 736 35332 776
rect 35372 736 35414 776
rect 35454 736 35496 776
rect 35536 736 41856 776
rect 1152 712 41856 736
<< via1 >>
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 35168 9808 35208 9848
rect 35250 9808 35290 9848
rect 35332 9808 35372 9848
rect 35414 9808 35454 9848
rect 35496 9808 35536 9848
rect 6412 9640 6452 9680
rect 7660 9640 7700 9680
rect 9004 9640 9044 9680
rect 9388 9640 9428 9680
rect 9772 9640 9812 9680
rect 10156 9640 10196 9680
rect 12652 9640 12692 9680
rect 13036 9640 13076 9680
rect 14764 9640 14804 9680
rect 18796 9640 18836 9680
rect 25036 9640 25076 9680
rect 27052 9640 27092 9680
rect 3244 9556 3284 9596
rect 22924 9556 22964 9596
rect 1612 9472 1652 9512
rect 2860 9472 2900 9512
rect 3436 9472 3476 9512
rect 4684 9472 4724 9512
rect 4876 9472 4916 9512
rect 4972 9472 5012 9512
rect 5068 9472 5108 9512
rect 5164 9472 5204 9512
rect 6220 9472 6260 9512
rect 6604 9472 6644 9512
rect 6700 9472 6740 9512
rect 6892 9472 6932 9512
rect 6988 9472 7028 9512
rect 7089 9472 7129 9512
rect 7372 9472 7412 9512
rect 7468 9472 7508 9512
rect 8140 9472 8180 9512
rect 8236 9472 8276 9512
rect 8332 9472 8372 9512
rect 8428 9472 8468 9512
rect 8716 9472 8756 9512
rect 8812 9472 8852 9512
rect 15148 9472 15188 9512
rect 16396 9472 16436 9512
rect 16780 9472 16820 9512
rect 18028 9472 18068 9512
rect 19468 9472 19508 9512
rect 20716 9472 20756 9512
rect 21196 9472 21236 9512
rect 21292 9472 21332 9512
rect 21676 9472 21716 9512
rect 22252 9472 22292 9512
rect 22732 9458 22772 9498
rect 23308 9472 23348 9512
rect 24556 9472 24596 9512
rect 25420 9472 25460 9512
rect 26668 9472 26708 9512
rect 29356 9472 29396 9512
rect 30604 9472 30644 9512
rect 31180 9472 31220 9512
rect 32428 9472 32468 9512
rect 32812 9472 32852 9512
rect 34060 9472 34100 9512
rect 34444 9472 34484 9512
rect 35692 9472 35732 9512
rect 36076 9472 36116 9512
rect 37324 9472 37364 9512
rect 37900 9472 37940 9512
rect 39148 9472 39188 9512
rect 39340 9472 39380 9512
rect 40588 9472 40628 9512
rect 9580 9388 9620 9428
rect 9964 9388 10004 9428
rect 10348 9388 10388 9428
rect 12844 9388 12884 9428
rect 13228 9388 13268 9428
rect 14956 9388 14996 9428
rect 18604 9388 18644 9428
rect 21772 9388 21812 9428
rect 25228 9388 25268 9428
rect 27244 9388 27284 9428
rect 40972 9388 41012 9428
rect 6220 9304 6260 9344
rect 26860 9304 26900 9344
rect 41356 9304 41396 9344
rect 3052 9220 3092 9260
rect 6604 9220 6644 9260
rect 16588 9220 16628 9260
rect 18220 9220 18260 9260
rect 20908 9220 20948 9260
rect 23116 9220 23156 9260
rect 30796 9220 30836 9260
rect 30988 9220 31028 9260
rect 32620 9220 32660 9260
rect 34252 9220 34292 9260
rect 37516 9220 37556 9260
rect 37708 9220 37748 9260
rect 40780 9220 40820 9260
rect 41164 9220 41204 9260
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 33928 9052 33968 9092
rect 34010 9052 34050 9092
rect 34092 9052 34132 9092
rect 34174 9052 34214 9092
rect 34256 9052 34296 9092
rect 9484 8884 9524 8924
rect 9868 8800 9908 8840
rect 10636 8800 10676 8840
rect 10828 8800 10868 8840
rect 11212 8800 11252 8840
rect 11788 8800 11828 8840
rect 12172 8800 12212 8840
rect 30028 8800 30068 8840
rect 9676 8716 9716 8756
rect 10060 8716 10100 8756
rect 10444 8716 10484 8756
rect 11020 8716 11060 8756
rect 11404 8716 11444 8756
rect 11596 8716 11636 8756
rect 11980 8716 12020 8756
rect 15244 8716 15284 8756
rect 18892 8716 18932 8756
rect 24364 8716 24404 8756
rect 26476 8716 26516 8756
rect 29452 8716 29492 8756
rect 29836 8716 29876 8756
rect 31468 8716 31508 8756
rect 32524 8716 32564 8756
rect 32908 8716 32948 8756
rect 35404 8716 35444 8756
rect 41356 8716 41396 8756
rect 1900 8632 1940 8672
rect 1996 8632 2036 8672
rect 2092 8632 2132 8672
rect 2476 8632 2516 8672
rect 2572 8632 2612 8672
rect 2860 8632 2900 8672
rect 2956 8632 2996 8672
rect 3340 8632 3380 8672
rect 3436 8632 3476 8672
rect 3916 8632 3956 8672
rect 4396 8637 4436 8677
rect 4780 8632 4820 8672
rect 6028 8632 6068 8672
rect 6796 8632 6836 8672
rect 6892 8632 6932 8672
rect 7276 8632 7316 8672
rect 7372 8632 7412 8672
rect 7852 8632 7892 8672
rect 8332 8637 8372 8677
rect 8812 8632 8852 8672
rect 9100 8632 9140 8672
rect 12364 8632 12404 8672
rect 13612 8632 13652 8672
rect 14140 8641 14180 8681
rect 14668 8632 14708 8672
rect 15148 8632 15188 8672
rect 15628 8632 15668 8672
rect 15724 8632 15764 8672
rect 16396 8632 16436 8672
rect 16492 8632 16532 8672
rect 16876 8632 16916 8672
rect 16972 8632 17012 8672
rect 17452 8632 17492 8672
rect 17932 8646 17972 8686
rect 18412 8632 18452 8672
rect 18508 8632 18548 8672
rect 18988 8632 19028 8672
rect 19468 8632 19508 8672
rect 19948 8637 19988 8677
rect 21772 8632 21812 8672
rect 21868 8632 21908 8672
rect 22252 8632 22292 8672
rect 22348 8632 22388 8672
rect 22828 8632 22868 8672
rect 23308 8646 23348 8686
rect 23884 8632 23924 8672
rect 23980 8632 24020 8672
rect 24460 8632 24500 8672
rect 24940 8632 24980 8672
rect 25468 8641 25508 8681
rect 25900 8632 25940 8672
rect 25996 8632 26036 8672
rect 26380 8632 26420 8672
rect 26956 8632 26996 8672
rect 27484 8641 27524 8681
rect 28012 8632 28052 8672
rect 29260 8632 29300 8672
rect 30508 8646 30548 8686
rect 30988 8632 31028 8672
rect 31564 8632 31604 8672
rect 31948 8612 31988 8652
rect 32044 8632 32084 8672
rect 33292 8632 33332 8672
rect 33388 8632 33428 8672
rect 33772 8632 33812 8672
rect 33868 8632 33908 8672
rect 34348 8632 34388 8672
rect 34828 8646 34868 8686
rect 35788 8632 35828 8672
rect 35884 8632 35924 8672
rect 36268 8632 36308 8672
rect 36364 8632 36404 8672
rect 36844 8632 36884 8672
rect 37372 8641 37412 8681
rect 37804 8632 37844 8672
rect 37900 8632 37940 8672
rect 38284 8632 38324 8672
rect 38380 8632 38420 8672
rect 38860 8632 38900 8672
rect 39340 8646 39380 8686
rect 39916 8632 39956 8672
rect 41164 8632 41204 8672
rect 8524 8548 8564 8588
rect 9196 8548 9236 8588
rect 18124 8548 18164 8588
rect 20140 8548 20180 8588
rect 25612 8548 25652 8588
rect 27628 8548 27668 8588
rect 30316 8548 30356 8588
rect 1804 8464 1844 8504
rect 2284 8464 2324 8504
rect 4588 8464 4628 8504
rect 6220 8464 6260 8504
rect 10252 8464 10292 8504
rect 13804 8464 13844 8504
rect 13996 8464 14036 8504
rect 20332 8464 20372 8504
rect 23500 8464 23540 8504
rect 27820 8464 27860 8504
rect 29644 8464 29684 8504
rect 32332 8464 32372 8504
rect 32716 8464 32756 8504
rect 35020 8464 35060 8504
rect 35212 8464 35252 8504
rect 37516 8464 37556 8504
rect 39532 8464 39572 8504
rect 39724 8464 39764 8504
rect 41548 8464 41588 8504
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 35168 8296 35208 8336
rect 35250 8296 35290 8336
rect 35332 8296 35372 8336
rect 35414 8296 35454 8336
rect 35496 8296 35536 8336
rect 4108 8170 4148 8210
rect 3340 8128 3380 8168
rect 8428 8128 8468 8168
rect 11116 8128 11156 8168
rect 13996 8128 14036 8168
rect 17740 8128 17780 8168
rect 19372 8128 19412 8168
rect 21004 8128 21044 8168
rect 23212 8128 23252 8168
rect 25516 8128 25556 8168
rect 25708 8128 25748 8168
rect 26284 8128 26324 8168
rect 30412 8128 30452 8168
rect 30796 8128 30836 8168
rect 33196 8128 33236 8168
rect 35692 8128 35732 8168
rect 37900 8128 37940 8168
rect 40684 8128 40724 8168
rect 10924 8044 10964 8084
rect 23020 8044 23060 8084
rect 28588 8044 28628 8084
rect 1900 7960 1940 8000
rect 3148 7960 3188 8000
rect 3820 7960 3860 8000
rect 3916 7961 3956 8001
rect 4300 7960 4340 8000
rect 4396 7960 4436 8000
rect 4492 7960 4532 8000
rect 4588 7960 4628 8000
rect 4780 7960 4820 8000
rect 6028 7960 6068 8000
rect 6700 7960 6740 8000
rect 6796 7960 6836 8000
rect 7756 7960 7796 8000
rect 8236 7946 8276 7986
rect 8620 7960 8660 8000
rect 8716 7960 8756 8000
rect 8812 7960 8852 8000
rect 8908 7960 8948 8000
rect 9100 7960 9140 8000
rect 9292 7960 9332 8000
rect 9484 7960 9524 8000
rect 10732 7960 10772 8000
rect 11260 7950 11300 7990
rect 11788 7960 11828 8000
rect 12268 7960 12308 8000
rect 12748 7960 12788 8000
rect 12844 7960 12884 8000
rect 14188 7960 14228 8000
rect 15436 7960 15476 8000
rect 16300 7960 16340 8000
rect 17548 7960 17588 8000
rect 17932 7960 17972 8000
rect 19180 7960 19220 8000
rect 19564 7960 19604 8000
rect 20812 7960 20852 8000
rect 21292 7960 21332 8000
rect 21388 7960 21428 8000
rect 21772 7960 21812 8000
rect 21868 7960 21908 8000
rect 22348 7960 22388 8000
rect 22828 7946 22868 7986
rect 24076 7960 24116 8000
rect 25324 7960 25364 8000
rect 26860 7960 26900 8000
rect 26956 7960 26996 8000
rect 27436 7960 27476 8000
rect 27916 7960 27956 8000
rect 28396 7955 28436 7995
rect 28780 7960 28820 8000
rect 30028 7960 30068 8000
rect 31468 7960 31508 8000
rect 31564 7960 31604 8000
rect 31948 7960 31988 8000
rect 32044 7960 32084 8000
rect 32524 7969 32564 8009
rect 33052 7950 33092 7990
rect 34060 7960 34100 8000
rect 35308 7960 35348 8000
rect 35884 7960 35924 8000
rect 37132 7960 37172 8000
rect 38956 7960 38996 8000
rect 39052 7960 39092 8000
rect 39436 7960 39476 8000
rect 39532 7960 39572 8000
rect 40012 7960 40052 8000
rect 40492 7946 40532 7986
rect 7180 7876 7220 7916
rect 7276 7876 7316 7916
rect 12364 7876 12404 7916
rect 23404 7876 23444 7916
rect 25900 7876 25940 7916
rect 26092 7865 26132 7905
rect 27340 7876 27380 7916
rect 30604 7876 30644 7916
rect 30988 7876 31028 7916
rect 33868 7876 33908 7916
rect 37516 7876 37556 7916
rect 37708 7876 37748 7916
rect 38284 7876 38324 7916
rect 38668 7876 38708 7916
rect 40876 7876 40916 7916
rect 41260 7876 41300 7916
rect 33676 7792 33716 7832
rect 41452 7792 41492 7832
rect 6220 7708 6260 7748
rect 9196 7708 9236 7748
rect 30220 7708 30260 7748
rect 35500 7708 35540 7748
rect 37324 7708 37364 7748
rect 38092 7708 38132 7748
rect 38476 7708 38516 7748
rect 41068 7708 41108 7748
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 33928 7540 33968 7580
rect 34010 7540 34050 7580
rect 34092 7540 34132 7580
rect 34174 7540 34214 7580
rect 34256 7540 34296 7580
rect 6028 7372 6068 7412
rect 6988 7372 7028 7412
rect 7372 7372 7412 7412
rect 7852 7372 7892 7412
rect 10444 7372 10484 7412
rect 10828 7372 10868 7412
rect 11020 7372 11060 7412
rect 12652 7372 12692 7412
rect 15724 7372 15764 7412
rect 22444 7372 22484 7412
rect 24076 7372 24116 7412
rect 26188 7372 26228 7412
rect 31852 7372 31892 7412
rect 33484 7372 33524 7412
rect 35404 7372 35444 7412
rect 41260 7372 41300 7412
rect 10252 7204 10292 7244
rect 10636 7204 10676 7244
rect 12844 7204 12884 7244
rect 13804 7204 13844 7244
rect 15532 7204 15572 7244
rect 18604 7204 18644 7244
rect 28300 7204 28340 7244
rect 28396 7204 28436 7244
rect 29836 7204 29876 7244
rect 35596 7204 35636 7244
rect 35788 7204 35828 7244
rect 36364 7204 36404 7244
rect 41452 7204 41492 7244
rect 1324 7120 1364 7160
rect 1516 7120 1556 7160
rect 1708 7120 1748 7160
rect 2956 7120 2996 7160
rect 3436 7120 3476 7160
rect 3532 7120 3572 7160
rect 3628 7120 3668 7160
rect 4108 7120 4148 7160
rect 4204 7120 4244 7160
rect 4588 7120 4628 7160
rect 5836 7120 5876 7160
rect 6316 7120 6356 7160
rect 6604 7120 6644 7160
rect 6700 7120 6740 7160
rect 7372 7120 7412 7160
rect 7564 7120 7604 7160
rect 7660 7120 7700 7160
rect 8044 7120 8084 7160
rect 9292 7120 9332 7160
rect 9484 7120 9524 7160
rect 9676 7120 9716 7160
rect 9772 7120 9812 7160
rect 10060 7120 10100 7160
rect 11212 7120 11252 7160
rect 12460 7120 12500 7160
rect 13324 7120 13364 7160
rect 13420 7120 13460 7160
rect 13900 7120 13940 7160
rect 14380 7120 14420 7160
rect 14860 7125 14900 7165
rect 15916 7120 15956 7160
rect 17164 7120 17204 7160
rect 18124 7120 18164 7160
rect 18220 7120 18260 7160
rect 18700 7120 18740 7160
rect 19180 7120 19220 7160
rect 19660 7125 19700 7165
rect 21004 7120 21044 7160
rect 22252 7120 22292 7160
rect 22636 7120 22676 7160
rect 23884 7120 23924 7160
rect 24748 7120 24788 7160
rect 25996 7120 26036 7160
rect 27820 7120 27860 7160
rect 27916 7120 27956 7160
rect 28876 7120 28916 7160
rect 29356 7125 29396 7165
rect 30220 7120 30260 7160
rect 31468 7120 31508 7160
rect 32044 7120 32084 7160
rect 33292 7120 33332 7160
rect 33676 7120 33716 7160
rect 34924 7120 34964 7160
rect 36556 7120 36596 7160
rect 37804 7120 37844 7160
rect 38380 7120 38420 7160
rect 39628 7120 39668 7160
rect 39820 7120 39860 7160
rect 41068 7120 41108 7160
rect 3148 7036 3188 7076
rect 15052 7036 15092 7076
rect 19852 7036 19892 7076
rect 1420 6952 1460 6992
rect 3724 6952 3764 6992
rect 3916 6952 3956 6992
rect 9580 6952 9620 6992
rect 9964 6952 10004 6992
rect 17356 6952 17396 6992
rect 29548 6952 29588 6992
rect 30028 6952 30068 6992
rect 31660 6952 31700 6992
rect 35980 6952 36020 6992
rect 36172 6952 36212 6992
rect 37996 6952 38036 6992
rect 38188 6952 38228 6992
rect 41644 6952 41684 6992
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 35168 6784 35208 6824
rect 35250 6784 35290 6824
rect 35332 6784 35372 6824
rect 35414 6784 35454 6824
rect 35496 6784 35536 6824
rect 4684 6616 4724 6656
rect 5164 6616 5204 6656
rect 5932 6616 5972 6656
rect 8428 6616 8468 6656
rect 10252 6616 10292 6656
rect 12460 6616 12500 6656
rect 14092 6616 14132 6656
rect 17740 6616 17780 6656
rect 25708 6616 25748 6656
rect 31564 6616 31604 6656
rect 31948 6616 31988 6656
rect 32524 6616 32564 6656
rect 34732 6616 34772 6656
rect 36844 6616 36884 6656
rect 37420 6616 37460 6656
rect 39436 6616 39476 6656
rect 41068 6616 41108 6656
rect 6508 6532 6548 6572
rect 15724 6532 15764 6572
rect 20620 6532 20660 6572
rect 23692 6532 23732 6572
rect 27532 6532 27572 6572
rect 29548 6532 29588 6572
rect 1228 6448 1268 6488
rect 2476 6448 2516 6488
rect 2956 6448 2996 6488
rect 3052 6448 3092 6488
rect 3436 6448 3476 6488
rect 4012 6448 4052 6488
rect 4492 6443 4532 6483
rect 4876 6448 4916 6488
rect 4972 6448 5012 6488
rect 5068 6448 5108 6488
rect 5356 6448 5396 6488
rect 5548 6448 5588 6488
rect 5740 6448 5780 6488
rect 5836 6448 5876 6488
rect 6028 6448 6068 6488
rect 6220 6448 6260 6488
rect 6316 6448 6356 6488
rect 6412 6448 6452 6488
rect 6700 6448 6740 6488
rect 6892 6448 6932 6488
rect 6988 6448 7028 6488
rect 7276 6448 7316 6488
rect 7564 6448 7604 6488
rect 7660 6448 7700 6488
rect 8140 6448 8180 6488
rect 8236 6448 8276 6488
rect 8332 6448 8372 6488
rect 8812 6448 8852 6488
rect 10060 6448 10100 6488
rect 10444 6448 10484 6488
rect 10636 6448 10676 6488
rect 10732 6448 10772 6488
rect 11020 6448 11060 6488
rect 12268 6448 12308 6488
rect 12652 6448 12692 6488
rect 13900 6448 13940 6488
rect 14284 6448 14324 6488
rect 15532 6448 15572 6488
rect 16012 6448 16052 6488
rect 16108 6448 16148 6488
rect 16492 6448 16532 6488
rect 17068 6448 17108 6488
rect 17548 6443 17588 6483
rect 18892 6448 18932 6488
rect 18988 6448 19028 6488
rect 19372 6448 19412 6488
rect 19468 6448 19508 6488
rect 19948 6448 19988 6488
rect 20428 6434 20468 6474
rect 22252 6448 22292 6488
rect 23500 6448 23540 6488
rect 23980 6448 24020 6488
rect 24076 6448 24116 6488
rect 24460 6448 24500 6488
rect 25036 6448 25076 6488
rect 25564 6438 25604 6478
rect 26092 6448 26132 6488
rect 27340 6448 27380 6488
rect 27820 6448 27860 6488
rect 27916 6448 27956 6488
rect 28396 6448 28436 6488
rect 28876 6448 28916 6488
rect 29356 6434 29396 6474
rect 29836 6448 29876 6488
rect 29932 6448 29972 6488
rect 30412 6448 30452 6488
rect 30892 6448 30932 6488
rect 31420 6438 31460 6478
rect 33004 6448 33044 6488
rect 33100 6448 33140 6488
rect 33580 6448 33620 6488
rect 34060 6448 34100 6488
rect 3532 6364 3572 6404
rect 16588 6364 16628 6404
rect 24556 6364 24596 6404
rect 28300 6364 28340 6404
rect 30316 6364 30356 6404
rect 31756 6364 31796 6404
rect 32140 6364 32180 6404
rect 32716 6364 32756 6404
rect 33484 6364 33524 6404
rect 34588 6406 34628 6446
rect 35116 6448 35156 6488
rect 35212 6448 35252 6488
rect 35596 6448 35636 6488
rect 36172 6448 36212 6488
rect 35692 6406 35732 6446
rect 36652 6434 36692 6474
rect 37708 6448 37748 6488
rect 37804 6448 37844 6488
rect 38188 6448 38228 6488
rect 38284 6448 38324 6488
rect 38764 6448 38804 6488
rect 39244 6443 39284 6483
rect 37228 6364 37268 6404
rect 39820 6364 39860 6404
rect 40396 6364 40436 6404
rect 40876 6364 40916 6404
rect 41260 6364 41300 6404
rect 2668 6280 2708 6320
rect 5452 6280 5492 6320
rect 40012 6280 40052 6320
rect 40204 6280 40244 6320
rect 41452 6280 41492 6320
rect 7948 6196 7988 6236
rect 10444 6196 10484 6236
rect 32332 6196 32372 6236
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 33928 6028 33968 6068
rect 34010 6028 34050 6068
rect 34092 6028 34132 6068
rect 34174 6028 34214 6068
rect 34256 6028 34296 6068
rect 2764 5860 2804 5900
rect 9772 5860 9812 5900
rect 10540 5860 10580 5900
rect 11500 5860 11540 5900
rect 11884 5860 11924 5900
rect 12268 5860 12308 5900
rect 13228 5860 13268 5900
rect 13804 5860 13844 5900
rect 17932 5860 17972 5900
rect 19564 5860 19604 5900
rect 21196 5860 21236 5900
rect 22828 5860 22868 5900
rect 25804 5860 25844 5900
rect 27532 5860 27572 5900
rect 27724 5860 27764 5900
rect 29356 5860 29396 5900
rect 31660 5860 31700 5900
rect 34924 5860 34964 5900
rect 37036 5860 37076 5900
rect 38188 5860 38228 5900
rect 38572 5860 38612 5900
rect 41068 5860 41108 5900
rect 11212 5776 11252 5816
rect 41452 5776 41492 5816
rect 11692 5692 11732 5732
rect 12076 5692 12116 5732
rect 12460 5692 12500 5732
rect 13420 5692 13460 5732
rect 13612 5692 13652 5732
rect 16300 5692 16340 5732
rect 31084 5692 31124 5732
rect 31468 5692 31508 5732
rect 35212 5692 35252 5732
rect 37420 5692 37460 5732
rect 37612 5692 37652 5732
rect 37996 5692 38036 5732
rect 38380 5692 38420 5732
rect 39340 5692 39380 5732
rect 39436 5692 39476 5732
rect 40876 5692 40916 5732
rect 41260 5692 41300 5732
rect 1324 5608 1364 5648
rect 2572 5608 2612 5648
rect 3244 5587 3284 5627
rect 3340 5608 3380 5648
rect 3436 5608 3476 5648
rect 3724 5608 3764 5648
rect 3820 5608 3860 5648
rect 3916 5608 3956 5648
rect 4012 5608 4052 5648
rect 4204 5608 4244 5648
rect 4300 5608 4340 5648
rect 4684 5608 4724 5648
rect 4780 5608 4820 5648
rect 4876 5608 4916 5648
rect 5164 5608 5204 5648
rect 6412 5608 6452 5648
rect 6796 5608 6836 5648
rect 8044 5608 8084 5648
rect 8524 5608 8564 5648
rect 8620 5608 8660 5648
rect 9100 5608 9140 5648
rect 9388 5608 9428 5648
rect 9998 5623 10038 5663
rect 10156 5608 10196 5648
rect 10252 5608 10292 5648
rect 10444 5608 10484 5648
rect 10540 5608 10580 5648
rect 10828 5608 10868 5648
rect 10924 5608 10964 5648
rect 13996 5608 14036 5648
rect 15244 5608 15284 5648
rect 16492 5608 16532 5648
rect 17740 5608 17780 5648
rect 18124 5608 18164 5648
rect 19372 5608 19412 5648
rect 19756 5608 19796 5648
rect 21004 5608 21044 5648
rect 21388 5608 21428 5648
rect 22636 5608 22676 5648
rect 24364 5608 24404 5648
rect 25612 5608 25652 5648
rect 26092 5608 26132 5648
rect 27340 5608 27380 5648
rect 27916 5608 27956 5648
rect 29164 5608 29204 5648
rect 29548 5608 29588 5648
rect 30796 5608 30836 5648
rect 31852 5608 31892 5648
rect 33100 5608 33140 5648
rect 33484 5608 33524 5648
rect 34732 5608 34772 5648
rect 35596 5608 35636 5648
rect 36844 5608 36884 5648
rect 38860 5608 38900 5648
rect 38956 5608 38996 5648
rect 39916 5608 39956 5648
rect 40396 5613 40436 5653
rect 8236 5524 8276 5564
rect 9484 5524 9524 5564
rect 40588 5524 40628 5564
rect 3532 5440 3572 5480
rect 4492 5440 4532 5480
rect 4972 5440 5012 5480
rect 6604 5440 6644 5480
rect 8812 5440 8852 5480
rect 15436 5440 15476 5480
rect 16108 5440 16148 5480
rect 31276 5440 31316 5480
rect 33292 5440 33332 5480
rect 35404 5440 35444 5480
rect 37228 5440 37268 5480
rect 37804 5440 37844 5480
rect 10732 5382 10772 5422
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 35168 5272 35208 5312
rect 35250 5272 35290 5312
rect 35332 5272 35372 5312
rect 35414 5272 35454 5312
rect 35496 5272 35536 5312
rect 4684 5104 4724 5144
rect 10444 5104 10484 5144
rect 20620 5104 20660 5144
rect 37228 5104 37268 5144
rect 40972 5104 41012 5144
rect 2668 5020 2708 5060
rect 9004 5020 9044 5060
rect 12076 5020 12116 5060
rect 14092 5020 14132 5060
rect 16492 5020 16532 5060
rect 16780 5020 16820 5060
rect 25516 5020 25556 5060
rect 30892 5020 30932 5060
rect 37420 5020 37460 5060
rect 1228 4936 1268 4976
rect 2476 4936 2516 4976
rect 2956 4936 2996 4976
rect 3052 4936 3092 4976
rect 4012 4936 4052 4976
rect 4492 4931 4532 4971
rect 5164 4936 5204 4976
rect 6412 4936 6452 4976
rect 6796 4936 6836 4976
rect 6988 4936 7028 4976
rect 7276 4936 7316 4976
rect 7372 4936 7412 4976
rect 8332 4936 8372 4976
rect 8812 4931 8852 4971
rect 9292 4936 9332 4976
rect 9580 4936 9620 4976
rect 9676 4936 9716 4976
rect 10156 4936 10196 4976
rect 10252 4936 10292 4976
rect 10636 4936 10676 4976
rect 11884 4936 11924 4976
rect 12364 4936 12404 4976
rect 12460 4936 12500 4976
rect 13420 4936 13460 4976
rect 13900 4922 13940 4962
rect 14764 4936 14804 4976
rect 14860 4936 14900 4976
rect 15340 4936 15380 4976
rect 15820 4936 15860 4976
rect 16300 4922 16340 4962
rect 16972 4922 17012 4962
rect 17452 4936 17492 4976
rect 17932 4936 17972 4976
rect 18412 4936 18452 4976
rect 18508 4936 18548 4976
rect 19180 4936 19220 4976
rect 20428 4936 20468 4976
rect 21676 4936 21716 4976
rect 22924 4936 22964 4976
rect 23788 4936 23828 4976
rect 23884 4936 23924 4976
rect 24268 4936 24308 4976
rect 24364 4936 24404 4976
rect 24844 4936 24884 4976
rect 25900 4936 25940 4976
rect 27148 4936 27188 4976
rect 27916 4936 27956 4976
rect 28876 4936 28916 4976
rect 29164 4936 29204 4976
rect 3436 4852 3476 4892
rect 3532 4852 3572 4892
rect 7756 4852 7796 4892
rect 7852 4852 7892 4892
rect 12844 4852 12884 4892
rect 12940 4852 12980 4892
rect 15244 4852 15284 4892
rect 25372 4894 25412 4934
rect 29260 4936 29300 4976
rect 29740 4936 29780 4976
rect 30220 4936 30260 4976
rect 30700 4922 30740 4962
rect 31276 4936 31316 4976
rect 32524 4936 32564 4976
rect 33292 4936 33332 4976
rect 34540 4936 34580 4976
rect 35500 4936 35540 4976
rect 35596 4936 35636 4976
rect 36556 4936 36596 4976
rect 37084 4926 37124 4966
rect 37612 4936 37652 4976
rect 38860 4936 38900 4976
rect 40780 4936 40820 4976
rect 18028 4852 18068 4892
rect 18796 4852 18836 4892
rect 23500 4852 23540 4892
rect 27436 4852 27476 4892
rect 29644 4852 29684 4892
rect 33100 4852 33140 4892
rect 35116 4852 35156 4892
rect 35980 4852 36020 4892
rect 39532 4894 39572 4934
rect 36076 4852 36116 4892
rect 39148 4852 39188 4892
rect 41164 4852 41204 4892
rect 41740 4852 41780 4892
rect 9964 4768 10004 4808
rect 18988 4768 19028 4808
rect 23308 4768 23348 4808
rect 25708 4768 25748 4808
rect 34924 4768 34964 4808
rect 39340 4768 39380 4808
rect 41356 4768 41396 4808
rect 6604 4684 6644 4724
rect 6796 4684 6836 4724
rect 23116 4684 23156 4724
rect 27628 4684 27668 4724
rect 32716 4684 32756 4724
rect 32908 4684 32948 4724
rect 34732 4684 34772 4724
rect 41548 4684 41588 4724
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 33928 4516 33968 4556
rect 34010 4516 34050 4556
rect 34092 4516 34132 4556
rect 34174 4516 34214 4556
rect 34256 4516 34296 4556
rect 2764 4348 2804 4388
rect 4876 4348 4916 4388
rect 5260 4348 5300 4388
rect 6892 4348 6932 4388
rect 7852 4348 7892 4388
rect 8812 4348 8852 4388
rect 9004 4348 9044 4388
rect 13612 4348 13652 4388
rect 16492 4348 16532 4388
rect 17068 4348 17108 4388
rect 18892 4348 18932 4388
rect 28588 4348 28628 4388
rect 30412 4348 30452 4388
rect 41548 4348 41588 4388
rect 14668 4180 14708 4220
rect 14764 4180 14804 4220
rect 16300 4180 16340 4220
rect 17260 4180 17300 4220
rect 20236 4180 20276 4220
rect 20332 4180 20372 4220
rect 21868 4180 21908 4220
rect 21964 4180 22004 4220
rect 1324 4096 1364 4136
rect 2572 4096 2612 4136
rect 2956 4096 2996 4136
rect 3052 4096 3092 4136
rect 3148 4096 3188 4136
rect 3436 4096 3476 4136
rect 4684 4096 4724 4136
rect 5068 4096 5108 4136
rect 5260 4096 5300 4136
rect 5356 4096 5396 4136
rect 5548 4096 5588 4136
rect 5644 4096 5684 4136
rect 5836 4096 5876 4136
rect 6220 4096 6260 4136
rect 6508 4096 6548 4136
rect 6604 4096 6644 4136
rect 7180 4096 7220 4136
rect 7468 4096 7508 4136
rect 7564 4096 7604 4136
rect 8140 4096 8180 4136
rect 8428 4096 8468 4136
rect 8524 4096 8564 4136
rect 9388 4096 9428 4136
rect 9676 4096 9716 4136
rect 10060 4096 10100 4136
rect 10348 4096 10388 4136
rect 10540 4096 10580 4136
rect 11788 4096 11828 4136
rect 12172 4096 12212 4136
rect 13420 4096 13460 4136
rect 14188 4096 14228 4136
rect 14284 4096 14324 4136
rect 15244 4096 15284 4136
rect 15724 4110 15764 4150
rect 17452 4096 17492 4136
rect 18700 4096 18740 4136
rect 19276 4101 19316 4141
rect 19756 4096 19796 4136
rect 20716 4096 20756 4136
rect 20812 4096 20852 4136
rect 21388 4096 21428 4136
rect 22972 4138 23012 4178
rect 25132 4180 25172 4220
rect 27148 4180 27188 4220
rect 27244 4180 27284 4220
rect 30220 4180 30260 4220
rect 31276 4180 31316 4220
rect 33292 4180 33332 4220
rect 21484 4096 21524 4136
rect 22444 4096 22484 4136
rect 24556 4096 24596 4136
rect 24652 4096 24692 4136
rect 25036 4096 25076 4136
rect 25612 4096 25652 4136
rect 26092 4101 26132 4141
rect 26668 4096 26708 4136
rect 26764 4096 26804 4136
rect 27724 4096 27764 4136
rect 28204 4101 28244 4141
rect 28780 4096 28820 4136
rect 30028 4096 30068 4136
rect 30700 4096 30740 4136
rect 30796 4096 30836 4136
rect 31180 4096 31220 4136
rect 31756 4096 31796 4136
rect 32236 4101 32276 4141
rect 32716 4096 32756 4136
rect 32812 4096 32852 4136
rect 34300 4138 34340 4178
rect 36460 4180 36500 4220
rect 36556 4180 36596 4220
rect 38092 4180 38132 4220
rect 38284 4180 38324 4220
rect 39532 4180 39572 4220
rect 39628 4180 39668 4220
rect 40972 4180 41012 4220
rect 41356 4180 41396 4220
rect 33196 4096 33236 4136
rect 33772 4096 33812 4136
rect 35596 4096 35636 4136
rect 35980 4096 36020 4136
rect 36076 4096 36116 4136
rect 37036 4096 37076 4136
rect 37564 4105 37604 4145
rect 39052 4096 39092 4136
rect 39148 4096 39188 4136
rect 40108 4096 40148 4136
rect 40588 4101 40628 4141
rect 9292 4012 9332 4052
rect 19084 4012 19124 4052
rect 23116 4012 23156 4052
rect 32428 4012 32468 4052
rect 34444 4012 34484 4052
rect 40780 4012 40820 4052
rect 3244 3928 3284 3968
rect 5740 3928 5780 3968
rect 10252 3928 10292 3968
rect 11980 3928 12020 3968
rect 15916 3928 15956 3968
rect 26284 3928 26324 3968
rect 28396 3928 28436 3968
rect 35116 3928 35156 3968
rect 37708 3928 37748 3968
rect 37900 3928 37940 3968
rect 38476 3928 38516 3968
rect 41164 3928 41204 3968
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 35168 3760 35208 3800
rect 35250 3760 35290 3800
rect 35332 3760 35372 3800
rect 35414 3760 35454 3800
rect 35496 3760 35536 3800
rect 2764 3592 2804 3632
rect 5260 3592 5300 3632
rect 8332 3592 8372 3632
rect 8908 3592 8948 3632
rect 12364 3592 12404 3632
rect 13996 3592 14036 3632
rect 14188 3592 14228 3632
rect 16204 3592 16244 3632
rect 16396 3592 16436 3632
rect 16780 3592 16820 3632
rect 19852 3592 19892 3632
rect 21484 3592 21524 3632
rect 21676 3592 21716 3632
rect 23980 3592 24020 3632
rect 26956 3592 26996 3632
rect 28588 3592 28628 3632
rect 28780 3592 28820 3632
rect 30412 3592 30452 3632
rect 32044 3592 32084 3632
rect 33676 3592 33716 3632
rect 35692 3592 35732 3632
rect 37612 3592 37652 3632
rect 39724 3592 39764 3632
rect 39916 3592 39956 3632
rect 4396 3508 4436 3548
rect 4684 3508 4724 3548
rect 7372 3508 7412 3548
rect 10924 3508 10964 3548
rect 1324 3424 1364 3464
rect 2572 3424 2612 3464
rect 2956 3424 2996 3464
rect 4204 3424 4244 3464
rect 4588 3424 4628 3464
rect 4780 3424 4820 3464
rect 4972 3424 5012 3464
rect 5068 3424 5108 3464
rect 5548 3424 5588 3464
rect 5932 3424 5972 3464
rect 6124 3424 6164 3464
rect 6220 3424 6260 3464
rect 6412 3424 6452 3464
rect 6700 3424 6740 3464
rect 6988 3424 7028 3464
rect 7276 3424 7316 3464
rect 7852 3424 7892 3464
rect 7948 3424 7988 3464
rect 8044 3424 8084 3464
rect 8140 3424 8180 3464
rect 8332 3424 8372 3464
rect 8524 3424 8564 3464
rect 8620 3424 8660 3464
rect 8812 3424 8852 3464
rect 9196 3424 9236 3464
rect 9292 3424 9332 3464
rect 10251 3433 10291 3473
rect 10732 3410 10772 3450
rect 11212 3424 11252 3464
rect 11500 3424 11540 3464
rect 11596 3424 11636 3464
rect 12076 3424 12116 3464
rect 12172 3424 12212 3464
rect 12556 3424 12596 3464
rect 14764 3424 14804 3464
rect 16012 3424 16052 3464
rect 16972 3424 17012 3464
rect 18220 3424 18260 3464
rect 18412 3424 18452 3464
rect 19660 3424 19700 3464
rect 20044 3424 20084 3464
rect 21292 3424 21332 3464
rect 22540 3424 22580 3464
rect 23788 3424 23828 3464
rect 25516 3424 25556 3464
rect 26764 3424 26804 3464
rect 27148 3424 27188 3464
rect 28396 3424 28436 3464
rect 28972 3424 29012 3464
rect 30220 3424 30260 3464
rect 30604 3424 30644 3464
rect 31852 3424 31892 3464
rect 32236 3424 32276 3464
rect 33484 3424 33524 3464
rect 34252 3424 34292 3464
rect 35500 3424 35540 3464
rect 36172 3424 36212 3464
rect 37420 3424 37460 3464
rect 38284 3424 38324 3464
rect 39532 3424 39572 3464
rect 40108 3424 40148 3464
rect 41356 3424 41396 3464
rect 9676 3340 9716 3380
rect 13804 3382 13844 3422
rect 9772 3340 9812 3380
rect 14380 3340 14420 3380
rect 16588 3340 16628 3380
rect 21868 3340 21908 3380
rect 24364 3340 24404 3380
rect 24748 3340 24788 3380
rect 25132 3340 25172 3380
rect 33868 3340 33908 3380
rect 38092 3340 38132 3380
rect 5548 3256 5588 3296
rect 11884 3256 11924 3296
rect 24940 3256 24980 3296
rect 25324 3256 25364 3296
rect 41548 3256 41588 3296
rect 2764 3172 2804 3212
rect 5740 3172 5780 3212
rect 5932 3172 5972 3212
rect 6700 3172 6740 3212
rect 7660 3172 7700 3212
rect 24556 3172 24596 3212
rect 37900 3172 37940 3212
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 33928 3004 33968 3044
rect 34010 3004 34050 3044
rect 34092 3004 34132 3044
rect 34174 3004 34214 3044
rect 34256 3004 34296 3044
rect 2956 2836 2996 2876
rect 6220 2836 6260 2876
rect 9964 2836 10004 2876
rect 13900 2836 13940 2876
rect 16300 2836 16340 2876
rect 26668 2836 26708 2876
rect 29548 2836 29588 2876
rect 30028 2836 30068 2876
rect 31660 2836 31700 2876
rect 32044 2836 32084 2876
rect 36364 2836 36404 2876
rect 36940 2836 36980 2876
rect 37612 2836 37652 2876
rect 6028 2752 6068 2792
rect 41644 2752 41684 2792
rect 4300 2668 4340 2708
rect 4396 2668 4436 2708
rect 1516 2584 1556 2624
rect 2764 2584 2804 2624
rect 3340 2589 3380 2629
rect 3820 2584 3860 2624
rect 4780 2584 4820 2624
rect 5644 2626 5684 2666
rect 7084 2668 7124 2708
rect 7180 2668 7220 2708
rect 10828 2668 10868 2708
rect 14668 2668 14708 2708
rect 14764 2668 14804 2708
rect 16108 2668 16148 2708
rect 17068 2668 17108 2708
rect 17164 2668 17204 2708
rect 19180 2668 19220 2708
rect 21196 2668 21236 2708
rect 21292 2668 21332 2708
rect 23788 2668 23828 2708
rect 23884 2668 23924 2708
rect 27052 2668 27092 2708
rect 28012 2668 28052 2708
rect 28108 2668 28148 2708
rect 29740 2668 29780 2708
rect 31852 2668 31892 2708
rect 32236 2668 32276 2708
rect 33292 2668 33332 2708
rect 33388 2668 33428 2708
rect 36556 2668 36596 2708
rect 37132 2668 37172 2708
rect 4876 2584 4916 2624
rect 5356 2584 5396 2624
rect 5740 2584 5780 2624
rect 6316 2584 6356 2624
rect 6604 2584 6644 2624
rect 6700 2584 6740 2624
rect 7660 2584 7700 2624
rect 8140 2589 8180 2629
rect 8524 2584 8564 2624
rect 9772 2584 9812 2624
rect 10252 2584 10292 2624
rect 10348 2584 10388 2624
rect 10732 2584 10772 2624
rect 11308 2584 11348 2624
rect 11788 2589 11828 2629
rect 12268 2584 12308 2624
rect 12460 2584 12500 2624
rect 13708 2584 13748 2624
rect 14188 2584 14228 2624
rect 14284 2584 14324 2624
rect 15244 2584 15284 2624
rect 15724 2589 15764 2629
rect 16588 2584 16628 2624
rect 16684 2584 16724 2624
rect 17644 2584 17684 2624
rect 18124 2589 18164 2629
rect 18700 2584 18740 2624
rect 18796 2584 18836 2624
rect 19276 2584 19316 2624
rect 19756 2584 19796 2624
rect 20284 2593 20324 2633
rect 20716 2584 20756 2624
rect 20812 2584 20852 2624
rect 21772 2584 21812 2624
rect 22300 2593 22340 2633
rect 23308 2584 23348 2624
rect 23404 2584 23444 2624
rect 24364 2584 24404 2624
rect 24844 2589 24884 2629
rect 25228 2584 25268 2624
rect 26476 2584 26516 2624
rect 27532 2584 27572 2624
rect 27628 2584 27668 2624
rect 28588 2584 28628 2624
rect 29116 2593 29156 2633
rect 30220 2584 30260 2624
rect 31468 2584 31508 2624
rect 32812 2584 32852 2624
rect 32908 2584 32948 2624
rect 33868 2584 33908 2624
rect 34396 2593 34436 2633
rect 34924 2584 34964 2624
rect 36172 2584 36212 2624
rect 38764 2584 38804 2624
rect 39628 2584 39668 2624
rect 40012 2584 40052 2624
rect 40204 2584 40244 2624
rect 41452 2584 41492 2624
rect 3148 2500 3188 2540
rect 15916 2500 15956 2540
rect 18316 2500 18356 2540
rect 25036 2500 25076 2540
rect 29260 2500 29300 2540
rect 8332 2416 8372 2456
rect 11980 2416 12020 2456
rect 12172 2416 12212 2456
rect 20428 2374 20468 2414
rect 22444 2416 22484 2456
rect 27244 2416 27284 2456
rect 34540 2416 34580 2456
rect 36748 2416 36788 2456
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 35168 2248 35208 2288
rect 35250 2248 35290 2288
rect 35332 2248 35372 2288
rect 35414 2248 35454 2288
rect 35496 2248 35536 2288
rect 2956 2080 2996 2120
rect 3532 2080 3572 2120
rect 5932 2080 5972 2120
rect 10924 2080 10964 2120
rect 14092 2080 14132 2120
rect 16012 2080 16052 2120
rect 17644 2080 17684 2120
rect 19276 2080 19316 2120
rect 21004 2080 21044 2120
rect 22636 2080 22676 2120
rect 24268 2080 24308 2120
rect 26284 2080 26324 2120
rect 30124 2080 30164 2120
rect 33196 2080 33236 2120
rect 36076 2080 36116 2120
rect 38956 2080 38996 2120
rect 41260 2080 41300 2120
rect 3244 1996 3284 2036
rect 8524 1996 8564 2036
rect 11884 1996 11924 2036
rect 26476 1996 26516 2036
rect 29932 1996 29972 2036
rect 33676 1996 33716 2036
rect 36556 1996 36596 2036
rect 1516 1912 1556 1952
rect 2764 1912 2804 1952
rect 3148 1912 3188 1952
rect 3340 1912 3380 1952
rect 3628 1912 3668 1952
rect 3724 1912 3764 1952
rect 3820 1912 3860 1952
rect 4204 1912 4244 1952
rect 5452 1912 5492 1952
rect 5740 1912 5780 1952
rect 5836 1912 5876 1952
rect 6028 1912 6068 1952
rect 6124 1912 6164 1952
rect 6281 1905 6321 1945
rect 6796 1912 6836 1952
rect 6892 1912 6932 1952
rect 7276 1912 7316 1952
rect 7372 1912 7412 1952
rect 7852 1912 7892 1952
rect 8332 1902 8372 1942
rect 9196 1912 9236 1952
rect 9292 1912 9332 1952
rect 9676 1912 9716 1952
rect 9772 1912 9812 1952
rect 10252 1912 10292 1952
rect 10732 1898 10772 1938
rect 11116 1912 11156 1952
rect 11212 1912 11252 1952
rect 11308 1912 11348 1952
rect 11404 1912 11444 1952
rect 11980 1912 12020 1952
rect 12268 1912 12308 1952
rect 12652 1912 12692 1952
rect 13900 1912 13940 1952
rect 14572 1912 14612 1952
rect 15820 1912 15860 1952
rect 16204 1912 16244 1952
rect 17452 1912 17492 1952
rect 17836 1912 17876 1952
rect 19084 1912 19124 1952
rect 19564 1912 19604 1952
rect 20812 1912 20852 1952
rect 21196 1912 21236 1952
rect 22444 1912 22484 1952
rect 22828 1912 22868 1952
rect 24076 1912 24116 1952
rect 24556 1912 24596 1952
rect 24652 1912 24692 1952
rect 25036 1912 25076 1952
rect 25132 1912 25172 1952
rect 25612 1912 25652 1952
rect 26092 1907 26132 1947
rect 26668 1912 26708 1952
rect 27916 1912 27956 1952
rect 28204 1912 28244 1952
rect 28300 1912 28340 1952
rect 28684 1912 28724 1952
rect 28780 1912 28820 1952
rect 29260 1912 29300 1952
rect 29740 1898 29780 1938
rect 30316 1912 30356 1952
rect 31564 1912 31604 1952
rect 31756 1912 31796 1952
rect 33004 1912 33044 1952
rect 34060 1912 34100 1952
rect 34924 1912 34964 1952
rect 36940 1912 36980 1952
rect 37804 1912 37844 1952
rect 39244 1912 39284 1952
rect 40780 1912 40820 1952
rect 4012 1660 4052 1700
rect 11596 1660 11636 1700
rect 39532 1660 39572 1700
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 33928 1492 33968 1532
rect 34010 1492 34050 1532
rect 34092 1492 34132 1532
rect 34174 1492 34214 1532
rect 34256 1492 34296 1532
rect 3340 1324 3380 1364
rect 11212 1324 11252 1364
rect 20908 1324 20948 1364
rect 24460 1324 24500 1364
rect 27916 1324 27956 1364
rect 29548 1324 29588 1364
rect 31564 1324 31604 1364
rect 41548 1324 41588 1364
rect 5260 1240 5300 1280
rect 7180 1240 7220 1280
rect 9580 1240 9620 1280
rect 11692 1240 11732 1280
rect 13612 1240 13652 1280
rect 15436 1240 15476 1280
rect 17356 1240 17396 1280
rect 19084 1240 19124 1280
rect 22540 1240 22580 1280
rect 24652 1240 24692 1280
rect 27724 1240 27764 1280
rect 32428 1240 32468 1280
rect 32812 1240 32852 1280
rect 34828 1240 34868 1280
rect 36268 1240 36308 1280
rect 36844 1240 36884 1280
rect 40204 1240 40244 1280
rect 40588 1240 40628 1280
rect 13804 1156 13844 1196
rect 32620 1156 32660 1196
rect 33004 1156 33044 1196
rect 35212 1156 35252 1196
rect 39628 1156 39668 1196
rect 40012 1156 40052 1196
rect 41164 1156 41204 1196
rect 41356 1156 41396 1196
rect 1516 1072 1556 1112
rect 1612 1072 1652 1112
rect 1708 1072 1748 1112
rect 1900 1072 1940 1112
rect 3148 1072 3188 1112
rect 3820 1072 3860 1112
rect 5068 1072 5108 1112
rect 5740 1072 5780 1112
rect 5836 1072 5876 1112
rect 6220 1072 6260 1112
rect 6316 1072 6356 1112
rect 6412 1072 6452 1112
rect 6700 1072 6740 1112
rect 6796 1072 6836 1112
rect 6892 1072 6932 1112
rect 6988 1072 7028 1112
rect 7468 1072 7508 1112
rect 7564 1072 7604 1112
rect 7852 1072 7892 1112
rect 8140 1072 8180 1112
rect 9388 1072 9428 1112
rect 9772 1072 9812 1112
rect 11020 1072 11060 1112
rect 11404 1072 11444 1112
rect 11500 1072 11540 1112
rect 11692 1072 11732 1112
rect 11884 1072 11924 1112
rect 11980 1072 12020 1112
rect 12076 1072 12116 1112
rect 12364 1072 12404 1112
rect 12460 1072 12500 1112
rect 12556 1072 12596 1112
rect 12652 1072 12692 1112
rect 12844 1072 12884 1112
rect 12940 1072 12980 1112
rect 13036 1072 13076 1112
rect 13132 1072 13172 1112
rect 13996 1072 14036 1112
rect 15244 1072 15284 1112
rect 15916 1072 15956 1112
rect 17164 1072 17204 1112
rect 17644 1072 17684 1112
rect 18892 1072 18932 1112
rect 19468 1072 19508 1112
rect 20716 1072 20756 1112
rect 21100 1072 21140 1112
rect 22348 1072 22388 1112
rect 23020 1072 23060 1112
rect 24268 1072 24308 1112
rect 24844 1072 24884 1112
rect 26092 1072 26132 1112
rect 26284 1072 26324 1112
rect 27532 1072 27572 1112
rect 28108 1072 28148 1112
rect 29356 1072 29396 1112
rect 29740 1072 29780 1112
rect 30988 1072 31028 1112
rect 31276 1072 31316 1112
rect 33388 1072 33428 1112
rect 34636 1072 34676 1112
rect 35596 1072 35636 1112
rect 36556 1072 36596 1112
rect 37996 1072 38036 1112
rect 38860 1072 38900 1112
rect 39244 1072 39284 1112
rect 1420 904 1460 944
rect 6028 904 6068 944
rect 6508 904 6548 944
rect 12172 904 12212 944
rect 35020 904 35060 944
rect 39436 904 39476 944
rect 39820 904 39860 944
rect 40972 904 41012 944
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 35168 736 35208 776
rect 35250 736 35290 776
rect 35332 736 35372 776
rect 35414 736 35454 776
rect 35496 736 35536 776
<< metal2 >>
rect 9464 10672 9544 10752
rect 9656 10672 9736 10752
rect 9848 10672 9928 10752
rect 10040 10672 10120 10752
rect 10232 10672 10312 10752
rect 10424 10672 10504 10752
rect 10616 10672 10696 10752
rect 10808 10672 10888 10752
rect 11000 10672 11080 10752
rect 11192 10672 11272 10752
rect 11384 10672 11464 10752
rect 11576 10672 11656 10752
rect 11768 10672 11848 10752
rect 11960 10672 12040 10752
rect 12152 10672 12232 10752
rect 12344 10672 12424 10752
rect 12536 10672 12616 10752
rect 12728 10672 12808 10752
rect 12920 10672 13000 10752
rect 13112 10672 13192 10752
rect 13304 10672 13384 10752
rect 13496 10672 13576 10752
rect 13688 10672 13768 10752
rect 13880 10672 13960 10752
rect 14072 10672 14152 10752
rect 14264 10672 14344 10752
rect 14456 10672 14536 10752
rect 14648 10672 14728 10752
rect 14840 10672 14920 10752
rect 15032 10672 15112 10752
rect 15224 10672 15304 10752
rect 15416 10672 15496 10752
rect 15608 10672 15688 10752
rect 15800 10672 15880 10752
rect 15992 10672 16072 10752
rect 16184 10672 16264 10752
rect 16376 10672 16456 10752
rect 16568 10672 16648 10752
rect 16760 10672 16840 10752
rect 16952 10672 17032 10752
rect 17144 10672 17224 10752
rect 17336 10672 17416 10752
rect 17528 10672 17608 10752
rect 17720 10672 17800 10752
rect 17912 10672 17992 10752
rect 18104 10672 18184 10752
rect 18296 10672 18376 10752
rect 18488 10672 18568 10752
rect 18680 10672 18760 10752
rect 18872 10672 18952 10752
rect 19064 10672 19144 10752
rect 19256 10672 19336 10752
rect 19448 10672 19528 10752
rect 19640 10672 19720 10752
rect 19832 10672 19912 10752
rect 20024 10672 20104 10752
rect 20216 10688 20296 10752
rect 20216 10672 20236 10688
rect 1707 10520 1749 10529
rect 1707 10480 1708 10520
rect 1748 10480 1749 10520
rect 1707 10471 1749 10480
rect 1611 10184 1653 10193
rect 1611 10144 1612 10184
rect 1652 10144 1653 10184
rect 1611 10135 1653 10144
rect 1612 9512 1652 10135
rect 1612 8933 1652 9472
rect 1611 8924 1653 8933
rect 1611 8884 1612 8924
rect 1652 8884 1653 8924
rect 1611 8875 1653 8884
rect 1708 8429 1748 10471
rect 4683 9848 4725 9857
rect 4683 9808 4684 9848
rect 4724 9808 4725 9848
rect 4683 9799 4725 9808
rect 4928 9848 5296 9857
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 4928 9799 5296 9808
rect 2860 9640 3188 9680
rect 2860 9512 2900 9640
rect 2860 9463 2900 9472
rect 2955 9512 2997 9521
rect 2955 9472 2956 9512
rect 2996 9472 2997 9512
rect 2955 9463 2997 9472
rect 2956 9008 2996 9463
rect 3148 9344 3188 9640
rect 3244 9596 3284 9607
rect 3244 9521 3284 9556
rect 3243 9512 3285 9521
rect 3436 9512 3476 9521
rect 3243 9472 3244 9512
rect 3284 9472 3285 9512
rect 3243 9463 3285 9472
rect 3340 9472 3436 9512
rect 3340 9344 3380 9472
rect 3436 9463 3476 9472
rect 4684 9512 4724 9799
rect 6412 9680 6452 9689
rect 7660 9680 7700 9689
rect 9004 9680 9044 9689
rect 6452 9640 6932 9680
rect 6412 9631 6452 9640
rect 4876 9512 4916 9521
rect 3148 9304 3380 9344
rect 3435 9344 3477 9353
rect 3435 9304 3436 9344
rect 3476 9304 3477 9344
rect 2860 8968 2996 9008
rect 3052 9260 3092 9269
rect 2860 8765 2900 8968
rect 2091 8756 2133 8765
rect 2091 8716 2092 8756
rect 2132 8716 2133 8756
rect 2091 8707 2133 8716
rect 2859 8756 2901 8765
rect 2859 8716 2860 8756
rect 2900 8716 2901 8756
rect 2859 8707 2901 8716
rect 1900 8672 1940 8681
rect 1804 8504 1844 8513
rect 1707 8420 1749 8429
rect 1707 8380 1708 8420
rect 1748 8380 1749 8420
rect 1707 8371 1749 8380
rect 1323 8168 1365 8177
rect 1323 8128 1324 8168
rect 1364 8128 1365 8168
rect 1323 8119 1365 8128
rect 1324 7328 1364 8119
rect 1708 7832 1748 8371
rect 1804 8009 1844 8464
rect 1900 8177 1940 8632
rect 1996 8672 2036 8681
rect 1996 8504 2036 8632
rect 2092 8672 2132 8707
rect 2092 8621 2132 8632
rect 2476 8672 2516 8681
rect 2284 8504 2324 8513
rect 1996 8464 2284 8504
rect 2284 8455 2324 8464
rect 1899 8168 1941 8177
rect 1899 8128 1900 8168
rect 1940 8128 1941 8168
rect 1899 8119 1941 8128
rect 1803 8000 1845 8009
rect 1803 7960 1804 8000
rect 1844 7960 1845 8000
rect 1803 7951 1845 7960
rect 1900 8000 1940 8009
rect 1900 7832 1940 7960
rect 1708 7792 1940 7832
rect 1707 7580 1749 7589
rect 1707 7540 1708 7580
rect 1748 7540 1749 7580
rect 1707 7531 1749 7540
rect 1228 7288 1364 7328
rect 1131 6488 1173 6497
rect 1131 6448 1132 6488
rect 1172 6448 1173 6488
rect 1131 6439 1173 6448
rect 1228 6488 1268 7288
rect 1228 6439 1268 6448
rect 1324 7160 1364 7169
rect 1132 5573 1172 6439
rect 1324 6320 1364 7120
rect 1516 7160 1556 7169
rect 1419 6992 1461 7001
rect 1419 6952 1420 6992
rect 1460 6952 1461 6992
rect 1419 6943 1461 6952
rect 1420 6858 1460 6943
rect 1516 6320 1556 7120
rect 1708 7160 1748 7531
rect 1803 7412 1845 7421
rect 1803 7372 1804 7412
rect 1844 7372 1845 7412
rect 1803 7363 1845 7372
rect 1708 7111 1748 7120
rect 1324 6280 1460 6320
rect 1516 6280 1748 6320
rect 1323 5984 1365 5993
rect 1323 5944 1324 5984
rect 1364 5944 1365 5984
rect 1323 5935 1365 5944
rect 1324 5648 1364 5935
rect 1324 5599 1364 5608
rect 1131 5564 1173 5573
rect 1131 5524 1132 5564
rect 1172 5524 1173 5564
rect 1131 5515 1173 5524
rect 1323 5480 1365 5489
rect 1323 5440 1324 5480
rect 1364 5440 1365 5480
rect 1323 5431 1365 5440
rect 1324 5237 1364 5431
rect 1323 5228 1365 5237
rect 1323 5188 1324 5228
rect 1364 5188 1365 5228
rect 1323 5179 1365 5188
rect 1228 4976 1268 4985
rect 1324 4976 1364 5179
rect 1268 4936 1364 4976
rect 1228 4927 1268 4936
rect 1131 4472 1173 4481
rect 1131 4432 1132 4472
rect 1172 4432 1173 4472
rect 1131 4423 1173 4432
rect 1132 2549 1172 4423
rect 1323 4136 1365 4145
rect 1323 4096 1324 4136
rect 1364 4096 1365 4136
rect 1323 4087 1365 4096
rect 1324 4002 1364 4087
rect 1420 3641 1460 6280
rect 1419 3632 1461 3641
rect 1419 3592 1420 3632
rect 1460 3592 1461 3632
rect 1419 3583 1461 3592
rect 1323 3464 1365 3473
rect 1323 3424 1324 3464
rect 1364 3424 1365 3464
rect 1323 3415 1365 3424
rect 1324 2801 1364 3415
rect 1323 2792 1365 2801
rect 1323 2752 1324 2792
rect 1364 2752 1365 2792
rect 1323 2743 1365 2752
rect 1131 2540 1173 2549
rect 1131 2500 1132 2540
rect 1172 2500 1173 2540
rect 1131 2491 1173 2500
rect 1420 1112 1460 3583
rect 1515 3380 1557 3389
rect 1515 3340 1516 3380
rect 1556 3340 1557 3380
rect 1515 3331 1557 3340
rect 1516 2624 1556 3331
rect 1556 2584 1652 2624
rect 1516 2575 1556 2584
rect 1515 2036 1557 2045
rect 1515 1996 1516 2036
rect 1556 1996 1557 2036
rect 1515 1987 1557 1996
rect 1516 1952 1556 1987
rect 1516 1901 1556 1912
rect 1612 1373 1652 2584
rect 1708 2129 1748 6280
rect 1804 5993 1844 7363
rect 2476 7085 2516 8632
rect 2571 8672 2613 8681
rect 2571 8632 2572 8672
rect 2612 8632 2613 8672
rect 2571 8623 2613 8632
rect 2860 8672 2900 8707
rect 3052 8681 3092 9220
rect 2572 8538 2612 8623
rect 2860 8622 2900 8632
rect 2956 8672 2996 8681
rect 2956 7748 2996 8632
rect 3051 8672 3093 8681
rect 3051 8632 3052 8672
rect 3092 8632 3093 8672
rect 3051 8623 3093 8632
rect 3148 8261 3188 9304
rect 3435 9295 3477 9304
rect 3340 8672 3380 8681
rect 3244 8632 3340 8672
rect 3147 8252 3189 8261
rect 3147 8212 3148 8252
rect 3188 8212 3189 8252
rect 3147 8203 3189 8212
rect 3148 8000 3188 8203
rect 3051 7748 3093 7757
rect 2956 7708 3052 7748
rect 3092 7708 3093 7748
rect 3051 7699 3093 7708
rect 2955 7328 2997 7337
rect 2955 7288 2956 7328
rect 2996 7288 2997 7328
rect 2955 7279 2997 7288
rect 2956 7160 2996 7279
rect 2956 7111 2996 7120
rect 2475 7076 2517 7085
rect 2475 7036 2476 7076
rect 2516 7036 2517 7076
rect 2475 7027 2517 7036
rect 2476 6488 2516 6497
rect 2955 6488 2997 6497
rect 1803 5984 1845 5993
rect 1803 5944 1804 5984
rect 1844 5944 1845 5984
rect 1803 5935 1845 5944
rect 2476 5648 2516 6448
rect 2764 6448 2956 6488
rect 2996 6448 2997 6488
rect 2667 6320 2709 6329
rect 2667 6280 2668 6320
rect 2708 6280 2709 6320
rect 2667 6271 2709 6280
rect 2668 6186 2708 6271
rect 2764 5900 2804 6448
rect 2955 6439 2997 6448
rect 3052 6488 3092 7699
rect 3148 7337 3188 7960
rect 3147 7328 3189 7337
rect 3147 7288 3148 7328
rect 3188 7288 3189 7328
rect 3147 7279 3189 7288
rect 3147 7160 3189 7169
rect 3147 7120 3148 7160
rect 3188 7120 3189 7160
rect 3147 7111 3189 7120
rect 3148 7076 3188 7111
rect 3148 7025 3188 7036
rect 2956 6354 2996 6439
rect 2764 5851 2804 5860
rect 2859 5732 2901 5741
rect 2859 5692 2860 5732
rect 2900 5692 2901 5732
rect 2859 5683 2901 5692
rect 2572 5648 2612 5657
rect 2476 5608 2572 5648
rect 2283 5396 2325 5405
rect 2283 5356 2284 5396
rect 2324 5356 2325 5396
rect 2283 5347 2325 5356
rect 2284 3137 2324 5347
rect 2476 4976 2516 5608
rect 2572 5599 2612 5608
rect 2668 5060 2708 5071
rect 2668 4985 2708 5020
rect 2476 4136 2516 4936
rect 2667 4976 2709 4985
rect 2667 4936 2668 4976
rect 2708 4936 2709 4976
rect 2667 4927 2709 4936
rect 2763 4892 2805 4901
rect 2763 4852 2764 4892
rect 2804 4852 2805 4892
rect 2763 4843 2805 4852
rect 2764 4388 2804 4843
rect 2764 4339 2804 4348
rect 2860 4220 2900 5683
rect 2956 5069 2996 5100
rect 2955 5060 2997 5069
rect 2955 5020 2956 5060
rect 2996 5020 2997 5060
rect 2955 5011 2997 5020
rect 2956 4976 2996 5011
rect 2956 4901 2996 4936
rect 3052 4976 3092 6448
rect 3244 6404 3284 8632
rect 3340 8623 3380 8632
rect 3436 8672 3476 9295
rect 3688 9092 4056 9101
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 3688 9043 4056 9052
rect 4684 9017 4724 9472
rect 4780 9472 4876 9512
rect 4683 9008 4725 9017
rect 4683 8968 4684 9008
rect 4724 8968 4725 9008
rect 4683 8959 4725 8968
rect 4780 8849 4820 9472
rect 4876 9463 4916 9472
rect 4971 9512 5013 9521
rect 4971 9472 4972 9512
rect 5012 9472 5013 9512
rect 4971 9463 5013 9472
rect 5068 9512 5108 9521
rect 4972 9378 5012 9463
rect 4875 9176 4917 9185
rect 4875 9136 4876 9176
rect 4916 9136 4917 9176
rect 4875 9127 4917 9136
rect 3819 8840 3861 8849
rect 3819 8800 3820 8840
rect 3860 8800 3861 8840
rect 3819 8791 3861 8800
rect 4779 8840 4821 8849
rect 4779 8800 4780 8840
rect 4820 8800 4821 8840
rect 4779 8791 4821 8800
rect 3339 8168 3381 8177
rect 3339 8128 3340 8168
rect 3380 8128 3381 8168
rect 3339 8119 3381 8128
rect 3340 8034 3380 8119
rect 3436 7328 3476 8632
rect 3820 8177 3860 8791
rect 4011 8756 4053 8765
rect 4011 8716 4012 8756
rect 4052 8716 4053 8756
rect 4011 8707 4053 8716
rect 3916 8672 3956 8683
rect 3916 8597 3956 8632
rect 3915 8588 3957 8597
rect 3915 8548 3916 8588
rect 3956 8548 3957 8588
rect 3915 8539 3957 8548
rect 3819 8168 3861 8177
rect 4012 8168 4052 8707
rect 4396 8681 4436 8686
rect 4395 8677 4437 8681
rect 4395 8632 4396 8677
rect 4436 8632 4437 8677
rect 4395 8623 4437 8632
rect 4780 8672 4820 8681
rect 4876 8672 4916 9127
rect 5068 8681 5108 9472
rect 5164 9512 5204 9521
rect 5164 9260 5204 9472
rect 5931 9512 5973 9521
rect 6220 9512 6260 9521
rect 6604 9512 6644 9521
rect 5931 9472 5932 9512
rect 5972 9472 5973 9512
rect 5931 9463 5973 9472
rect 6124 9472 6220 9512
rect 5164 9220 5492 9260
rect 4820 8632 4916 8672
rect 5067 8672 5109 8681
rect 5067 8632 5068 8672
rect 5108 8632 5109 8672
rect 4780 8623 4820 8632
rect 5067 8623 5109 8632
rect 4396 8542 4436 8623
rect 4588 8504 4628 8513
rect 4628 8464 4724 8504
rect 4588 8455 4628 8464
rect 3819 8128 3820 8168
rect 3860 8128 3861 8168
rect 3819 8119 3861 8128
rect 3915 8128 4052 8168
rect 4108 8210 4148 8219
rect 4108 8168 4148 8170
rect 4108 8128 4532 8168
rect 3915 8010 3955 8128
rect 3819 8000 3861 8009
rect 3819 7960 3820 8000
rect 3860 7960 3861 8000
rect 3915 8001 3956 8010
rect 3915 7961 3916 8001
rect 3915 7960 3956 7961
rect 3819 7951 3861 7960
rect 3916 7952 3956 7960
rect 4299 8000 4341 8009
rect 4299 7960 4300 8000
rect 4340 7960 4341 8000
rect 4299 7951 4341 7960
rect 4396 8000 4436 8009
rect 3820 7866 3860 7951
rect 4300 7866 4340 7951
rect 4396 7832 4436 7960
rect 4492 8000 4532 8128
rect 4588 8009 4628 8094
rect 4492 7951 4532 7960
rect 4587 8000 4629 8009
rect 4587 7960 4588 8000
rect 4628 7960 4629 8000
rect 4587 7951 4629 7960
rect 4684 7832 4724 8464
rect 4928 8336 5296 8345
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 4928 8287 5296 8296
rect 4779 8084 4821 8093
rect 4779 8044 4780 8084
rect 4820 8044 4821 8084
rect 4779 8035 4821 8044
rect 4780 8000 4820 8035
rect 4780 7949 4820 7960
rect 4396 7792 4724 7832
rect 3688 7580 4056 7589
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 3688 7531 4056 7540
rect 4587 7580 4629 7589
rect 4587 7540 4588 7580
rect 4628 7540 4629 7580
rect 4587 7531 4629 7540
rect 3340 7288 3476 7328
rect 3819 7328 3861 7337
rect 4203 7328 4245 7337
rect 3819 7288 3820 7328
rect 3860 7288 3861 7328
rect 3340 6740 3380 7288
rect 3819 7279 3861 7288
rect 4108 7288 4204 7328
rect 4244 7288 4245 7328
rect 3436 7160 3476 7169
rect 3436 6917 3476 7120
rect 3531 7160 3573 7169
rect 3531 7120 3532 7160
rect 3572 7120 3573 7160
rect 3531 7111 3573 7120
rect 3628 7160 3668 7169
rect 3532 7026 3572 7111
rect 3435 6908 3477 6917
rect 3435 6868 3436 6908
rect 3476 6868 3477 6908
rect 3435 6859 3477 6868
rect 3340 6700 3572 6740
rect 3436 6488 3476 6497
rect 3339 6404 3381 6413
rect 3436 6404 3476 6448
rect 3244 6364 3340 6404
rect 3380 6364 3476 6404
rect 3532 6404 3572 6700
rect 3628 6497 3668 7120
rect 3820 7085 3860 7279
rect 4108 7160 4148 7288
rect 4203 7279 4245 7288
rect 4108 7111 4148 7120
rect 4203 7160 4245 7169
rect 4588 7160 4628 7531
rect 4203 7120 4204 7160
rect 4244 7120 4532 7160
rect 4203 7111 4245 7120
rect 3819 7076 3861 7085
rect 3819 7036 3820 7076
rect 3860 7036 3861 7076
rect 3819 7027 3861 7036
rect 3724 6992 3764 7001
rect 3627 6488 3669 6497
rect 3627 6448 3628 6488
rect 3668 6448 3669 6488
rect 3627 6439 3669 6448
rect 3339 6355 3381 6364
rect 3532 6320 3572 6364
rect 3436 6280 3572 6320
rect 3436 5825 3476 6280
rect 3628 6236 3668 6439
rect 3724 6245 3764 6952
rect 3820 6413 3860 7027
rect 4204 7026 4244 7111
rect 3916 6992 3956 7001
rect 3819 6404 3861 6413
rect 3819 6364 3820 6404
rect 3860 6364 3861 6404
rect 3819 6355 3861 6364
rect 3532 6196 3668 6236
rect 3723 6236 3765 6245
rect 3723 6196 3724 6236
rect 3764 6196 3765 6236
rect 3916 6236 3956 6952
rect 4011 6488 4053 6497
rect 4011 6448 4012 6488
rect 4052 6448 4053 6488
rect 4011 6439 4053 6448
rect 4492 6483 4532 7120
rect 4588 7111 4628 7120
rect 5355 6992 5397 7001
rect 5355 6952 5356 6992
rect 5396 6952 5397 6992
rect 5355 6943 5397 6952
rect 4928 6824 5296 6833
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 4928 6775 5296 6784
rect 4684 6656 4724 6665
rect 5163 6656 5205 6665
rect 4724 6616 5012 6656
rect 4684 6607 4724 6616
rect 4012 6354 4052 6439
rect 4492 6434 4532 6443
rect 4876 6488 4916 6499
rect 4876 6413 4916 6448
rect 4972 6488 5012 6616
rect 5163 6616 5164 6656
rect 5204 6616 5205 6656
rect 5163 6607 5205 6616
rect 5164 6522 5204 6607
rect 4972 6439 5012 6448
rect 5068 6488 5108 6497
rect 4875 6404 4917 6413
rect 4875 6364 4876 6404
rect 4916 6364 4917 6404
rect 4875 6355 4917 6364
rect 5068 6329 5108 6448
rect 5356 6488 5396 6943
rect 5452 6497 5492 9220
rect 5932 8849 5972 9463
rect 6124 9353 6164 9472
rect 6220 9463 6260 9472
rect 6508 9472 6604 9512
rect 6123 9344 6165 9353
rect 6123 9304 6124 9344
rect 6164 9304 6165 9344
rect 6123 9295 6165 9304
rect 6220 9344 6260 9353
rect 6220 8849 6260 9304
rect 5931 8840 5973 8849
rect 5931 8800 5932 8840
rect 5972 8800 5973 8840
rect 5931 8791 5973 8800
rect 6219 8840 6261 8849
rect 6219 8800 6220 8840
rect 6260 8800 6261 8840
rect 6219 8791 6261 8800
rect 6028 8672 6068 8681
rect 6028 8177 6068 8632
rect 6411 8672 6453 8681
rect 6411 8632 6412 8672
rect 6452 8632 6453 8672
rect 6411 8623 6453 8632
rect 6219 8504 6261 8513
rect 6219 8464 6220 8504
rect 6260 8464 6261 8504
rect 6219 8455 6261 8464
rect 6220 8370 6260 8455
rect 5835 8168 5877 8177
rect 5835 8128 5836 8168
rect 5876 8128 5877 8168
rect 5835 8119 5877 8128
rect 6027 8168 6069 8177
rect 6027 8128 6028 8168
rect 6068 8128 6069 8168
rect 6027 8119 6069 8128
rect 5739 7664 5781 7673
rect 5739 7624 5740 7664
rect 5780 7624 5781 7664
rect 5739 7615 5781 7624
rect 5547 7496 5589 7505
rect 5547 7456 5548 7496
rect 5588 7456 5589 7496
rect 5547 7447 5589 7456
rect 5356 6439 5396 6448
rect 5451 6488 5493 6497
rect 5451 6448 5452 6488
rect 5492 6448 5493 6488
rect 5451 6439 5493 6448
rect 5548 6488 5588 7447
rect 5548 6439 5588 6448
rect 5740 6488 5780 7615
rect 5836 7169 5876 8119
rect 6028 8000 6068 8119
rect 6028 7951 6068 7960
rect 6123 8000 6165 8009
rect 6123 7960 6124 8000
rect 6164 7960 6165 8000
rect 6123 7951 6165 7960
rect 6315 8000 6357 8009
rect 6315 7960 6316 8000
rect 6356 7960 6357 8000
rect 6315 7951 6357 7960
rect 6124 7832 6164 7951
rect 6028 7792 6164 7832
rect 6028 7673 6068 7792
rect 6220 7748 6260 7757
rect 6124 7708 6220 7748
rect 6027 7664 6069 7673
rect 6027 7624 6028 7664
rect 6068 7624 6069 7664
rect 6027 7615 6069 7624
rect 6028 7412 6068 7615
rect 6124 7589 6164 7708
rect 6220 7699 6260 7708
rect 6123 7580 6165 7589
rect 6123 7540 6124 7580
rect 6164 7540 6165 7580
rect 6123 7531 6165 7540
rect 6028 7363 6068 7372
rect 5835 7160 5877 7169
rect 5835 7120 5836 7160
rect 5876 7120 5877 7160
rect 5835 7111 5877 7120
rect 5836 7026 5876 7111
rect 5932 6665 5972 6750
rect 5931 6656 5973 6665
rect 5931 6616 5932 6656
rect 5972 6616 5973 6656
rect 5931 6607 5973 6616
rect 5740 6439 5780 6448
rect 5836 6488 5876 6497
rect 6028 6488 6068 6497
rect 5876 6448 5972 6488
rect 5836 6439 5876 6448
rect 5163 6404 5205 6413
rect 5163 6364 5164 6404
rect 5204 6364 5205 6404
rect 5163 6355 5205 6364
rect 4203 6320 4245 6329
rect 4203 6280 4204 6320
rect 4244 6280 4245 6320
rect 4203 6271 4245 6280
rect 4491 6320 4533 6329
rect 4491 6280 4492 6320
rect 4532 6280 4533 6320
rect 4491 6271 4533 6280
rect 5067 6320 5109 6329
rect 5067 6280 5068 6320
rect 5108 6280 5109 6320
rect 5067 6271 5109 6280
rect 3916 6196 4148 6236
rect 3532 5900 3572 6196
rect 3723 6187 3765 6196
rect 3688 6068 4056 6077
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 3688 6019 4056 6028
rect 4108 5900 4148 6196
rect 3532 5860 3764 5900
rect 3147 5816 3189 5825
rect 3147 5776 3148 5816
rect 3188 5776 3189 5816
rect 3147 5767 3189 5776
rect 3435 5816 3477 5825
rect 3435 5776 3436 5816
rect 3476 5776 3477 5816
rect 3435 5767 3477 5776
rect 3052 4927 3092 4936
rect 2955 4892 2997 4901
rect 2955 4852 2956 4892
rect 2996 4852 2997 4892
rect 2955 4843 2997 4852
rect 3148 4808 3188 5767
rect 3340 5657 3380 5742
rect 3339 5648 3381 5657
rect 3244 5627 3284 5636
rect 3339 5608 3340 5648
rect 3380 5608 3381 5648
rect 3339 5599 3381 5608
rect 3436 5648 3476 5657
rect 3244 4985 3284 5587
rect 3436 5153 3476 5608
rect 3724 5648 3764 5860
rect 3724 5599 3764 5608
rect 3820 5860 4148 5900
rect 3820 5648 3860 5860
rect 4204 5816 4244 6271
rect 4299 6236 4341 6245
rect 4299 6196 4300 6236
rect 4340 6196 4341 6236
rect 4299 6187 4341 6196
rect 3820 5599 3860 5608
rect 3916 5776 4244 5816
rect 3916 5648 3956 5776
rect 3916 5599 3956 5608
rect 4012 5648 4052 5657
rect 4204 5648 4244 5657
rect 4052 5608 4204 5648
rect 4012 5599 4052 5608
rect 4204 5599 4244 5608
rect 4300 5648 4340 6187
rect 4300 5599 4340 5608
rect 3532 5480 3572 5489
rect 3532 5321 3572 5440
rect 3627 5480 3669 5489
rect 3627 5440 3628 5480
rect 3668 5440 3669 5480
rect 3627 5431 3669 5440
rect 4107 5480 4149 5489
rect 4107 5440 4108 5480
rect 4148 5440 4149 5480
rect 4107 5431 4149 5440
rect 4492 5480 4532 6271
rect 4971 6236 5013 6245
rect 4971 6196 4972 6236
rect 5012 6196 5013 6236
rect 4971 6187 5013 6196
rect 4972 5741 5012 6187
rect 4971 5732 5013 5741
rect 4971 5692 4972 5732
rect 5012 5692 5013 5732
rect 4971 5683 5013 5692
rect 4684 5648 4724 5657
rect 4492 5431 4532 5440
rect 4588 5608 4684 5648
rect 3531 5312 3573 5321
rect 3531 5272 3532 5312
rect 3572 5272 3573 5312
rect 3531 5263 3573 5272
rect 3435 5144 3477 5153
rect 3435 5104 3436 5144
rect 3476 5104 3477 5144
rect 3435 5095 3477 5104
rect 3243 4976 3285 4985
rect 3628 4976 3668 5431
rect 3723 5312 3765 5321
rect 3723 5272 3724 5312
rect 3764 5272 3765 5312
rect 3723 5263 3765 5272
rect 3724 5069 3764 5263
rect 3723 5060 3765 5069
rect 3723 5020 3724 5060
rect 3764 5020 3765 5060
rect 3723 5011 3765 5020
rect 3243 4936 3244 4976
rect 3284 4936 3285 4976
rect 3243 4927 3285 4936
rect 3532 4936 3668 4976
rect 4012 4976 4052 4985
rect 3436 4892 3476 4901
rect 3148 4768 3284 4808
rect 2764 4180 2900 4220
rect 2572 4136 2612 4145
rect 2476 4096 2572 4136
rect 2572 3464 2612 4096
rect 2764 3893 2804 4180
rect 2956 4136 2996 4145
rect 2860 4096 2956 4136
rect 2763 3884 2805 3893
rect 2763 3844 2764 3884
rect 2804 3844 2805 3884
rect 2763 3835 2805 3844
rect 2763 3632 2805 3641
rect 2763 3592 2764 3632
rect 2804 3592 2805 3632
rect 2763 3583 2805 3592
rect 2764 3498 2804 3583
rect 1803 3128 1845 3137
rect 1803 3088 1804 3128
rect 1844 3088 1845 3128
rect 1803 3079 1845 3088
rect 2283 3128 2325 3137
rect 2283 3088 2284 3128
rect 2324 3088 2325 3128
rect 2283 3079 2325 3088
rect 1707 2120 1749 2129
rect 1707 2080 1708 2120
rect 1748 2080 1749 2120
rect 1707 2071 1749 2080
rect 1611 1364 1653 1373
rect 1611 1324 1612 1364
rect 1652 1324 1653 1364
rect 1611 1315 1653 1324
rect 1516 1112 1556 1121
rect 1420 1072 1516 1112
rect 1516 1063 1556 1072
rect 1612 1112 1652 1121
rect 1419 944 1461 953
rect 1419 904 1420 944
rect 1460 904 1461 944
rect 1612 944 1652 1072
rect 1708 1112 1748 2071
rect 1804 2045 1844 3079
rect 1995 2876 2037 2885
rect 1995 2836 1996 2876
rect 2036 2836 2037 2876
rect 1995 2827 2037 2836
rect 1803 2036 1845 2045
rect 1803 1996 1804 2036
rect 1844 1996 1845 2036
rect 1803 1987 1845 1996
rect 1899 1952 1941 1961
rect 1899 1912 1900 1952
rect 1940 1912 1941 1952
rect 1899 1903 1941 1912
rect 1900 1457 1940 1903
rect 1899 1448 1941 1457
rect 1899 1408 1900 1448
rect 1940 1408 1941 1448
rect 1899 1399 1941 1408
rect 1708 1063 1748 1072
rect 1900 1112 1940 1399
rect 1900 1063 1940 1072
rect 1996 944 2036 2827
rect 2572 2633 2612 3424
rect 2667 3464 2709 3473
rect 2667 3424 2668 3464
rect 2708 3424 2709 3464
rect 2667 3415 2709 3424
rect 2571 2624 2613 2633
rect 2571 2584 2572 2624
rect 2612 2584 2613 2624
rect 2571 2575 2613 2584
rect 2668 1793 2708 3415
rect 2763 3212 2805 3221
rect 2763 3172 2764 3212
rect 2804 3172 2805 3212
rect 2763 3163 2805 3172
rect 2764 3078 2804 3163
rect 2860 3128 2900 4096
rect 2956 4087 2996 4096
rect 3052 4136 3092 4145
rect 2955 3464 2997 3473
rect 2955 3424 2956 3464
rect 2996 3424 2997 3464
rect 2955 3415 2997 3424
rect 2956 3330 2996 3415
rect 2955 3128 2997 3137
rect 2860 3088 2956 3128
rect 2996 3088 2997 3128
rect 2955 3079 2997 3088
rect 2859 2960 2901 2969
rect 2859 2920 2860 2960
rect 2900 2920 2901 2960
rect 2859 2911 2901 2920
rect 2763 2624 2805 2633
rect 2763 2584 2764 2624
rect 2804 2584 2805 2624
rect 2763 2575 2805 2584
rect 2764 1952 2804 2575
rect 2667 1784 2709 1793
rect 2667 1744 2668 1784
rect 2708 1744 2709 1784
rect 2667 1735 2709 1744
rect 2764 1205 2804 1912
rect 2860 1280 2900 2911
rect 2956 2876 2996 3079
rect 2956 2827 2996 2836
rect 3052 2540 3092 4096
rect 3147 4136 3189 4145
rect 3147 4096 3148 4136
rect 3188 4096 3189 4136
rect 3244 4136 3284 4768
rect 3436 4733 3476 4852
rect 3532 4892 3572 4936
rect 3435 4724 3477 4733
rect 3435 4684 3436 4724
rect 3476 4684 3477 4724
rect 3435 4675 3477 4684
rect 3532 4388 3572 4852
rect 4012 4733 4052 4936
rect 4011 4724 4053 4733
rect 4011 4684 4012 4724
rect 4052 4684 4053 4724
rect 4011 4675 4053 4684
rect 3688 4556 4056 4565
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 3688 4507 4056 4516
rect 3532 4348 3668 4388
rect 3436 4136 3476 4145
rect 3244 4096 3436 4136
rect 3147 4087 3189 4096
rect 3436 4087 3476 4096
rect 3148 4002 3188 4087
rect 3244 3968 3284 3977
rect 3147 3884 3189 3893
rect 3147 3844 3148 3884
rect 3188 3844 3189 3884
rect 3147 3835 3189 3844
rect 3148 2969 3188 3835
rect 3147 2960 3189 2969
rect 3147 2920 3148 2960
rect 3188 2920 3189 2960
rect 3147 2911 3189 2920
rect 3244 2549 3284 3928
rect 3531 3968 3573 3977
rect 3531 3928 3532 3968
rect 3572 3928 3573 3968
rect 3531 3919 3573 3928
rect 3340 2629 3380 2638
rect 3148 2540 3188 2549
rect 3052 2500 3148 2540
rect 3148 2491 3188 2500
rect 3243 2540 3285 2549
rect 3243 2500 3244 2540
rect 3284 2500 3285 2540
rect 3243 2491 3285 2500
rect 3340 2213 3380 2589
rect 3435 2624 3477 2633
rect 3435 2584 3436 2624
rect 3476 2584 3477 2624
rect 3435 2575 3477 2584
rect 2955 2204 2997 2213
rect 2955 2164 2956 2204
rect 2996 2164 2997 2204
rect 2955 2155 2997 2164
rect 3339 2204 3381 2213
rect 3339 2164 3340 2204
rect 3380 2164 3381 2204
rect 3339 2155 3381 2164
rect 2956 2120 2996 2155
rect 2956 2069 2996 2080
rect 3243 2120 3285 2129
rect 3243 2080 3244 2120
rect 3284 2080 3285 2120
rect 3243 2071 3285 2080
rect 3244 2036 3284 2071
rect 3244 1985 3284 1996
rect 3147 1952 3189 1961
rect 3147 1912 3148 1952
rect 3188 1912 3189 1952
rect 3147 1903 3189 1912
rect 3340 1952 3380 1961
rect 3436 1952 3476 2575
rect 3532 2540 3572 3919
rect 3628 3473 3668 4348
rect 3627 3464 3669 3473
rect 3627 3424 3628 3464
rect 3668 3424 3669 3464
rect 3627 3415 3669 3424
rect 3688 3044 4056 3053
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 3688 2995 4056 3004
rect 3915 2876 3957 2885
rect 3915 2836 3916 2876
rect 3956 2836 3957 2876
rect 3915 2827 3957 2836
rect 3819 2792 3861 2801
rect 3819 2752 3820 2792
rect 3860 2752 3861 2792
rect 3819 2743 3861 2752
rect 3820 2624 3860 2743
rect 3820 2575 3860 2584
rect 3532 2500 3668 2540
rect 3628 2297 3668 2500
rect 3627 2288 3669 2297
rect 3627 2248 3628 2288
rect 3668 2248 3669 2288
rect 3627 2239 3669 2248
rect 3531 2204 3573 2213
rect 3531 2164 3532 2204
rect 3572 2164 3573 2204
rect 3531 2155 3573 2164
rect 3532 2120 3572 2155
rect 3532 2069 3572 2080
rect 3380 1912 3476 1952
rect 3628 1952 3668 1961
rect 3148 1818 3188 1903
rect 3340 1364 3380 1912
rect 3628 1709 3668 1912
rect 3724 1952 3764 1961
rect 3724 1793 3764 1912
rect 3820 1952 3860 1961
rect 3916 1952 3956 2827
rect 3860 1912 3956 1952
rect 3820 1903 3860 1912
rect 3723 1784 3765 1793
rect 3723 1744 3724 1784
rect 3764 1744 3765 1784
rect 3723 1735 3765 1744
rect 4012 1709 4052 1794
rect 3627 1700 3669 1709
rect 3627 1660 3628 1700
rect 3668 1660 3669 1700
rect 3627 1651 3669 1660
rect 4011 1700 4053 1709
rect 4011 1660 4012 1700
rect 4052 1660 4053 1700
rect 4011 1651 4053 1660
rect 3688 1532 4056 1541
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 3688 1483 4056 1492
rect 4108 1448 4148 5431
rect 4299 5144 4341 5153
rect 4299 5104 4300 5144
rect 4340 5104 4341 5144
rect 4299 5095 4341 5104
rect 4300 4472 4340 5095
rect 4491 4976 4533 4985
rect 4491 4931 4492 4976
rect 4532 4931 4533 4976
rect 4491 4927 4533 4931
rect 4492 4841 4532 4927
rect 4588 4556 4628 5608
rect 4684 5599 4724 5608
rect 4780 5648 4820 5657
rect 4684 5144 4724 5153
rect 4780 5144 4820 5608
rect 4875 5648 4917 5657
rect 4875 5608 4876 5648
rect 4916 5608 4917 5648
rect 4875 5599 4917 5608
rect 5164 5648 5204 6355
rect 5451 6320 5493 6329
rect 5451 6280 5452 6320
rect 5492 6280 5493 6320
rect 5451 6271 5493 6280
rect 5452 6186 5492 6271
rect 5164 5599 5204 5608
rect 5355 5648 5397 5657
rect 5355 5608 5356 5648
rect 5396 5608 5397 5648
rect 5355 5599 5397 5608
rect 4876 5514 4916 5599
rect 4972 5489 5012 5574
rect 4971 5480 5013 5489
rect 4971 5440 4972 5480
rect 5012 5440 5013 5480
rect 4971 5431 5013 5440
rect 4928 5312 5296 5321
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 4928 5263 5296 5272
rect 4724 5104 4820 5144
rect 4684 5095 4724 5104
rect 5067 5060 5109 5069
rect 5259 5060 5301 5069
rect 5067 5020 5068 5060
rect 5108 5020 5109 5060
rect 5067 5011 5109 5020
rect 5164 5020 5260 5060
rect 5300 5020 5301 5060
rect 4588 4516 4916 4556
rect 4300 4432 4628 4472
rect 4203 4388 4245 4397
rect 4203 4348 4204 4388
rect 4244 4348 4245 4388
rect 4203 4339 4245 4348
rect 4204 3464 4244 4339
rect 4588 4313 4628 4432
rect 4683 4388 4725 4397
rect 4683 4348 4684 4388
rect 4724 4348 4725 4388
rect 4683 4339 4725 4348
rect 4876 4388 4916 4516
rect 5068 4472 5108 5011
rect 5164 4976 5204 5020
rect 5259 5011 5301 5020
rect 5164 4927 5204 4936
rect 5068 4432 5204 4472
rect 4916 4348 5108 4388
rect 4876 4339 4916 4348
rect 4587 4304 4629 4313
rect 4587 4264 4588 4304
rect 4628 4264 4629 4304
rect 4587 4255 4629 4264
rect 4395 3548 4437 3557
rect 4395 3508 4396 3548
rect 4436 3508 4437 3548
rect 4395 3499 4437 3508
rect 4204 3415 4244 3424
rect 4396 3414 4436 3499
rect 4491 3464 4533 3473
rect 4491 3424 4492 3464
rect 4532 3424 4533 3464
rect 4491 3415 4533 3424
rect 4588 3464 4628 4255
rect 4684 4136 4724 4339
rect 4684 4087 4724 4096
rect 5068 4136 5108 4348
rect 5164 4136 5204 4432
rect 5260 4388 5300 4397
rect 5356 4388 5396 5599
rect 5300 4348 5396 4388
rect 5260 4339 5300 4348
rect 5260 4136 5300 4145
rect 5164 4096 5260 4136
rect 5068 4087 5108 4096
rect 5260 4087 5300 4096
rect 5356 4136 5396 4145
rect 5548 4136 5588 4145
rect 4779 3968 4821 3977
rect 4779 3928 4780 3968
rect 4820 3928 4821 3968
rect 4779 3919 4821 3928
rect 4683 3884 4725 3893
rect 4683 3844 4684 3884
rect 4724 3844 4725 3884
rect 4683 3835 4725 3844
rect 4684 3548 4724 3835
rect 4684 3499 4724 3508
rect 4299 3380 4341 3389
rect 4299 3340 4300 3380
rect 4340 3340 4341 3380
rect 4299 3331 4341 3340
rect 4300 2885 4340 3331
rect 4299 2876 4341 2885
rect 4299 2836 4300 2876
rect 4340 2836 4341 2876
rect 4299 2827 4341 2836
rect 4299 2708 4341 2717
rect 4299 2668 4300 2708
rect 4340 2668 4341 2708
rect 4299 2659 4341 2668
rect 4396 2708 4436 2717
rect 4492 2708 4532 3415
rect 4436 2668 4532 2708
rect 4396 2659 4436 2668
rect 4300 2574 4340 2659
rect 4588 1961 4628 3424
rect 4780 3464 4820 3919
rect 5356 3893 5396 4096
rect 5452 4096 5548 4136
rect 5355 3884 5397 3893
rect 5355 3844 5356 3884
rect 5396 3844 5397 3884
rect 5355 3835 5397 3844
rect 4928 3800 5296 3809
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 4928 3751 5296 3760
rect 5260 3632 5300 3641
rect 5452 3632 5492 4096
rect 5548 4087 5588 4096
rect 5644 4136 5684 4145
rect 5300 3592 5492 3632
rect 5260 3583 5300 3592
rect 5548 3473 5588 3558
rect 4780 3415 4820 3424
rect 4972 3464 5012 3473
rect 4972 3305 5012 3424
rect 5068 3464 5108 3473
rect 4971 3296 5013 3305
rect 4971 3256 4972 3296
rect 5012 3256 5013 3296
rect 4971 3247 5013 3256
rect 4875 3212 4917 3221
rect 4875 3172 4876 3212
rect 4916 3172 4917 3212
rect 4875 3163 4917 3172
rect 4780 2624 4820 2635
rect 4780 2549 4820 2584
rect 4876 2624 4916 3163
rect 4972 2633 5012 3247
rect 5068 2969 5108 3424
rect 5547 3464 5589 3473
rect 5547 3424 5548 3464
rect 5588 3424 5589 3464
rect 5547 3415 5589 3424
rect 5451 3296 5493 3305
rect 5548 3296 5588 3305
rect 5451 3256 5452 3296
rect 5492 3256 5548 3296
rect 5451 3247 5493 3256
rect 5548 3247 5588 3256
rect 5644 3128 5684 4096
rect 5836 4136 5876 4145
rect 5932 4136 5972 6448
rect 6028 6320 6068 6448
rect 6124 6320 6164 7531
rect 6316 7160 6356 7951
rect 6219 6824 6261 6833
rect 6219 6784 6220 6824
rect 6260 6784 6261 6824
rect 6219 6775 6261 6784
rect 6220 6497 6260 6775
rect 6316 6740 6356 7120
rect 6412 6917 6452 8623
rect 6508 8513 6548 9472
rect 6604 9463 6644 9472
rect 6699 9512 6741 9521
rect 6699 9472 6700 9512
rect 6740 9472 6741 9512
rect 6699 9463 6741 9472
rect 6892 9512 6932 9640
rect 7180 9640 7508 9680
rect 6892 9463 6932 9472
rect 6988 9512 7028 9521
rect 7089 9512 7129 9521
rect 6700 9378 6740 9463
rect 6603 9260 6645 9269
rect 6603 9220 6604 9260
rect 6644 9220 6645 9260
rect 6603 9211 6645 9220
rect 6604 9126 6644 9211
rect 6795 8840 6837 8849
rect 6795 8800 6796 8840
rect 6836 8800 6837 8840
rect 6795 8791 6837 8800
rect 6796 8672 6836 8791
rect 6700 8632 6796 8672
rect 6507 8504 6549 8513
rect 6507 8464 6508 8504
rect 6548 8464 6549 8504
rect 6507 8455 6549 8464
rect 6700 8009 6740 8632
rect 6796 8623 6836 8632
rect 6891 8672 6933 8681
rect 6891 8632 6892 8672
rect 6932 8632 6933 8672
rect 6891 8623 6933 8632
rect 6892 8538 6932 8623
rect 6891 8168 6933 8177
rect 6891 8128 6892 8168
rect 6932 8128 6933 8168
rect 6891 8119 6933 8128
rect 6699 8000 6741 8009
rect 6699 7960 6700 8000
rect 6740 7960 6741 8000
rect 6699 7951 6741 7960
rect 6796 8000 6836 8009
rect 6700 7866 6740 7951
rect 6699 7496 6741 7505
rect 6699 7456 6700 7496
rect 6740 7456 6741 7496
rect 6699 7447 6741 7456
rect 6604 7160 6644 7171
rect 6604 7085 6644 7120
rect 6700 7160 6740 7447
rect 6700 7111 6740 7120
rect 6603 7076 6645 7085
rect 6603 7036 6604 7076
rect 6644 7036 6645 7076
rect 6603 7027 6645 7036
rect 6796 6917 6836 7960
rect 6411 6908 6453 6917
rect 6411 6868 6412 6908
rect 6452 6868 6453 6908
rect 6411 6859 6453 6868
rect 6795 6908 6837 6917
rect 6795 6868 6796 6908
rect 6836 6868 6837 6908
rect 6795 6859 6837 6868
rect 6316 6700 6740 6740
rect 6219 6488 6261 6497
rect 6219 6448 6220 6488
rect 6260 6448 6261 6488
rect 6219 6439 6261 6448
rect 6316 6488 6356 6700
rect 6507 6572 6549 6581
rect 6507 6532 6508 6572
rect 6548 6532 6549 6572
rect 6507 6523 6549 6532
rect 6316 6439 6356 6448
rect 6412 6488 6452 6497
rect 6412 6320 6452 6448
rect 6508 6438 6548 6523
rect 6700 6488 6740 6700
rect 6892 6656 6932 8119
rect 6988 7589 7028 9472
rect 7084 9472 7089 9512
rect 7084 9463 7129 9472
rect 6987 7580 7029 7589
rect 6987 7540 6988 7580
rect 7028 7540 7029 7580
rect 6987 7531 7029 7540
rect 6988 7412 7028 7421
rect 7084 7412 7124 9463
rect 7180 8597 7220 9640
rect 7372 9512 7412 9521
rect 7276 9472 7372 9512
rect 7276 8849 7316 9472
rect 7372 9463 7412 9472
rect 7468 9512 7508 9640
rect 7468 9463 7508 9472
rect 7275 8840 7317 8849
rect 7275 8800 7276 8840
rect 7316 8800 7317 8840
rect 7275 8791 7317 8800
rect 7467 8840 7509 8849
rect 7467 8800 7468 8840
rect 7508 8800 7509 8840
rect 7467 8791 7509 8800
rect 7276 8672 7316 8681
rect 7179 8588 7221 8597
rect 7179 8548 7180 8588
rect 7220 8548 7221 8588
rect 7179 8539 7221 8548
rect 7276 8177 7316 8632
rect 7372 8672 7412 8681
rect 7275 8168 7317 8177
rect 7275 8128 7276 8168
rect 7316 8128 7317 8168
rect 7275 8119 7317 8128
rect 7028 7372 7124 7412
rect 7180 7916 7220 7925
rect 6988 7363 7028 7372
rect 7083 6908 7125 6917
rect 7083 6868 7084 6908
rect 7124 6868 7125 6908
rect 7083 6859 7125 6868
rect 6700 6439 6740 6448
rect 6796 6616 6932 6656
rect 6796 6320 6836 6616
rect 6891 6488 6933 6497
rect 6891 6448 6892 6488
rect 6932 6448 6933 6488
rect 6891 6439 6933 6448
rect 6988 6488 7028 6497
rect 6892 6354 6932 6439
rect 6028 6280 6452 6320
rect 6508 6280 6836 6320
rect 6315 6152 6357 6161
rect 6315 6112 6316 6152
rect 6356 6112 6357 6152
rect 6315 6103 6357 6112
rect 6219 4724 6261 4733
rect 6219 4684 6220 4724
rect 6260 4684 6261 4724
rect 6219 4675 6261 4684
rect 6220 4136 6260 4675
rect 6316 4304 6356 6103
rect 6412 5648 6452 5657
rect 6412 5321 6452 5608
rect 6411 5312 6453 5321
rect 6411 5272 6412 5312
rect 6452 5272 6453 5312
rect 6411 5263 6453 5272
rect 6412 4976 6452 5263
rect 6412 4481 6452 4936
rect 6411 4472 6453 4481
rect 6411 4432 6412 4472
rect 6452 4432 6453 4472
rect 6411 4423 6453 4432
rect 6508 4388 6548 6280
rect 6988 6236 7028 6448
rect 6700 6196 7028 6236
rect 6604 5480 6644 5489
rect 6604 5069 6644 5440
rect 6603 5060 6645 5069
rect 6603 5020 6604 5060
rect 6644 5020 6645 5060
rect 6603 5011 6645 5020
rect 6603 4724 6645 4733
rect 6603 4684 6604 4724
rect 6644 4684 6645 4724
rect 6603 4675 6645 4684
rect 6604 4590 6644 4675
rect 6700 4649 6740 6196
rect 6891 6068 6933 6077
rect 6891 6028 6892 6068
rect 6932 6028 6933 6068
rect 6891 6019 6933 6028
rect 6796 5648 6836 5657
rect 6796 5573 6836 5608
rect 6795 5564 6837 5573
rect 6795 5524 6796 5564
rect 6836 5524 6837 5564
rect 6795 5515 6837 5524
rect 6796 5153 6836 5515
rect 6892 5237 6932 6019
rect 6891 5228 6933 5237
rect 6891 5188 6892 5228
rect 6932 5188 6933 5228
rect 6891 5179 6933 5188
rect 6795 5144 6837 5153
rect 6795 5104 6796 5144
rect 6836 5104 6837 5144
rect 6795 5095 6837 5104
rect 6795 4976 6837 4985
rect 6795 4936 6796 4976
rect 6836 4936 6837 4976
rect 6795 4927 6837 4936
rect 6987 4976 7029 4985
rect 6987 4936 6988 4976
rect 7028 4936 7029 4976
rect 6987 4927 7029 4936
rect 6796 4842 6836 4927
rect 6988 4842 7028 4927
rect 7084 4808 7124 6859
rect 7180 6656 7220 7876
rect 7275 7916 7317 7925
rect 7275 7876 7276 7916
rect 7316 7876 7317 7916
rect 7275 7867 7317 7876
rect 7276 7757 7316 7867
rect 7275 7748 7317 7757
rect 7275 7708 7276 7748
rect 7316 7708 7317 7748
rect 7275 7699 7317 7708
rect 7372 7673 7412 8632
rect 7371 7664 7413 7673
rect 7371 7624 7372 7664
rect 7412 7624 7413 7664
rect 7371 7615 7413 7624
rect 7275 7580 7317 7589
rect 7275 7540 7276 7580
rect 7316 7540 7317 7580
rect 7275 7531 7317 7540
rect 7276 7160 7316 7531
rect 7372 7412 7412 7421
rect 7468 7412 7508 8791
rect 7563 7748 7605 7757
rect 7563 7708 7564 7748
rect 7604 7708 7605 7748
rect 7563 7699 7605 7708
rect 7412 7372 7508 7412
rect 7372 7363 7412 7372
rect 7372 7160 7412 7169
rect 7276 7120 7372 7160
rect 7372 7111 7412 7120
rect 7564 7160 7604 7699
rect 7564 7111 7604 7120
rect 7660 7160 7700 9640
rect 7948 9640 8756 9680
rect 7852 8672 7892 8681
rect 7756 8000 7796 8011
rect 7756 7925 7796 7960
rect 7755 7916 7797 7925
rect 7755 7876 7756 7916
rect 7796 7876 7797 7916
rect 7755 7867 7797 7876
rect 7852 7580 7892 8632
rect 7660 7111 7700 7120
rect 7756 7540 7892 7580
rect 7563 6656 7605 6665
rect 7180 6616 7508 6656
rect 7276 6488 7316 6497
rect 7180 6448 7276 6488
rect 7180 4985 7220 6448
rect 7276 6439 7316 6448
rect 7276 5069 7316 5100
rect 7275 5060 7317 5069
rect 7275 5020 7276 5060
rect 7316 5020 7317 5060
rect 7275 5011 7317 5020
rect 7179 4976 7221 4985
rect 7179 4936 7180 4976
rect 7220 4936 7221 4976
rect 7179 4927 7221 4936
rect 7276 4976 7316 5011
rect 7276 4901 7316 4936
rect 7372 4976 7412 4985
rect 7275 4892 7317 4901
rect 7275 4852 7276 4892
rect 7316 4852 7317 4892
rect 7275 4843 7317 4852
rect 7084 4768 7220 4808
rect 6796 4724 6836 4733
rect 7180 4724 7220 4768
rect 7180 4684 7316 4724
rect 6699 4640 6741 4649
rect 6699 4600 6700 4640
rect 6740 4600 6741 4640
rect 6699 4591 6741 4600
rect 6508 4348 6644 4388
rect 6316 4264 6548 4304
rect 5932 4096 6164 4136
rect 5836 4052 5876 4096
rect 5836 4012 6068 4052
rect 5740 3968 5780 3977
rect 5740 3389 5780 3928
rect 6028 3557 6068 4012
rect 6027 3548 6069 3557
rect 6027 3508 6028 3548
rect 6068 3508 6069 3548
rect 6027 3499 6069 3508
rect 5932 3464 5972 3473
rect 5739 3380 5781 3389
rect 5739 3340 5740 3380
rect 5780 3340 5781 3380
rect 5932 3380 5972 3424
rect 6028 3380 6068 3499
rect 5932 3340 6068 3380
rect 5739 3331 5781 3340
rect 5739 3212 5781 3221
rect 5932 3212 5972 3221
rect 5739 3172 5740 3212
rect 5780 3172 5781 3212
rect 5739 3163 5781 3172
rect 5836 3172 5932 3212
rect 5452 3088 5684 3128
rect 5067 2960 5109 2969
rect 5067 2920 5068 2960
rect 5108 2920 5109 2960
rect 5067 2911 5109 2920
rect 5356 2633 5396 2718
rect 4876 2575 4916 2584
rect 4971 2624 5013 2633
rect 4971 2584 4972 2624
rect 5012 2584 5013 2624
rect 4971 2575 5013 2584
rect 5355 2624 5397 2633
rect 5355 2584 5356 2624
rect 5396 2584 5397 2624
rect 5355 2575 5397 2584
rect 4779 2540 4821 2549
rect 4779 2500 4780 2540
rect 4820 2500 4821 2540
rect 4779 2491 4821 2500
rect 5355 2456 5397 2465
rect 5355 2416 5356 2456
rect 5396 2416 5397 2456
rect 5355 2407 5397 2416
rect 4779 2288 4821 2297
rect 4779 2248 4780 2288
rect 4820 2248 4821 2288
rect 4779 2239 4821 2248
rect 4928 2288 5296 2297
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 4928 2239 5296 2248
rect 4780 2045 4820 2239
rect 4779 2036 4821 2045
rect 4779 1996 4780 2036
rect 4820 1996 4821 2036
rect 4779 1987 4821 1996
rect 4204 1952 4244 1961
rect 4587 1952 4629 1961
rect 4244 1912 4340 1952
rect 4204 1903 4244 1912
rect 4108 1408 4244 1448
rect 3340 1315 3380 1324
rect 4107 1280 4149 1289
rect 2860 1240 2996 1280
rect 2763 1196 2805 1205
rect 2763 1156 2764 1196
rect 2804 1156 2805 1196
rect 2763 1147 2805 1156
rect 1612 904 2036 944
rect 1419 895 1461 904
rect 1420 810 1460 895
rect 2956 80 2996 1240
rect 4107 1240 4108 1280
rect 4148 1240 4149 1280
rect 4107 1231 4149 1240
rect 3147 1196 3189 1205
rect 3147 1156 3148 1196
rect 3188 1156 3189 1196
rect 3147 1147 3189 1156
rect 3148 1112 3188 1147
rect 3148 1061 3188 1072
rect 3819 1112 3861 1121
rect 3819 1072 3820 1112
rect 3860 1072 3861 1112
rect 3819 1063 3861 1072
rect 3820 978 3860 1063
rect 4108 80 4148 1231
rect 4204 869 4244 1408
rect 4300 1121 4340 1912
rect 4587 1912 4588 1952
rect 4628 1912 4629 1952
rect 4587 1903 4629 1912
rect 5260 1280 5300 1291
rect 5260 1205 5300 1240
rect 5259 1196 5301 1205
rect 5259 1156 5260 1196
rect 5300 1156 5301 1196
rect 5259 1147 5301 1156
rect 4299 1112 4341 1121
rect 4299 1072 4300 1112
rect 4340 1072 4341 1112
rect 4299 1063 4341 1072
rect 5067 1112 5109 1121
rect 5067 1072 5068 1112
rect 5108 1072 5109 1112
rect 5067 1063 5109 1072
rect 5068 978 5108 1063
rect 4203 860 4245 869
rect 4203 820 4204 860
rect 4244 820 4245 860
rect 4203 811 4245 820
rect 4928 776 5296 785
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 4928 727 5296 736
rect 5356 608 5396 2407
rect 5452 2129 5492 3088
rect 5740 3078 5780 3163
rect 5547 2960 5589 2969
rect 5547 2920 5548 2960
rect 5588 2920 5589 2960
rect 5547 2911 5589 2920
rect 5548 2540 5588 2911
rect 5643 2792 5685 2801
rect 5643 2752 5644 2792
rect 5684 2752 5685 2792
rect 5643 2743 5685 2752
rect 5644 2666 5684 2743
rect 5644 2617 5684 2626
rect 5740 2624 5780 2633
rect 5740 2540 5780 2584
rect 5548 2500 5780 2540
rect 5547 2372 5589 2381
rect 5547 2332 5548 2372
rect 5588 2332 5589 2372
rect 5547 2323 5589 2332
rect 5451 2120 5493 2129
rect 5451 2080 5452 2120
rect 5492 2080 5493 2120
rect 5451 2071 5493 2080
rect 5452 1952 5492 1961
rect 5548 1952 5588 2323
rect 5740 1952 5780 1961
rect 5492 1912 5588 1952
rect 5644 1912 5740 1952
rect 5452 1457 5492 1912
rect 5451 1448 5493 1457
rect 5451 1408 5452 1448
rect 5492 1408 5493 1448
rect 5451 1399 5493 1408
rect 5644 1205 5684 1912
rect 5740 1903 5780 1912
rect 5836 1952 5876 3172
rect 5932 3163 5972 3172
rect 6028 2969 6068 3340
rect 6124 3464 6164 4096
rect 6220 4087 6260 4096
rect 6508 4136 6548 4264
rect 6027 2960 6069 2969
rect 6027 2920 6028 2960
rect 6068 2920 6069 2960
rect 6027 2911 6069 2920
rect 6124 2876 6164 3424
rect 6220 3464 6260 3473
rect 6412 3464 6452 3473
rect 6260 3424 6412 3464
rect 6220 3305 6260 3424
rect 6412 3415 6452 3424
rect 6219 3296 6261 3305
rect 6219 3256 6220 3296
rect 6260 3256 6261 3296
rect 6219 3247 6261 3256
rect 6508 3221 6548 4096
rect 6604 4136 6644 4348
rect 6604 3473 6644 4096
rect 6603 3464 6645 3473
rect 6603 3424 6604 3464
rect 6644 3424 6645 3464
rect 6603 3415 6645 3424
rect 6700 3464 6740 4591
rect 6796 3977 6836 4684
rect 6891 4556 6933 4565
rect 6891 4516 6892 4556
rect 6932 4516 6933 4556
rect 6891 4507 6933 4516
rect 6892 4388 6932 4507
rect 6892 4339 6932 4348
rect 7180 4136 7220 4147
rect 7180 4061 7220 4096
rect 6987 4052 7029 4061
rect 6987 4012 6988 4052
rect 7028 4012 7029 4052
rect 6987 4003 7029 4012
rect 7179 4052 7221 4061
rect 7179 4012 7180 4052
rect 7220 4012 7221 4052
rect 7179 4003 7221 4012
rect 6795 3968 6837 3977
rect 6795 3928 6796 3968
rect 6836 3928 6837 3968
rect 6795 3919 6837 3928
rect 6700 3415 6740 3424
rect 6988 3464 7028 4003
rect 7083 3884 7125 3893
rect 7083 3844 7084 3884
rect 7124 3844 7125 3884
rect 7083 3835 7125 3844
rect 6988 3415 7028 3424
rect 6603 3296 6645 3305
rect 6603 3256 6604 3296
rect 6644 3256 6645 3296
rect 6603 3247 6645 3256
rect 6507 3212 6549 3221
rect 6507 3172 6508 3212
rect 6548 3172 6549 3212
rect 6507 3163 6549 3172
rect 6220 2876 6260 2885
rect 6124 2836 6220 2876
rect 6220 2827 6260 2836
rect 6028 2792 6068 2801
rect 6068 2752 6164 2792
rect 6028 2743 6068 2752
rect 6124 2708 6164 2752
rect 6315 2708 6357 2717
rect 6124 2668 6260 2708
rect 5931 2624 5973 2633
rect 5931 2584 5932 2624
rect 5972 2584 5973 2624
rect 5931 2575 5973 2584
rect 5932 2120 5972 2575
rect 6220 2456 6260 2668
rect 6315 2668 6316 2708
rect 6356 2668 6357 2708
rect 6315 2659 6357 2668
rect 6316 2624 6356 2659
rect 6316 2573 6356 2584
rect 6604 2624 6644 3247
rect 6700 3212 6740 3221
rect 6987 3212 7029 3221
rect 6740 3172 6836 3212
rect 6700 3163 6740 3172
rect 6220 2416 6356 2456
rect 6123 2372 6165 2381
rect 6123 2332 6124 2372
rect 6164 2332 6165 2372
rect 6123 2323 6165 2332
rect 5932 2071 5972 2080
rect 6027 2120 6069 2129
rect 6027 2080 6028 2120
rect 6068 2080 6069 2120
rect 6027 2071 6069 2080
rect 5836 1903 5876 1912
rect 6028 1952 6068 2071
rect 6124 1961 6164 2323
rect 6316 2288 6356 2416
rect 6281 2248 6356 2288
rect 6028 1903 6068 1912
rect 6123 1952 6165 1961
rect 6123 1912 6124 1952
rect 6164 1912 6165 1952
rect 6123 1903 6165 1912
rect 6281 1945 6321 2248
rect 6124 1818 6164 1903
rect 6281 1896 6321 1905
rect 6411 1952 6453 1961
rect 6411 1912 6412 1952
rect 6452 1912 6453 1952
rect 6411 1903 6453 1912
rect 6219 1784 6261 1793
rect 6219 1744 6220 1784
rect 6260 1744 6261 1784
rect 6219 1735 6261 1744
rect 5739 1700 5781 1709
rect 5739 1660 5740 1700
rect 5780 1660 5781 1700
rect 5739 1651 5781 1660
rect 5643 1196 5685 1205
rect 5643 1156 5644 1196
rect 5684 1156 5685 1196
rect 5643 1147 5685 1156
rect 5451 1112 5493 1121
rect 5451 1072 5452 1112
rect 5492 1072 5493 1112
rect 5451 1063 5493 1072
rect 5740 1112 5780 1651
rect 6027 1616 6069 1625
rect 6027 1576 6028 1616
rect 6068 1576 6069 1616
rect 6027 1567 6069 1576
rect 5740 1063 5780 1072
rect 5835 1112 5877 1121
rect 5835 1072 5836 1112
rect 5876 1072 5877 1112
rect 5835 1063 5877 1072
rect 5452 785 5492 1063
rect 5836 978 5876 1063
rect 6028 944 6068 1567
rect 6123 1532 6165 1541
rect 6123 1492 6124 1532
rect 6164 1492 6165 1532
rect 6123 1483 6165 1492
rect 6028 895 6068 904
rect 5451 776 5493 785
rect 5451 736 5452 776
rect 5492 736 5493 776
rect 5451 727 5493 736
rect 5260 568 5396 608
rect 5260 80 5300 568
rect 6124 449 6164 1483
rect 6220 1112 6260 1735
rect 6315 1700 6357 1709
rect 6315 1660 6316 1700
rect 6356 1660 6357 1700
rect 6315 1651 6357 1660
rect 6220 1063 6260 1072
rect 6316 1112 6356 1651
rect 6316 1063 6356 1072
rect 6412 1112 6452 1903
rect 6604 1709 6644 2584
rect 6700 2624 6740 2633
rect 6700 2381 6740 2584
rect 6699 2372 6741 2381
rect 6699 2332 6700 2372
rect 6740 2332 6741 2372
rect 6699 2323 6741 2332
rect 6796 2120 6836 3172
rect 6987 3172 6988 3212
rect 7028 3172 7029 3212
rect 6987 3163 7029 3172
rect 6988 2708 7028 3163
rect 6700 2080 6836 2120
rect 6892 2668 7028 2708
rect 7084 2708 7124 3835
rect 7179 3632 7221 3641
rect 7179 3592 7180 3632
rect 7220 3592 7221 3632
rect 7179 3583 7221 3592
rect 6603 1700 6645 1709
rect 6603 1660 6604 1700
rect 6644 1660 6645 1700
rect 6603 1651 6645 1660
rect 6412 1063 6452 1072
rect 6700 1112 6740 2080
rect 6796 1952 6836 1961
rect 6796 1709 6836 1912
rect 6892 1952 6932 2668
rect 7084 2659 7124 2668
rect 7180 2708 7220 3583
rect 7180 2659 7220 2668
rect 7276 3464 7316 4684
rect 7372 4565 7412 4936
rect 7371 4556 7413 4565
rect 7371 4516 7372 4556
rect 7412 4516 7413 4556
rect 7371 4507 7413 4516
rect 7468 4304 7508 6616
rect 7563 6616 7564 6656
rect 7604 6616 7605 6656
rect 7563 6607 7605 6616
rect 7564 6488 7604 6607
rect 7564 6439 7604 6448
rect 7660 6488 7700 6497
rect 7660 6161 7700 6448
rect 7659 6152 7701 6161
rect 7659 6112 7660 6152
rect 7700 6112 7701 6152
rect 7659 6103 7701 6112
rect 7756 5069 7796 7540
rect 7852 7412 7892 7421
rect 7948 7412 7988 9640
rect 8140 9512 8180 9521
rect 8140 8849 8180 9472
rect 8236 9512 8276 9521
rect 8139 8840 8181 8849
rect 8139 8800 8140 8840
rect 8180 8800 8181 8840
rect 8139 8791 8181 8800
rect 8139 8672 8181 8681
rect 8139 8632 8140 8672
rect 8180 8632 8181 8672
rect 8139 8623 8181 8632
rect 8140 8000 8180 8623
rect 8236 8084 8276 9472
rect 8332 9512 8372 9640
rect 8332 9463 8372 9472
rect 8428 9512 8468 9521
rect 8716 9512 8756 9640
rect 8908 9640 9004 9680
rect 8468 9472 8660 9512
rect 8428 9463 8468 9472
rect 8427 9260 8469 9269
rect 8427 9220 8428 9260
rect 8468 9220 8469 9260
rect 8427 9211 8469 9220
rect 8332 8681 8372 8767
rect 8331 8677 8373 8681
rect 8331 8632 8332 8677
rect 8372 8632 8373 8677
rect 8331 8623 8373 8632
rect 8331 8504 8373 8513
rect 8331 8464 8332 8504
rect 8372 8464 8373 8504
rect 8331 8455 8373 8464
rect 8332 8336 8372 8455
rect 8428 8420 8468 9211
rect 8620 8756 8660 9472
rect 8716 9463 8756 9472
rect 8811 9512 8853 9521
rect 8811 9472 8812 9512
rect 8852 9472 8853 9512
rect 8811 9463 8853 9472
rect 8812 9378 8852 9463
rect 8811 8756 8853 8765
rect 8620 8716 8756 8756
rect 8523 8672 8565 8681
rect 8523 8632 8524 8672
rect 8564 8632 8565 8672
rect 8523 8623 8565 8632
rect 8524 8588 8564 8623
rect 8524 8537 8564 8548
rect 8428 8380 8660 8420
rect 8332 8296 8564 8336
rect 8427 8168 8469 8177
rect 8427 8128 8428 8168
rect 8468 8128 8469 8168
rect 8427 8119 8469 8128
rect 8236 8044 8372 8084
rect 8140 7986 8276 8000
rect 8140 7960 8236 7986
rect 8236 7589 8276 7946
rect 8235 7580 8277 7589
rect 8235 7540 8236 7580
rect 8276 7540 8277 7580
rect 8235 7531 8277 7540
rect 7892 7372 7988 7412
rect 8139 7412 8181 7421
rect 8139 7372 8140 7412
rect 8180 7372 8181 7412
rect 7852 7363 7892 7372
rect 8139 7363 8181 7372
rect 8043 7160 8085 7169
rect 8043 7120 8044 7160
rect 8084 7120 8085 7160
rect 8043 7111 8085 7120
rect 7851 6656 7893 6665
rect 7851 6616 7852 6656
rect 7892 6616 7893 6656
rect 7851 6607 7893 6616
rect 7563 5060 7605 5069
rect 7563 5020 7564 5060
rect 7604 5020 7605 5060
rect 7563 5011 7605 5020
rect 7755 5060 7797 5069
rect 7755 5020 7756 5060
rect 7796 5020 7797 5060
rect 7852 5060 7892 6607
rect 7948 6236 7988 6245
rect 7948 5237 7988 6196
rect 8044 5648 8084 7111
rect 8140 6665 8180 7363
rect 8139 6656 8181 6665
rect 8139 6616 8140 6656
rect 8180 6616 8181 6656
rect 8332 6656 8372 8044
rect 8428 8034 8468 8119
rect 8428 6656 8468 6665
rect 8332 6616 8428 6656
rect 8139 6607 8181 6616
rect 8428 6607 8468 6616
rect 8235 6572 8277 6581
rect 8235 6532 8236 6572
rect 8276 6532 8277 6572
rect 8235 6523 8277 6532
rect 8139 6488 8181 6497
rect 8139 6448 8140 6488
rect 8180 6448 8181 6488
rect 8139 6439 8181 6448
rect 8236 6488 8276 6523
rect 8140 6354 8180 6439
rect 8236 6437 8276 6448
rect 8332 6488 8372 6497
rect 8524 6488 8564 8296
rect 8620 8000 8660 8380
rect 8620 7951 8660 7960
rect 8716 8000 8756 8716
rect 8811 8716 8812 8756
rect 8852 8716 8853 8756
rect 8811 8707 8853 8716
rect 8812 8672 8852 8707
rect 8812 8621 8852 8632
rect 8908 8504 8948 9640
rect 9004 9631 9044 9640
rect 9388 9680 9428 9689
rect 9484 9680 9524 10672
rect 9428 9640 9524 9680
rect 9676 9680 9716 10672
rect 9772 9680 9812 9689
rect 9676 9640 9772 9680
rect 9868 9680 9908 10672
rect 10060 9848 10100 10672
rect 10252 10025 10292 10672
rect 10251 10016 10293 10025
rect 10251 9976 10252 10016
rect 10292 9976 10293 10016
rect 10251 9967 10293 9976
rect 10060 9808 10292 9848
rect 10156 9680 10196 9689
rect 9868 9640 10156 9680
rect 9388 9631 9428 9640
rect 9772 9631 9812 9640
rect 10156 9631 10196 9640
rect 9099 9596 9141 9605
rect 9099 9556 9100 9596
rect 9140 9556 9141 9596
rect 9099 9547 9141 9556
rect 9100 9101 9140 9547
rect 9483 9512 9525 9521
rect 9483 9472 9484 9512
rect 9524 9472 9525 9512
rect 9483 9463 9525 9472
rect 10155 9512 10197 9521
rect 10155 9472 10156 9512
rect 10196 9472 10197 9512
rect 10155 9463 10197 9472
rect 9099 9092 9141 9101
rect 9099 9052 9100 9092
rect 9140 9052 9141 9092
rect 9099 9043 9141 9052
rect 9387 9092 9429 9101
rect 9387 9052 9388 9092
rect 9428 9052 9429 9092
rect 9387 9043 9429 9052
rect 9099 8672 9141 8681
rect 9099 8632 9100 8672
rect 9140 8632 9141 8672
rect 9099 8623 9141 8632
rect 9100 8538 9140 8623
rect 9196 8588 9236 8597
rect 8716 7951 8756 7960
rect 8812 8464 8948 8504
rect 8812 8000 8852 8464
rect 9196 8177 9236 8548
rect 9195 8168 9237 8177
rect 9195 8128 9196 8168
rect 9236 8128 9237 8168
rect 9195 8119 9237 8128
rect 8812 7951 8852 7960
rect 8908 8000 8948 8009
rect 9099 8000 9141 8009
rect 8948 7960 9044 8000
rect 8908 7951 8948 7960
rect 8811 7664 8853 7673
rect 8811 7624 8812 7664
rect 8852 7624 8853 7664
rect 8811 7615 8853 7624
rect 8812 7085 8852 7615
rect 8811 7076 8853 7085
rect 8811 7036 8812 7076
rect 8852 7036 8853 7076
rect 8811 7027 8853 7036
rect 8372 6448 8564 6488
rect 8811 6488 8853 6497
rect 8811 6448 8812 6488
rect 8852 6448 8853 6488
rect 8332 6439 8372 6448
rect 8811 6439 8853 6448
rect 8812 6354 8852 6439
rect 8427 6320 8469 6329
rect 8427 6280 8428 6320
rect 8468 6280 8469 6320
rect 8427 6271 8469 6280
rect 8044 5321 8084 5608
rect 8235 5564 8277 5573
rect 8235 5524 8236 5564
rect 8276 5524 8277 5564
rect 8235 5515 8277 5524
rect 8236 5430 8276 5515
rect 8043 5312 8085 5321
rect 8043 5272 8044 5312
rect 8084 5272 8085 5312
rect 8043 5263 8085 5272
rect 7947 5228 7989 5237
rect 7947 5188 7948 5228
rect 7988 5188 7989 5228
rect 7947 5179 7989 5188
rect 7852 5020 7988 5060
rect 7755 5011 7797 5020
rect 7372 4264 7508 4304
rect 7372 3893 7412 4264
rect 7468 4136 7508 4147
rect 7468 4061 7508 4096
rect 7564 4136 7604 5011
rect 7467 4052 7509 4061
rect 7467 4012 7468 4052
rect 7508 4012 7509 4052
rect 7467 4003 7509 4012
rect 7371 3884 7413 3893
rect 7371 3844 7372 3884
rect 7412 3844 7413 3884
rect 7371 3835 7413 3844
rect 7372 3548 7412 3835
rect 7372 3499 7412 3508
rect 7083 2540 7125 2549
rect 7083 2500 7084 2540
rect 7124 2500 7125 2540
rect 7083 2491 7125 2500
rect 7084 1952 7124 2491
rect 7276 2381 7316 3424
rect 7371 3380 7413 3389
rect 7371 3340 7372 3380
rect 7412 3340 7413 3380
rect 7371 3331 7413 3340
rect 7372 2549 7412 3331
rect 7371 2540 7413 2549
rect 7371 2500 7372 2540
rect 7412 2500 7413 2540
rect 7371 2491 7413 2500
rect 7275 2372 7317 2381
rect 7275 2332 7276 2372
rect 7316 2332 7317 2372
rect 7275 2323 7317 2332
rect 7276 1952 7316 1961
rect 7084 1912 7276 1952
rect 6892 1903 6932 1912
rect 7276 1903 7316 1912
rect 7372 1952 7412 1961
rect 7468 1952 7508 4003
rect 7564 3977 7604 4096
rect 7756 4892 7796 4901
rect 7563 3968 7605 3977
rect 7563 3928 7564 3968
rect 7604 3928 7605 3968
rect 7563 3919 7605 3928
rect 7563 3464 7605 3473
rect 7563 3424 7564 3464
rect 7604 3424 7605 3464
rect 7563 3415 7605 3424
rect 7564 2372 7604 3415
rect 7660 3212 7700 3221
rect 7756 3212 7796 4852
rect 7852 4892 7892 4901
rect 7852 4388 7892 4852
rect 7852 4339 7892 4348
rect 7948 3641 7988 5020
rect 8044 4733 8084 5263
rect 8331 5228 8373 5237
rect 8331 5188 8332 5228
rect 8372 5188 8373 5228
rect 8331 5179 8373 5188
rect 8332 4976 8372 5179
rect 8332 4927 8372 4936
rect 8428 4808 8468 6271
rect 8524 5648 8564 5657
rect 8524 5573 8564 5608
rect 8620 5648 8660 5657
rect 8660 5608 8948 5648
rect 8620 5599 8660 5608
rect 8523 5564 8565 5573
rect 8523 5524 8524 5564
rect 8564 5524 8565 5564
rect 8523 5515 8565 5524
rect 8524 5069 8564 5515
rect 8811 5480 8853 5489
rect 8811 5440 8812 5480
rect 8852 5440 8853 5480
rect 8811 5431 8853 5440
rect 8812 5346 8852 5431
rect 8523 5060 8565 5069
rect 8523 5020 8524 5060
rect 8564 5020 8565 5060
rect 8523 5011 8565 5020
rect 8811 4976 8853 4985
rect 8811 4931 8812 4976
rect 8852 4931 8853 4976
rect 8811 4927 8853 4931
rect 8812 4841 8852 4927
rect 8428 4768 8660 4808
rect 8043 4724 8085 4733
rect 8043 4684 8044 4724
rect 8084 4684 8085 4724
rect 8043 4675 8085 4684
rect 8427 4472 8469 4481
rect 8427 4432 8428 4472
rect 8468 4432 8469 4472
rect 8427 4423 8469 4432
rect 8139 4220 8181 4229
rect 8139 4180 8140 4220
rect 8180 4180 8181 4220
rect 8139 4171 8181 4180
rect 8140 4136 8180 4171
rect 8140 4085 8180 4096
rect 8331 4136 8373 4145
rect 8331 4096 8332 4136
rect 8372 4096 8373 4136
rect 8331 4087 8373 4096
rect 8428 4136 8468 4423
rect 8523 4304 8565 4313
rect 8523 4264 8524 4304
rect 8564 4264 8565 4304
rect 8523 4255 8565 4264
rect 8428 4087 8468 4096
rect 8524 4136 8564 4255
rect 8524 4087 8564 4096
rect 7947 3632 7989 3641
rect 7947 3592 7948 3632
rect 7988 3592 7989 3632
rect 7947 3583 7989 3592
rect 8332 3632 8372 4087
rect 8427 3800 8469 3809
rect 8427 3760 8428 3800
rect 8468 3760 8469 3800
rect 8427 3751 8469 3760
rect 8332 3583 8372 3592
rect 7700 3172 7796 3212
rect 7852 3464 7892 3473
rect 7660 3163 7700 3172
rect 7659 2792 7701 2801
rect 7659 2752 7660 2792
rect 7700 2752 7701 2792
rect 7659 2743 7701 2752
rect 7660 2624 7700 2743
rect 7852 2633 7892 3424
rect 7948 3464 7988 3473
rect 7660 2575 7700 2584
rect 7851 2624 7893 2633
rect 7851 2584 7852 2624
rect 7892 2584 7893 2624
rect 7851 2575 7893 2584
rect 7851 2456 7893 2465
rect 7851 2416 7852 2456
rect 7892 2416 7893 2456
rect 7851 2407 7893 2416
rect 7564 2332 7700 2372
rect 7563 2204 7605 2213
rect 7563 2164 7564 2204
rect 7604 2164 7605 2204
rect 7563 2155 7605 2164
rect 7412 1912 7508 1952
rect 7372 1903 7412 1912
rect 6987 1868 7029 1877
rect 6987 1828 6988 1868
rect 7028 1828 7029 1868
rect 6987 1819 7029 1828
rect 6795 1700 6837 1709
rect 6795 1660 6796 1700
rect 6836 1660 6837 1700
rect 6795 1651 6837 1660
rect 6891 1196 6933 1205
rect 6891 1156 6892 1196
rect 6932 1156 6933 1196
rect 6891 1147 6933 1156
rect 6700 1063 6740 1072
rect 6796 1112 6836 1121
rect 6508 944 6548 953
rect 6796 944 6836 1072
rect 6892 1112 6932 1147
rect 6892 1061 6932 1072
rect 6988 1112 7028 1819
rect 7564 1616 7604 2155
rect 7660 1709 7700 2332
rect 7852 1952 7892 2407
rect 7948 2297 7988 3424
rect 8043 3464 8085 3473
rect 8043 3424 8044 3464
rect 8084 3424 8085 3464
rect 8043 3415 8085 3424
rect 8140 3464 8180 3473
rect 8044 3330 8084 3415
rect 8140 2960 8180 3424
rect 8332 3464 8372 3473
rect 8332 3137 8372 3424
rect 8331 3128 8373 3137
rect 8331 3088 8332 3128
rect 8372 3088 8373 3128
rect 8331 3079 8373 3088
rect 8044 2920 8180 2960
rect 7947 2288 7989 2297
rect 7947 2248 7948 2288
rect 7988 2248 7989 2288
rect 7947 2239 7989 2248
rect 7852 1903 7892 1912
rect 7755 1784 7797 1793
rect 7755 1744 7756 1784
rect 7796 1744 7797 1784
rect 7755 1735 7797 1744
rect 7659 1700 7701 1709
rect 7659 1660 7660 1700
rect 7700 1660 7701 1700
rect 7659 1651 7701 1660
rect 7468 1576 7604 1616
rect 7180 1280 7220 1289
rect 7180 1121 7220 1240
rect 6988 1063 7028 1072
rect 7179 1112 7221 1121
rect 7179 1072 7180 1112
rect 7220 1072 7221 1112
rect 7179 1063 7221 1072
rect 7468 1112 7508 1576
rect 7468 1063 7508 1072
rect 7564 1112 7604 1121
rect 7756 1112 7796 1735
rect 8044 1289 8084 2920
rect 8140 2629 8180 2638
rect 8140 2465 8180 2589
rect 8428 2540 8468 3751
rect 8524 3464 8564 3473
rect 8524 2960 8564 3424
rect 8620 3464 8660 4768
rect 8811 4388 8853 4397
rect 8811 4348 8812 4388
rect 8852 4348 8853 4388
rect 8908 4388 8948 5608
rect 9004 5573 9044 7960
rect 9099 7960 9100 8000
rect 9140 7960 9141 8000
rect 9099 7951 9141 7960
rect 9292 8000 9332 8009
rect 9100 7866 9140 7951
rect 9195 7748 9237 7757
rect 9195 7708 9196 7748
rect 9236 7708 9237 7748
rect 9195 7699 9237 7708
rect 9196 7614 9236 7699
rect 9292 7328 9332 7960
rect 9196 7288 9332 7328
rect 9100 5648 9140 5657
rect 9003 5564 9045 5573
rect 9003 5524 9004 5564
rect 9044 5524 9045 5564
rect 9003 5515 9045 5524
rect 9003 5060 9045 5069
rect 9003 5020 9004 5060
rect 9044 5020 9045 5060
rect 9003 5011 9045 5020
rect 9004 4926 9044 5011
rect 9100 4976 9140 5608
rect 9196 5228 9236 7288
rect 9292 7160 9332 7169
rect 9388 7160 9428 9043
rect 9484 8924 9524 9463
rect 9579 9428 9621 9437
rect 9579 9388 9580 9428
rect 9620 9388 9621 9428
rect 9579 9379 9621 9388
rect 9964 9428 10004 9437
rect 9580 9294 9620 9379
rect 9675 9344 9717 9353
rect 9675 9304 9676 9344
rect 9716 9304 9717 9344
rect 9675 9295 9717 9304
rect 9579 9008 9621 9017
rect 9676 9008 9716 9295
rect 9579 8968 9580 9008
rect 9620 8968 9716 9008
rect 9579 8959 9621 8968
rect 9484 8875 9524 8884
rect 9484 8000 9524 8009
rect 9580 8000 9620 8959
rect 9867 8840 9909 8849
rect 9867 8800 9868 8840
rect 9908 8800 9909 8840
rect 9867 8791 9909 8800
rect 9524 7960 9620 8000
rect 9676 8756 9716 8765
rect 9484 7951 9524 7960
rect 9676 7925 9716 8716
rect 9868 8706 9908 8791
rect 9964 8345 10004 9388
rect 10060 8756 10100 8765
rect 9963 8336 10005 8345
rect 9963 8296 9964 8336
rect 10004 8296 10005 8336
rect 9963 8287 10005 8296
rect 9675 7916 9717 7925
rect 9675 7876 9676 7916
rect 9716 7876 9717 7916
rect 9675 7867 9717 7876
rect 10060 7580 10100 8716
rect 10156 8000 10196 9463
rect 10252 8849 10292 9808
rect 10348 9428 10388 9437
rect 10348 9269 10388 9388
rect 10347 9260 10389 9269
rect 10347 9220 10348 9260
rect 10388 9220 10389 9260
rect 10347 9211 10389 9220
rect 10444 8924 10484 10672
rect 10539 10016 10581 10025
rect 10539 9976 10540 10016
rect 10580 9976 10581 10016
rect 10539 9967 10581 9976
rect 10348 8884 10484 8924
rect 10251 8840 10293 8849
rect 10251 8800 10252 8840
rect 10292 8800 10293 8840
rect 10251 8791 10293 8800
rect 10252 8504 10292 8513
rect 10348 8504 10388 8884
rect 10292 8464 10388 8504
rect 10444 8756 10484 8765
rect 10252 8455 10292 8464
rect 10444 8177 10484 8716
rect 10540 8513 10580 9967
rect 10636 8840 10676 10672
rect 10731 9008 10773 9017
rect 10731 8968 10732 9008
rect 10772 8968 10773 9008
rect 10731 8959 10773 8968
rect 10636 8791 10676 8800
rect 10539 8504 10581 8513
rect 10539 8464 10540 8504
rect 10580 8464 10581 8504
rect 10539 8455 10581 8464
rect 10443 8168 10485 8177
rect 10443 8128 10444 8168
rect 10484 8128 10485 8168
rect 10732 8168 10772 8959
rect 10828 8840 10868 10672
rect 10923 9428 10965 9437
rect 10923 9388 10924 9428
rect 10964 9388 10965 9428
rect 10923 9379 10965 9388
rect 10828 8791 10868 8800
rect 10924 8588 10964 9379
rect 11020 9008 11060 10672
rect 11212 9680 11252 10672
rect 11404 9857 11444 10672
rect 11403 9848 11445 9857
rect 11403 9808 11404 9848
rect 11444 9808 11445 9848
rect 11403 9799 11445 9808
rect 11212 9640 11540 9680
rect 11211 9344 11253 9353
rect 11211 9304 11212 9344
rect 11252 9304 11253 9344
rect 11211 9295 11253 9304
rect 11212 9101 11252 9295
rect 11211 9092 11253 9101
rect 11211 9052 11212 9092
rect 11252 9052 11253 9092
rect 11211 9043 11253 9052
rect 11020 8968 11156 9008
rect 11020 8765 11060 8850
rect 11116 8840 11156 8968
rect 11212 8840 11252 8849
rect 11116 8800 11212 8840
rect 11212 8791 11252 8800
rect 11019 8756 11061 8765
rect 11019 8716 11020 8756
rect 11060 8716 11061 8756
rect 11019 8707 11061 8716
rect 11404 8756 11444 8765
rect 10924 8548 11156 8588
rect 11116 8168 11156 8548
rect 10732 8128 10868 8168
rect 10443 8119 10485 8128
rect 10635 8084 10677 8093
rect 10635 8044 10636 8084
rect 10676 8044 10677 8084
rect 10635 8035 10677 8044
rect 10156 7960 10484 8000
rect 10060 7540 10388 7580
rect 10251 7412 10293 7421
rect 10251 7372 10252 7412
rect 10292 7372 10293 7412
rect 10251 7363 10293 7372
rect 10252 7244 10292 7363
rect 10252 7195 10292 7204
rect 9332 7120 9428 7160
rect 9483 7160 9525 7169
rect 9483 7120 9484 7160
rect 9524 7120 9525 7160
rect 9292 7111 9332 7120
rect 9483 7111 9525 7120
rect 9676 7160 9716 7169
rect 9484 7026 9524 7111
rect 9676 7001 9716 7120
rect 9772 7160 9812 7169
rect 10060 7160 10100 7169
rect 9812 7120 9908 7160
rect 9772 7111 9812 7120
rect 9580 6992 9620 7001
rect 9387 6824 9429 6833
rect 9387 6784 9388 6824
rect 9428 6784 9429 6824
rect 9387 6775 9429 6784
rect 9388 5648 9428 6775
rect 9580 5741 9620 6952
rect 9675 6992 9717 7001
rect 9675 6952 9676 6992
rect 9716 6952 9717 6992
rect 9675 6943 9717 6952
rect 9579 5732 9621 5741
rect 9579 5692 9580 5732
rect 9620 5692 9621 5732
rect 9579 5683 9621 5692
rect 9388 5599 9428 5608
rect 9484 5564 9524 5573
rect 9196 5188 9428 5228
rect 9292 4976 9332 4985
rect 9100 4936 9292 4976
rect 9004 4388 9044 4397
rect 8908 4348 9004 4388
rect 8811 4339 8853 4348
rect 9004 4339 9044 4348
rect 8812 4254 8852 4339
rect 9100 4229 9140 4936
rect 9292 4927 9332 4936
rect 9388 4565 9428 5188
rect 9484 4649 9524 5524
rect 9676 5144 9716 6943
rect 9771 6488 9813 6497
rect 9771 6448 9772 6488
rect 9812 6448 9813 6488
rect 9771 6439 9813 6448
rect 9772 5900 9812 6439
rect 9772 5851 9812 5860
rect 9676 5104 9812 5144
rect 9772 4985 9812 5104
rect 9580 4976 9620 4985
rect 9483 4640 9525 4649
rect 9483 4600 9484 4640
rect 9524 4600 9525 4640
rect 9483 4591 9525 4600
rect 9387 4556 9429 4565
rect 9387 4516 9388 4556
rect 9428 4516 9429 4556
rect 9387 4507 9429 4516
rect 9388 4313 9428 4507
rect 9387 4304 9429 4313
rect 9580 4304 9620 4936
rect 9676 4976 9716 4985
rect 9676 4640 9716 4936
rect 9771 4976 9813 4985
rect 9771 4936 9772 4976
rect 9812 4936 9813 4976
rect 9771 4927 9813 4936
rect 9868 4808 9908 7120
rect 10100 7120 10196 7160
rect 10060 7111 10100 7120
rect 9964 6992 10004 7001
rect 9964 5909 10004 6952
rect 10156 6656 10196 7120
rect 10252 6656 10292 6665
rect 10156 6616 10252 6656
rect 10348 6656 10388 7540
rect 10444 7412 10484 7960
rect 10636 7580 10676 8035
rect 10732 8000 10772 8009
rect 10732 7757 10772 7960
rect 10731 7748 10773 7757
rect 10731 7708 10732 7748
rect 10772 7708 10773 7748
rect 10731 7699 10773 7708
rect 10636 7540 10772 7580
rect 10444 7363 10484 7372
rect 10635 7244 10677 7253
rect 10635 7204 10636 7244
rect 10676 7204 10677 7244
rect 10732 7244 10772 7540
rect 10828 7412 10868 8128
rect 11116 8119 11156 8128
rect 10923 8084 10965 8093
rect 10923 8044 10924 8084
rect 10964 8044 10965 8084
rect 10923 8035 10965 8044
rect 10924 7950 10964 8035
rect 11020 7990 11300 8000
rect 11020 7960 11260 7990
rect 10923 7664 10965 7673
rect 10923 7624 10924 7664
rect 10964 7624 10965 7664
rect 10923 7615 10965 7624
rect 10828 7363 10868 7372
rect 10732 7204 10868 7244
rect 10635 7195 10677 7204
rect 10636 7110 10676 7195
rect 10635 6992 10677 7001
rect 10635 6952 10636 6992
rect 10676 6952 10677 6992
rect 10635 6943 10677 6952
rect 10348 6616 10580 6656
rect 10252 6607 10292 6616
rect 10060 6488 10100 6497
rect 10444 6488 10484 6497
rect 10060 6329 10100 6448
rect 10348 6448 10444 6488
rect 10059 6320 10101 6329
rect 10059 6280 10060 6320
rect 10100 6280 10101 6320
rect 10059 6271 10101 6280
rect 9963 5900 10005 5909
rect 9963 5860 9964 5900
rect 10004 5860 10005 5900
rect 9963 5851 10005 5860
rect 9997 5732 10039 5741
rect 9997 5692 9998 5732
rect 10038 5692 10039 5732
rect 9997 5683 10039 5692
rect 9998 5663 10038 5683
rect 9998 5597 10038 5623
rect 10156 5648 10196 5657
rect 10156 5489 10196 5608
rect 10252 5648 10292 5657
rect 10155 5480 10197 5489
rect 10155 5440 10156 5480
rect 10196 5440 10197 5480
rect 10155 5431 10197 5440
rect 10059 5228 10101 5237
rect 10059 5188 10060 5228
rect 10100 5188 10101 5228
rect 10059 5179 10101 5188
rect 9964 4808 10004 4817
rect 9868 4768 9964 4808
rect 9964 4759 10004 4768
rect 10060 4640 10100 5179
rect 10252 5144 10292 5608
rect 10348 5312 10388 6448
rect 10444 6439 10484 6448
rect 10444 6236 10484 6245
rect 10444 5648 10484 6196
rect 10540 6161 10580 6616
rect 10636 6488 10676 6943
rect 10636 6439 10676 6448
rect 10731 6488 10773 6497
rect 10731 6448 10732 6488
rect 10772 6448 10773 6488
rect 10731 6439 10773 6448
rect 10732 6354 10772 6439
rect 10828 6329 10868 7204
rect 10827 6320 10869 6329
rect 10827 6280 10828 6320
rect 10868 6280 10869 6320
rect 10827 6271 10869 6280
rect 10539 6152 10581 6161
rect 10539 6112 10540 6152
rect 10580 6112 10581 6152
rect 10539 6103 10581 6112
rect 10540 5909 10580 5994
rect 10924 5984 10964 7615
rect 11020 7412 11060 7960
rect 11260 7941 11300 7950
rect 11115 7832 11157 7841
rect 11115 7792 11116 7832
rect 11156 7792 11157 7832
rect 11115 7783 11157 7792
rect 11020 7363 11060 7372
rect 11019 6656 11061 6665
rect 11019 6616 11020 6656
rect 11060 6616 11061 6656
rect 11019 6607 11061 6616
rect 11020 6488 11060 6607
rect 11116 6488 11156 7783
rect 11307 7748 11349 7757
rect 11307 7708 11308 7748
rect 11348 7708 11349 7748
rect 11307 7699 11349 7708
rect 11212 7160 11252 7169
rect 11308 7160 11348 7699
rect 11252 7120 11348 7160
rect 11212 7111 11252 7120
rect 11404 6581 11444 8716
rect 11403 6572 11445 6581
rect 11403 6532 11404 6572
rect 11444 6532 11445 6572
rect 11403 6523 11445 6532
rect 11116 6448 11348 6488
rect 11020 5993 11060 6448
rect 11115 6320 11157 6329
rect 11115 6280 11116 6320
rect 11156 6280 11157 6320
rect 11115 6271 11157 6280
rect 11116 6068 11156 6271
rect 11308 6236 11348 6448
rect 11308 6196 11360 6236
rect 11320 6152 11360 6196
rect 11320 6112 11444 6152
rect 11116 6028 11348 6068
rect 10636 5944 10964 5984
rect 11019 5984 11061 5993
rect 11019 5944 11020 5984
rect 11060 5944 11061 5984
rect 10539 5900 10581 5909
rect 10539 5860 10540 5900
rect 10580 5860 10581 5900
rect 10539 5851 10581 5860
rect 10539 5732 10581 5741
rect 10539 5692 10540 5732
rect 10580 5692 10581 5732
rect 10539 5683 10581 5692
rect 10444 5599 10484 5608
rect 10540 5648 10580 5683
rect 10540 5597 10580 5608
rect 10348 5272 10580 5312
rect 10444 5144 10484 5153
rect 10252 5104 10444 5144
rect 10444 5095 10484 5104
rect 10155 4976 10197 4985
rect 10155 4936 10156 4976
rect 10196 4936 10197 4976
rect 10155 4927 10197 4936
rect 10252 4976 10292 4985
rect 10156 4842 10196 4927
rect 9676 4600 10100 4640
rect 9387 4264 9388 4304
rect 9428 4264 9429 4304
rect 9387 4255 9429 4264
rect 9484 4264 9620 4304
rect 9099 4220 9141 4229
rect 9099 4180 9100 4220
rect 9140 4180 9141 4220
rect 9099 4171 9141 4180
rect 9388 4136 9428 4145
rect 9292 4052 9332 4061
rect 8811 3800 8853 3809
rect 8811 3760 8812 3800
rect 8852 3760 8853 3800
rect 8811 3751 8853 3760
rect 8715 3632 8757 3641
rect 8715 3592 8716 3632
rect 8756 3592 8757 3632
rect 8715 3583 8757 3592
rect 8620 3415 8660 3424
rect 8716 3137 8756 3583
rect 8812 3464 8852 3751
rect 8907 3632 8949 3641
rect 9292 3632 9332 4012
rect 8907 3592 8908 3632
rect 8948 3592 8949 3632
rect 8907 3583 8949 3592
rect 9100 3592 9332 3632
rect 8908 3498 8948 3583
rect 9100 3473 9140 3592
rect 9388 3557 9428 4096
rect 9387 3548 9429 3557
rect 9387 3508 9388 3548
rect 9428 3508 9429 3548
rect 9387 3499 9429 3508
rect 8812 3415 8852 3424
rect 9099 3464 9141 3473
rect 9099 3424 9100 3464
rect 9140 3424 9141 3464
rect 9099 3415 9141 3424
rect 9196 3464 9236 3473
rect 8715 3128 8757 3137
rect 8715 3088 8716 3128
rect 8756 3088 8757 3128
rect 8715 3079 8757 3088
rect 8524 2920 8756 2960
rect 8524 2624 8564 2633
rect 8524 2540 8564 2584
rect 8428 2500 8564 2540
rect 8139 2456 8181 2465
rect 8332 2456 8372 2465
rect 8139 2416 8140 2456
rect 8180 2416 8276 2456
rect 8139 2407 8181 2416
rect 8236 1952 8276 2416
rect 8332 2213 8372 2416
rect 8524 2213 8564 2500
rect 8331 2204 8373 2213
rect 8331 2164 8332 2204
rect 8372 2164 8373 2204
rect 8331 2155 8373 2164
rect 8523 2204 8565 2213
rect 8523 2164 8524 2204
rect 8564 2164 8565 2204
rect 8523 2155 8565 2164
rect 8524 2036 8564 2045
rect 8236 1942 8372 1952
rect 8236 1912 8332 1942
rect 8332 1893 8372 1902
rect 8139 1868 8181 1877
rect 8139 1828 8140 1868
rect 8180 1828 8181 1868
rect 8139 1819 8181 1828
rect 8140 1457 8180 1819
rect 8524 1793 8564 1996
rect 8523 1784 8565 1793
rect 8523 1744 8524 1784
rect 8564 1744 8565 1784
rect 8523 1735 8565 1744
rect 8139 1448 8181 1457
rect 8139 1408 8140 1448
rect 8180 1408 8181 1448
rect 8139 1399 8181 1408
rect 8043 1280 8085 1289
rect 8043 1240 8044 1280
rect 8084 1240 8085 1280
rect 8043 1231 8085 1240
rect 7604 1072 7796 1112
rect 7851 1112 7893 1121
rect 7851 1072 7852 1112
rect 7892 1072 7893 1112
rect 7564 1063 7604 1072
rect 7851 1063 7893 1072
rect 8140 1112 8180 1399
rect 8140 1063 8180 1072
rect 7852 978 7892 1063
rect 8716 1028 8756 2920
rect 9100 2717 9140 3415
rect 9099 2708 9141 2717
rect 9099 2668 9100 2708
rect 9140 2668 9141 2708
rect 9099 2659 9141 2668
rect 9196 2465 9236 3424
rect 9292 3464 9332 3473
rect 9292 3221 9332 3424
rect 9291 3212 9333 3221
rect 9291 3172 9292 3212
rect 9332 3172 9333 3212
rect 9291 3163 9333 3172
rect 9292 2969 9332 3163
rect 9291 2960 9333 2969
rect 9291 2920 9292 2960
rect 9332 2920 9333 2960
rect 9291 2911 9333 2920
rect 9388 2633 9428 3499
rect 9484 2885 9524 4264
rect 9675 4220 9717 4229
rect 9675 4180 9676 4220
rect 9716 4180 9717 4220
rect 9675 4171 9717 4180
rect 9579 4136 9621 4145
rect 9579 4096 9580 4136
rect 9620 4096 9621 4136
rect 9579 4087 9621 4096
rect 9676 4136 9716 4171
rect 9580 3893 9620 4087
rect 9676 4085 9716 4096
rect 9771 4052 9813 4061
rect 9771 4012 9772 4052
rect 9812 4012 9813 4052
rect 9771 4003 9813 4012
rect 9579 3884 9621 3893
rect 9579 3844 9580 3884
rect 9620 3844 9621 3884
rect 9579 3835 9621 3844
rect 9483 2876 9525 2885
rect 9483 2836 9484 2876
rect 9524 2836 9525 2876
rect 9483 2827 9525 2836
rect 9387 2624 9429 2633
rect 9387 2584 9388 2624
rect 9428 2584 9429 2624
rect 9387 2575 9429 2584
rect 9195 2456 9237 2465
rect 9195 2416 9196 2456
rect 9236 2416 9237 2456
rect 9195 2407 9237 2416
rect 9196 1952 9236 2407
rect 9291 2372 9333 2381
rect 9291 2332 9292 2372
rect 9332 2332 9333 2372
rect 9291 2323 9333 2332
rect 9483 2372 9525 2381
rect 9483 2332 9484 2372
rect 9524 2332 9525 2372
rect 9483 2323 9525 2332
rect 9196 1903 9236 1912
rect 9292 1952 9332 2323
rect 9292 1903 9332 1912
rect 8620 988 8756 1028
rect 9388 1112 9428 1121
rect 9484 1112 9524 2323
rect 9580 1952 9620 3835
rect 9772 3632 9812 4003
rect 9867 3716 9909 3725
rect 9867 3676 9868 3716
rect 9908 3676 9909 3716
rect 9867 3667 9909 3676
rect 9772 3592 9816 3632
rect 9676 3380 9716 3391
rect 9776 3389 9816 3592
rect 9676 3305 9716 3340
rect 9772 3380 9816 3389
rect 9812 3340 9816 3380
rect 9772 3331 9812 3340
rect 9675 3296 9717 3305
rect 9675 3256 9676 3296
rect 9716 3256 9717 3296
rect 9675 3247 9717 3256
rect 9771 3212 9813 3221
rect 9771 3172 9772 3212
rect 9812 3172 9813 3212
rect 9771 3163 9813 3172
rect 9675 3128 9717 3137
rect 9675 3088 9676 3128
rect 9716 3088 9717 3128
rect 9675 3079 9717 3088
rect 9676 2204 9716 3079
rect 9772 2624 9812 3163
rect 9772 2381 9812 2584
rect 9771 2372 9813 2381
rect 9771 2332 9772 2372
rect 9812 2332 9813 2372
rect 9771 2323 9813 2332
rect 9676 2164 9812 2204
rect 9676 1952 9716 1961
rect 9580 1912 9676 1952
rect 9676 1903 9716 1912
rect 9772 1952 9812 2164
rect 9772 1903 9812 1912
rect 9579 1280 9621 1289
rect 9579 1240 9580 1280
rect 9620 1240 9621 1280
rect 9579 1231 9621 1240
rect 9580 1146 9620 1231
rect 9428 1072 9524 1112
rect 9771 1112 9813 1121
rect 9771 1072 9772 1112
rect 9812 1072 9813 1112
rect 6548 904 6836 944
rect 7563 944 7605 953
rect 7563 904 7564 944
rect 7604 904 7605 944
rect 6508 895 6548 904
rect 7563 895 7605 904
rect 6123 440 6165 449
rect 6123 400 6124 440
rect 6164 400 6165 440
rect 6123 391 6165 400
rect 6411 188 6453 197
rect 6411 148 6412 188
rect 6452 148 6453 188
rect 6411 139 6453 148
rect 6412 80 6452 139
rect 7564 80 7604 895
rect 8620 701 8660 988
rect 8715 860 8757 869
rect 8715 820 8716 860
rect 8756 820 8757 860
rect 8715 811 8757 820
rect 8619 692 8661 701
rect 8619 652 8620 692
rect 8660 652 8661 692
rect 8619 643 8661 652
rect 8716 80 8756 811
rect 9388 785 9428 1072
rect 9771 1063 9813 1072
rect 9772 978 9812 1063
rect 9387 776 9429 785
rect 9387 736 9388 776
rect 9428 736 9429 776
rect 9387 727 9429 736
rect 9868 80 9908 3667
rect 9964 3137 10004 4600
rect 10252 4397 10292 4936
rect 10443 4808 10485 4817
rect 10443 4768 10444 4808
rect 10484 4768 10485 4808
rect 10443 4759 10485 4768
rect 10347 4640 10389 4649
rect 10347 4600 10348 4640
rect 10388 4600 10389 4640
rect 10347 4591 10389 4600
rect 10251 4388 10293 4397
rect 10251 4348 10252 4388
rect 10292 4348 10293 4388
rect 10251 4339 10293 4348
rect 10348 4313 10388 4591
rect 10347 4304 10389 4313
rect 10347 4264 10348 4304
rect 10388 4264 10389 4304
rect 10347 4255 10389 4264
rect 10060 4136 10100 4145
rect 9963 3128 10005 3137
rect 9963 3088 9964 3128
rect 10004 3088 10005 3128
rect 9963 3079 10005 3088
rect 9964 2876 10004 2885
rect 10060 2876 10100 4096
rect 10348 4136 10388 4255
rect 10444 4136 10484 4759
rect 10540 4304 10580 5272
rect 10636 5237 10676 5944
rect 11019 5935 11061 5944
rect 10923 5816 10965 5825
rect 11212 5816 11252 5825
rect 10923 5776 10924 5816
rect 10964 5776 10965 5816
rect 10923 5767 10965 5776
rect 11020 5776 11212 5816
rect 10827 5732 10869 5741
rect 10827 5692 10828 5732
rect 10868 5692 10869 5732
rect 10827 5683 10869 5692
rect 10828 5648 10868 5683
rect 10828 5597 10868 5608
rect 10924 5648 10964 5767
rect 10924 5599 10964 5608
rect 10732 5422 10772 5431
rect 10635 5228 10677 5237
rect 10635 5188 10636 5228
rect 10676 5188 10677 5228
rect 10635 5179 10677 5188
rect 10732 5069 10772 5382
rect 10731 5060 10773 5069
rect 10731 5020 10732 5060
rect 10772 5020 10773 5060
rect 10731 5011 10773 5020
rect 10635 4976 10677 4985
rect 10635 4936 10636 4976
rect 10676 4936 10677 4976
rect 10635 4927 10677 4936
rect 10636 4842 10676 4927
rect 10731 4472 10773 4481
rect 10731 4432 10732 4472
rect 10772 4432 10773 4472
rect 10731 4423 10773 4432
rect 10540 4264 10676 4304
rect 10540 4136 10580 4145
rect 10444 4096 10540 4136
rect 10348 4087 10388 4096
rect 10155 3968 10197 3977
rect 10155 3928 10156 3968
rect 10196 3928 10197 3968
rect 10155 3919 10197 3928
rect 10252 3968 10292 3977
rect 10292 3928 10484 3968
rect 10252 3919 10292 3928
rect 10156 3548 10196 3919
rect 10347 3800 10389 3809
rect 10347 3760 10348 3800
rect 10388 3760 10389 3800
rect 10347 3751 10389 3760
rect 10251 3548 10293 3557
rect 10156 3508 10252 3548
rect 10292 3508 10293 3548
rect 10251 3499 10293 3508
rect 10251 3473 10291 3499
rect 10251 3414 10291 3433
rect 10348 3296 10388 3751
rect 10004 2836 10100 2876
rect 9964 2827 10004 2836
rect 10060 2465 10100 2836
rect 10156 3256 10388 3296
rect 10156 2717 10196 3256
rect 10251 2792 10293 2801
rect 10251 2752 10252 2792
rect 10292 2752 10293 2792
rect 10251 2743 10293 2752
rect 10155 2708 10197 2717
rect 10155 2668 10156 2708
rect 10196 2668 10197 2708
rect 10155 2659 10197 2668
rect 10059 2456 10101 2465
rect 10059 2416 10060 2456
rect 10100 2416 10101 2456
rect 10059 2407 10101 2416
rect 10060 2045 10100 2407
rect 10059 2036 10101 2045
rect 10059 1996 10060 2036
rect 10100 1996 10101 2036
rect 10059 1987 10101 1996
rect 10156 1952 10196 2659
rect 10252 2624 10292 2743
rect 10348 2633 10388 2718
rect 10252 2120 10292 2584
rect 10347 2624 10389 2633
rect 10347 2584 10348 2624
rect 10388 2584 10389 2624
rect 10347 2575 10389 2584
rect 10252 2080 10388 2120
rect 10252 1952 10292 1961
rect 10156 1912 10252 1952
rect 10252 1903 10292 1912
rect 10348 1289 10388 2080
rect 10347 1280 10389 1289
rect 10347 1240 10348 1280
rect 10388 1240 10389 1280
rect 10347 1231 10389 1240
rect 10444 869 10484 3928
rect 10540 3893 10580 4096
rect 10539 3884 10581 3893
rect 10539 3844 10540 3884
rect 10580 3844 10581 3884
rect 10539 3835 10581 3844
rect 10636 3641 10676 4264
rect 10732 3977 10772 4423
rect 10731 3968 10773 3977
rect 10731 3928 10732 3968
rect 10772 3928 10773 3968
rect 10731 3919 10773 3928
rect 10635 3632 10677 3641
rect 10635 3592 10636 3632
rect 10676 3592 10677 3632
rect 10635 3583 10677 3592
rect 10923 3548 10965 3557
rect 10923 3508 10924 3548
rect 10964 3508 10965 3548
rect 10923 3499 10965 3508
rect 10827 3464 10869 3473
rect 10732 3450 10772 3459
rect 10827 3424 10828 3464
rect 10868 3424 10869 3464
rect 10827 3415 10869 3424
rect 10635 3212 10677 3221
rect 10635 3172 10636 3212
rect 10676 3172 10677 3212
rect 10635 3163 10677 3172
rect 10636 2885 10676 3163
rect 10635 2876 10677 2885
rect 10635 2836 10636 2876
rect 10676 2836 10677 2876
rect 10635 2827 10677 2836
rect 10636 2624 10676 2827
rect 10732 2801 10772 3410
rect 10828 3053 10868 3415
rect 10924 3414 10964 3499
rect 10827 3044 10869 3053
rect 10827 3004 10828 3044
rect 10868 3004 10869 3044
rect 10827 2995 10869 3004
rect 10731 2792 10773 2801
rect 10731 2752 10732 2792
rect 10772 2752 10773 2792
rect 10731 2743 10773 2752
rect 10828 2708 10868 2995
rect 10828 2659 10868 2668
rect 10732 2624 10772 2633
rect 10636 2584 10732 2624
rect 10732 2575 10772 2584
rect 10923 2540 10965 2549
rect 10828 2500 10924 2540
rect 10964 2500 10965 2540
rect 10828 2456 10868 2500
rect 10923 2491 10965 2500
rect 10732 2416 10868 2456
rect 10732 1938 10772 2416
rect 10923 2120 10965 2129
rect 10923 2080 10924 2120
rect 10964 2080 10965 2120
rect 10923 2071 10965 2080
rect 10924 1986 10964 2071
rect 10732 1289 10772 1898
rect 10731 1280 10773 1289
rect 10731 1240 10732 1280
rect 10772 1240 10773 1280
rect 11020 1280 11060 5776
rect 11212 5767 11252 5776
rect 11308 5321 11348 6028
rect 11307 5312 11349 5321
rect 11307 5272 11308 5312
rect 11348 5272 11349 5312
rect 11307 5263 11349 5272
rect 11404 5144 11444 6112
rect 11500 5900 11540 9640
rect 11596 8924 11636 10672
rect 11788 9017 11828 10672
rect 11883 10352 11925 10361
rect 11883 10312 11884 10352
rect 11924 10312 11925 10352
rect 11883 10303 11925 10312
rect 11787 9008 11829 9017
rect 11787 8968 11788 9008
rect 11828 8968 11829 9008
rect 11787 8959 11829 8968
rect 11596 8884 11732 8924
rect 11596 8756 11636 8765
rect 11596 8513 11636 8716
rect 11595 8504 11637 8513
rect 11595 8464 11596 8504
rect 11636 8464 11637 8504
rect 11595 8455 11637 8464
rect 11692 8168 11732 8884
rect 11788 8840 11828 8849
rect 11884 8840 11924 10303
rect 11980 8924 12020 10672
rect 12172 10361 12212 10672
rect 12267 10604 12309 10613
rect 12267 10564 12268 10604
rect 12308 10564 12309 10604
rect 12267 10555 12309 10564
rect 12171 10352 12213 10361
rect 12171 10312 12172 10352
rect 12212 10312 12213 10352
rect 12171 10303 12213 10312
rect 12171 10184 12213 10193
rect 12171 10144 12172 10184
rect 12212 10144 12213 10184
rect 12171 10135 12213 10144
rect 11980 8884 12116 8924
rect 11828 8800 11924 8840
rect 11788 8791 11828 8800
rect 11979 8756 12021 8765
rect 11979 8716 11980 8756
rect 12020 8716 12021 8756
rect 11979 8707 12021 8716
rect 11980 8622 12020 8707
rect 11692 8128 11924 8168
rect 11788 8000 11828 8009
rect 11788 7505 11828 7960
rect 11787 7496 11829 7505
rect 11787 7456 11788 7496
rect 11828 7456 11829 7496
rect 11787 7447 11829 7456
rect 11595 6740 11637 6749
rect 11595 6700 11596 6740
rect 11636 6700 11637 6740
rect 11595 6691 11637 6700
rect 11500 5851 11540 5860
rect 11596 5564 11636 6691
rect 11692 5741 11732 5826
rect 11691 5732 11733 5741
rect 11691 5692 11692 5732
rect 11732 5692 11733 5732
rect 11691 5683 11733 5692
rect 11596 5524 11732 5564
rect 11595 5228 11637 5237
rect 11595 5188 11596 5228
rect 11636 5188 11637 5228
rect 11595 5179 11637 5188
rect 11308 5104 11444 5144
rect 11212 3464 11252 3473
rect 11116 3424 11212 3464
rect 11116 1952 11156 3424
rect 11212 3415 11252 3424
rect 11211 3128 11253 3137
rect 11211 3088 11212 3128
rect 11252 3088 11253 3128
rect 11211 3079 11253 3088
rect 11212 2624 11252 3079
rect 11308 2801 11348 5104
rect 11596 3725 11636 5179
rect 11595 3716 11637 3725
rect 11595 3676 11596 3716
rect 11636 3676 11637 3716
rect 11595 3667 11637 3676
rect 11499 3464 11541 3473
rect 11499 3424 11500 3464
rect 11540 3424 11541 3464
rect 11499 3415 11541 3424
rect 11596 3464 11636 3473
rect 11403 3380 11445 3389
rect 11403 3340 11404 3380
rect 11444 3340 11445 3380
rect 11403 3331 11445 3340
rect 11307 2792 11349 2801
rect 11307 2752 11308 2792
rect 11348 2752 11349 2792
rect 11307 2743 11349 2752
rect 11308 2624 11348 2633
rect 11212 2584 11308 2624
rect 11308 2575 11348 2584
rect 11211 2456 11253 2465
rect 11404 2456 11444 3331
rect 11500 3330 11540 3415
rect 11211 2416 11212 2456
rect 11252 2416 11253 2456
rect 11211 2407 11253 2416
rect 11308 2416 11444 2456
rect 11116 1700 11156 1912
rect 11212 1952 11252 2407
rect 11212 1903 11252 1912
rect 11308 1952 11348 2416
rect 11596 2129 11636 3424
rect 11595 2120 11637 2129
rect 11595 2080 11596 2120
rect 11636 2080 11637 2120
rect 11595 2071 11637 2080
rect 11308 1903 11348 1912
rect 11403 1952 11445 1961
rect 11403 1912 11404 1952
rect 11444 1912 11445 1952
rect 11403 1903 11445 1912
rect 11404 1818 11444 1903
rect 11596 1700 11636 1709
rect 11116 1660 11252 1700
rect 11212 1364 11252 1660
rect 11212 1289 11252 1324
rect 11404 1660 11596 1700
rect 11211 1280 11253 1289
rect 11020 1240 11156 1280
rect 10731 1231 10773 1240
rect 11020 1112 11060 1121
rect 10924 1072 11020 1112
rect 10443 860 10485 869
rect 10443 820 10444 860
rect 10484 820 10485 860
rect 10443 811 10485 820
rect 10924 785 10964 1072
rect 11020 1063 11060 1072
rect 11116 944 11156 1240
rect 11211 1240 11212 1280
rect 11252 1240 11253 1280
rect 11211 1231 11253 1240
rect 11212 1200 11252 1231
rect 11404 1112 11444 1660
rect 11596 1651 11636 1660
rect 11692 1448 11732 5524
rect 11788 5237 11828 7447
rect 11884 5900 11924 8128
rect 12076 7589 12116 8884
rect 12172 8840 12212 10135
rect 12172 8791 12212 8800
rect 12171 8420 12213 8429
rect 12171 8380 12172 8420
rect 12212 8380 12213 8420
rect 12171 8371 12213 8380
rect 12075 7580 12117 7589
rect 12075 7540 12076 7580
rect 12116 7540 12117 7580
rect 12075 7531 12117 7540
rect 11979 6320 12021 6329
rect 11979 6280 11980 6320
rect 12020 6280 12021 6320
rect 11979 6271 12021 6280
rect 11884 5851 11924 5860
rect 11787 5228 11829 5237
rect 11787 5188 11788 5228
rect 11828 5188 11829 5228
rect 11787 5179 11829 5188
rect 11884 4976 11924 4985
rect 11980 4976 12020 6271
rect 12172 5900 12212 8371
rect 12268 8000 12308 10555
rect 12364 10016 12404 10672
rect 12556 10193 12596 10672
rect 12555 10184 12597 10193
rect 12555 10144 12556 10184
rect 12596 10144 12597 10184
rect 12555 10135 12597 10144
rect 12748 10016 12788 10672
rect 12940 10100 12980 10672
rect 13132 10184 13172 10672
rect 13132 10144 13268 10184
rect 12940 10060 13172 10100
rect 12364 9976 12692 10016
rect 12748 9976 13076 10016
rect 12652 9680 12692 9976
rect 12652 9631 12692 9640
rect 13036 9680 13076 9976
rect 13036 9631 13076 9640
rect 13035 9512 13077 9521
rect 13035 9472 13036 9512
rect 13076 9472 13077 9512
rect 13035 9463 13077 9472
rect 12844 9428 12884 9437
rect 12884 9388 12980 9428
rect 12844 9379 12884 9388
rect 12459 9344 12501 9353
rect 12459 9304 12460 9344
rect 12500 9304 12501 9344
rect 12459 9295 12501 9304
rect 12363 9008 12405 9017
rect 12363 8968 12364 9008
rect 12404 8968 12405 9008
rect 12363 8959 12405 8968
rect 12364 8672 12404 8959
rect 12364 8623 12404 8632
rect 12268 7951 12308 7960
rect 12364 7916 12404 7925
rect 12268 6488 12308 6497
rect 12268 6329 12308 6448
rect 12267 6320 12309 6329
rect 12267 6280 12268 6320
rect 12308 6280 12309 6320
rect 12267 6271 12309 6280
rect 12364 6245 12404 7876
rect 12460 7160 12500 9295
rect 12747 9092 12789 9101
rect 12747 9052 12748 9092
rect 12788 9052 12789 9092
rect 12747 9043 12789 9052
rect 12748 8000 12788 9043
rect 12748 7951 12788 7960
rect 12843 8000 12885 8009
rect 12843 7960 12844 8000
rect 12884 7960 12885 8000
rect 12843 7951 12885 7960
rect 12844 7866 12884 7951
rect 12651 7580 12693 7589
rect 12651 7540 12652 7580
rect 12692 7540 12693 7580
rect 12651 7531 12693 7540
rect 12652 7412 12692 7531
rect 12652 7363 12692 7372
rect 12843 7244 12885 7253
rect 12843 7204 12844 7244
rect 12884 7204 12885 7244
rect 12843 7195 12885 7204
rect 12460 7111 12500 7120
rect 12844 7110 12884 7195
rect 12747 6908 12789 6917
rect 12747 6868 12748 6908
rect 12788 6868 12789 6908
rect 12747 6859 12789 6868
rect 12459 6656 12501 6665
rect 12459 6616 12460 6656
rect 12500 6616 12501 6656
rect 12459 6607 12501 6616
rect 12460 6522 12500 6607
rect 12651 6488 12693 6497
rect 12651 6448 12652 6488
rect 12692 6448 12693 6488
rect 12651 6439 12693 6448
rect 12363 6236 12405 6245
rect 12363 6196 12364 6236
rect 12404 6196 12405 6236
rect 12363 6187 12405 6196
rect 12652 6077 12692 6439
rect 12651 6068 12693 6077
rect 12651 6028 12652 6068
rect 12692 6028 12693 6068
rect 12651 6019 12693 6028
rect 12268 5900 12308 5909
rect 12172 5860 12268 5900
rect 12268 5851 12308 5860
rect 12076 5732 12116 5741
rect 12076 5237 12116 5692
rect 12460 5732 12500 5741
rect 12500 5692 12596 5732
rect 12460 5683 12500 5692
rect 12075 5228 12117 5237
rect 12075 5188 12076 5228
rect 12116 5188 12117 5228
rect 12075 5179 12117 5188
rect 12076 5060 12116 5069
rect 12116 5020 12404 5060
rect 12076 5011 12116 5020
rect 11924 4936 12020 4976
rect 11884 4927 11924 4936
rect 11980 4808 12020 4936
rect 12364 4976 12404 5020
rect 12364 4927 12404 4936
rect 12460 4976 12500 4985
rect 11980 4768 12308 4808
rect 11979 4640 12021 4649
rect 11979 4600 11980 4640
rect 12020 4600 12021 4640
rect 11979 4591 12021 4600
rect 11980 4229 12020 4591
rect 11979 4220 12021 4229
rect 11979 4180 11980 4220
rect 12020 4180 12021 4220
rect 11979 4171 12021 4180
rect 12171 4220 12213 4229
rect 12171 4180 12172 4220
rect 12212 4180 12213 4220
rect 12171 4171 12213 4180
rect 11787 4136 11829 4145
rect 11787 4096 11788 4136
rect 11828 4096 11829 4136
rect 11787 4087 11829 4096
rect 12172 4136 12212 4171
rect 11788 4002 11828 4087
rect 12172 4085 12212 4096
rect 12268 3977 12308 4768
rect 12460 4724 12500 4936
rect 12364 4684 12500 4724
rect 11883 3968 11925 3977
rect 11883 3928 11884 3968
rect 11924 3928 11925 3968
rect 11883 3919 11925 3928
rect 11980 3968 12020 3977
rect 12267 3968 12309 3977
rect 12020 3928 12116 3968
rect 11980 3919 12020 3928
rect 11884 3716 11924 3919
rect 11788 3676 11924 3716
rect 11788 2960 11828 3676
rect 12076 3473 12116 3928
rect 12267 3928 12268 3968
rect 12308 3928 12309 3968
rect 12267 3919 12309 3928
rect 12364 3809 12404 4684
rect 12459 4556 12501 4565
rect 12459 4516 12460 4556
rect 12500 4516 12501 4556
rect 12459 4507 12501 4516
rect 12363 3800 12405 3809
rect 12363 3760 12364 3800
rect 12404 3760 12405 3800
rect 12363 3751 12405 3760
rect 12364 3632 12404 3641
rect 12268 3592 12364 3632
rect 12075 3464 12117 3473
rect 12075 3424 12076 3464
rect 12116 3424 12117 3464
rect 12075 3415 12117 3424
rect 12172 3464 12212 3473
rect 11884 3296 11924 3305
rect 12172 3296 12212 3424
rect 11924 3256 12212 3296
rect 11884 3247 11924 3256
rect 12268 3044 12308 3592
rect 12364 3583 12404 3592
rect 12460 3212 12500 4507
rect 12556 4145 12596 5692
rect 12748 4229 12788 6859
rect 12940 5573 12980 9388
rect 12939 5564 12981 5573
rect 12939 5524 12940 5564
rect 12980 5524 12981 5564
rect 12939 5515 12981 5524
rect 12844 4892 12884 4901
rect 12844 4649 12884 4852
rect 12940 4892 12980 4901
rect 12843 4640 12885 4649
rect 12843 4600 12844 4640
rect 12884 4600 12885 4640
rect 12843 4591 12885 4600
rect 12747 4220 12789 4229
rect 12747 4180 12748 4220
rect 12788 4180 12789 4220
rect 12747 4171 12789 4180
rect 12555 4136 12597 4145
rect 12555 4096 12556 4136
rect 12596 4096 12597 4136
rect 12555 4087 12597 4096
rect 12940 4061 12980 4852
rect 12939 4052 12981 4061
rect 12939 4012 12940 4052
rect 12980 4012 12981 4052
rect 12939 4003 12981 4012
rect 13036 3641 13076 9463
rect 13132 5900 13172 10060
rect 13228 9605 13268 10144
rect 13227 9596 13269 9605
rect 13227 9556 13228 9596
rect 13268 9556 13269 9596
rect 13227 9547 13269 9556
rect 13227 9428 13269 9437
rect 13227 9388 13228 9428
rect 13268 9388 13269 9428
rect 13227 9379 13269 9388
rect 13228 9294 13268 9379
rect 13324 7328 13364 10672
rect 13516 8849 13556 10672
rect 13708 8849 13748 10672
rect 13900 9941 13940 10672
rect 13899 9932 13941 9941
rect 13899 9892 13900 9932
rect 13940 9892 13941 9932
rect 13899 9883 13941 9892
rect 14092 9521 14132 10672
rect 14091 9512 14133 9521
rect 14091 9472 14092 9512
rect 14132 9472 14133 9512
rect 14091 9463 14133 9472
rect 13803 8924 13845 8933
rect 13803 8884 13804 8924
rect 13844 8884 13845 8924
rect 13803 8875 13845 8884
rect 13515 8840 13557 8849
rect 13515 8800 13516 8840
rect 13556 8800 13557 8840
rect 13515 8791 13557 8800
rect 13707 8840 13749 8849
rect 13707 8800 13708 8840
rect 13748 8800 13749 8840
rect 13707 8791 13749 8800
rect 13612 8672 13652 8681
rect 13804 8672 13844 8875
rect 14284 8849 14324 10672
rect 14476 9680 14516 10672
rect 14668 10613 14708 10672
rect 14667 10604 14709 10613
rect 14667 10564 14668 10604
rect 14708 10564 14709 10604
rect 14667 10555 14709 10564
rect 14860 9773 14900 10672
rect 14955 10604 14997 10613
rect 14955 10564 14956 10604
rect 14996 10564 14997 10604
rect 14955 10555 14997 10564
rect 14859 9764 14901 9773
rect 14859 9724 14860 9764
rect 14900 9724 14901 9764
rect 14859 9715 14901 9724
rect 14764 9680 14804 9689
rect 14476 9640 14764 9680
rect 14764 9631 14804 9640
rect 14956 9596 14996 10555
rect 14860 9556 14996 9596
rect 14283 8840 14325 8849
rect 14283 8800 14284 8840
rect 14324 8800 14325 8840
rect 14283 8791 14325 8800
rect 14140 8681 14180 8690
rect 13612 7757 13652 8632
rect 13708 8632 13844 8672
rect 14092 8641 14140 8672
rect 14092 8632 14180 8641
rect 14668 8672 14708 8681
rect 13611 7748 13653 7757
rect 13611 7708 13612 7748
rect 13652 7708 13653 7748
rect 13611 7699 13653 7708
rect 13324 7288 13556 7328
rect 13324 7160 13364 7169
rect 13324 6665 13364 7120
rect 13420 7160 13460 7169
rect 13420 7085 13460 7120
rect 13419 7076 13461 7085
rect 13419 7036 13420 7076
rect 13460 7036 13461 7076
rect 13419 7027 13461 7036
rect 13420 6917 13460 7027
rect 13419 6908 13461 6917
rect 13419 6868 13420 6908
rect 13460 6868 13461 6908
rect 13419 6859 13461 6868
rect 13323 6656 13365 6665
rect 13323 6616 13324 6656
rect 13364 6616 13365 6656
rect 13323 6607 13365 6616
rect 13228 5900 13268 5909
rect 13132 5860 13228 5900
rect 13228 5851 13268 5860
rect 13420 5732 13460 5741
rect 13324 5692 13420 5732
rect 13324 4985 13364 5692
rect 13420 5683 13460 5692
rect 13323 4976 13365 4985
rect 13323 4936 13324 4976
rect 13364 4936 13365 4976
rect 13323 4927 13365 4936
rect 13420 4976 13460 4985
rect 13420 4304 13460 4936
rect 13324 4264 13460 4304
rect 13227 4220 13269 4229
rect 13227 4180 13228 4220
rect 13268 4180 13269 4220
rect 13227 4171 13269 4180
rect 13035 3632 13077 3641
rect 13035 3592 13036 3632
rect 13076 3592 13077 3632
rect 13035 3583 13077 3592
rect 12555 3464 12597 3473
rect 12555 3424 12556 3464
rect 12596 3424 12597 3464
rect 12555 3415 12597 3424
rect 12556 3330 12596 3415
rect 12460 3172 12596 3212
rect 12076 3004 12308 3044
rect 11883 2960 11925 2969
rect 11788 2920 11884 2960
rect 11924 2920 11925 2960
rect 11883 2911 11925 2920
rect 11788 2629 11828 2638
rect 11788 2129 11828 2589
rect 11884 2204 11924 2911
rect 11979 2456 12021 2465
rect 11979 2416 11980 2456
rect 12020 2416 12021 2456
rect 11979 2407 12021 2416
rect 11980 2322 12020 2407
rect 11884 2164 12020 2204
rect 11787 2120 11829 2129
rect 11787 2080 11788 2120
rect 11828 2080 11829 2120
rect 11787 2071 11829 2080
rect 11883 2036 11925 2045
rect 11883 1996 11884 2036
rect 11924 1996 11925 2036
rect 11883 1987 11925 1996
rect 11884 1902 11924 1987
rect 11980 1952 12020 2164
rect 11980 1903 12020 1912
rect 11787 1868 11829 1877
rect 11787 1828 11788 1868
rect 11828 1828 11829 1868
rect 11787 1819 11829 1828
rect 11788 1532 11828 1819
rect 11788 1492 12020 1532
rect 11596 1408 11732 1448
rect 11499 1196 11541 1205
rect 11499 1156 11500 1196
rect 11540 1156 11541 1196
rect 11499 1147 11541 1156
rect 11404 1063 11444 1072
rect 11500 1112 11540 1147
rect 11500 1061 11540 1072
rect 11020 904 11156 944
rect 10923 776 10965 785
rect 10923 736 10924 776
rect 10964 736 10965 776
rect 10923 727 10965 736
rect 11020 80 11060 904
rect 2936 0 3016 80
rect 4088 0 4168 80
rect 5240 0 5320 80
rect 6392 0 6472 80
rect 7544 0 7624 80
rect 8696 0 8776 80
rect 9848 0 9928 80
rect 11000 0 11080 80
rect 11596 60 11636 1408
rect 11692 1280 11732 1289
rect 11732 1240 11924 1280
rect 11692 1231 11732 1240
rect 11691 1112 11733 1121
rect 11691 1072 11692 1112
rect 11732 1072 11733 1112
rect 11691 1063 11733 1072
rect 11884 1112 11924 1240
rect 11884 1063 11924 1072
rect 11980 1112 12020 1492
rect 11980 1063 12020 1072
rect 12076 1112 12116 3004
rect 12268 2633 12308 2718
rect 12267 2624 12309 2633
rect 12267 2584 12268 2624
rect 12308 2584 12309 2624
rect 12267 2575 12309 2584
rect 12460 2624 12500 2633
rect 12172 2456 12212 2465
rect 12172 1205 12212 2416
rect 12267 1952 12309 1961
rect 12267 1912 12268 1952
rect 12308 1912 12309 1952
rect 12267 1903 12309 1912
rect 12268 1818 12308 1903
rect 12460 1877 12500 2584
rect 12556 2045 12596 3172
rect 12939 2624 12981 2633
rect 12939 2584 12940 2624
rect 12980 2584 12981 2624
rect 12939 2575 12981 2584
rect 12651 2372 12693 2381
rect 12651 2332 12652 2372
rect 12692 2332 12693 2372
rect 12651 2323 12693 2332
rect 12555 2036 12597 2045
rect 12555 1996 12556 2036
rect 12596 1996 12597 2036
rect 12555 1987 12597 1996
rect 12652 1952 12692 2323
rect 12747 2204 12789 2213
rect 12747 2164 12748 2204
rect 12788 2164 12789 2204
rect 12747 2155 12789 2164
rect 12459 1868 12501 1877
rect 12459 1828 12460 1868
rect 12500 1828 12501 1868
rect 12459 1819 12501 1828
rect 12460 1532 12500 1819
rect 12268 1492 12500 1532
rect 12171 1196 12213 1205
rect 12171 1156 12172 1196
rect 12212 1156 12213 1196
rect 12171 1147 12213 1156
rect 12076 1063 12116 1072
rect 11692 978 11732 1063
rect 12171 944 12213 953
rect 12171 904 12172 944
rect 12212 904 12213 944
rect 12171 895 12213 904
rect 12172 810 12212 895
rect 12268 281 12308 1492
rect 12652 1457 12692 1912
rect 12651 1448 12693 1457
rect 12651 1408 12652 1448
rect 12692 1408 12693 1448
rect 12651 1399 12693 1408
rect 12748 1289 12788 2155
rect 12459 1280 12501 1289
rect 12459 1240 12460 1280
rect 12500 1240 12501 1280
rect 12459 1231 12501 1240
rect 12747 1280 12789 1289
rect 12747 1240 12748 1280
rect 12788 1240 12789 1280
rect 12747 1231 12789 1240
rect 12363 1112 12405 1121
rect 12363 1072 12364 1112
rect 12404 1072 12405 1112
rect 12363 1063 12405 1072
rect 12460 1112 12500 1231
rect 12460 1063 12500 1072
rect 12555 1112 12597 1121
rect 12555 1072 12556 1112
rect 12596 1072 12597 1112
rect 12555 1063 12597 1072
rect 12652 1112 12692 1121
rect 12364 978 12404 1063
rect 12556 978 12596 1063
rect 12652 869 12692 1072
rect 12843 1112 12885 1121
rect 12843 1072 12844 1112
rect 12884 1072 12885 1112
rect 12843 1063 12885 1072
rect 12940 1112 12980 2575
rect 13035 1952 13077 1961
rect 13035 1912 13036 1952
rect 13076 1912 13077 1952
rect 13035 1903 13077 1912
rect 12940 1063 12980 1072
rect 13036 1112 13076 1903
rect 13036 1063 13076 1072
rect 13132 1112 13172 1121
rect 13228 1112 13268 4171
rect 13324 2801 13364 4264
rect 13420 4136 13460 4145
rect 13420 3977 13460 4096
rect 13419 3968 13461 3977
rect 13419 3928 13420 3968
rect 13460 3928 13461 3968
rect 13419 3919 13461 3928
rect 13323 2792 13365 2801
rect 13323 2752 13324 2792
rect 13364 2752 13365 2792
rect 13323 2743 13365 2752
rect 13172 1072 13268 1112
rect 13132 1063 13172 1072
rect 12844 978 12884 1063
rect 12651 860 12693 869
rect 12651 820 12652 860
rect 12692 820 12693 860
rect 12651 811 12693 820
rect 12267 272 12309 281
rect 12267 232 12268 272
rect 12308 232 12309 272
rect 12267 223 12309 232
rect 11980 148 12217 188
rect 11980 60 12020 148
rect 12177 104 12217 148
rect 12172 80 12217 104
rect 13324 80 13364 2743
rect 13516 1280 13556 7288
rect 13708 5900 13748 8632
rect 13899 8588 13941 8597
rect 13804 8548 13900 8588
rect 13940 8548 13941 8588
rect 13804 8504 13844 8548
rect 13899 8539 13941 8548
rect 13804 8455 13844 8464
rect 13996 8504 14036 8513
rect 13996 8345 14036 8464
rect 13995 8336 14037 8345
rect 13995 8296 13996 8336
rect 14036 8296 14037 8336
rect 13995 8287 14037 8296
rect 13996 8168 14036 8177
rect 14092 8168 14132 8632
rect 14668 8345 14708 8632
rect 14667 8336 14709 8345
rect 14667 8296 14668 8336
rect 14708 8296 14709 8336
rect 14667 8287 14709 8296
rect 14036 8128 14132 8168
rect 13996 8119 14036 8128
rect 14188 8000 14228 8009
rect 14188 7757 14228 7960
rect 14187 7748 14229 7757
rect 14187 7708 14188 7748
rect 14228 7708 14229 7748
rect 14187 7699 14229 7708
rect 14379 7496 14421 7505
rect 14379 7456 14380 7496
rect 14420 7456 14421 7496
rect 14379 7447 14421 7456
rect 13803 7328 13845 7337
rect 13803 7288 13804 7328
rect 13844 7288 13845 7328
rect 13803 7279 13845 7288
rect 13804 7244 13844 7279
rect 13804 7193 13844 7204
rect 13899 7160 13941 7169
rect 13899 7120 13900 7160
rect 13940 7120 13941 7160
rect 13899 7111 13941 7120
rect 14380 7160 14420 7447
rect 14860 7328 14900 9556
rect 14955 9428 14997 9437
rect 14955 9388 14956 9428
rect 14996 9388 14997 9428
rect 14955 9379 14997 9388
rect 14956 9294 14996 9379
rect 15052 8849 15092 10672
rect 15244 10193 15284 10672
rect 15243 10184 15285 10193
rect 15243 10144 15244 10184
rect 15284 10144 15285 10184
rect 15243 10135 15285 10144
rect 15243 10016 15285 10025
rect 15243 9976 15244 10016
rect 15284 9976 15285 10016
rect 15243 9967 15285 9976
rect 15147 9680 15189 9689
rect 15147 9640 15148 9680
rect 15188 9640 15189 9680
rect 15147 9631 15189 9640
rect 15148 9512 15188 9631
rect 15148 9463 15188 9472
rect 15244 9101 15284 9967
rect 15339 9428 15381 9437
rect 15339 9388 15340 9428
rect 15380 9388 15381 9428
rect 15339 9379 15381 9388
rect 15243 9092 15285 9101
rect 15243 9052 15244 9092
rect 15284 9052 15285 9092
rect 15243 9043 15285 9052
rect 15051 8840 15093 8849
rect 15051 8800 15052 8840
rect 15092 8800 15093 8840
rect 15051 8791 15093 8800
rect 15244 8756 15284 9043
rect 15244 8707 15284 8716
rect 15147 8672 15189 8681
rect 15147 8632 15148 8672
rect 15188 8632 15189 8672
rect 15147 8623 15189 8632
rect 14860 7288 14996 7328
rect 14380 7111 14420 7120
rect 14860 7165 14900 7174
rect 13900 7001 13940 7111
rect 13899 6992 13941 7001
rect 13899 6952 13900 6992
rect 13940 6952 13941 6992
rect 13899 6943 13941 6952
rect 14860 6740 14900 7125
rect 14092 6700 14900 6740
rect 14092 6656 14132 6700
rect 14092 6607 14132 6616
rect 13900 6488 13940 6497
rect 13900 6329 13940 6448
rect 14283 6488 14325 6497
rect 14283 6448 14284 6488
rect 14324 6448 14325 6488
rect 14283 6439 14325 6448
rect 13899 6320 13941 6329
rect 13899 6280 13900 6320
rect 13940 6280 13941 6320
rect 13899 6271 13941 6280
rect 13804 5900 13844 5909
rect 13708 5860 13804 5900
rect 13804 5851 13844 5860
rect 13995 5816 14037 5825
rect 13995 5776 13996 5816
rect 14036 5776 14037 5816
rect 13995 5767 14037 5776
rect 13612 5732 13652 5741
rect 13612 5069 13652 5692
rect 13996 5648 14036 5767
rect 14284 5657 14324 6439
rect 13996 5405 14036 5608
rect 14283 5648 14325 5657
rect 14283 5608 14284 5648
rect 14324 5608 14325 5648
rect 14283 5599 14325 5608
rect 14475 5480 14517 5489
rect 14475 5440 14476 5480
rect 14516 5440 14517 5480
rect 14475 5431 14517 5440
rect 13995 5396 14037 5405
rect 13995 5356 13996 5396
rect 14036 5356 14037 5396
rect 13995 5347 14037 5356
rect 13611 5060 13653 5069
rect 13611 5020 13612 5060
rect 13652 5020 13653 5060
rect 13611 5011 13653 5020
rect 14091 5060 14133 5069
rect 14091 5020 14092 5060
rect 14132 5020 14133 5060
rect 14091 5011 14133 5020
rect 13900 4962 13940 4971
rect 14092 4926 14132 5011
rect 13900 4472 13940 4922
rect 13612 4432 13940 4472
rect 13612 4388 13652 4432
rect 13995 4388 14037 4397
rect 13612 4339 13652 4348
rect 13900 4348 13996 4388
rect 14036 4348 14037 4388
rect 13803 3968 13845 3977
rect 13803 3928 13804 3968
rect 13844 3928 13845 3968
rect 13803 3919 13845 3928
rect 13804 3557 13844 3919
rect 13803 3548 13845 3557
rect 13803 3508 13804 3548
rect 13844 3508 13845 3548
rect 13803 3499 13845 3508
rect 13804 3422 13844 3499
rect 13708 2624 13748 2633
rect 13804 2624 13844 3382
rect 13900 2876 13940 4348
rect 13995 4339 14037 4348
rect 14283 4220 14325 4229
rect 14283 4180 14284 4220
rect 14324 4180 14325 4220
rect 14283 4171 14325 4180
rect 14188 4136 14228 4145
rect 13996 4096 14188 4136
rect 13996 3632 14036 4096
rect 14188 4087 14228 4096
rect 14284 4136 14324 4171
rect 14284 4085 14324 4096
rect 13996 3583 14036 3592
rect 14187 3632 14229 3641
rect 14187 3592 14188 3632
rect 14228 3592 14229 3632
rect 14187 3583 14229 3592
rect 14188 3498 14228 3583
rect 14379 3380 14421 3389
rect 14379 3340 14380 3380
rect 14420 3340 14421 3380
rect 14379 3331 14421 3340
rect 14380 3246 14420 3331
rect 14283 3128 14325 3137
rect 14283 3088 14284 3128
rect 14324 3088 14325 3128
rect 14283 3079 14325 3088
rect 13900 2827 13940 2836
rect 14284 2717 14324 3079
rect 14283 2708 14325 2717
rect 14283 2668 14284 2708
rect 14324 2668 14325 2708
rect 14283 2659 14325 2668
rect 14188 2624 14228 2633
rect 13748 2584 13940 2624
rect 13708 2575 13748 2584
rect 13900 1952 13940 2584
rect 14092 2120 14132 2129
rect 14188 2120 14228 2584
rect 14284 2624 14324 2659
rect 14284 2574 14324 2584
rect 14132 2080 14228 2120
rect 14092 2071 14132 2080
rect 13900 1903 13940 1912
rect 13612 1280 13652 1289
rect 13516 1240 13612 1280
rect 13612 1231 13652 1240
rect 13803 1196 13845 1205
rect 13803 1156 13804 1196
rect 13844 1156 13845 1196
rect 13803 1147 13845 1156
rect 13804 1062 13844 1147
rect 13995 1112 14037 1121
rect 13995 1072 13996 1112
rect 14036 1072 14037 1112
rect 13995 1063 14037 1072
rect 13996 978 14036 1063
rect 14476 80 14516 5431
rect 14764 4976 14804 4985
rect 14764 4397 14804 4936
rect 14860 4976 14900 4985
rect 14860 4817 14900 4936
rect 14859 4808 14901 4817
rect 14859 4768 14860 4808
rect 14900 4768 14901 4808
rect 14859 4759 14901 4768
rect 14763 4388 14805 4397
rect 14763 4348 14764 4388
rect 14804 4348 14805 4388
rect 14763 4339 14805 4348
rect 14667 4304 14709 4313
rect 14667 4264 14668 4304
rect 14708 4264 14709 4304
rect 14667 4255 14709 4264
rect 14668 4220 14708 4255
rect 14668 4169 14708 4180
rect 14764 4220 14804 4229
rect 14860 4220 14900 4759
rect 14804 4180 14900 4220
rect 14764 4171 14804 4180
rect 14956 4052 14996 7288
rect 15051 7244 15093 7253
rect 15051 7204 15052 7244
rect 15092 7204 15093 7244
rect 15051 7195 15093 7204
rect 15052 7076 15092 7195
rect 15052 7027 15092 7036
rect 15148 6665 15188 8623
rect 15243 8336 15285 8345
rect 15243 8296 15244 8336
rect 15284 8296 15285 8336
rect 15243 8287 15285 8296
rect 15147 6656 15189 6665
rect 15147 6616 15148 6656
rect 15188 6616 15189 6656
rect 15147 6607 15189 6616
rect 15244 6474 15284 8287
rect 15340 7085 15380 9379
rect 15436 8849 15476 10672
rect 15628 9428 15668 10672
rect 15820 10529 15860 10672
rect 15819 10520 15861 10529
rect 15819 10480 15820 10520
rect 15860 10480 15861 10520
rect 15819 10471 15861 10480
rect 15915 10100 15957 10109
rect 15915 10060 15916 10100
rect 15956 10060 15957 10100
rect 15915 10051 15957 10060
rect 15532 9388 15668 9428
rect 15435 8840 15477 8849
rect 15435 8800 15436 8840
rect 15476 8800 15477 8840
rect 15435 8791 15477 8800
rect 15532 8177 15572 9388
rect 15819 8840 15861 8849
rect 15819 8800 15820 8840
rect 15860 8800 15861 8840
rect 15819 8791 15861 8800
rect 15628 8672 15668 8681
rect 15531 8168 15573 8177
rect 15531 8128 15532 8168
rect 15572 8128 15573 8168
rect 15531 8119 15573 8128
rect 15628 8093 15668 8632
rect 15724 8672 15764 8683
rect 15724 8597 15764 8632
rect 15723 8588 15765 8597
rect 15723 8548 15724 8588
rect 15764 8548 15765 8588
rect 15723 8539 15765 8548
rect 15627 8084 15669 8093
rect 15627 8044 15628 8084
rect 15668 8044 15669 8084
rect 15627 8035 15669 8044
rect 15435 8000 15477 8009
rect 15435 7960 15436 8000
rect 15476 7960 15477 8000
rect 15435 7951 15477 7960
rect 15436 7866 15476 7951
rect 15723 7496 15765 7505
rect 15723 7456 15724 7496
rect 15764 7456 15765 7496
rect 15723 7447 15765 7456
rect 15724 7412 15764 7447
rect 15724 7361 15764 7372
rect 15531 7244 15573 7253
rect 15531 7204 15532 7244
rect 15572 7204 15573 7244
rect 15531 7195 15573 7204
rect 15532 7110 15572 7195
rect 15339 7076 15381 7085
rect 15339 7036 15340 7076
rect 15380 7036 15381 7076
rect 15339 7027 15381 7036
rect 15531 6992 15573 7001
rect 15531 6952 15532 6992
rect 15572 6952 15573 6992
rect 15531 6943 15573 6952
rect 15339 6656 15381 6665
rect 15339 6616 15340 6656
rect 15380 6616 15381 6656
rect 15339 6607 15381 6616
rect 15148 6434 15284 6474
rect 15148 5069 15188 6434
rect 15243 6320 15285 6329
rect 15243 6280 15244 6320
rect 15284 6280 15285 6320
rect 15243 6271 15285 6280
rect 15244 5648 15284 6271
rect 15244 5599 15284 5608
rect 15147 5060 15189 5069
rect 15147 5020 15148 5060
rect 15188 5020 15189 5060
rect 15147 5011 15189 5020
rect 14668 4012 14996 4052
rect 14668 3221 14708 4012
rect 15148 3968 15188 5011
rect 15340 4976 15380 6607
rect 15532 6488 15572 6943
rect 15820 6740 15860 8791
rect 15916 7328 15956 10051
rect 16012 7412 16052 10672
rect 16204 7496 16244 10672
rect 16396 9689 16436 10672
rect 16491 9848 16533 9857
rect 16491 9808 16492 9848
rect 16532 9808 16533 9848
rect 16491 9799 16533 9808
rect 16395 9680 16437 9689
rect 16395 9640 16396 9680
rect 16436 9640 16437 9680
rect 16395 9631 16437 9640
rect 16299 9596 16341 9605
rect 16299 9556 16300 9596
rect 16340 9556 16341 9596
rect 16299 9547 16341 9556
rect 16300 9353 16340 9547
rect 16396 9512 16436 9521
rect 16492 9512 16532 9799
rect 16588 9521 16628 10672
rect 16780 9680 16820 10672
rect 16875 10352 16917 10361
rect 16875 10312 16876 10352
rect 16916 10312 16917 10352
rect 16875 10303 16917 10312
rect 16684 9640 16820 9680
rect 16436 9472 16532 9512
rect 16587 9512 16629 9521
rect 16587 9472 16588 9512
rect 16628 9472 16629 9512
rect 16396 9463 16436 9472
rect 16587 9463 16629 9472
rect 16299 9344 16341 9353
rect 16299 9304 16300 9344
rect 16340 9304 16341 9344
rect 16299 9295 16341 9304
rect 16300 8000 16340 9295
rect 16588 9260 16628 9269
rect 16396 9220 16588 9260
rect 16396 8672 16436 9220
rect 16588 9211 16628 9220
rect 16491 9092 16533 9101
rect 16491 9052 16492 9092
rect 16532 9052 16533 9092
rect 16491 9043 16533 9052
rect 16396 8623 16436 8632
rect 16492 8672 16532 9043
rect 16300 7951 16340 7960
rect 16204 7456 16340 7496
rect 16012 7372 16244 7412
rect 15916 7288 16148 7328
rect 15916 7160 15956 7169
rect 15916 6749 15956 7120
rect 15532 6439 15572 6448
rect 15628 6700 15860 6740
rect 15915 6740 15957 6749
rect 15915 6700 15916 6740
rect 15956 6700 15957 6740
rect 15628 5564 15668 6700
rect 15915 6691 15957 6700
rect 15724 6572 15764 6581
rect 15764 6532 16052 6572
rect 15724 6523 15764 6532
rect 16012 6488 16052 6532
rect 16012 6439 16052 6448
rect 16108 6488 16148 7288
rect 16108 5984 16148 6448
rect 16012 5944 16148 5984
rect 15628 5524 15956 5564
rect 15436 5480 15476 5489
rect 15476 5440 15764 5480
rect 15436 5431 15476 5440
rect 15627 5312 15669 5321
rect 15627 5272 15628 5312
rect 15668 5272 15669 5312
rect 15627 5263 15669 5272
rect 15243 4892 15285 4901
rect 15243 4852 15244 4892
rect 15284 4852 15285 4892
rect 15243 4843 15285 4852
rect 15244 4758 15284 4843
rect 15244 4136 15284 4145
rect 15340 4136 15380 4936
rect 15284 4096 15380 4136
rect 15244 4087 15284 4096
rect 15148 3928 15284 3968
rect 15147 3548 15189 3557
rect 15147 3508 15148 3548
rect 15188 3508 15189 3548
rect 15147 3499 15189 3508
rect 14763 3464 14805 3473
rect 14763 3424 14764 3464
rect 14804 3424 14805 3464
rect 14763 3415 14805 3424
rect 14764 3330 14804 3415
rect 14667 3212 14709 3221
rect 14667 3172 14668 3212
rect 14708 3172 14709 3212
rect 14667 3163 14709 3172
rect 14668 2708 14708 3163
rect 14763 2960 14805 2969
rect 14763 2920 14764 2960
rect 14804 2920 14805 2960
rect 14763 2911 14805 2920
rect 14668 2659 14708 2668
rect 14764 2708 14804 2911
rect 14764 2659 14804 2668
rect 14572 1952 14612 1963
rect 14572 1877 14612 1912
rect 14571 1868 14613 1877
rect 14571 1828 14572 1868
rect 14612 1828 14613 1868
rect 14571 1819 14613 1828
rect 14572 1541 14612 1819
rect 14571 1532 14613 1541
rect 14571 1492 14572 1532
rect 14612 1492 14613 1532
rect 14571 1483 14613 1492
rect 15148 1112 15188 3499
rect 15244 2624 15284 3928
rect 15531 3800 15573 3809
rect 15531 3760 15532 3800
rect 15572 3760 15573 3800
rect 15531 3751 15573 3760
rect 15532 3305 15572 3751
rect 15531 3296 15573 3305
rect 15531 3256 15532 3296
rect 15572 3256 15573 3296
rect 15531 3247 15573 3256
rect 15628 3212 15668 5263
rect 15724 4150 15764 5440
rect 15819 5060 15861 5069
rect 15819 5020 15820 5060
rect 15860 5020 15861 5060
rect 15819 5011 15861 5020
rect 15820 4976 15860 5011
rect 15820 4925 15860 4936
rect 15916 4220 15956 5524
rect 15724 4101 15764 4110
rect 15820 4180 15956 4220
rect 15820 3296 15860 4180
rect 15915 3968 15957 3977
rect 15915 3928 15916 3968
rect 15956 3928 15957 3968
rect 15915 3919 15957 3928
rect 15916 3834 15956 3919
rect 16012 3809 16052 5944
rect 16108 5480 16148 5489
rect 16204 5480 16244 7372
rect 16300 6320 16340 7456
rect 16492 6488 16532 8632
rect 16300 6280 16436 6320
rect 16148 5440 16244 5480
rect 16300 5732 16340 5741
rect 16108 5431 16148 5440
rect 16300 5060 16340 5692
rect 16396 5228 16436 6280
rect 16492 5825 16532 6448
rect 16587 6404 16629 6413
rect 16587 6364 16588 6404
rect 16628 6364 16629 6404
rect 16587 6355 16629 6364
rect 16588 6270 16628 6355
rect 16491 5816 16533 5825
rect 16491 5776 16492 5816
rect 16532 5776 16533 5816
rect 16491 5767 16533 5776
rect 16491 5648 16533 5657
rect 16491 5608 16492 5648
rect 16532 5608 16533 5648
rect 16491 5599 16533 5608
rect 16492 5405 16532 5599
rect 16491 5396 16533 5405
rect 16491 5356 16492 5396
rect 16532 5356 16533 5396
rect 16491 5347 16533 5356
rect 16396 5188 16628 5228
rect 16492 5060 16532 5069
rect 16300 5020 16492 5060
rect 16492 5011 16532 5020
rect 16300 4962 16340 4971
rect 16300 4388 16340 4922
rect 16588 4892 16628 5188
rect 16204 4348 16340 4388
rect 16396 4852 16628 4892
rect 16011 3800 16053 3809
rect 16011 3760 16012 3800
rect 16052 3760 16053 3800
rect 16011 3751 16053 3760
rect 16204 3632 16244 4348
rect 16300 4220 16340 4229
rect 16300 3977 16340 4180
rect 16299 3968 16341 3977
rect 16299 3928 16300 3968
rect 16340 3928 16341 3968
rect 16299 3919 16341 3928
rect 16204 3583 16244 3592
rect 16396 3632 16436 4852
rect 16684 4397 16724 9640
rect 16780 9512 16820 9523
rect 16780 9437 16820 9472
rect 16779 9428 16821 9437
rect 16779 9388 16780 9428
rect 16820 9388 16821 9428
rect 16779 9379 16821 9388
rect 16779 9092 16821 9101
rect 16876 9092 16916 10303
rect 16972 9101 17012 10672
rect 17067 9680 17109 9689
rect 17067 9640 17068 9680
rect 17108 9640 17109 9680
rect 17067 9631 17109 9640
rect 16779 9052 16780 9092
rect 16820 9052 16916 9092
rect 16971 9092 17013 9101
rect 16971 9052 16972 9092
rect 17012 9052 17013 9092
rect 16779 9043 16821 9052
rect 16971 9043 17013 9052
rect 16875 8672 16917 8681
rect 16875 8632 16876 8672
rect 16916 8632 16917 8672
rect 16875 8623 16917 8632
rect 16972 8672 17012 8681
rect 16876 8538 16916 8623
rect 16972 8513 17012 8632
rect 16971 8504 17013 8513
rect 16971 8464 16972 8504
rect 17012 8464 17013 8504
rect 16971 8455 17013 8464
rect 16779 6740 16821 6749
rect 16779 6700 16780 6740
rect 16820 6700 16821 6740
rect 16779 6691 16821 6700
rect 16780 6077 16820 6691
rect 17068 6656 17108 9631
rect 17164 8849 17204 10672
rect 17259 9848 17301 9857
rect 17259 9808 17260 9848
rect 17300 9808 17301 9848
rect 17259 9799 17301 9808
rect 17163 8840 17205 8849
rect 17163 8800 17164 8840
rect 17204 8800 17205 8840
rect 17163 8791 17205 8800
rect 17163 8000 17205 8009
rect 17163 7960 17164 8000
rect 17204 7960 17205 8000
rect 17163 7951 17205 7960
rect 17164 7160 17204 7951
rect 17164 7001 17204 7120
rect 17163 6992 17205 7001
rect 17163 6952 17164 6992
rect 17204 6952 17205 6992
rect 17163 6943 17205 6952
rect 17068 6616 17204 6656
rect 17067 6488 17109 6497
rect 17067 6448 17068 6488
rect 17108 6448 17109 6488
rect 17067 6439 17109 6448
rect 17068 6354 17108 6439
rect 16779 6068 16821 6077
rect 16779 6028 16780 6068
rect 16820 6028 16821 6068
rect 16779 6019 16821 6028
rect 17067 5816 17109 5825
rect 17067 5776 17068 5816
rect 17108 5776 17109 5816
rect 17067 5767 17109 5776
rect 16780 5069 16820 5154
rect 16779 5060 16821 5069
rect 16779 5020 16780 5060
rect 16820 5020 16821 5060
rect 16779 5011 16821 5020
rect 16972 4962 17012 4971
rect 16972 4733 17012 4922
rect 17068 4817 17108 5767
rect 17067 4808 17109 4817
rect 17067 4768 17068 4808
rect 17108 4768 17109 4808
rect 17067 4759 17109 4768
rect 16779 4724 16821 4733
rect 16779 4684 16780 4724
rect 16820 4684 16821 4724
rect 16779 4675 16821 4684
rect 16971 4724 17013 4733
rect 16971 4684 16972 4724
rect 17012 4684 17013 4724
rect 16971 4675 17013 4684
rect 16491 4388 16533 4397
rect 16491 4348 16492 4388
rect 16532 4348 16533 4388
rect 16491 4339 16533 4348
rect 16683 4388 16725 4397
rect 16683 4348 16684 4388
rect 16724 4348 16725 4388
rect 16683 4339 16725 4348
rect 16492 4254 16532 4339
rect 16396 3583 16436 3592
rect 16780 3632 16820 4675
rect 17164 4640 17204 6616
rect 17260 6329 17300 9799
rect 17356 9521 17396 10672
rect 17355 9512 17397 9521
rect 17355 9472 17356 9512
rect 17396 9472 17397 9512
rect 17355 9463 17397 9472
rect 17452 8672 17492 8683
rect 17452 8597 17492 8632
rect 17451 8588 17493 8597
rect 17451 8548 17452 8588
rect 17492 8548 17493 8588
rect 17451 8539 17493 8548
rect 17548 8420 17588 10672
rect 17643 9680 17685 9689
rect 17643 9640 17644 9680
rect 17684 9640 17685 9680
rect 17643 9631 17685 9640
rect 17644 9437 17684 9631
rect 17643 9428 17685 9437
rect 17643 9388 17644 9428
rect 17684 9388 17685 9428
rect 17643 9379 17685 9388
rect 17452 8380 17588 8420
rect 17452 7505 17492 8380
rect 17547 8000 17589 8009
rect 17547 7960 17548 8000
rect 17588 7960 17589 8000
rect 17644 8000 17684 9379
rect 17740 8933 17780 10672
rect 17932 9605 17972 10672
rect 18124 10529 18164 10672
rect 18123 10520 18165 10529
rect 18123 10480 18124 10520
rect 18164 10480 18165 10520
rect 18123 10471 18165 10480
rect 18027 9848 18069 9857
rect 18027 9808 18028 9848
rect 18068 9808 18069 9848
rect 18027 9799 18069 9808
rect 17931 9596 17973 9605
rect 17931 9556 17932 9596
rect 17972 9556 17973 9596
rect 17931 9547 17973 9556
rect 18028 9512 18068 9799
rect 18316 9596 18356 10672
rect 18508 9857 18548 10672
rect 18507 9848 18549 9857
rect 18507 9808 18508 9848
rect 18548 9808 18549 9848
rect 18507 9799 18549 9808
rect 18700 9680 18740 10672
rect 18796 9680 18836 9689
rect 18700 9640 18796 9680
rect 18796 9631 18836 9640
rect 18316 9556 18740 9596
rect 18028 9463 18068 9472
rect 18604 9428 18644 9437
rect 17835 9260 17877 9269
rect 18220 9260 18260 9269
rect 17835 9220 17836 9260
rect 17876 9220 17877 9260
rect 17835 9211 17877 9220
rect 18028 9220 18220 9260
rect 17739 8924 17781 8933
rect 17739 8884 17740 8924
rect 17780 8884 17781 8924
rect 17739 8875 17781 8884
rect 17836 8429 17876 9211
rect 18028 8840 18068 9220
rect 18220 9211 18260 9220
rect 18604 8924 18644 9388
rect 17932 8800 18068 8840
rect 18124 8884 18644 8924
rect 17932 8686 17972 8800
rect 17932 8637 17972 8646
rect 18124 8588 18164 8884
rect 18412 8672 18452 8681
rect 18124 8539 18164 8548
rect 18220 8632 18412 8672
rect 17835 8420 17877 8429
rect 17835 8380 17836 8420
rect 17876 8380 17877 8420
rect 17835 8371 17877 8380
rect 18220 8252 18260 8632
rect 18412 8623 18452 8632
rect 18508 8672 18548 8681
rect 18315 8504 18357 8513
rect 18315 8464 18316 8504
rect 18356 8464 18357 8504
rect 18315 8455 18357 8464
rect 17740 8212 18260 8252
rect 17740 8168 17780 8212
rect 17740 8119 17780 8128
rect 17932 8000 17972 8009
rect 17644 7960 17932 8000
rect 17547 7951 17589 7960
rect 17932 7951 17972 7960
rect 17548 7866 17588 7951
rect 17835 7580 17877 7589
rect 17835 7540 17836 7580
rect 17876 7540 17877 7580
rect 17835 7531 17877 7540
rect 17451 7496 17493 7505
rect 17451 7456 17452 7496
rect 17492 7456 17493 7496
rect 17451 7447 17493 7456
rect 17739 7412 17781 7421
rect 17739 7372 17740 7412
rect 17780 7372 17781 7412
rect 17739 7363 17781 7372
rect 17643 7160 17685 7169
rect 17643 7120 17644 7160
rect 17684 7120 17685 7160
rect 17643 7111 17685 7120
rect 17644 7001 17684 7111
rect 17356 6992 17396 7001
rect 17643 6992 17685 7001
rect 17396 6952 17588 6992
rect 17356 6943 17396 6952
rect 17355 6824 17397 6833
rect 17355 6784 17356 6824
rect 17396 6784 17397 6824
rect 17355 6775 17397 6784
rect 17259 6320 17301 6329
rect 17259 6280 17260 6320
rect 17300 6280 17301 6320
rect 17259 6271 17301 6280
rect 17356 5144 17396 6775
rect 17451 6488 17493 6497
rect 17451 6448 17452 6488
rect 17492 6448 17493 6488
rect 17451 6439 17493 6448
rect 17548 6483 17588 6952
rect 17643 6952 17644 6992
rect 17684 6952 17685 6992
rect 17643 6943 17685 6952
rect 17740 6656 17780 7363
rect 17836 6833 17876 7531
rect 18316 7169 18356 8455
rect 18411 8420 18453 8429
rect 18411 8380 18412 8420
rect 18452 8380 18453 8420
rect 18411 8371 18453 8380
rect 18124 7160 18164 7169
rect 17932 7120 18124 7160
rect 17835 6824 17877 6833
rect 17835 6784 17836 6824
rect 17876 6784 17877 6824
rect 17835 6775 17877 6784
rect 17740 6607 17780 6616
rect 17068 4600 17204 4640
rect 17260 5104 17396 5144
rect 16971 4472 17013 4481
rect 16971 4432 16972 4472
rect 17012 4432 17013 4472
rect 16971 4423 17013 4432
rect 16972 4229 17012 4423
rect 17068 4388 17108 4600
rect 17260 4388 17300 5104
rect 17355 4976 17397 4985
rect 17355 4936 17356 4976
rect 17396 4936 17397 4976
rect 17355 4927 17397 4936
rect 17452 4976 17492 6439
rect 17548 6434 17588 6443
rect 17547 6320 17589 6329
rect 17547 6280 17548 6320
rect 17588 6280 17589 6320
rect 17547 6271 17589 6280
rect 17548 5069 17588 6271
rect 17739 5900 17781 5909
rect 17739 5860 17740 5900
rect 17780 5860 17781 5900
rect 17739 5851 17781 5860
rect 17740 5648 17780 5851
rect 17644 5608 17740 5648
rect 17547 5060 17589 5069
rect 17547 5020 17548 5060
rect 17588 5020 17589 5060
rect 17547 5011 17589 5020
rect 17452 4927 17492 4936
rect 17068 4339 17108 4348
rect 17164 4348 17300 4388
rect 16971 4220 17013 4229
rect 17164 4220 17204 4348
rect 16971 4180 16972 4220
rect 17012 4180 17013 4220
rect 16971 4171 17013 4180
rect 17068 4180 17204 4220
rect 17260 4220 17300 4229
rect 16780 3583 16820 3592
rect 16011 3548 16053 3557
rect 16011 3508 16012 3548
rect 16052 3508 16053 3548
rect 16011 3499 16053 3508
rect 16012 3464 16052 3499
rect 16012 3413 16052 3424
rect 16971 3464 17013 3473
rect 16971 3424 16972 3464
rect 17012 3424 17013 3464
rect 16971 3415 17013 3424
rect 16588 3380 16628 3389
rect 16628 3340 16820 3380
rect 16588 3331 16628 3340
rect 15820 3256 16340 3296
rect 15628 3172 15860 3212
rect 15244 2575 15284 2584
rect 15724 2629 15764 2638
rect 15339 2288 15381 2297
rect 15339 2248 15340 2288
rect 15380 2248 15381 2288
rect 15339 2239 15381 2248
rect 15244 1112 15284 1121
rect 15148 1072 15244 1112
rect 15244 953 15284 1072
rect 15243 944 15285 953
rect 15243 904 15244 944
rect 15284 904 15285 944
rect 15243 895 15285 904
rect 15340 188 15380 2239
rect 15724 1784 15764 2589
rect 15820 2129 15860 3172
rect 16300 2876 16340 3256
rect 16300 2827 16340 2836
rect 16683 2876 16725 2885
rect 16683 2836 16684 2876
rect 16724 2836 16725 2876
rect 16683 2827 16725 2836
rect 16108 2708 16148 2717
rect 15916 2540 15956 2549
rect 16108 2540 16148 2668
rect 16588 2633 16628 2718
rect 16684 2717 16724 2827
rect 16683 2708 16725 2717
rect 16683 2668 16684 2708
rect 16724 2668 16725 2708
rect 16683 2659 16725 2668
rect 16203 2624 16245 2633
rect 16203 2584 16204 2624
rect 16244 2584 16245 2624
rect 16203 2575 16245 2584
rect 16587 2624 16629 2633
rect 16587 2584 16588 2624
rect 16628 2584 16629 2624
rect 16587 2575 16629 2584
rect 16684 2624 16724 2659
rect 15956 2500 16148 2540
rect 15916 2491 15956 2500
rect 15819 2120 15861 2129
rect 15819 2080 15820 2120
rect 15860 2080 15861 2120
rect 15819 2071 15861 2080
rect 16012 2120 16052 2129
rect 16204 2120 16244 2575
rect 16684 2574 16724 2584
rect 16299 2540 16341 2549
rect 16299 2500 16300 2540
rect 16340 2500 16341 2540
rect 16299 2491 16341 2500
rect 16052 2080 16244 2120
rect 16012 2071 16052 2080
rect 16300 2036 16340 2491
rect 16780 2045 16820 3340
rect 16204 1996 16340 2036
rect 16779 2036 16821 2045
rect 16779 1996 16780 2036
rect 16820 1996 16821 2036
rect 15436 1744 15764 1784
rect 15820 1952 15860 1961
rect 15436 1280 15476 1744
rect 15436 1231 15476 1240
rect 15820 1205 15860 1912
rect 15915 1952 15957 1961
rect 15915 1912 15916 1952
rect 15956 1912 15957 1952
rect 15915 1903 15957 1912
rect 16204 1952 16244 1996
rect 16779 1987 16821 1996
rect 15916 1541 15956 1903
rect 16204 1877 16244 1912
rect 16203 1868 16245 1877
rect 16203 1828 16204 1868
rect 16244 1828 16245 1868
rect 16203 1819 16245 1828
rect 16204 1788 16244 1819
rect 15915 1532 15957 1541
rect 15915 1492 15916 1532
rect 15956 1492 15957 1532
rect 15915 1483 15957 1492
rect 15819 1196 15861 1205
rect 15819 1156 15820 1196
rect 15860 1156 15861 1196
rect 15819 1147 15861 1156
rect 15820 785 15860 1147
rect 15916 1112 15956 1483
rect 16779 1280 16821 1289
rect 16779 1240 16780 1280
rect 16820 1240 16821 1280
rect 16779 1231 16821 1240
rect 15916 1063 15956 1072
rect 15819 776 15861 785
rect 15819 736 15820 776
rect 15860 736 15861 776
rect 15819 727 15861 736
rect 15340 148 15668 188
rect 15628 80 15668 148
rect 16780 80 16820 1231
rect 16972 1112 17012 3415
rect 17068 2708 17108 4180
rect 17260 3977 17300 4180
rect 17259 3968 17301 3977
rect 17259 3928 17260 3968
rect 17300 3928 17301 3968
rect 17259 3919 17301 3928
rect 17163 2876 17205 2885
rect 17163 2836 17164 2876
rect 17204 2836 17205 2876
rect 17163 2827 17205 2836
rect 17068 2659 17108 2668
rect 17164 2708 17204 2827
rect 17164 2659 17204 2668
rect 17356 1280 17396 4927
rect 17548 4901 17588 5011
rect 17547 4892 17589 4901
rect 17547 4852 17548 4892
rect 17588 4852 17589 4892
rect 17547 4843 17589 4852
rect 17452 4136 17492 4145
rect 17452 2381 17492 4096
rect 17644 3800 17684 5608
rect 17740 5599 17780 5608
rect 17836 5564 17876 6775
rect 17932 5900 17972 7120
rect 18124 7111 18164 7120
rect 18220 7160 18260 7169
rect 18315 7160 18357 7169
rect 18260 7120 18316 7160
rect 18356 7120 18357 7160
rect 18220 7111 18260 7120
rect 18315 7111 18357 7120
rect 18316 7026 18356 7111
rect 18123 6068 18165 6077
rect 18123 6028 18124 6068
rect 18164 6028 18165 6068
rect 18123 6019 18165 6028
rect 17932 5851 17972 5860
rect 18124 5648 18164 6019
rect 18412 5993 18452 8371
rect 18508 7673 18548 8632
rect 18700 8261 18740 9556
rect 18892 9269 18932 10672
rect 18891 9260 18933 9269
rect 18891 9220 18892 9260
rect 18932 9220 18933 9260
rect 19084 9260 19124 10672
rect 19276 9437 19316 10672
rect 19371 10436 19413 10445
rect 19371 10396 19372 10436
rect 19412 10396 19413 10436
rect 19371 10387 19413 10396
rect 19275 9428 19317 9437
rect 19275 9388 19276 9428
rect 19316 9388 19317 9428
rect 19275 9379 19317 9388
rect 19084 9220 19316 9260
rect 18891 9211 18933 9220
rect 18808 9092 19176 9101
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 18808 9043 19176 9052
rect 18891 8840 18933 8849
rect 18891 8800 18892 8840
rect 18932 8800 18933 8840
rect 18891 8791 18933 8800
rect 18892 8756 18932 8791
rect 18699 8252 18741 8261
rect 18699 8212 18700 8252
rect 18740 8212 18741 8252
rect 18699 8203 18741 8212
rect 18892 7748 18932 8716
rect 18988 8672 19028 8681
rect 18988 8513 19028 8632
rect 18987 8504 19029 8513
rect 18987 8464 18988 8504
rect 19028 8464 19029 8504
rect 18987 8455 19029 8464
rect 19179 8000 19221 8009
rect 19179 7960 19180 8000
rect 19220 7960 19221 8000
rect 19179 7951 19221 7960
rect 19180 7757 19220 7951
rect 18700 7708 18932 7748
rect 19179 7748 19221 7757
rect 19179 7708 19180 7748
rect 19220 7708 19221 7748
rect 18507 7664 18549 7673
rect 18507 7624 18508 7664
rect 18548 7624 18549 7664
rect 18507 7615 18549 7624
rect 18700 7580 18740 7708
rect 19179 7699 19221 7708
rect 18604 7540 18740 7580
rect 18808 7580 19176 7589
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 18604 7253 18644 7540
rect 18808 7531 19176 7540
rect 19179 7412 19221 7421
rect 19179 7372 19180 7412
rect 19220 7372 19221 7412
rect 19179 7363 19221 7372
rect 18603 7244 18645 7253
rect 18603 7204 18604 7244
rect 18644 7204 18645 7244
rect 18603 7195 18645 7204
rect 18604 7110 18644 7195
rect 18700 7160 18740 7169
rect 18700 6992 18740 7120
rect 18604 6952 18740 6992
rect 19180 7160 19220 7363
rect 18604 6665 18644 6952
rect 19180 6833 19220 7120
rect 19179 6824 19221 6833
rect 19179 6784 19180 6824
rect 19220 6784 19221 6824
rect 19179 6775 19221 6784
rect 18603 6656 18645 6665
rect 18603 6616 18604 6656
rect 18644 6616 18645 6656
rect 18603 6607 18645 6616
rect 18604 6245 18644 6607
rect 18892 6488 18932 6497
rect 18603 6236 18645 6245
rect 18892 6236 18932 6448
rect 18988 6488 19028 6499
rect 18988 6413 19028 6448
rect 18987 6404 19029 6413
rect 18987 6364 18988 6404
rect 19028 6364 19029 6404
rect 18987 6355 19029 6364
rect 18603 6196 18604 6236
rect 18644 6196 18645 6236
rect 18603 6187 18645 6196
rect 18700 6196 18932 6236
rect 18411 5984 18453 5993
rect 18411 5944 18412 5984
rect 18452 5944 18453 5984
rect 18411 5935 18453 5944
rect 18124 5573 18164 5608
rect 18123 5564 18165 5573
rect 17836 5524 18068 5564
rect 18028 5228 18068 5524
rect 18123 5524 18124 5564
rect 18164 5524 18165 5564
rect 18123 5515 18165 5524
rect 17932 5188 18068 5228
rect 17932 5144 17972 5188
rect 17548 3760 17684 3800
rect 17740 5104 17972 5144
rect 17548 3473 17588 3760
rect 17547 3464 17589 3473
rect 17547 3424 17548 3464
rect 17588 3424 17589 3464
rect 17547 3415 17589 3424
rect 17644 2624 17684 2633
rect 17740 2624 17780 5104
rect 18027 5060 18069 5069
rect 17932 5020 18028 5060
rect 18068 5020 18069 5060
rect 17932 4976 17972 5020
rect 18027 5011 18069 5020
rect 17932 4927 17972 4936
rect 18412 4976 18452 4985
rect 17835 4892 17877 4901
rect 17835 4852 17836 4892
rect 17876 4852 17877 4892
rect 17835 4843 17877 4852
rect 18028 4892 18068 4903
rect 17684 2584 17780 2624
rect 17644 2575 17684 2584
rect 17836 2465 17876 4843
rect 18028 4817 18068 4852
rect 18315 4892 18357 4901
rect 18315 4852 18316 4892
rect 18356 4852 18357 4892
rect 18315 4843 18357 4852
rect 18027 4808 18069 4817
rect 18027 4768 18028 4808
rect 18068 4768 18069 4808
rect 18027 4759 18069 4768
rect 18219 3464 18261 3473
rect 18219 3424 18220 3464
rect 18260 3424 18261 3464
rect 18219 3415 18261 3424
rect 18220 3330 18260 3415
rect 18124 2629 18164 2638
rect 17835 2456 17877 2465
rect 17835 2416 17836 2456
rect 17876 2416 17877 2456
rect 17835 2407 17877 2416
rect 17451 2372 17493 2381
rect 17451 2332 17452 2372
rect 17492 2332 17493 2372
rect 17451 2323 17493 2332
rect 17644 2120 17684 2129
rect 18124 2120 18164 2589
rect 18316 2540 18356 4843
rect 18412 4145 18452 4936
rect 18507 4976 18549 4985
rect 18507 4936 18508 4976
rect 18548 4936 18549 4976
rect 18507 4927 18549 4936
rect 18508 4842 18548 4927
rect 18700 4388 18740 6196
rect 18808 6068 19176 6077
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 18808 6019 19176 6028
rect 19179 5732 19221 5741
rect 19179 5692 19180 5732
rect 19220 5692 19221 5732
rect 19179 5683 19221 5692
rect 19180 5405 19220 5683
rect 19179 5396 19221 5405
rect 19179 5356 19180 5396
rect 19220 5356 19221 5396
rect 19179 5347 19221 5356
rect 19180 4985 19220 5070
rect 19179 4976 19221 4985
rect 19179 4936 19180 4976
rect 19220 4936 19221 4976
rect 19179 4927 19221 4936
rect 18795 4892 18837 4901
rect 18795 4852 18796 4892
rect 18836 4852 18837 4892
rect 18795 4843 18837 4852
rect 18796 4758 18836 4843
rect 18988 4808 19028 4817
rect 19276 4808 19316 9220
rect 19372 8849 19412 10387
rect 19468 9689 19508 10672
rect 19467 9680 19509 9689
rect 19467 9640 19468 9680
rect 19508 9640 19509 9680
rect 19467 9631 19509 9640
rect 19467 9512 19509 9521
rect 19467 9472 19468 9512
rect 19508 9472 19509 9512
rect 19467 9463 19509 9472
rect 19468 9378 19508 9463
rect 19660 8849 19700 10672
rect 19371 8840 19413 8849
rect 19371 8800 19372 8840
rect 19412 8800 19413 8840
rect 19371 8791 19413 8800
rect 19659 8840 19701 8849
rect 19659 8800 19660 8840
rect 19700 8800 19701 8840
rect 19659 8791 19701 8800
rect 19468 8672 19508 8681
rect 19371 8336 19413 8345
rect 19371 8296 19372 8336
rect 19412 8296 19413 8336
rect 19371 8287 19413 8296
rect 19372 8168 19412 8287
rect 19372 8119 19412 8128
rect 19371 7916 19413 7925
rect 19371 7876 19372 7916
rect 19412 7876 19413 7916
rect 19371 7867 19413 7876
rect 19372 7169 19412 7867
rect 19468 7841 19508 8632
rect 19852 8252 19892 10672
rect 20044 10025 20084 10672
rect 20235 10648 20236 10672
rect 20276 10672 20296 10688
rect 20408 10672 20488 10752
rect 20600 10672 20680 10752
rect 20792 10672 20872 10752
rect 20984 10672 21064 10752
rect 21176 10672 21256 10752
rect 21368 10672 21448 10752
rect 21560 10672 21640 10752
rect 21752 10672 21832 10752
rect 21944 10672 22024 10752
rect 22136 10672 22216 10752
rect 22328 10672 22408 10752
rect 22520 10672 22600 10752
rect 22712 10672 22792 10752
rect 22904 10672 22984 10752
rect 23096 10672 23176 10752
rect 23288 10672 23368 10752
rect 23480 10672 23560 10752
rect 23672 10672 23752 10752
rect 23864 10672 23944 10752
rect 24056 10672 24136 10752
rect 24248 10672 24328 10752
rect 24440 10672 24520 10752
rect 24632 10672 24712 10752
rect 24824 10672 24904 10752
rect 25016 10672 25096 10752
rect 25208 10672 25288 10752
rect 25400 10688 25480 10752
rect 25400 10672 25420 10688
rect 20276 10648 20277 10672
rect 20235 10639 20277 10648
rect 20236 10025 20276 10639
rect 20043 10016 20085 10025
rect 20043 9976 20044 10016
rect 20084 9976 20085 10016
rect 20043 9967 20085 9976
rect 20235 10016 20277 10025
rect 20235 9976 20236 10016
rect 20276 9976 20277 10016
rect 20428 10016 20468 10672
rect 20620 10109 20660 10672
rect 20619 10100 20661 10109
rect 20619 10060 20620 10100
rect 20660 10060 20661 10100
rect 20619 10051 20661 10060
rect 20428 9976 20564 10016
rect 20235 9967 20277 9976
rect 20048 9848 20416 9857
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20048 9799 20416 9808
rect 20331 9680 20373 9689
rect 20331 9640 20332 9680
rect 20372 9640 20373 9680
rect 20331 9631 20373 9640
rect 20139 8756 20181 8765
rect 20139 8716 20140 8756
rect 20180 8716 20181 8756
rect 20139 8707 20181 8716
rect 19948 8677 19988 8686
rect 19948 8345 19988 8637
rect 20140 8588 20180 8707
rect 20140 8539 20180 8548
rect 20332 8504 20372 9631
rect 20524 9596 20564 9976
rect 20812 9857 20852 10672
rect 20811 9848 20853 9857
rect 20811 9808 20812 9848
rect 20852 9808 20853 9848
rect 20811 9799 20853 9808
rect 20428 9556 20564 9596
rect 20428 8513 20468 9556
rect 20716 9521 20756 9606
rect 21004 9596 21044 10672
rect 21196 9689 21236 10672
rect 21291 9932 21333 9941
rect 21291 9892 21292 9932
rect 21332 9892 21333 9932
rect 21291 9883 21333 9892
rect 21195 9680 21237 9689
rect 21195 9640 21196 9680
rect 21236 9640 21237 9680
rect 21195 9631 21237 9640
rect 20812 9556 21044 9596
rect 20715 9512 20757 9521
rect 20524 9472 20716 9512
rect 20756 9472 20757 9512
rect 20332 8455 20372 8464
rect 20427 8504 20469 8513
rect 20427 8464 20428 8504
rect 20468 8464 20469 8504
rect 20427 8455 20469 8464
rect 19947 8336 19989 8345
rect 19947 8296 19948 8336
rect 19988 8296 19989 8336
rect 19947 8287 19989 8296
rect 20048 8336 20416 8345
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20048 8287 20416 8296
rect 19756 8212 19892 8252
rect 19756 8093 19796 8212
rect 19755 8084 19797 8093
rect 19755 8044 19756 8084
rect 19796 8044 19797 8084
rect 19755 8035 19797 8044
rect 19563 8000 19605 8009
rect 19563 7960 19564 8000
rect 19604 7960 19605 8000
rect 19563 7951 19605 7960
rect 19564 7866 19604 7951
rect 19467 7832 19509 7841
rect 19467 7792 19468 7832
rect 19508 7792 19509 7832
rect 19467 7783 19509 7792
rect 19563 7580 19605 7589
rect 19563 7540 19564 7580
rect 19604 7540 19605 7580
rect 19563 7531 19605 7540
rect 19467 7244 19509 7253
rect 19467 7204 19468 7244
rect 19508 7204 19509 7244
rect 19467 7195 19509 7204
rect 19371 7160 19413 7169
rect 19371 7120 19372 7160
rect 19412 7120 19413 7160
rect 19371 7111 19413 7120
rect 19372 6488 19412 7111
rect 19372 6439 19412 6448
rect 19468 6488 19508 7195
rect 19468 6439 19508 6448
rect 19564 6413 19604 7531
rect 19660 7165 19700 7174
rect 19563 6404 19605 6413
rect 19563 6364 19564 6404
rect 19604 6364 19605 6404
rect 19563 6355 19605 6364
rect 19467 5984 19509 5993
rect 19467 5944 19468 5984
rect 19508 5944 19509 5984
rect 19467 5935 19509 5944
rect 19371 5900 19413 5909
rect 19371 5860 19372 5900
rect 19412 5860 19413 5900
rect 19371 5851 19413 5860
rect 19372 5648 19412 5851
rect 19372 5599 19412 5608
rect 19028 4768 19316 4808
rect 18988 4759 19028 4768
rect 19468 4724 19508 5935
rect 19564 5900 19604 5909
rect 19660 5900 19700 7125
rect 19756 6824 19796 8035
rect 19947 7832 19989 7841
rect 19947 7792 19948 7832
rect 19988 7792 19989 7832
rect 19947 7783 19989 7792
rect 19851 7076 19893 7085
rect 19851 7036 19852 7076
rect 19892 7036 19893 7076
rect 19851 7027 19893 7036
rect 19852 6942 19892 7027
rect 19756 6784 19892 6824
rect 19755 6404 19797 6413
rect 19755 6364 19756 6404
rect 19796 6364 19797 6404
rect 19755 6355 19797 6364
rect 19604 5860 19700 5900
rect 19564 5851 19604 5860
rect 19756 5816 19796 6355
rect 19276 4684 19508 4724
rect 19660 5776 19796 5816
rect 18808 4556 19176 4565
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 18808 4507 19176 4516
rect 18892 4388 18932 4397
rect 19276 4388 19316 4684
rect 19371 4556 19413 4565
rect 19371 4516 19372 4556
rect 19412 4516 19413 4556
rect 19371 4507 19413 4516
rect 18700 4348 18892 4388
rect 18892 4339 18932 4348
rect 19180 4348 19316 4388
rect 18411 4136 18453 4145
rect 18411 4096 18412 4136
rect 18452 4096 18453 4136
rect 18411 4087 18453 4096
rect 18700 4136 18740 4145
rect 18412 3968 18452 4087
rect 18412 3928 18548 3968
rect 18411 3464 18453 3473
rect 18411 3424 18412 3464
rect 18452 3424 18453 3464
rect 18411 3415 18453 3424
rect 18412 3330 18452 3415
rect 18508 3053 18548 3928
rect 18603 3800 18645 3809
rect 18603 3760 18604 3800
rect 18644 3760 18645 3800
rect 18603 3751 18645 3760
rect 18507 3044 18549 3053
rect 18507 3004 18508 3044
rect 18548 3004 18549 3044
rect 18507 2995 18549 3004
rect 18604 2876 18644 3751
rect 18700 3557 18740 4096
rect 19084 4052 19124 4061
rect 19180 4052 19220 4348
rect 19124 4012 19220 4052
rect 19276 4141 19316 4150
rect 19084 4003 19124 4012
rect 18891 3884 18933 3893
rect 19276 3884 19316 4101
rect 18891 3844 18892 3884
rect 18932 3844 18933 3884
rect 18891 3835 18933 3844
rect 19084 3844 19316 3884
rect 18699 3548 18741 3557
rect 18699 3508 18700 3548
rect 18740 3508 18741 3548
rect 18699 3499 18741 3508
rect 18892 3473 18932 3835
rect 19084 3641 19124 3844
rect 19179 3716 19221 3725
rect 19179 3676 19180 3716
rect 19220 3676 19221 3716
rect 19179 3667 19221 3676
rect 19083 3632 19125 3641
rect 19083 3592 19084 3632
rect 19124 3592 19125 3632
rect 19083 3583 19125 3592
rect 18891 3464 18933 3473
rect 18891 3424 18892 3464
rect 18932 3424 18933 3464
rect 18891 3415 18933 3424
rect 19180 3221 19220 3667
rect 19275 3548 19317 3557
rect 19275 3508 19276 3548
rect 19316 3508 19317 3548
rect 19275 3499 19317 3508
rect 19179 3212 19221 3221
rect 19179 3172 19180 3212
rect 19220 3172 19221 3212
rect 19179 3163 19221 3172
rect 18808 3044 19176 3053
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 18808 2995 19176 3004
rect 19276 2876 19316 3499
rect 18604 2836 18836 2876
rect 18316 2491 18356 2500
rect 18700 2624 18740 2633
rect 17684 2080 18164 2120
rect 17644 2071 17684 2080
rect 17356 1231 17396 1240
rect 17452 1952 17492 1961
rect 17452 1205 17492 1912
rect 17835 1952 17877 1961
rect 17835 1912 17836 1952
rect 17876 1912 17877 1952
rect 17835 1903 17877 1912
rect 17836 1818 17876 1903
rect 18700 1373 18740 2584
rect 18796 2624 18836 2836
rect 18796 2575 18836 2584
rect 19084 2836 19316 2876
rect 19084 1952 19124 2836
rect 19372 2792 19412 4507
rect 19660 3893 19700 5776
rect 19756 5648 19796 5657
rect 19756 5573 19796 5608
rect 19755 5564 19797 5573
rect 19755 5524 19756 5564
rect 19796 5524 19797 5564
rect 19755 5515 19797 5524
rect 19756 5237 19796 5515
rect 19755 5228 19797 5237
rect 19755 5188 19756 5228
rect 19796 5188 19797 5228
rect 19755 5179 19797 5188
rect 19852 4229 19892 6784
rect 19948 6488 19988 7783
rect 20048 6824 20416 6833
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20048 6775 20416 6784
rect 19948 6439 19988 6448
rect 20428 6474 20468 6483
rect 20428 5648 20468 6434
rect 20524 5909 20564 9472
rect 20715 9463 20757 9472
rect 20812 9344 20852 9556
rect 21196 9512 21236 9521
rect 20716 9304 20852 9344
rect 21004 9472 21196 9512
rect 20619 8840 20661 8849
rect 20619 8800 20620 8840
rect 20660 8800 20661 8840
rect 20619 8791 20661 8800
rect 20620 6740 20660 8791
rect 20716 7589 20756 9304
rect 20907 9260 20949 9269
rect 20907 9220 20908 9260
rect 20948 9220 20949 9260
rect 20907 9211 20949 9220
rect 20908 9126 20948 9211
rect 20907 8504 20949 8513
rect 20907 8464 20908 8504
rect 20948 8464 20949 8504
rect 20907 8455 20949 8464
rect 20812 8000 20852 8009
rect 20812 7757 20852 7960
rect 20811 7748 20853 7757
rect 20811 7708 20812 7748
rect 20852 7708 20853 7748
rect 20811 7699 20853 7708
rect 20715 7580 20757 7589
rect 20715 7540 20716 7580
rect 20756 7540 20757 7580
rect 20715 7531 20757 7540
rect 20620 6700 20756 6740
rect 20619 6572 20661 6581
rect 20619 6532 20620 6572
rect 20660 6532 20661 6572
rect 20619 6523 20661 6532
rect 20620 6438 20660 6523
rect 20523 5900 20565 5909
rect 20523 5860 20524 5900
rect 20564 5860 20565 5900
rect 20523 5851 20565 5860
rect 20428 5608 20660 5648
rect 20048 5312 20416 5321
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20048 5263 20416 5272
rect 20427 5144 20469 5153
rect 20427 5104 20428 5144
rect 20468 5104 20469 5144
rect 20427 5095 20469 5104
rect 20620 5144 20660 5608
rect 20620 5095 20660 5104
rect 20428 4976 20468 5095
rect 20428 4927 20468 4936
rect 20235 4808 20277 4817
rect 20235 4768 20236 4808
rect 20276 4768 20277 4808
rect 20235 4759 20277 4768
rect 20236 4388 20276 4759
rect 20236 4348 20468 4388
rect 19851 4220 19893 4229
rect 19851 4180 19852 4220
rect 19892 4180 19893 4220
rect 19851 4171 19893 4180
rect 20236 4220 20276 4348
rect 20236 4171 20276 4180
rect 20331 4220 20373 4229
rect 20331 4180 20332 4220
rect 20372 4180 20373 4220
rect 20331 4171 20373 4180
rect 19756 4136 19796 4145
rect 19659 3884 19701 3893
rect 19659 3844 19660 3884
rect 19700 3844 19701 3884
rect 19659 3835 19701 3844
rect 19756 3800 19796 4096
rect 20332 4086 20372 4171
rect 20428 4061 20468 4348
rect 20716 4136 20756 6700
rect 20812 5489 20852 7699
rect 20811 5480 20853 5489
rect 20811 5440 20812 5480
rect 20852 5440 20853 5480
rect 20811 5431 20853 5440
rect 20812 5153 20852 5431
rect 20811 5144 20853 5153
rect 20811 5104 20812 5144
rect 20852 5104 20853 5144
rect 20811 5095 20853 5104
rect 20908 4220 20948 8455
rect 21004 8168 21044 9472
rect 21196 9463 21236 9472
rect 21292 9512 21332 9883
rect 21292 8849 21332 9472
rect 21291 8840 21333 8849
rect 21291 8800 21292 8840
rect 21332 8800 21333 8840
rect 21291 8791 21333 8800
rect 21004 8119 21044 8128
rect 21292 8000 21332 8009
rect 21003 7160 21045 7169
rect 21003 7120 21004 7160
rect 21044 7120 21045 7160
rect 21003 7111 21045 7120
rect 21004 7026 21044 7111
rect 21196 5900 21236 5909
rect 21292 5900 21332 7960
rect 21236 5860 21332 5900
rect 21388 8000 21428 10672
rect 21580 10025 21620 10672
rect 21675 10100 21717 10109
rect 21675 10060 21676 10100
rect 21716 10060 21717 10100
rect 21675 10051 21717 10060
rect 21579 10016 21621 10025
rect 21579 9976 21580 10016
rect 21620 9976 21621 10016
rect 21579 9967 21621 9976
rect 21483 9848 21525 9857
rect 21676 9848 21716 10051
rect 21483 9808 21484 9848
rect 21524 9808 21525 9848
rect 21483 9799 21525 9808
rect 21580 9808 21716 9848
rect 21196 5851 21236 5860
rect 21388 5816 21428 7960
rect 21292 5776 21428 5816
rect 21195 5732 21237 5741
rect 21195 5692 21196 5732
rect 21236 5692 21237 5732
rect 21195 5683 21237 5692
rect 21004 5648 21044 5657
rect 21004 5489 21044 5608
rect 21003 5480 21045 5489
rect 21003 5440 21004 5480
rect 21044 5440 21045 5480
rect 21003 5431 21045 5440
rect 20908 4180 21044 4220
rect 20427 4052 20469 4061
rect 20427 4012 20428 4052
rect 20468 4012 20469 4052
rect 20427 4003 20469 4012
rect 20716 3968 20756 4096
rect 20812 4136 20852 4145
rect 20852 4096 20948 4136
rect 20812 4087 20852 4096
rect 20716 3928 20852 3968
rect 19947 3800 19989 3809
rect 19756 3760 19948 3800
rect 19988 3760 19989 3800
rect 19659 3548 19701 3557
rect 19659 3508 19660 3548
rect 19700 3508 19701 3548
rect 19659 3499 19701 3508
rect 19660 3464 19700 3499
rect 19660 3413 19700 3424
rect 19467 3212 19509 3221
rect 19467 3172 19468 3212
rect 19508 3172 19509 3212
rect 19467 3163 19509 3172
rect 19180 2752 19412 2792
rect 19180 2708 19220 2752
rect 19468 2708 19508 3163
rect 19756 2801 19796 3760
rect 19947 3751 19989 3760
rect 20048 3800 20416 3809
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20048 3751 20416 3760
rect 19851 3632 19893 3641
rect 19851 3592 19852 3632
rect 19892 3592 19893 3632
rect 19851 3583 19893 3592
rect 19852 3498 19892 3583
rect 20043 3464 20085 3473
rect 20043 3424 20044 3464
rect 20084 3424 20085 3464
rect 20043 3415 20085 3424
rect 20044 3330 20084 3415
rect 19755 2792 19797 2801
rect 19755 2752 19756 2792
rect 19796 2752 19797 2792
rect 19755 2743 19797 2752
rect 19180 2659 19220 2668
rect 19276 2668 19508 2708
rect 19276 2624 19316 2668
rect 19276 2575 19316 2584
rect 19756 2624 19796 2743
rect 20284 2633 20324 2642
rect 20324 2593 20564 2633
rect 20284 2584 20324 2593
rect 19756 2575 19796 2584
rect 20427 2540 20469 2549
rect 20427 2500 20428 2540
rect 20468 2500 20469 2540
rect 20427 2491 20469 2500
rect 20428 2414 20468 2491
rect 19275 2372 19317 2381
rect 19275 2332 19276 2372
rect 19316 2332 19317 2372
rect 20428 2365 20468 2374
rect 19275 2323 19317 2332
rect 19276 2120 19316 2323
rect 20048 2288 20416 2297
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20048 2239 20416 2248
rect 19276 2071 19316 2080
rect 19563 1952 19605 1961
rect 19084 1903 19124 1912
rect 19468 1912 19564 1952
rect 19604 1912 19605 1952
rect 18808 1532 19176 1541
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 18808 1483 19176 1492
rect 18699 1364 18741 1373
rect 18699 1324 18700 1364
rect 18740 1324 18741 1364
rect 18699 1315 18741 1324
rect 19083 1364 19125 1373
rect 19083 1324 19084 1364
rect 19124 1324 19125 1364
rect 19083 1315 19125 1324
rect 19084 1280 19124 1315
rect 19084 1229 19124 1240
rect 17451 1196 17493 1205
rect 17451 1156 17452 1196
rect 17492 1156 17493 1196
rect 17451 1147 17493 1156
rect 17931 1196 17973 1205
rect 17931 1156 17932 1196
rect 17972 1156 17973 1196
rect 17931 1147 17973 1156
rect 18891 1196 18933 1205
rect 18891 1156 18892 1196
rect 18932 1156 18933 1196
rect 18891 1147 18933 1156
rect 17164 1112 17204 1121
rect 16972 1072 17164 1112
rect 17164 869 17204 1072
rect 17643 1112 17685 1121
rect 17643 1072 17644 1112
rect 17684 1072 17685 1112
rect 17643 1063 17685 1072
rect 17644 978 17684 1063
rect 17163 860 17205 869
rect 17163 820 17164 860
rect 17204 820 17205 860
rect 17163 811 17205 820
rect 17932 80 17972 1147
rect 18892 1112 18932 1147
rect 18892 1061 18932 1072
rect 19468 1112 19508 1912
rect 19563 1903 19605 1912
rect 19564 1818 19604 1903
rect 20524 1373 20564 2593
rect 20716 2624 20756 2633
rect 20716 2120 20756 2584
rect 20812 2624 20852 3928
rect 20812 2575 20852 2584
rect 20908 2381 20948 4096
rect 21004 3809 21044 4180
rect 21003 3800 21045 3809
rect 21003 3760 21004 3800
rect 21044 3760 21045 3800
rect 21003 3751 21045 3760
rect 21004 2717 21044 3751
rect 21099 3548 21141 3557
rect 21099 3508 21100 3548
rect 21140 3508 21141 3548
rect 21099 3499 21141 3508
rect 21100 3053 21140 3499
rect 21099 3044 21141 3053
rect 21099 3004 21100 3044
rect 21140 3004 21141 3044
rect 21099 2995 21141 3004
rect 21003 2708 21045 2717
rect 21003 2668 21004 2708
rect 21044 2668 21045 2708
rect 21003 2659 21045 2668
rect 20907 2372 20949 2381
rect 20907 2332 20908 2372
rect 20948 2332 20949 2372
rect 20907 2323 20949 2332
rect 21004 2120 21044 2129
rect 20716 2080 21004 2120
rect 21004 2071 21044 2080
rect 20812 1952 20852 1961
rect 21100 1952 21140 2995
rect 21196 2708 21236 5683
rect 21292 4733 21332 5776
rect 21388 5648 21428 5657
rect 21388 5405 21428 5608
rect 21387 5396 21429 5405
rect 21387 5356 21388 5396
rect 21428 5356 21429 5396
rect 21387 5347 21429 5356
rect 21291 4724 21333 4733
rect 21291 4684 21292 4724
rect 21332 4684 21333 4724
rect 21291 4675 21333 4684
rect 21484 4145 21524 9799
rect 21388 4136 21428 4145
rect 21388 3800 21428 4096
rect 21483 4136 21525 4145
rect 21483 4096 21484 4136
rect 21524 4096 21525 4136
rect 21483 4087 21525 4096
rect 21484 4002 21524 4087
rect 21388 3760 21524 3800
rect 21484 3632 21524 3760
rect 21484 3583 21524 3592
rect 21292 3464 21332 3473
rect 21332 3424 21428 3464
rect 21292 3415 21332 3424
rect 21291 3128 21333 3137
rect 21291 3088 21292 3128
rect 21332 3088 21333 3128
rect 21291 3079 21333 3088
rect 21196 2659 21236 2668
rect 21292 2708 21332 3079
rect 21292 2659 21332 2668
rect 21388 2381 21428 3424
rect 21580 3221 21620 9808
rect 21675 9680 21717 9689
rect 21675 9640 21676 9680
rect 21716 9640 21717 9680
rect 21675 9631 21717 9640
rect 21676 9512 21716 9631
rect 21772 9596 21812 10672
rect 21964 10109 22004 10672
rect 21963 10100 22005 10109
rect 21963 10060 21964 10100
rect 22004 10060 22005 10100
rect 21963 10051 22005 10060
rect 22156 9857 22196 10672
rect 22348 10613 22388 10672
rect 22347 10604 22389 10613
rect 22347 10564 22348 10604
rect 22388 10564 22389 10604
rect 22347 10555 22389 10564
rect 22348 9857 22388 10555
rect 22155 9848 22197 9857
rect 22155 9808 22156 9848
rect 22196 9808 22197 9848
rect 22155 9799 22197 9808
rect 22347 9848 22389 9857
rect 22347 9808 22348 9848
rect 22388 9808 22389 9848
rect 22347 9799 22389 9808
rect 22155 9680 22197 9689
rect 22155 9640 22156 9680
rect 22196 9640 22197 9680
rect 22155 9631 22197 9640
rect 21772 9556 22100 9596
rect 21676 9463 21716 9472
rect 21772 9428 21812 9437
rect 21812 9388 21908 9428
rect 21772 9379 21812 9388
rect 21771 9260 21813 9269
rect 21771 9220 21772 9260
rect 21812 9220 21813 9260
rect 21771 9211 21813 9220
rect 21675 9092 21717 9101
rect 21675 9052 21676 9092
rect 21716 9052 21717 9092
rect 21675 9043 21717 9052
rect 21676 7337 21716 9043
rect 21772 8672 21812 9211
rect 21868 8933 21908 9388
rect 21867 8924 21909 8933
rect 21867 8884 21868 8924
rect 21908 8884 21909 8924
rect 21867 8875 21909 8884
rect 21868 8681 21908 8875
rect 21772 8623 21812 8632
rect 21867 8672 21909 8681
rect 21867 8632 21868 8672
rect 21908 8632 21909 8672
rect 21867 8623 21909 8632
rect 21868 8504 21908 8623
rect 21772 8464 21908 8504
rect 21772 8000 21812 8464
rect 21867 8336 21909 8345
rect 21867 8296 21868 8336
rect 21908 8296 21909 8336
rect 21867 8287 21909 8296
rect 21772 7951 21812 7960
rect 21868 8000 21908 8287
rect 22060 8009 22100 9556
rect 22156 8840 22196 9631
rect 22252 9512 22292 9521
rect 22292 9472 22484 9512
rect 22252 9463 22292 9472
rect 22156 8800 22292 8840
rect 22252 8672 22292 8800
rect 22444 8765 22484 9472
rect 22443 8756 22485 8765
rect 22443 8716 22444 8756
rect 22484 8716 22485 8756
rect 22443 8707 22485 8716
rect 22252 8345 22292 8632
rect 22348 8672 22388 8683
rect 22348 8597 22388 8632
rect 22347 8588 22389 8597
rect 22347 8548 22348 8588
rect 22388 8548 22389 8588
rect 22347 8539 22389 8548
rect 22251 8336 22293 8345
rect 22251 8296 22252 8336
rect 22292 8296 22293 8336
rect 22251 8287 22293 8296
rect 21868 7951 21908 7960
rect 22059 8000 22101 8009
rect 22059 7960 22060 8000
rect 22100 7960 22101 8000
rect 22059 7951 22101 7960
rect 22348 8000 22388 8009
rect 22444 8000 22484 8707
rect 22388 7960 22484 8000
rect 22348 7951 22388 7960
rect 22059 7748 22101 7757
rect 22059 7708 22060 7748
rect 22100 7708 22101 7748
rect 22059 7699 22101 7708
rect 21867 7664 21909 7673
rect 21867 7624 21868 7664
rect 21908 7624 21909 7664
rect 21867 7615 21909 7624
rect 21675 7328 21717 7337
rect 21675 7288 21676 7328
rect 21716 7288 21717 7328
rect 21675 7279 21717 7288
rect 21676 4976 21716 4985
rect 21676 4397 21716 4936
rect 21675 4388 21717 4397
rect 21675 4348 21676 4388
rect 21716 4348 21717 4388
rect 21675 4339 21717 4348
rect 21868 4220 21908 7615
rect 21868 4171 21908 4180
rect 21963 4220 22005 4229
rect 21963 4180 21964 4220
rect 22004 4180 22005 4220
rect 21963 4171 22005 4180
rect 21964 4086 22004 4171
rect 21867 3884 21909 3893
rect 21772 3844 21868 3884
rect 21908 3844 21909 3884
rect 21675 3800 21717 3809
rect 21675 3760 21676 3800
rect 21716 3760 21717 3800
rect 21675 3751 21717 3760
rect 21676 3632 21716 3751
rect 21676 3583 21716 3592
rect 21579 3212 21621 3221
rect 21579 3172 21580 3212
rect 21620 3172 21621 3212
rect 21579 3163 21621 3172
rect 21772 2624 21812 3844
rect 21867 3835 21909 3844
rect 21868 3380 21908 3389
rect 21868 2633 21908 3340
rect 21772 2575 21812 2584
rect 21867 2624 21909 2633
rect 21867 2584 21868 2624
rect 21908 2584 21909 2624
rect 21867 2575 21909 2584
rect 22060 2540 22100 7699
rect 22540 7673 22580 10672
rect 22732 9596 22772 10672
rect 22924 9941 22964 10672
rect 22923 9932 22965 9941
rect 22923 9892 22924 9932
rect 22964 9892 22965 9932
rect 22923 9883 22965 9892
rect 22924 9596 22964 9605
rect 22732 9556 22868 9596
rect 22732 9498 22772 9507
rect 22539 7664 22581 7673
rect 22539 7624 22540 7664
rect 22580 7624 22581 7664
rect 22539 7615 22581 7624
rect 22444 7412 22484 7421
rect 22732 7412 22772 9458
rect 22828 8849 22868 9556
rect 22827 8840 22869 8849
rect 22827 8800 22828 8840
rect 22868 8800 22869 8840
rect 22827 8791 22869 8800
rect 22827 8672 22869 8681
rect 22827 8632 22828 8672
rect 22868 8632 22869 8672
rect 22827 8623 22869 8632
rect 22828 8429 22868 8623
rect 22924 8513 22964 9556
rect 23116 9428 23156 10672
rect 23308 9680 23348 10672
rect 23308 9640 23444 9680
rect 23307 9512 23349 9521
rect 23307 9472 23308 9512
rect 23348 9472 23349 9512
rect 23307 9463 23349 9472
rect 23020 9388 23156 9428
rect 22923 8504 22965 8513
rect 22923 8464 22924 8504
rect 22964 8464 22965 8504
rect 22923 8455 22965 8464
rect 22827 8420 22869 8429
rect 22827 8380 22828 8420
rect 22868 8380 22869 8420
rect 22827 8371 22869 8380
rect 23020 8336 23060 9388
rect 23308 9378 23348 9463
rect 23116 9260 23156 9269
rect 23156 9220 23348 9260
rect 23116 9211 23156 9220
rect 23211 8840 23253 8849
rect 23211 8800 23212 8840
rect 23252 8800 23253 8840
rect 23211 8791 23253 8800
rect 23212 8513 23252 8791
rect 23308 8686 23348 9220
rect 23308 8637 23348 8646
rect 23211 8504 23253 8513
rect 23404 8504 23444 9640
rect 23500 8849 23540 10672
rect 23692 10361 23732 10672
rect 23691 10352 23733 10361
rect 23691 10312 23692 10352
rect 23732 10312 23733 10352
rect 23691 10303 23733 10312
rect 23499 8840 23541 8849
rect 23884 8840 23924 10672
rect 23499 8800 23500 8840
rect 23540 8800 23541 8840
rect 23499 8791 23541 8800
rect 23788 8800 23924 8840
rect 23211 8464 23212 8504
rect 23252 8464 23253 8504
rect 23211 8455 23253 8464
rect 23308 8464 23444 8504
rect 23500 8504 23540 8513
rect 22924 8296 23060 8336
rect 22484 7372 22772 7412
rect 22828 7986 22868 7995
rect 22444 7363 22484 7372
rect 22347 7328 22389 7337
rect 22347 7288 22348 7328
rect 22388 7288 22389 7328
rect 22347 7279 22389 7288
rect 22155 7160 22197 7169
rect 22155 7120 22156 7160
rect 22196 7120 22197 7160
rect 22155 7111 22197 7120
rect 22252 7160 22292 7169
rect 22156 6488 22196 7111
rect 22252 6833 22292 7120
rect 22251 6824 22293 6833
rect 22251 6784 22252 6824
rect 22292 6784 22293 6824
rect 22251 6775 22293 6784
rect 22252 6488 22292 6497
rect 22156 6448 22252 6488
rect 22252 6439 22292 6448
rect 22348 4817 22388 7279
rect 22635 7160 22677 7169
rect 22635 7120 22636 7160
rect 22676 7120 22677 7160
rect 22635 7111 22677 7120
rect 22636 7026 22676 7111
rect 22635 6824 22677 6833
rect 22635 6784 22636 6824
rect 22676 6784 22677 6824
rect 22635 6775 22677 6784
rect 22539 5984 22581 5993
rect 22539 5944 22540 5984
rect 22580 5944 22581 5984
rect 22539 5935 22581 5944
rect 22540 5405 22580 5935
rect 22636 5648 22676 6775
rect 22828 5900 22868 7946
rect 22924 7085 22964 8296
rect 23211 8168 23253 8177
rect 23211 8128 23212 8168
rect 23252 8128 23253 8168
rect 23211 8119 23253 8128
rect 23019 8084 23061 8093
rect 23019 8044 23020 8084
rect 23060 8044 23061 8084
rect 23019 8035 23061 8044
rect 23020 7950 23060 8035
rect 23212 8034 23252 8119
rect 23308 7165 23348 8464
rect 23404 7916 23444 7925
rect 23500 7916 23540 8464
rect 23444 7876 23540 7916
rect 23404 7867 23444 7876
rect 23788 7589 23828 8800
rect 23884 8672 23924 8681
rect 23884 7832 23924 8632
rect 23980 8672 24020 8681
rect 24076 8672 24116 10672
rect 24268 9941 24308 10672
rect 24363 10016 24405 10025
rect 24363 9976 24364 10016
rect 24404 9976 24405 10016
rect 24363 9967 24405 9976
rect 24267 9932 24309 9941
rect 24267 9892 24268 9932
rect 24308 9892 24309 9932
rect 24267 9883 24309 9892
rect 24364 9428 24404 9967
rect 24268 9388 24404 9428
rect 24171 8840 24213 8849
rect 24171 8800 24172 8840
rect 24212 8800 24213 8840
rect 24171 8791 24213 8800
rect 24020 8632 24116 8672
rect 23980 8093 24020 8632
rect 23979 8084 24021 8093
rect 23979 8044 23980 8084
rect 24020 8044 24021 8084
rect 23979 8035 24021 8044
rect 24076 8009 24116 8094
rect 24075 8000 24117 8009
rect 24075 7960 24076 8000
rect 24116 7960 24117 8000
rect 24075 7951 24117 7960
rect 23884 7792 24116 7832
rect 23883 7664 23925 7673
rect 23883 7624 23884 7664
rect 23924 7624 23925 7664
rect 23883 7615 23925 7624
rect 23787 7580 23829 7589
rect 23787 7540 23788 7580
rect 23828 7540 23829 7580
rect 23787 7531 23829 7540
rect 23212 7125 23348 7165
rect 23884 7160 23924 7615
rect 24076 7412 24116 7792
rect 24076 7363 24116 7372
rect 22923 7076 22965 7085
rect 22923 7036 22924 7076
rect 22964 7036 22965 7076
rect 22923 7027 22965 7036
rect 22828 5851 22868 5860
rect 22924 5732 22964 7027
rect 23212 6749 23252 7125
rect 23500 7120 23884 7160
rect 23211 6740 23253 6749
rect 23211 6700 23212 6740
rect 23252 6700 23253 6740
rect 23211 6691 23253 6700
rect 22636 5489 22676 5608
rect 22828 5692 22964 5732
rect 22635 5480 22677 5489
rect 22635 5440 22636 5480
rect 22676 5440 22677 5480
rect 22635 5431 22677 5440
rect 22539 5396 22581 5405
rect 22539 5356 22540 5396
rect 22580 5356 22581 5396
rect 22539 5347 22581 5356
rect 22636 5060 22676 5431
rect 22636 5020 22772 5060
rect 22732 4901 22772 5020
rect 22731 4892 22773 4901
rect 22731 4852 22732 4892
rect 22772 4852 22773 4892
rect 22731 4843 22773 4852
rect 22347 4808 22389 4817
rect 22347 4768 22348 4808
rect 22388 4768 22389 4808
rect 22347 4759 22389 4768
rect 22828 4565 22868 5692
rect 22923 5144 22965 5153
rect 22923 5104 22924 5144
rect 22964 5104 22965 5144
rect 22923 5095 22965 5104
rect 22924 4976 22964 5095
rect 22924 4927 22964 4936
rect 23116 4724 23156 4733
rect 22827 4556 22869 4565
rect 22827 4516 22828 4556
rect 22868 4516 22869 4556
rect 22827 4507 22869 4516
rect 23116 4220 23156 4684
rect 23212 4313 23252 6691
rect 23500 6488 23540 7120
rect 23884 7111 23924 7120
rect 23692 6572 23732 6581
rect 23732 6532 24020 6572
rect 23692 6523 23732 6532
rect 23307 6404 23349 6413
rect 23307 6364 23308 6404
rect 23348 6364 23349 6404
rect 23307 6355 23349 6364
rect 23308 4808 23348 6355
rect 23500 5153 23540 6448
rect 23980 6488 24020 6532
rect 23980 6439 24020 6448
rect 24076 6488 24116 6497
rect 24172 6488 24212 8791
rect 24116 6448 24212 6488
rect 24076 6439 24116 6448
rect 23499 5144 23541 5153
rect 24075 5144 24117 5153
rect 23499 5104 23500 5144
rect 23540 5104 23636 5144
rect 23499 5095 23541 5104
rect 23308 4759 23348 4768
rect 23500 4892 23540 4901
rect 23211 4304 23253 4313
rect 23211 4264 23212 4304
rect 23252 4264 23253 4304
rect 23211 4255 23253 4264
rect 22972 4180 23156 4220
rect 22972 4178 23012 4180
rect 22444 4136 22484 4145
rect 22972 4129 23012 4138
rect 22444 3893 22484 4096
rect 23116 4052 23156 4061
rect 23500 4052 23540 4852
rect 23156 4012 23540 4052
rect 23116 4003 23156 4012
rect 22443 3884 22485 3893
rect 22443 3844 22444 3884
rect 22484 3844 22485 3884
rect 22443 3835 22485 3844
rect 23596 3800 23636 5104
rect 24075 5104 24076 5144
rect 24116 5104 24117 5144
rect 24075 5095 24117 5104
rect 23788 4976 23828 4985
rect 23691 4892 23733 4901
rect 23691 4852 23692 4892
rect 23732 4852 23733 4892
rect 23691 4843 23733 4852
rect 23500 3760 23636 3800
rect 22539 3632 22581 3641
rect 22539 3592 22540 3632
rect 22580 3592 22581 3632
rect 22539 3583 22581 3592
rect 22540 3464 22580 3583
rect 22540 3415 22580 3424
rect 22443 3296 22485 3305
rect 22443 3256 22444 3296
rect 22484 3256 22485 3296
rect 22443 3247 22485 3256
rect 22300 2633 22340 2642
rect 22340 2624 22375 2633
rect 22340 2593 22388 2624
rect 22300 2584 22388 2593
rect 22060 2500 22196 2540
rect 21387 2372 21429 2381
rect 21292 2332 21388 2372
rect 21428 2332 21429 2372
rect 20852 1912 21140 1952
rect 20812 1903 20852 1912
rect 20523 1364 20565 1373
rect 20523 1324 20524 1364
rect 20564 1324 20565 1364
rect 20523 1315 20565 1324
rect 20907 1364 20949 1373
rect 20907 1324 20908 1364
rect 20948 1324 20949 1364
rect 20907 1315 20949 1324
rect 20908 1230 20948 1315
rect 21100 1280 21140 1912
rect 21195 1952 21237 1961
rect 21195 1912 21196 1952
rect 21236 1912 21237 1952
rect 21195 1903 21237 1912
rect 21196 1818 21236 1903
rect 21100 1240 21236 1280
rect 21003 1196 21045 1205
rect 21003 1156 21004 1196
rect 21044 1156 21045 1196
rect 21003 1147 21045 1156
rect 19083 944 19125 953
rect 19083 904 19084 944
rect 19124 904 19125 944
rect 19083 895 19125 904
rect 19084 80 19124 895
rect 19468 533 19508 1072
rect 20716 1112 20756 1121
rect 20716 1028 20756 1072
rect 21004 1028 21044 1147
rect 21099 1112 21141 1121
rect 21099 1072 21100 1112
rect 21140 1072 21141 1112
rect 21099 1063 21141 1072
rect 20716 988 21044 1028
rect 21100 978 21140 1063
rect 21196 1037 21236 1240
rect 21195 1028 21237 1037
rect 21195 988 21196 1028
rect 21236 988 21237 1028
rect 21195 979 21237 988
rect 21292 953 21332 2332
rect 21387 2323 21429 2332
rect 21387 1028 21429 1037
rect 21387 988 21388 1028
rect 21428 988 21429 1028
rect 21387 979 21429 988
rect 21291 944 21333 953
rect 21291 904 21292 944
rect 21332 904 21333 944
rect 21291 895 21333 904
rect 19947 860 19989 869
rect 19947 820 19948 860
rect 19988 820 19989 860
rect 19947 811 19989 820
rect 19467 524 19509 533
rect 19467 484 19468 524
rect 19508 484 19509 524
rect 19467 475 19509 484
rect 19948 113 19988 811
rect 20048 776 20416 785
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20048 727 20416 736
rect 19947 104 19989 113
rect 11596 20 12020 60
rect 12152 0 12232 80
rect 13304 0 13384 80
rect 14456 0 14536 80
rect 15608 0 15688 80
rect 16760 0 16840 80
rect 17912 0 17992 80
rect 19064 0 19144 80
rect 19947 64 19948 104
rect 19988 64 19989 104
rect 20235 104 20277 113
rect 20235 80 20236 104
rect 19947 55 19989 64
rect 20216 64 20236 80
rect 20276 80 20277 104
rect 21388 80 21428 979
rect 20276 64 20296 80
rect 20216 0 20296 64
rect 21368 0 21448 80
rect 22156 60 22196 2500
rect 22348 2120 22388 2584
rect 22444 2456 22484 3247
rect 23403 3212 23445 3221
rect 23403 3172 23404 3212
rect 23444 3172 23445 3212
rect 23403 3163 23445 3172
rect 23308 2633 23348 2718
rect 22635 2624 22677 2633
rect 22635 2584 22636 2624
rect 22676 2584 22677 2624
rect 22635 2575 22677 2584
rect 23307 2624 23349 2633
rect 23307 2584 23308 2624
rect 23348 2584 23349 2624
rect 23307 2575 23349 2584
rect 23404 2624 23444 3163
rect 23404 2575 23444 2584
rect 22444 2407 22484 2416
rect 22636 2120 22676 2575
rect 23500 2381 23540 3760
rect 23692 3464 23732 4843
rect 23788 3632 23828 4936
rect 23884 4976 23924 4985
rect 23884 3809 23924 4936
rect 24076 4229 24116 5095
rect 24172 4976 24212 6448
rect 24268 5228 24308 9388
rect 24363 9260 24405 9269
rect 24363 9220 24364 9260
rect 24404 9220 24405 9260
rect 24363 9211 24405 9220
rect 24364 9017 24404 9211
rect 24460 9101 24500 10672
rect 24652 9605 24692 10672
rect 24747 9932 24789 9941
rect 24747 9892 24748 9932
rect 24788 9892 24789 9932
rect 24747 9883 24789 9892
rect 24651 9596 24693 9605
rect 24651 9556 24652 9596
rect 24692 9556 24693 9596
rect 24651 9547 24693 9556
rect 24556 9512 24596 9521
rect 24556 9353 24596 9472
rect 24555 9344 24597 9353
rect 24555 9304 24556 9344
rect 24596 9304 24597 9344
rect 24555 9295 24597 9304
rect 24459 9092 24501 9101
rect 24459 9052 24460 9092
rect 24500 9052 24501 9092
rect 24459 9043 24501 9052
rect 24556 9017 24596 9295
rect 24363 9008 24405 9017
rect 24363 8968 24364 9008
rect 24404 8968 24405 9008
rect 24363 8959 24405 8968
rect 24555 9008 24597 9017
rect 24555 8968 24556 9008
rect 24596 8968 24597 9008
rect 24555 8959 24597 8968
rect 24364 8849 24404 8880
rect 24363 8840 24405 8849
rect 24363 8800 24364 8840
rect 24404 8800 24405 8840
rect 24363 8791 24405 8800
rect 24555 8840 24597 8849
rect 24555 8800 24556 8840
rect 24596 8800 24597 8840
rect 24555 8791 24597 8800
rect 24364 8756 24404 8791
rect 24364 8707 24404 8716
rect 24460 8672 24500 8681
rect 24556 8672 24596 8791
rect 24500 8632 24596 8672
rect 24460 8623 24500 8632
rect 24459 7580 24501 7589
rect 24459 7540 24460 7580
rect 24500 7540 24501 7580
rect 24459 7531 24501 7540
rect 24460 6488 24500 7531
rect 24748 7421 24788 9883
rect 24844 8849 24884 10672
rect 25036 10613 25076 10672
rect 25035 10604 25077 10613
rect 25035 10564 25036 10604
rect 25076 10564 25077 10604
rect 25035 10555 25077 10564
rect 25228 10529 25268 10672
rect 25419 10648 25420 10672
rect 25460 10672 25480 10688
rect 25592 10672 25672 10752
rect 25784 10672 25864 10752
rect 25976 10672 26056 10752
rect 26168 10672 26248 10752
rect 26360 10672 26440 10752
rect 26552 10672 26632 10752
rect 26744 10672 26824 10752
rect 26936 10672 27016 10752
rect 27128 10672 27208 10752
rect 27320 10672 27400 10752
rect 27512 10672 27592 10752
rect 27704 10672 27784 10752
rect 27896 10672 27976 10752
rect 28088 10672 28168 10752
rect 28280 10672 28360 10752
rect 28472 10672 28552 10752
rect 28664 10672 28744 10752
rect 28856 10672 28936 10752
rect 29048 10672 29128 10752
rect 29240 10672 29320 10752
rect 29432 10672 29512 10752
rect 29624 10672 29704 10752
rect 29816 10672 29896 10752
rect 30008 10672 30088 10752
rect 30200 10672 30280 10752
rect 30392 10672 30472 10752
rect 30584 10672 30664 10752
rect 30776 10672 30856 10752
rect 30968 10672 31048 10752
rect 31160 10672 31240 10752
rect 31352 10672 31432 10752
rect 31544 10672 31624 10752
rect 31736 10672 31816 10752
rect 31928 10672 32008 10752
rect 32120 10672 32200 10752
rect 32312 10672 32392 10752
rect 32504 10672 32584 10752
rect 32696 10672 32776 10752
rect 32888 10672 32968 10752
rect 33080 10672 33160 10752
rect 33272 10672 33352 10752
rect 33464 10672 33544 10752
rect 39627 10688 39669 10697
rect 25460 10648 25461 10672
rect 25419 10639 25461 10648
rect 24939 10520 24981 10529
rect 24939 10480 24940 10520
rect 24980 10480 24981 10520
rect 24939 10471 24981 10480
rect 25227 10520 25269 10529
rect 25227 10480 25228 10520
rect 25268 10480 25269 10520
rect 25227 10471 25269 10480
rect 24940 9680 24980 10471
rect 25036 9680 25076 9689
rect 24940 9640 25036 9680
rect 25036 9631 25076 9640
rect 25419 9512 25461 9521
rect 25419 9472 25420 9512
rect 25460 9472 25461 9512
rect 25419 9463 25461 9472
rect 25228 9428 25268 9437
rect 25228 9008 25268 9388
rect 25420 9269 25460 9463
rect 25419 9260 25461 9269
rect 25419 9220 25420 9260
rect 25460 9220 25461 9260
rect 25419 9211 25461 9220
rect 25612 9092 25652 10672
rect 25804 9101 25844 10672
rect 25803 9092 25845 9101
rect 25612 9052 25748 9092
rect 25228 8968 25652 9008
rect 24843 8840 24885 8849
rect 24843 8800 24844 8840
rect 24884 8800 24885 8840
rect 24843 8791 24885 8800
rect 24844 7757 24884 8791
rect 25468 8681 25508 8690
rect 24940 8672 24980 8681
rect 25508 8641 25556 8672
rect 25468 8632 25556 8641
rect 24940 8177 24980 8632
rect 25323 8420 25365 8429
rect 25323 8380 25324 8420
rect 25364 8380 25365 8420
rect 25323 8371 25365 8380
rect 24939 8168 24981 8177
rect 24939 8128 24940 8168
rect 24980 8128 24981 8168
rect 24939 8119 24981 8128
rect 24843 7748 24885 7757
rect 24843 7708 24844 7748
rect 24884 7708 24885 7748
rect 24843 7699 24885 7708
rect 24555 7412 24597 7421
rect 24555 7372 24556 7412
rect 24596 7372 24597 7412
rect 24555 7363 24597 7372
rect 24747 7412 24789 7421
rect 24747 7372 24748 7412
rect 24788 7372 24789 7412
rect 24747 7363 24789 7372
rect 24363 5648 24405 5657
rect 24363 5608 24364 5648
rect 24404 5608 24405 5648
rect 24363 5599 24405 5608
rect 24364 5514 24404 5599
rect 24268 5188 24404 5228
rect 24268 4985 24308 5070
rect 24267 4976 24309 4985
rect 24172 4936 24268 4976
rect 24308 4936 24309 4976
rect 24267 4927 24309 4936
rect 24364 4976 24404 5188
rect 24460 5153 24500 6448
rect 24556 6404 24596 7363
rect 24747 7160 24789 7169
rect 24747 7120 24748 7160
rect 24788 7120 24789 7160
rect 24747 7111 24789 7120
rect 24651 6824 24693 6833
rect 24651 6784 24652 6824
rect 24692 6784 24693 6824
rect 24651 6775 24693 6784
rect 24556 6161 24596 6364
rect 24555 6152 24597 6161
rect 24555 6112 24556 6152
rect 24596 6112 24597 6152
rect 24555 6103 24597 6112
rect 24459 5144 24501 5153
rect 24459 5104 24460 5144
rect 24500 5104 24501 5144
rect 24652 5144 24692 6775
rect 24748 6413 24788 7111
rect 24940 6833 24980 8119
rect 25324 8000 25364 8371
rect 25516 8168 25556 8632
rect 25612 8588 25652 8968
rect 25612 8539 25652 8548
rect 25708 8420 25748 9052
rect 25803 9052 25804 9092
rect 25844 9052 25845 9092
rect 25803 9043 25845 9052
rect 25516 8119 25556 8128
rect 25612 8380 25748 8420
rect 25900 8672 25940 8681
rect 25324 7673 25364 7960
rect 25323 7664 25365 7673
rect 25323 7624 25324 7664
rect 25364 7624 25460 7664
rect 25323 7615 25365 7624
rect 24939 6824 24981 6833
rect 24939 6784 24940 6824
rect 24980 6784 24981 6824
rect 24939 6775 24981 6784
rect 25035 6656 25077 6665
rect 25035 6616 25036 6656
rect 25076 6616 25077 6656
rect 25035 6607 25077 6616
rect 25036 6488 25076 6607
rect 25076 6448 25268 6488
rect 25036 6439 25076 6448
rect 24747 6404 24789 6413
rect 24747 6364 24748 6404
rect 24788 6364 24789 6404
rect 24747 6355 24789 6364
rect 24843 6236 24885 6245
rect 24843 6196 24844 6236
rect 24884 6196 24885 6236
rect 24843 6187 24885 6196
rect 24652 5104 24788 5144
rect 24459 5095 24501 5104
rect 24364 4808 24404 4936
rect 24651 4976 24693 4985
rect 24651 4936 24652 4976
rect 24692 4936 24693 4976
rect 24651 4927 24693 4936
rect 24172 4768 24404 4808
rect 24075 4220 24117 4229
rect 24075 4180 24076 4220
rect 24116 4180 24117 4220
rect 24075 4171 24117 4180
rect 24076 4061 24116 4171
rect 24075 4052 24117 4061
rect 24075 4012 24076 4052
rect 24116 4012 24117 4052
rect 24075 4003 24117 4012
rect 23883 3800 23925 3809
rect 23883 3760 23884 3800
rect 23924 3760 23925 3800
rect 23883 3751 23925 3760
rect 24172 3716 24212 4768
rect 24459 4724 24501 4733
rect 24459 4684 24460 4724
rect 24500 4684 24501 4724
rect 24459 4675 24501 4684
rect 24267 4304 24309 4313
rect 24267 4264 24268 4304
rect 24308 4264 24309 4304
rect 24267 4255 24309 4264
rect 24076 3676 24212 3716
rect 23980 3632 24020 3641
rect 23788 3592 23980 3632
rect 23980 3583 24020 3592
rect 23788 3464 23828 3473
rect 23692 3424 23788 3464
rect 23692 3053 23732 3424
rect 23788 3415 23828 3424
rect 24076 3053 24116 3676
rect 24171 3548 24213 3557
rect 24171 3508 24172 3548
rect 24212 3508 24213 3548
rect 24171 3499 24213 3508
rect 23691 3044 23733 3053
rect 23691 3004 23692 3044
rect 23732 3004 23733 3044
rect 23691 2995 23733 3004
rect 23883 3044 23925 3053
rect 23883 3004 23884 3044
rect 23924 3004 23925 3044
rect 23883 2995 23925 3004
rect 24075 3044 24117 3053
rect 24075 3004 24076 3044
rect 24116 3004 24117 3044
rect 24075 2995 24117 3004
rect 23787 2708 23829 2717
rect 23787 2668 23788 2708
rect 23828 2668 23829 2708
rect 23787 2659 23829 2668
rect 23884 2708 23924 2995
rect 23884 2659 23924 2668
rect 23788 2574 23828 2659
rect 23499 2372 23541 2381
rect 23499 2332 23500 2372
rect 23540 2332 23541 2372
rect 23499 2323 23541 2332
rect 22348 2080 22580 2120
rect 22444 1952 22484 1961
rect 22348 1112 22388 1123
rect 22348 1037 22388 1072
rect 22347 1028 22389 1037
rect 22347 988 22348 1028
rect 22388 988 22389 1028
rect 22347 979 22389 988
rect 22444 869 22484 1912
rect 22540 1280 22580 2080
rect 22636 2071 22676 2080
rect 22827 1952 22869 1961
rect 22827 1912 22828 1952
rect 22868 1912 22869 1952
rect 22827 1903 22869 1912
rect 22828 1373 22868 1903
rect 23500 1877 23540 2323
rect 24075 1952 24117 1961
rect 24075 1912 24076 1952
rect 24116 1912 24117 1952
rect 24075 1903 24117 1912
rect 23019 1868 23061 1877
rect 23019 1828 23020 1868
rect 23060 1828 23061 1868
rect 23019 1819 23061 1828
rect 23499 1868 23541 1877
rect 23499 1828 23500 1868
rect 23540 1828 23541 1868
rect 23499 1819 23541 1828
rect 23020 1457 23060 1819
rect 24076 1818 24116 1903
rect 24172 1541 24212 3499
rect 24268 2120 24308 4255
rect 24364 3380 24404 3389
rect 24364 2801 24404 3340
rect 24363 2792 24405 2801
rect 24363 2752 24364 2792
rect 24404 2752 24405 2792
rect 24363 2743 24405 2752
rect 24364 2624 24404 2633
rect 24460 2624 24500 4675
rect 24555 4304 24597 4313
rect 24555 4264 24556 4304
rect 24596 4264 24597 4304
rect 24555 4255 24597 4264
rect 24556 4136 24596 4255
rect 24556 4087 24596 4096
rect 24652 4136 24692 4927
rect 24555 3212 24597 3221
rect 24555 3172 24556 3212
rect 24596 3172 24597 3212
rect 24555 3163 24597 3172
rect 24556 3078 24596 3163
rect 24555 2792 24597 2801
rect 24555 2752 24556 2792
rect 24596 2752 24597 2792
rect 24555 2743 24597 2752
rect 24404 2584 24500 2624
rect 24364 2575 24404 2584
rect 24556 2540 24596 2743
rect 24652 2717 24692 4096
rect 24748 3893 24788 5104
rect 24844 4976 24884 6187
rect 25131 6152 25173 6161
rect 25131 6112 25132 6152
rect 25172 6112 25173 6152
rect 25131 6103 25173 6112
rect 24939 5480 24981 5489
rect 24939 5440 24940 5480
rect 24980 5440 24981 5480
rect 24939 5431 24981 5440
rect 24844 4733 24884 4936
rect 24843 4724 24885 4733
rect 24843 4684 24844 4724
rect 24884 4684 24885 4724
rect 24843 4675 24885 4684
rect 24747 3884 24789 3893
rect 24747 3844 24748 3884
rect 24788 3844 24789 3884
rect 24747 3835 24789 3844
rect 24940 3800 24980 5431
rect 25132 4220 25172 6103
rect 25132 4171 25172 4180
rect 25036 4136 25076 4147
rect 25228 4136 25268 6448
rect 25420 6152 25460 7624
rect 25612 6665 25652 8380
rect 25707 8252 25749 8261
rect 25707 8212 25708 8252
rect 25748 8212 25749 8252
rect 25707 8203 25749 8212
rect 25708 8168 25748 8203
rect 25708 8117 25748 8128
rect 25900 8084 25940 8632
rect 25996 8672 26036 10672
rect 26188 9176 26228 10672
rect 26380 9941 26420 10672
rect 26572 10025 26612 10672
rect 26571 10016 26613 10025
rect 26571 9976 26572 10016
rect 26612 9976 26613 10016
rect 26571 9967 26613 9976
rect 26379 9932 26421 9941
rect 26379 9892 26380 9932
rect 26420 9892 26421 9932
rect 26379 9883 26421 9892
rect 26668 9512 26708 9521
rect 26572 9472 26668 9512
rect 26572 9353 26612 9472
rect 26668 9463 26708 9472
rect 26571 9344 26613 9353
rect 26764 9344 26804 10672
rect 26956 9932 26996 10672
rect 27148 10445 27188 10672
rect 27147 10436 27189 10445
rect 27147 10396 27148 10436
rect 27188 10396 27189 10436
rect 27147 10387 27189 10396
rect 26956 9892 27188 9932
rect 27051 9764 27093 9773
rect 27051 9724 27052 9764
rect 27092 9724 27093 9764
rect 27051 9715 27093 9724
rect 27052 9680 27092 9715
rect 27052 9629 27092 9640
rect 26571 9304 26572 9344
rect 26612 9304 26613 9344
rect 26571 9295 26613 9304
rect 26668 9304 26804 9344
rect 26860 9344 26900 9353
rect 26900 9304 27092 9344
rect 26092 9136 26228 9176
rect 26092 9008 26132 9136
rect 26092 8968 26228 9008
rect 25996 8623 26036 8632
rect 25900 8044 26036 8084
rect 25900 7916 25940 7925
rect 25804 7876 25900 7916
rect 25611 6656 25653 6665
rect 25611 6616 25612 6656
rect 25652 6616 25653 6656
rect 25611 6607 25653 6616
rect 25708 6656 25748 6665
rect 25804 6656 25844 7876
rect 25900 7867 25940 7876
rect 25996 7673 26036 8044
rect 26092 7905 26132 7914
rect 25995 7664 26037 7673
rect 25995 7624 25996 7664
rect 26036 7624 26037 7664
rect 25995 7615 26037 7624
rect 25748 6616 25844 6656
rect 25996 7160 26036 7169
rect 25708 6607 25748 6616
rect 25564 6478 25604 6487
rect 25604 6438 25844 6474
rect 25564 6434 25844 6438
rect 25564 6429 25604 6434
rect 25420 6112 25652 6152
rect 25612 5648 25652 6112
rect 25804 5900 25844 6434
rect 25804 5851 25844 5860
rect 25996 5657 26036 7120
rect 26092 6656 26132 7865
rect 26188 7832 26228 8968
rect 26283 8924 26325 8933
rect 26283 8884 26284 8924
rect 26324 8884 26325 8924
rect 26283 8875 26325 8884
rect 26284 8168 26324 8875
rect 26476 8849 26516 8851
rect 26475 8840 26517 8849
rect 26475 8800 26476 8840
rect 26516 8800 26517 8840
rect 26475 8791 26517 8800
rect 26476 8756 26516 8791
rect 26476 8707 26516 8716
rect 26380 8672 26420 8681
rect 26380 8588 26420 8632
rect 26571 8588 26613 8597
rect 26380 8548 26572 8588
rect 26612 8548 26613 8588
rect 26571 8539 26613 8548
rect 26379 8336 26421 8345
rect 26379 8296 26380 8336
rect 26420 8296 26421 8336
rect 26379 8287 26421 8296
rect 26284 8119 26324 8128
rect 26188 7792 26324 7832
rect 26187 7664 26229 7673
rect 26187 7624 26188 7664
rect 26228 7624 26229 7664
rect 26187 7615 26229 7624
rect 26188 7412 26228 7615
rect 26188 7363 26228 7372
rect 26092 6616 26228 6656
rect 26092 6488 26132 6499
rect 26092 6413 26132 6448
rect 26091 6404 26133 6413
rect 26091 6364 26092 6404
rect 26132 6364 26133 6404
rect 26091 6355 26133 6364
rect 25612 5599 25652 5608
rect 25995 5648 26037 5657
rect 25995 5608 25996 5648
rect 26036 5608 26037 5648
rect 25995 5599 26037 5608
rect 26092 5648 26132 5657
rect 26092 5405 26132 5608
rect 26091 5396 26133 5405
rect 26091 5356 26092 5396
rect 26132 5356 26133 5396
rect 26091 5347 26133 5356
rect 25515 5060 25557 5069
rect 25515 5020 25516 5060
rect 25556 5020 25557 5060
rect 25515 5011 25557 5020
rect 25372 4934 25412 4943
rect 25516 4926 25556 5011
rect 25899 4976 25941 4985
rect 25899 4936 25900 4976
rect 25940 4936 25941 4976
rect 25899 4927 25941 4936
rect 25372 4892 25412 4894
rect 25372 4852 25460 4892
rect 25420 4808 25460 4852
rect 25900 4842 25940 4927
rect 25708 4808 25748 4817
rect 25420 4768 25708 4808
rect 25708 4759 25748 4768
rect 25612 4136 25652 4145
rect 26092 4141 26132 4150
rect 25228 4096 25612 4136
rect 25652 4096 25748 4136
rect 25036 4061 25076 4096
rect 25612 4087 25652 4096
rect 25035 4052 25077 4061
rect 25035 4012 25036 4052
rect 25076 4012 25077 4052
rect 25035 4003 25077 4012
rect 25611 3884 25653 3893
rect 25611 3844 25612 3884
rect 25652 3844 25653 3884
rect 25611 3835 25653 3844
rect 24940 3760 25172 3800
rect 24747 3716 24789 3725
rect 24747 3676 24748 3716
rect 24788 3676 24789 3716
rect 24747 3667 24789 3676
rect 24748 3380 24788 3667
rect 24940 3557 24980 3760
rect 24939 3548 24981 3557
rect 24939 3508 24940 3548
rect 24980 3508 24981 3548
rect 24939 3499 24981 3508
rect 24748 3331 24788 3340
rect 25035 3380 25077 3389
rect 25035 3340 25036 3380
rect 25076 3340 25077 3380
rect 25035 3331 25077 3340
rect 25132 3380 25172 3760
rect 25515 3464 25557 3473
rect 25515 3424 25516 3464
rect 25556 3424 25557 3464
rect 25515 3415 25557 3424
rect 25132 3331 25172 3340
rect 25227 3380 25269 3389
rect 25227 3340 25228 3380
rect 25268 3340 25269 3380
rect 25227 3331 25269 3340
rect 24939 3296 24981 3305
rect 24939 3256 24940 3296
rect 24980 3256 24981 3296
rect 24939 3247 24981 3256
rect 24940 3162 24980 3247
rect 24939 3044 24981 3053
rect 24939 3004 24940 3044
rect 24980 3004 24981 3044
rect 24939 2995 24981 3004
rect 24651 2708 24693 2717
rect 24651 2668 24652 2708
rect 24692 2668 24693 2708
rect 24651 2659 24693 2668
rect 24268 2071 24308 2080
rect 24460 2500 24596 2540
rect 24267 1952 24309 1961
rect 24267 1912 24268 1952
rect 24308 1912 24309 1952
rect 24267 1903 24309 1912
rect 24171 1532 24213 1541
rect 24171 1492 24172 1532
rect 24212 1492 24213 1532
rect 24171 1483 24213 1492
rect 23019 1448 23061 1457
rect 23019 1408 23020 1448
rect 23060 1408 23061 1448
rect 23019 1399 23061 1408
rect 22827 1364 22869 1373
rect 22827 1324 22828 1364
rect 22868 1324 22869 1364
rect 22827 1315 22869 1324
rect 22540 1231 22580 1240
rect 23020 1112 23060 1399
rect 23020 1063 23060 1072
rect 24268 1112 24308 1903
rect 24460 1625 24500 2500
rect 24556 1952 24596 1961
rect 24459 1616 24501 1625
rect 24459 1576 24460 1616
rect 24500 1576 24501 1616
rect 24459 1567 24501 1576
rect 24460 1364 24500 1373
rect 24556 1364 24596 1912
rect 24652 1952 24692 2659
rect 24844 2629 24884 2638
rect 24747 2120 24789 2129
rect 24747 2080 24748 2120
rect 24788 2080 24789 2120
rect 24747 2071 24789 2080
rect 24652 1903 24692 1912
rect 24748 1793 24788 2071
rect 24747 1784 24789 1793
rect 24747 1744 24748 1784
rect 24788 1744 24789 1784
rect 24747 1735 24789 1744
rect 24500 1324 24596 1364
rect 24460 1315 24500 1324
rect 24652 1280 24692 1289
rect 24844 1280 24884 2589
rect 24940 1952 24980 2995
rect 25036 2540 25076 3331
rect 25131 3128 25173 3137
rect 25131 3088 25132 3128
rect 25172 3088 25173 3128
rect 25131 3079 25173 3088
rect 25036 2491 25076 2500
rect 25036 1952 25076 1961
rect 24940 1912 25036 1952
rect 25036 1903 25076 1912
rect 25132 1952 25172 3079
rect 25132 1903 25172 1912
rect 25228 2624 25268 3331
rect 25323 3296 25365 3305
rect 25323 3256 25324 3296
rect 25364 3256 25365 3296
rect 25323 3247 25365 3256
rect 25324 3162 25364 3247
rect 25516 2969 25556 3415
rect 25515 2960 25557 2969
rect 25515 2920 25516 2960
rect 25556 2920 25557 2960
rect 25515 2911 25557 2920
rect 25228 1541 25268 2584
rect 25612 1952 25652 3835
rect 25612 1903 25652 1912
rect 25708 1877 25748 4096
rect 26092 2885 26132 4101
rect 26091 2876 26133 2885
rect 26091 2836 26092 2876
rect 26132 2836 26133 2876
rect 26091 2827 26133 2836
rect 26091 2036 26133 2045
rect 26091 1996 26092 2036
rect 26132 1996 26133 2036
rect 26091 1987 26133 1996
rect 26092 1947 26132 1987
rect 26092 1898 26132 1907
rect 25707 1868 25749 1877
rect 25707 1828 25708 1868
rect 25748 1828 25749 1868
rect 25707 1819 25749 1828
rect 25899 1616 25941 1625
rect 25899 1576 25900 1616
rect 25940 1576 25941 1616
rect 25899 1567 25941 1576
rect 25227 1532 25269 1541
rect 25227 1492 25228 1532
rect 25268 1492 25269 1532
rect 25227 1483 25269 1492
rect 25900 1289 25940 1567
rect 24692 1240 24884 1280
rect 25899 1280 25941 1289
rect 25899 1240 25900 1280
rect 25940 1240 25941 1280
rect 24652 1231 24692 1240
rect 25899 1231 25941 1240
rect 26091 1280 26133 1289
rect 26091 1240 26092 1280
rect 26132 1240 26133 1280
rect 26091 1231 26133 1240
rect 26092 1121 26132 1231
rect 26188 1205 26228 6616
rect 26284 4565 26324 7792
rect 26283 4556 26325 4565
rect 26283 4516 26284 4556
rect 26324 4516 26325 4556
rect 26283 4507 26325 4516
rect 26283 3968 26325 3977
rect 26283 3928 26284 3968
rect 26324 3928 26325 3968
rect 26283 3919 26325 3928
rect 26284 3834 26324 3919
rect 26380 3800 26420 8287
rect 26668 6497 26708 9304
rect 26860 9295 26900 9304
rect 26955 9176 26997 9185
rect 26860 9136 26956 9176
rect 26996 9136 26997 9176
rect 26860 9092 26900 9136
rect 26955 9127 26997 9136
rect 26764 9052 26900 9092
rect 26764 7832 26804 9052
rect 27052 9008 27092 9304
rect 26860 8968 27092 9008
rect 26860 8000 26900 8968
rect 26955 8672 26997 8681
rect 26955 8632 26956 8672
rect 26996 8632 27092 8672
rect 26955 8623 26997 8632
rect 26956 8538 26996 8623
rect 26860 7951 26900 7960
rect 26956 8000 26996 8009
rect 26956 7832 26996 7960
rect 26764 7792 26996 7832
rect 27052 7169 27092 8632
rect 27148 8084 27188 9892
rect 27243 9428 27285 9437
rect 27243 9388 27244 9428
rect 27284 9388 27285 9428
rect 27243 9379 27285 9388
rect 27244 9294 27284 9379
rect 27340 8261 27380 10672
rect 27532 9689 27572 10672
rect 27531 9680 27573 9689
rect 27531 9640 27532 9680
rect 27572 9640 27573 9680
rect 27531 9631 27573 9640
rect 27627 9428 27669 9437
rect 27627 9388 27628 9428
rect 27668 9388 27669 9428
rect 27627 9379 27669 9388
rect 27484 8681 27524 8690
rect 27524 8641 27572 8672
rect 27484 8632 27572 8641
rect 27339 8252 27381 8261
rect 27339 8212 27340 8252
rect 27380 8212 27381 8252
rect 27339 8203 27381 8212
rect 27148 8044 27476 8084
rect 27051 7160 27093 7169
rect 27051 7120 27052 7160
rect 27092 7120 27093 7160
rect 27051 7111 27093 7120
rect 26763 6908 26805 6917
rect 26763 6868 26764 6908
rect 26804 6868 26805 6908
rect 26763 6859 26805 6868
rect 26667 6488 26709 6497
rect 26667 6448 26668 6488
rect 26708 6448 26709 6488
rect 26667 6439 26709 6448
rect 26571 5732 26613 5741
rect 26571 5692 26572 5732
rect 26612 5692 26613 5732
rect 26571 5683 26613 5692
rect 26572 4985 26612 5683
rect 26571 4976 26613 4985
rect 26571 4936 26572 4976
rect 26612 4936 26613 4976
rect 26571 4927 26613 4936
rect 26380 3760 26480 3800
rect 26440 3716 26480 3760
rect 26440 3676 26516 3716
rect 26476 3389 26516 3676
rect 26572 3473 26612 4927
rect 26668 4136 26708 4145
rect 26668 3632 26708 4096
rect 26764 4136 26804 6859
rect 27147 6740 27189 6749
rect 27147 6700 27148 6740
rect 27188 6700 27189 6740
rect 27147 6691 27189 6700
rect 27148 6497 27188 6691
rect 27147 6488 27189 6497
rect 27147 6448 27148 6488
rect 27188 6448 27189 6488
rect 27147 6439 27189 6448
rect 27147 4976 27189 4985
rect 27147 4936 27148 4976
rect 27188 4936 27189 4976
rect 27147 4927 27189 4936
rect 27148 4842 27188 4927
rect 27244 4229 27284 8044
rect 27436 8000 27476 8044
rect 27436 7951 27476 7960
rect 27340 7916 27380 7925
rect 27340 7589 27380 7876
rect 27339 7580 27381 7589
rect 27339 7540 27340 7580
rect 27380 7540 27381 7580
rect 27339 7531 27381 7540
rect 27532 7076 27572 8632
rect 27628 8588 27668 9379
rect 27628 8539 27668 8548
rect 27724 7589 27764 10672
rect 27916 10109 27956 10672
rect 27915 10100 27957 10109
rect 27915 10060 27916 10100
rect 27956 10060 27957 10100
rect 27915 10051 27957 10060
rect 28108 8840 28148 10672
rect 28300 9008 28340 10672
rect 28300 8968 28436 9008
rect 28108 8800 28244 8840
rect 28012 8765 28052 8767
rect 28011 8756 28053 8765
rect 28011 8716 28012 8756
rect 28052 8716 28053 8756
rect 28011 8707 28053 8716
rect 28012 8672 28052 8707
rect 28204 8677 28244 8800
rect 28299 8756 28341 8765
rect 28299 8716 28300 8756
rect 28340 8716 28341 8756
rect 28299 8707 28341 8716
rect 28012 8623 28052 8632
rect 28108 8637 28244 8677
rect 27820 8504 27860 8513
rect 27820 8009 27860 8464
rect 27915 8336 27957 8345
rect 27915 8296 27916 8336
rect 27956 8296 27957 8336
rect 27915 8287 27957 8296
rect 27819 8000 27861 8009
rect 27819 7960 27820 8000
rect 27860 7960 27861 8000
rect 27819 7951 27861 7960
rect 27916 8000 27956 8287
rect 27916 7951 27956 7960
rect 28108 7673 28148 8637
rect 28300 7841 28340 8707
rect 28396 8681 28436 8968
rect 28492 8924 28532 10672
rect 28492 8884 28628 8924
rect 28395 8672 28437 8681
rect 28395 8632 28396 8672
rect 28436 8632 28437 8672
rect 28395 8623 28437 8632
rect 28588 8345 28628 8884
rect 28684 8765 28724 10672
rect 28683 8756 28725 8765
rect 28683 8716 28684 8756
rect 28724 8716 28725 8756
rect 28683 8707 28725 8716
rect 28876 8681 28916 10672
rect 28971 9092 29013 9101
rect 28971 9052 28972 9092
rect 29012 9052 29013 9092
rect 28971 9043 29013 9052
rect 28875 8672 28917 8681
rect 28875 8632 28876 8672
rect 28916 8632 28917 8672
rect 28875 8623 28917 8632
rect 28779 8504 28821 8513
rect 28779 8464 28780 8504
rect 28820 8464 28821 8504
rect 28779 8455 28821 8464
rect 28587 8336 28629 8345
rect 28587 8296 28588 8336
rect 28628 8296 28724 8336
rect 28587 8287 28629 8296
rect 28491 8252 28533 8261
rect 28491 8212 28492 8252
rect 28532 8212 28533 8252
rect 28491 8203 28533 8212
rect 28395 8000 28437 8009
rect 28395 7955 28396 8000
rect 28436 7955 28437 8000
rect 28395 7951 28437 7955
rect 28396 7865 28436 7951
rect 28299 7832 28341 7841
rect 28299 7792 28300 7832
rect 28340 7792 28341 7832
rect 28299 7783 28341 7792
rect 28107 7664 28149 7673
rect 28107 7624 28108 7664
rect 28148 7624 28149 7664
rect 28107 7615 28149 7624
rect 27723 7580 27765 7589
rect 27723 7540 27724 7580
rect 27764 7540 27765 7580
rect 27723 7531 27765 7540
rect 28203 7580 28245 7589
rect 28203 7540 28204 7580
rect 28244 7540 28245 7580
rect 28203 7531 28245 7540
rect 27436 7036 27572 7076
rect 27820 7160 27860 7169
rect 27340 6488 27380 6497
rect 27340 5816 27380 6448
rect 27436 5900 27476 7036
rect 27820 6740 27860 7120
rect 27916 7160 27956 7169
rect 27916 7001 27956 7120
rect 27915 6992 27957 7001
rect 27915 6952 27916 6992
rect 27956 6952 27957 6992
rect 27915 6943 27957 6952
rect 27820 6700 28052 6740
rect 27532 6572 27572 6581
rect 27572 6532 27860 6572
rect 27532 6523 27572 6532
rect 27820 6488 27860 6532
rect 27916 6497 27956 6582
rect 27820 6439 27860 6448
rect 27915 6488 27957 6497
rect 27915 6448 27916 6488
rect 27956 6448 27957 6488
rect 27915 6439 27957 6448
rect 27627 6320 27669 6329
rect 28012 6320 28052 6700
rect 27627 6280 27628 6320
rect 27668 6280 27669 6320
rect 27627 6271 27669 6280
rect 27724 6280 28052 6320
rect 27532 5900 27572 5909
rect 27436 5860 27532 5900
rect 27532 5851 27572 5860
rect 27340 5776 27466 5816
rect 27426 5741 27466 5776
rect 27426 5732 27477 5741
rect 27426 5692 27436 5732
rect 27476 5692 27477 5732
rect 27435 5683 27477 5692
rect 27339 5648 27381 5657
rect 27339 5608 27340 5648
rect 27380 5608 27381 5648
rect 27339 5599 27381 5608
rect 27051 4220 27093 4229
rect 27148 4220 27188 4229
rect 27051 4180 27052 4220
rect 27092 4180 27148 4220
rect 27051 4171 27093 4180
rect 27148 4171 27188 4180
rect 27243 4220 27285 4229
rect 27243 4180 27244 4220
rect 27284 4180 27285 4220
rect 27243 4171 27285 4180
rect 26764 4087 26804 4096
rect 27244 4086 27284 4171
rect 27147 3884 27189 3893
rect 27147 3844 27148 3884
rect 27188 3844 27189 3884
rect 27147 3835 27189 3844
rect 26956 3632 26996 3641
rect 26668 3592 26956 3632
rect 26956 3583 26996 3592
rect 26571 3464 26613 3473
rect 26571 3424 26572 3464
rect 26612 3424 26613 3464
rect 26571 3415 26613 3424
rect 26763 3464 26805 3473
rect 26763 3424 26764 3464
rect 26804 3424 26805 3464
rect 26763 3415 26805 3424
rect 27148 3464 27188 3835
rect 27148 3415 27188 3424
rect 26475 3380 26517 3389
rect 26475 3340 26476 3380
rect 26516 3340 26517 3380
rect 26475 3331 26517 3340
rect 26764 3330 26804 3415
rect 27051 3044 27093 3053
rect 27051 3004 27052 3044
rect 27092 3004 27093 3044
rect 27051 2995 27093 3004
rect 26667 2876 26709 2885
rect 26667 2836 26668 2876
rect 26708 2836 26709 2876
rect 26667 2827 26709 2836
rect 26668 2742 26708 2827
rect 27052 2717 27092 2995
rect 27051 2708 27093 2717
rect 27051 2668 27052 2708
rect 27092 2668 27093 2708
rect 27051 2659 27093 2668
rect 26476 2624 26516 2633
rect 26476 2540 26516 2584
rect 27052 2574 27092 2659
rect 26476 2500 26708 2540
rect 26283 2120 26325 2129
rect 26283 2080 26284 2120
rect 26324 2080 26325 2120
rect 26283 2071 26325 2080
rect 26284 1986 26324 2071
rect 26475 2036 26517 2045
rect 26475 1996 26476 2036
rect 26516 1996 26517 2036
rect 26475 1987 26517 1996
rect 26476 1902 26516 1987
rect 26668 1961 26708 2500
rect 27244 2456 27284 2465
rect 27244 2213 27284 2416
rect 27243 2204 27285 2213
rect 27243 2164 27244 2204
rect 27284 2164 27285 2204
rect 27243 2155 27285 2164
rect 26667 1952 26709 1961
rect 26667 1912 26668 1952
rect 26708 1912 26709 1952
rect 26667 1903 26709 1912
rect 26668 1818 26708 1903
rect 26283 1364 26325 1373
rect 26283 1324 26284 1364
rect 26324 1324 26325 1364
rect 26283 1315 26325 1324
rect 26187 1196 26229 1205
rect 26187 1156 26188 1196
rect 26228 1156 26229 1196
rect 26187 1147 26229 1156
rect 26284 1121 26324 1315
rect 24268 1063 24308 1072
rect 24844 1112 24884 1121
rect 24844 869 24884 1072
rect 26091 1112 26133 1121
rect 26091 1072 26092 1112
rect 26132 1072 26133 1112
rect 26091 1063 26133 1072
rect 26283 1112 26325 1121
rect 26283 1072 26284 1112
rect 26324 1072 26325 1112
rect 26283 1063 26325 1072
rect 25995 1028 26037 1037
rect 25995 988 25996 1028
rect 26036 988 26037 1028
rect 25995 979 26037 988
rect 22443 860 22485 869
rect 22443 820 22444 860
rect 22484 820 22485 860
rect 22443 811 22485 820
rect 24843 860 24885 869
rect 24843 820 24844 860
rect 24884 820 24885 860
rect 24843 811 24885 820
rect 23691 272 23733 281
rect 23691 232 23692 272
rect 23732 232 23733 272
rect 23691 223 23733 232
rect 22348 80 22580 104
rect 23692 80 23732 223
rect 24843 188 24885 197
rect 24843 148 24844 188
rect 24884 148 24885 188
rect 24843 139 24885 148
rect 24844 80 24884 139
rect 25996 80 26036 979
rect 26092 978 26132 1063
rect 26284 978 26324 1063
rect 27147 944 27189 953
rect 27147 904 27148 944
rect 27188 904 27189 944
rect 27147 895 27189 904
rect 27148 80 27188 895
rect 27340 869 27380 5599
rect 27435 5564 27477 5573
rect 27435 5524 27436 5564
rect 27476 5524 27477 5564
rect 27435 5515 27477 5524
rect 27436 5153 27476 5515
rect 27628 5321 27668 6271
rect 27724 5900 27764 6280
rect 27724 5851 27764 5860
rect 27915 5732 27957 5741
rect 27915 5692 27916 5732
rect 27956 5692 27957 5732
rect 27915 5683 27957 5692
rect 27916 5648 27956 5683
rect 27916 5597 27956 5608
rect 28011 5480 28053 5489
rect 28011 5440 28012 5480
rect 28052 5440 28053 5480
rect 28011 5431 28053 5440
rect 27627 5312 27669 5321
rect 27627 5272 27628 5312
rect 27668 5272 27669 5312
rect 27627 5263 27669 5272
rect 27915 5312 27957 5321
rect 27915 5272 27916 5312
rect 27956 5272 27957 5312
rect 27915 5263 27957 5272
rect 27435 5144 27477 5153
rect 27435 5104 27436 5144
rect 27476 5104 27477 5144
rect 27435 5095 27477 5104
rect 27436 4892 27476 5095
rect 27916 4985 27956 5263
rect 27915 4976 27957 4985
rect 27915 4936 27916 4976
rect 27956 4936 27957 4976
rect 27915 4927 27957 4936
rect 27436 4843 27476 4852
rect 27916 4842 27956 4927
rect 27627 4724 27669 4733
rect 27627 4684 27628 4724
rect 27668 4684 27669 4724
rect 27627 4675 27669 4684
rect 27628 4590 27668 4675
rect 27723 4640 27765 4649
rect 27723 4600 27724 4640
rect 27764 4600 27765 4640
rect 27723 4591 27765 4600
rect 27531 4472 27573 4481
rect 27531 4432 27532 4472
rect 27572 4432 27573 4472
rect 27531 4423 27573 4432
rect 27435 4136 27477 4145
rect 27435 4096 27436 4136
rect 27476 4096 27477 4136
rect 27435 4087 27477 4096
rect 27436 3893 27476 4087
rect 27532 3968 27572 4423
rect 27627 4304 27669 4313
rect 27627 4264 27628 4304
rect 27668 4264 27669 4304
rect 27627 4255 27669 4264
rect 27628 4145 27668 4255
rect 27627 4136 27669 4145
rect 27627 4096 27628 4136
rect 27668 4096 27669 4136
rect 27627 4087 27669 4096
rect 27724 4136 27764 4591
rect 27819 4304 27861 4313
rect 27819 4264 27820 4304
rect 27860 4264 27861 4304
rect 27819 4255 27861 4264
rect 27724 4087 27764 4096
rect 27820 3968 27860 4255
rect 28012 3968 28052 5431
rect 28204 4901 28244 7531
rect 28299 7412 28341 7421
rect 28299 7372 28300 7412
rect 28340 7372 28341 7412
rect 28299 7363 28341 7372
rect 28300 7244 28340 7363
rect 28300 7195 28340 7204
rect 28396 7244 28436 7253
rect 28492 7244 28532 8203
rect 28587 8084 28629 8093
rect 28587 8044 28588 8084
rect 28628 8044 28629 8084
rect 28587 8035 28629 8044
rect 28588 7950 28628 8035
rect 28587 7748 28629 7757
rect 28587 7708 28588 7748
rect 28628 7708 28629 7748
rect 28587 7699 28629 7708
rect 28436 7204 28532 7244
rect 28396 7195 28436 7204
rect 28588 7076 28628 7699
rect 28396 7036 28628 7076
rect 28396 6488 28436 7036
rect 28588 6917 28628 7036
rect 28587 6908 28629 6917
rect 28587 6868 28588 6908
rect 28628 6868 28629 6908
rect 28684 6908 28724 8296
rect 28780 8177 28820 8455
rect 28779 8168 28821 8177
rect 28779 8128 28780 8168
rect 28820 8128 28821 8168
rect 28779 8119 28821 8128
rect 28779 8000 28821 8009
rect 28779 7960 28780 8000
rect 28820 7960 28821 8000
rect 28779 7951 28821 7960
rect 28780 7866 28820 7951
rect 28779 7664 28821 7673
rect 28779 7624 28780 7664
rect 28820 7624 28821 7664
rect 28779 7615 28821 7624
rect 28780 6992 28820 7615
rect 28876 7160 28916 8623
rect 28876 7111 28916 7120
rect 28780 6952 28916 6992
rect 28684 6868 28820 6908
rect 28587 6859 28629 6868
rect 28683 6740 28725 6749
rect 28683 6700 28684 6740
rect 28724 6700 28725 6740
rect 28683 6691 28725 6700
rect 28587 6656 28629 6665
rect 28587 6616 28588 6656
rect 28628 6616 28629 6656
rect 28587 6607 28629 6616
rect 28299 6404 28341 6413
rect 28299 6364 28300 6404
rect 28340 6364 28341 6404
rect 28299 6355 28341 6364
rect 28300 6270 28340 6355
rect 28203 4892 28245 4901
rect 28203 4852 28204 4892
rect 28244 4852 28245 4892
rect 28203 4843 28245 4852
rect 28396 4313 28436 6448
rect 28491 6488 28533 6497
rect 28491 6448 28492 6488
rect 28532 6448 28533 6488
rect 28491 6439 28533 6448
rect 28395 4304 28437 4313
rect 28395 4264 28396 4304
rect 28436 4264 28437 4304
rect 28395 4255 28437 4264
rect 27532 3928 27668 3968
rect 27435 3884 27477 3893
rect 27435 3844 27436 3884
rect 27476 3844 27477 3884
rect 27435 3835 27477 3844
rect 27435 3464 27477 3473
rect 27435 3424 27436 3464
rect 27476 3424 27477 3464
rect 27435 3415 27477 3424
rect 27436 1112 27476 3415
rect 27532 2624 27572 2633
rect 27532 1364 27572 2584
rect 27628 2624 27668 3928
rect 27724 3928 27860 3968
rect 27916 3928 28052 3968
rect 28204 4141 28244 4150
rect 27724 2885 27764 3928
rect 27916 3884 27956 3928
rect 27820 3844 27956 3884
rect 27723 2876 27765 2885
rect 27723 2836 27724 2876
rect 27764 2836 27765 2876
rect 27723 2827 27765 2836
rect 27628 2575 27668 2584
rect 27820 1952 27860 3844
rect 28204 3725 28244 4101
rect 28395 3968 28437 3977
rect 28395 3928 28396 3968
rect 28436 3928 28437 3968
rect 28395 3919 28437 3928
rect 28396 3834 28436 3919
rect 28203 3716 28245 3725
rect 28203 3676 28204 3716
rect 28244 3676 28245 3716
rect 28203 3667 28245 3676
rect 28395 3464 28437 3473
rect 28395 3424 28396 3464
rect 28436 3424 28437 3464
rect 28395 3415 28437 3424
rect 28299 3380 28341 3389
rect 28299 3340 28300 3380
rect 28340 3340 28341 3380
rect 28299 3331 28341 3340
rect 28011 2876 28053 2885
rect 28011 2836 28012 2876
rect 28052 2836 28053 2876
rect 28011 2827 28053 2836
rect 28012 2708 28052 2827
rect 28012 2659 28052 2668
rect 28107 2708 28149 2717
rect 28107 2668 28108 2708
rect 28148 2668 28149 2708
rect 28107 2659 28149 2668
rect 28108 2574 28148 2659
rect 27916 1952 27956 1961
rect 28204 1952 28244 1961
rect 27820 1912 27916 1952
rect 27532 1324 27668 1364
rect 27628 1280 27668 1324
rect 27820 1289 27860 1912
rect 27916 1903 27956 1912
rect 28012 1912 28204 1952
rect 27916 1364 27956 1373
rect 28012 1364 28052 1912
rect 28204 1903 28244 1912
rect 28300 1952 28340 3331
rect 28396 3330 28436 3415
rect 28492 2624 28532 6439
rect 28588 6245 28628 6607
rect 28587 6236 28629 6245
rect 28587 6196 28588 6236
rect 28628 6196 28629 6236
rect 28587 6187 28629 6196
rect 28587 4388 28629 4397
rect 28587 4348 28588 4388
rect 28628 4348 28629 4388
rect 28587 4339 28629 4348
rect 28588 4254 28628 4339
rect 28587 3716 28629 3725
rect 28587 3676 28588 3716
rect 28628 3676 28629 3716
rect 28587 3667 28629 3676
rect 28588 3632 28628 3667
rect 28684 3632 28724 6691
rect 28780 4733 28820 6868
rect 28876 6665 28916 6952
rect 28875 6656 28917 6665
rect 28875 6616 28876 6656
rect 28916 6616 28917 6656
rect 28875 6607 28917 6616
rect 28875 6488 28917 6497
rect 28972 6488 29012 9043
rect 29068 8849 29108 10672
rect 29163 9764 29205 9773
rect 29163 9724 29164 9764
rect 29204 9724 29205 9764
rect 29163 9715 29205 9724
rect 29164 9269 29204 9715
rect 29260 9437 29300 10672
rect 29356 9512 29396 9521
rect 29259 9428 29301 9437
rect 29259 9388 29260 9428
rect 29300 9388 29301 9428
rect 29259 9379 29301 9388
rect 29356 9353 29396 9472
rect 29355 9344 29397 9353
rect 29355 9304 29356 9344
rect 29396 9304 29397 9344
rect 29355 9295 29397 9304
rect 29163 9260 29205 9269
rect 29163 9220 29164 9260
rect 29204 9220 29205 9260
rect 29163 9211 29205 9220
rect 29067 8840 29109 8849
rect 29067 8800 29068 8840
rect 29108 8800 29109 8840
rect 29067 8791 29109 8800
rect 29164 8756 29204 9211
rect 29452 9101 29492 10672
rect 29451 9092 29493 9101
rect 29451 9052 29452 9092
rect 29492 9052 29493 9092
rect 29451 9043 29493 9052
rect 29452 8756 29492 8765
rect 29164 8716 29300 8756
rect 29260 8672 29300 8716
rect 29260 8623 29300 8632
rect 29452 7757 29492 8716
rect 29644 8672 29684 10672
rect 29739 9428 29781 9437
rect 29739 9388 29740 9428
rect 29780 9388 29781 9428
rect 29739 9379 29781 9388
rect 29548 8632 29684 8672
rect 29451 7748 29493 7757
rect 29451 7708 29452 7748
rect 29492 7708 29493 7748
rect 29451 7699 29493 7708
rect 29067 7244 29109 7253
rect 29067 7204 29068 7244
rect 29108 7204 29109 7244
rect 29067 7195 29109 7204
rect 28875 6448 28876 6488
rect 28916 6448 29012 6488
rect 28875 6439 28917 6448
rect 28876 6354 28916 6439
rect 28876 4976 28916 4985
rect 28779 4724 28821 4733
rect 28779 4684 28780 4724
rect 28820 4684 28821 4724
rect 28779 4675 28821 4684
rect 28780 4136 28820 4145
rect 28780 3977 28820 4096
rect 28779 3968 28821 3977
rect 28779 3928 28780 3968
rect 28820 3928 28821 3968
rect 28779 3919 28821 3928
rect 28780 3632 28820 3641
rect 28684 3592 28780 3632
rect 28588 3581 28628 3592
rect 28780 3583 28820 3592
rect 28588 2624 28628 2633
rect 28492 2584 28588 2624
rect 28628 2584 28820 2624
rect 28588 2575 28628 2584
rect 28300 1903 28340 1912
rect 28683 1952 28725 1961
rect 28683 1912 28684 1952
rect 28724 1912 28725 1952
rect 28683 1903 28725 1912
rect 28780 1952 28820 2584
rect 28780 1903 28820 1912
rect 28684 1818 28724 1903
rect 27956 1324 28052 1364
rect 27916 1315 27956 1324
rect 28876 1289 28916 4936
rect 28971 3968 29013 3977
rect 28971 3928 28972 3968
rect 29012 3928 29013 3968
rect 28971 3919 29013 3928
rect 28972 3473 29012 3919
rect 28971 3464 29013 3473
rect 28971 3424 28972 3464
rect 29012 3424 29013 3464
rect 28971 3415 29013 3424
rect 29068 3296 29108 7195
rect 29356 7165 29396 7174
rect 29548 7160 29588 8632
rect 29643 8504 29685 8513
rect 29643 8464 29644 8504
rect 29684 8464 29685 8504
rect 29643 8455 29685 8464
rect 29644 8370 29684 8455
rect 29356 6749 29396 7125
rect 29452 7120 29588 7160
rect 29355 6740 29397 6749
rect 29355 6700 29356 6740
rect 29396 6700 29397 6740
rect 29355 6691 29397 6700
rect 29356 6474 29396 6483
rect 29356 5900 29396 6434
rect 29356 5851 29396 5860
rect 29164 5648 29204 5659
rect 29164 5573 29204 5608
rect 29163 5564 29205 5573
rect 29163 5524 29164 5564
rect 29204 5524 29205 5564
rect 29163 5515 29205 5524
rect 29164 4976 29204 4985
rect 29164 4397 29204 4936
rect 29260 4976 29300 4985
rect 29260 4817 29300 4936
rect 29259 4808 29301 4817
rect 29259 4768 29260 4808
rect 29300 4768 29301 4808
rect 29259 4759 29301 4768
rect 29163 4388 29205 4397
rect 29163 4348 29164 4388
rect 29204 4348 29205 4388
rect 29163 4339 29205 4348
rect 28972 3256 29108 3296
rect 28972 2381 29012 3256
rect 29355 3212 29397 3221
rect 29355 3172 29356 3212
rect 29396 3172 29397 3212
rect 29355 3163 29397 3172
rect 29356 2801 29396 3163
rect 29452 2876 29492 7120
rect 29548 6992 29588 7001
rect 29548 6833 29588 6952
rect 29547 6824 29589 6833
rect 29547 6784 29548 6824
rect 29588 6784 29589 6824
rect 29547 6775 29589 6784
rect 29548 6572 29588 6581
rect 29588 6532 29684 6572
rect 29548 6523 29588 6532
rect 29547 5648 29589 5657
rect 29547 5608 29548 5648
rect 29588 5608 29589 5648
rect 29547 5599 29589 5608
rect 29548 5514 29588 5599
rect 29644 5060 29684 6532
rect 29740 6329 29780 9379
rect 29836 8933 29876 10672
rect 29835 8924 29877 8933
rect 29835 8884 29836 8924
rect 29876 8884 29877 8924
rect 29835 8875 29877 8884
rect 30028 8840 30068 10672
rect 30123 9596 30165 9605
rect 30123 9556 30124 9596
rect 30164 9556 30165 9596
rect 30123 9547 30165 9556
rect 30124 9176 30164 9547
rect 30220 9260 30260 10672
rect 30412 9689 30452 10672
rect 30411 9680 30453 9689
rect 30604 9680 30644 10672
rect 30411 9640 30412 9680
rect 30452 9640 30453 9680
rect 30411 9631 30453 9640
rect 30508 9640 30644 9680
rect 30220 9220 30452 9260
rect 30124 9136 30260 9176
rect 30028 8791 30068 8800
rect 29835 8756 29877 8765
rect 29835 8716 29836 8756
rect 29876 8716 29877 8756
rect 29835 8707 29877 8716
rect 29836 8429 29876 8707
rect 29835 8420 29877 8429
rect 29835 8380 29836 8420
rect 29876 8380 29877 8420
rect 29835 8371 29877 8380
rect 30027 8000 30069 8009
rect 30027 7960 30028 8000
rect 30068 7960 30069 8000
rect 30027 7951 30069 7960
rect 30028 7866 30068 7951
rect 30220 7916 30260 9136
rect 30315 8588 30357 8597
rect 30315 8548 30316 8588
rect 30356 8548 30357 8588
rect 30315 8539 30357 8548
rect 30316 8454 30356 8539
rect 30412 8168 30452 9220
rect 30508 9092 30548 9640
rect 30796 9605 30836 10672
rect 30891 9680 30933 9689
rect 30891 9640 30892 9680
rect 30932 9640 30933 9680
rect 30891 9631 30933 9640
rect 30795 9596 30837 9605
rect 30795 9556 30796 9596
rect 30836 9556 30837 9596
rect 30795 9547 30837 9556
rect 30604 9512 30644 9523
rect 30604 9437 30644 9472
rect 30603 9428 30645 9437
rect 30603 9388 30604 9428
rect 30644 9388 30645 9428
rect 30603 9379 30645 9388
rect 30795 9260 30837 9269
rect 30795 9220 30796 9260
rect 30836 9220 30837 9260
rect 30795 9211 30837 9220
rect 30796 9126 30836 9211
rect 30508 9052 30644 9092
rect 30507 8924 30549 8933
rect 30507 8884 30508 8924
rect 30548 8884 30549 8924
rect 30507 8875 30549 8884
rect 30508 8686 30548 8875
rect 30508 8637 30548 8646
rect 30604 8513 30644 9052
rect 30892 9008 30932 9631
rect 30988 9428 31028 10672
rect 31180 9680 31220 10672
rect 31180 9640 31316 9680
rect 31180 9512 31220 9521
rect 31180 9437 31220 9472
rect 31179 9428 31221 9437
rect 30988 9388 31124 9428
rect 30796 8968 30932 9008
rect 30988 9260 31028 9269
rect 30699 8840 30741 8849
rect 30699 8800 30700 8840
rect 30740 8800 30741 8840
rect 30699 8791 30741 8800
rect 30603 8504 30645 8513
rect 30603 8464 30604 8504
rect 30644 8464 30645 8504
rect 30603 8455 30645 8464
rect 30412 8119 30452 8128
rect 30604 7916 30644 7925
rect 30220 7876 30452 7916
rect 30220 7748 30260 7757
rect 29932 7708 30220 7748
rect 29836 7253 29876 7338
rect 29835 7244 29877 7253
rect 29835 7204 29836 7244
rect 29876 7204 29877 7244
rect 29835 7195 29877 7204
rect 29932 7076 29972 7708
rect 30220 7699 30260 7708
rect 30219 7160 30261 7169
rect 30219 7120 30220 7160
rect 30260 7120 30261 7160
rect 30219 7111 30261 7120
rect 29836 7036 29972 7076
rect 29836 6488 29876 7036
rect 30220 7026 30260 7111
rect 30028 6992 30068 7001
rect 29931 6908 29973 6917
rect 29931 6868 29932 6908
rect 29972 6868 29973 6908
rect 29931 6859 29973 6868
rect 29836 6439 29876 6448
rect 29932 6488 29972 6859
rect 29932 6439 29972 6448
rect 29739 6320 29781 6329
rect 29739 6280 29740 6320
rect 29780 6280 29781 6320
rect 29739 6271 29781 6280
rect 30028 5825 30068 6952
rect 30123 6824 30165 6833
rect 30123 6784 30124 6824
rect 30164 6784 30165 6824
rect 30123 6775 30165 6784
rect 30027 5816 30069 5825
rect 30027 5776 30028 5816
rect 30068 5776 30069 5816
rect 30027 5767 30069 5776
rect 30124 5405 30164 6775
rect 30412 6488 30452 7876
rect 30604 7757 30644 7876
rect 30603 7748 30645 7757
rect 30603 7708 30604 7748
rect 30644 7708 30645 7748
rect 30603 7699 30645 7708
rect 30316 6404 30356 6413
rect 30219 6320 30261 6329
rect 30219 6280 30220 6320
rect 30260 6280 30261 6320
rect 30219 6271 30261 6280
rect 30123 5396 30165 5405
rect 30123 5356 30124 5396
rect 30164 5356 30165 5396
rect 30123 5347 30165 5356
rect 30220 5321 30260 6271
rect 30219 5312 30261 5321
rect 30219 5272 30220 5312
rect 30260 5272 30261 5312
rect 30219 5263 30261 5272
rect 29548 5020 29684 5060
rect 29548 4556 29588 5020
rect 29740 4976 29780 4985
rect 29643 4892 29685 4901
rect 29643 4852 29644 4892
rect 29684 4852 29685 4892
rect 29643 4843 29685 4852
rect 29644 4758 29684 4843
rect 29740 4817 29780 4936
rect 30220 4976 30260 5263
rect 30220 4927 30260 4936
rect 30316 4817 30356 6364
rect 30412 4901 30452 6448
rect 30700 5732 30740 8791
rect 30796 8168 30836 8968
rect 30988 8933 31028 9220
rect 30987 8924 31029 8933
rect 30987 8884 30988 8924
rect 31028 8884 31029 8924
rect 30987 8875 31029 8884
rect 30987 8672 31029 8681
rect 30987 8632 30988 8672
rect 31028 8632 31029 8672
rect 30987 8623 31029 8632
rect 30988 8538 31028 8623
rect 30796 8119 30836 8128
rect 30987 8000 31029 8009
rect 30987 7960 30988 8000
rect 31028 7960 31029 8000
rect 30987 7951 31029 7960
rect 30988 7916 31028 7951
rect 30988 7253 31028 7876
rect 30987 7244 31029 7253
rect 30987 7204 30988 7244
rect 31028 7204 31029 7244
rect 30987 7195 31029 7204
rect 30892 6488 30932 6497
rect 30796 6448 30892 6488
rect 30796 6329 30836 6448
rect 30892 6439 30932 6448
rect 30795 6320 30837 6329
rect 31084 6320 31124 9388
rect 31179 9388 31180 9428
rect 31220 9388 31221 9428
rect 31179 9379 31221 9388
rect 31180 8009 31220 9379
rect 31179 8000 31221 8009
rect 31179 7960 31180 8000
rect 31220 7960 31221 8000
rect 31179 7951 31221 7960
rect 30795 6280 30796 6320
rect 30836 6280 30837 6320
rect 30795 6271 30837 6280
rect 30892 6280 31124 6320
rect 31179 6320 31221 6329
rect 31179 6280 31180 6320
rect 31220 6280 31221 6320
rect 30604 5692 30740 5732
rect 30411 4892 30453 4901
rect 30411 4852 30412 4892
rect 30452 4852 30453 4892
rect 30411 4843 30453 4852
rect 29739 4808 29781 4817
rect 29739 4768 29740 4808
rect 29780 4768 29781 4808
rect 29739 4759 29781 4768
rect 30315 4808 30357 4817
rect 30315 4768 30316 4808
rect 30356 4768 30357 4808
rect 30315 4759 30357 4768
rect 29548 4516 29684 4556
rect 29548 2876 29588 2885
rect 29452 2836 29548 2876
rect 29548 2827 29588 2836
rect 29355 2792 29397 2801
rect 29355 2752 29356 2792
rect 29396 2752 29397 2792
rect 29355 2743 29397 2752
rect 29116 2633 29156 2642
rect 29260 2633 29300 2635
rect 29259 2624 29301 2633
rect 29156 2593 29204 2624
rect 29116 2584 29204 2593
rect 28971 2372 29013 2381
rect 28971 2332 28972 2372
rect 29012 2332 29013 2372
rect 28971 2323 29013 2332
rect 29164 2129 29204 2584
rect 29259 2584 29260 2624
rect 29300 2584 29301 2624
rect 29259 2575 29301 2584
rect 29260 2540 29300 2575
rect 29260 2491 29300 2500
rect 29163 2120 29205 2129
rect 29163 2080 29164 2120
rect 29204 2080 29205 2120
rect 29163 2071 29205 2080
rect 29260 1952 29300 1961
rect 29356 1952 29396 2743
rect 29547 2624 29589 2633
rect 29547 2584 29548 2624
rect 29588 2584 29589 2624
rect 29547 2575 29589 2584
rect 29300 1912 29396 1952
rect 29260 1903 29300 1912
rect 29548 1625 29588 2575
rect 29644 2297 29684 4516
rect 30412 4388 30452 4397
rect 30604 4388 30644 5692
rect 30796 5648 30836 5657
rect 30700 5608 30796 5648
rect 30700 5237 30740 5608
rect 30796 5599 30836 5608
rect 30892 5480 30932 6280
rect 31179 6271 31221 6280
rect 31084 5732 31124 5741
rect 30796 5440 30932 5480
rect 30988 5692 31084 5732
rect 30699 5228 30741 5237
rect 30699 5188 30700 5228
rect 30740 5188 30741 5228
rect 30699 5179 30741 5188
rect 30452 4348 30644 4388
rect 30700 4962 30740 4971
rect 30412 4339 30452 4348
rect 30700 4304 30740 4922
rect 30796 4892 30836 5440
rect 30892 5069 30932 5154
rect 30891 5060 30933 5069
rect 30891 5020 30892 5060
rect 30932 5020 30933 5060
rect 30891 5011 30933 5020
rect 30796 4852 30932 4892
rect 30795 4640 30837 4649
rect 30795 4600 30796 4640
rect 30836 4600 30837 4640
rect 30795 4591 30837 4600
rect 30508 4264 30740 4304
rect 30220 4220 30260 4229
rect 30124 4180 30220 4220
rect 30028 4136 30068 4145
rect 29932 4096 30028 4136
rect 29932 3557 29972 4096
rect 30028 4087 30068 4096
rect 30027 3800 30069 3809
rect 30027 3760 30028 3800
rect 30068 3760 30069 3800
rect 30027 3751 30069 3760
rect 29931 3548 29973 3557
rect 29931 3508 29932 3548
rect 29972 3508 29973 3548
rect 29931 3499 29973 3508
rect 29835 3380 29877 3389
rect 29835 3340 29836 3380
rect 29876 3340 29877 3380
rect 29835 3331 29877 3340
rect 29740 2708 29780 2717
rect 29740 2540 29780 2668
rect 29836 2624 29876 3331
rect 29932 3053 29972 3499
rect 29931 3044 29973 3053
rect 29931 3004 29932 3044
rect 29972 3004 29973 3044
rect 29931 2995 29973 3004
rect 30028 2876 30068 3751
rect 30028 2827 30068 2836
rect 29931 2624 29973 2633
rect 29836 2584 29932 2624
rect 29972 2584 29973 2624
rect 29931 2575 29973 2584
rect 29740 2500 29876 2540
rect 29643 2288 29685 2297
rect 29643 2248 29644 2288
rect 29684 2248 29685 2288
rect 29643 2239 29685 2248
rect 29740 1938 29780 1947
rect 29547 1616 29589 1625
rect 29547 1576 29548 1616
rect 29588 1576 29589 1616
rect 29547 1567 29589 1576
rect 29355 1532 29397 1541
rect 29355 1492 29356 1532
rect 29396 1492 29397 1532
rect 29355 1483 29397 1492
rect 27724 1280 27764 1289
rect 27628 1240 27724 1280
rect 27724 1231 27764 1240
rect 27819 1280 27861 1289
rect 27819 1240 27820 1280
rect 27860 1240 27861 1280
rect 27819 1231 27861 1240
rect 28875 1280 28917 1289
rect 28875 1240 28876 1280
rect 28916 1240 28917 1280
rect 28875 1231 28917 1240
rect 28299 1196 28341 1205
rect 28299 1156 28300 1196
rect 28340 1156 28341 1196
rect 28299 1147 28341 1156
rect 27532 1112 27572 1121
rect 27436 1072 27532 1112
rect 27532 1063 27572 1072
rect 28108 1112 28148 1121
rect 28108 869 28148 1072
rect 27339 860 27381 869
rect 27339 820 27340 860
rect 27380 820 27381 860
rect 27339 811 27381 820
rect 28107 860 28149 869
rect 28107 820 28108 860
rect 28148 820 28149 860
rect 28107 811 28149 820
rect 28300 80 28340 1147
rect 29356 1112 29396 1483
rect 29740 1448 29780 1898
rect 29548 1408 29780 1448
rect 29548 1364 29588 1408
rect 29836 1373 29876 2500
rect 30124 2288 30164 4180
rect 30220 4171 30260 4180
rect 30412 3632 30452 3641
rect 30508 3632 30548 4264
rect 30700 4136 30740 4145
rect 30700 3809 30740 4096
rect 30796 4136 30836 4591
rect 30796 4087 30836 4096
rect 30699 3800 30741 3809
rect 30699 3760 30700 3800
rect 30740 3760 30741 3800
rect 30699 3751 30741 3760
rect 30452 3592 30548 3632
rect 30412 3583 30452 3592
rect 30220 3464 30260 3475
rect 30220 3389 30260 3424
rect 30315 3464 30357 3473
rect 30315 3424 30316 3464
rect 30356 3424 30357 3464
rect 30315 3415 30357 3424
rect 30603 3464 30645 3473
rect 30603 3424 30604 3464
rect 30644 3424 30645 3464
rect 30603 3415 30645 3424
rect 30219 3380 30261 3389
rect 30219 3340 30220 3380
rect 30260 3340 30261 3380
rect 30219 3331 30261 3340
rect 30219 3044 30261 3053
rect 30219 3004 30220 3044
rect 30260 3004 30261 3044
rect 30219 2995 30261 3004
rect 30028 2248 30164 2288
rect 30220 2624 30260 2995
rect 29931 2036 29973 2045
rect 29931 1996 29932 2036
rect 29972 1996 29973 2036
rect 29931 1987 29973 1996
rect 29932 1902 29972 1987
rect 29548 1315 29588 1324
rect 29835 1364 29877 1373
rect 29835 1324 29836 1364
rect 29876 1324 29877 1364
rect 29835 1315 29877 1324
rect 29356 1063 29396 1072
rect 29740 1112 29780 1121
rect 29740 869 29780 1072
rect 29739 860 29781 869
rect 29739 820 29740 860
rect 29780 820 29781 860
rect 29739 811 29781 820
rect 30028 113 30068 2248
rect 30123 2120 30165 2129
rect 30123 2080 30124 2120
rect 30164 2080 30165 2120
rect 30123 2071 30165 2080
rect 30124 1986 30164 2071
rect 30220 869 30260 2584
rect 30316 1952 30356 3415
rect 30604 3330 30644 3415
rect 30316 1903 30356 1912
rect 30892 869 30932 4852
rect 30988 2381 31028 5692
rect 31084 5683 31124 5692
rect 31180 5480 31220 6271
rect 31276 5900 31316 9640
rect 31372 9185 31412 10672
rect 31371 9176 31413 9185
rect 31371 9136 31372 9176
rect 31412 9136 31413 9176
rect 31371 9127 31413 9136
rect 31564 9008 31604 10672
rect 31756 9176 31796 10672
rect 31851 9596 31893 9605
rect 31851 9556 31852 9596
rect 31892 9556 31893 9596
rect 31851 9547 31893 9556
rect 31852 9344 31892 9547
rect 31948 9428 31988 10672
rect 32140 9512 32180 10672
rect 32332 9689 32372 10672
rect 32331 9680 32373 9689
rect 32331 9640 32332 9680
rect 32372 9640 32373 9680
rect 32331 9631 32373 9640
rect 32428 9512 32468 9521
rect 32140 9472 32372 9512
rect 31948 9388 32276 9428
rect 31852 9304 31988 9344
rect 31756 9136 31892 9176
rect 31564 8968 31796 9008
rect 31756 8924 31796 8968
rect 31852 8933 31892 9136
rect 31851 8924 31893 8933
rect 31756 8884 31799 8924
rect 31759 8840 31799 8884
rect 31851 8884 31852 8924
rect 31892 8884 31893 8924
rect 31851 8875 31893 8884
rect 31756 8800 31799 8840
rect 31468 8756 31508 8765
rect 31372 8716 31468 8756
rect 31372 8597 31412 8716
rect 31468 8707 31508 8716
rect 31563 8672 31605 8681
rect 31563 8632 31564 8672
rect 31604 8632 31605 8672
rect 31563 8623 31605 8632
rect 31371 8588 31413 8597
rect 31371 8548 31372 8588
rect 31412 8548 31413 8588
rect 31371 8539 31413 8548
rect 31372 7505 31412 8539
rect 31564 8261 31604 8623
rect 31659 8420 31701 8429
rect 31659 8380 31660 8420
rect 31700 8380 31701 8420
rect 31659 8371 31701 8380
rect 31563 8252 31605 8261
rect 31563 8212 31564 8252
rect 31604 8212 31605 8252
rect 31563 8203 31605 8212
rect 31468 8000 31508 8009
rect 31371 7496 31413 7505
rect 31371 7456 31372 7496
rect 31412 7456 31413 7496
rect 31371 7447 31413 7456
rect 31468 7421 31508 7960
rect 31564 8000 31604 8009
rect 31660 8000 31700 8371
rect 31604 7960 31700 8000
rect 31564 7951 31604 7960
rect 31467 7412 31509 7421
rect 31467 7372 31468 7412
rect 31508 7372 31509 7412
rect 31467 7363 31509 7372
rect 31467 7244 31509 7253
rect 31467 7204 31468 7244
rect 31508 7204 31509 7244
rect 31467 7195 31509 7204
rect 31468 7160 31508 7195
rect 31468 7109 31508 7120
rect 31660 6992 31700 7001
rect 31468 6952 31660 6992
rect 31468 6488 31508 6952
rect 31660 6943 31700 6952
rect 31659 6740 31701 6749
rect 31659 6700 31660 6740
rect 31700 6700 31701 6740
rect 31659 6691 31701 6700
rect 31563 6656 31605 6665
rect 31563 6616 31564 6656
rect 31604 6616 31605 6656
rect 31563 6607 31605 6616
rect 31564 6522 31604 6607
rect 31420 6478 31508 6488
rect 31460 6448 31508 6478
rect 31420 6429 31460 6438
rect 31660 5900 31700 6691
rect 31756 6572 31796 8800
rect 31948 8756 31988 9304
rect 32043 9260 32085 9269
rect 32043 9220 32044 9260
rect 32084 9220 32085 9260
rect 32043 9211 32085 9220
rect 31852 8716 31988 8756
rect 31852 7673 31892 8716
rect 32044 8672 32084 9211
rect 32139 9092 32181 9101
rect 32139 9052 32140 9092
rect 32180 9052 32181 9092
rect 32139 9043 32181 9052
rect 31948 8652 31988 8661
rect 32044 8623 32084 8632
rect 31948 8177 31988 8612
rect 32043 8504 32085 8513
rect 32043 8464 32044 8504
rect 32084 8464 32085 8504
rect 32043 8455 32085 8464
rect 31947 8168 31989 8177
rect 31947 8128 31948 8168
rect 31988 8128 31989 8168
rect 31947 8119 31989 8128
rect 31947 8000 31989 8009
rect 31947 7960 31948 8000
rect 31988 7960 31989 8000
rect 31947 7951 31989 7960
rect 32044 8000 32084 8455
rect 32044 7951 32084 7960
rect 31948 7866 31988 7951
rect 32043 7748 32085 7757
rect 32043 7708 32044 7748
rect 32084 7708 32085 7748
rect 32043 7699 32085 7708
rect 31851 7664 31893 7673
rect 31851 7624 31852 7664
rect 31892 7624 31893 7664
rect 31851 7615 31893 7624
rect 31947 7496 31989 7505
rect 31947 7456 31948 7496
rect 31988 7456 31989 7496
rect 31947 7447 31989 7456
rect 31851 7412 31893 7421
rect 31851 7372 31852 7412
rect 31892 7372 31893 7412
rect 31851 7363 31893 7372
rect 31852 7278 31892 7363
rect 31948 6992 31988 7447
rect 32044 7421 32084 7699
rect 32043 7412 32085 7421
rect 32043 7372 32044 7412
rect 32084 7372 32085 7412
rect 32043 7363 32085 7372
rect 32044 7160 32084 7363
rect 32044 7111 32084 7120
rect 31948 6952 32084 6992
rect 31947 6656 31989 6665
rect 31947 6616 31948 6656
rect 31988 6616 31989 6656
rect 31947 6607 31989 6616
rect 31756 6532 31892 6572
rect 31276 5860 31604 5900
rect 31468 5732 31508 5741
rect 31372 5692 31468 5732
rect 31276 5480 31316 5489
rect 31180 5440 31276 5480
rect 31276 5431 31316 5440
rect 31083 5396 31125 5405
rect 31083 5356 31084 5396
rect 31124 5356 31125 5396
rect 31083 5347 31125 5356
rect 30987 2372 31029 2381
rect 30987 2332 30988 2372
rect 31028 2332 31029 2372
rect 30987 2323 31029 2332
rect 30987 1112 31029 1121
rect 30987 1072 30988 1112
rect 31028 1072 31029 1112
rect 30987 1063 31029 1072
rect 30988 978 31028 1063
rect 30219 860 30261 869
rect 30219 820 30220 860
rect 30260 820 30261 860
rect 30219 811 30261 820
rect 30891 860 30933 869
rect 30891 820 30892 860
rect 30932 820 30933 860
rect 30891 811 30933 820
rect 29451 104 29493 113
rect 29451 80 29452 104
rect 22348 64 22600 80
rect 22348 60 22388 64
rect 22156 20 22388 60
rect 22520 0 22600 64
rect 23672 0 23752 80
rect 24824 0 24904 80
rect 25976 0 26056 80
rect 27128 0 27208 80
rect 28280 0 28360 80
rect 29432 64 29452 80
rect 29492 80 29493 104
rect 30027 104 30069 113
rect 29492 64 29512 80
rect 29432 0 29512 64
rect 30027 64 30028 104
rect 30068 64 30069 104
rect 30603 104 30645 113
rect 30603 80 30604 104
rect 30027 55 30069 64
rect 30584 64 30604 80
rect 30644 80 30645 104
rect 30795 104 30837 113
rect 30644 64 30664 80
rect 30584 0 30664 64
rect 30795 64 30796 104
rect 30836 64 30837 104
rect 30795 60 30837 64
rect 31084 60 31124 5347
rect 31179 5312 31221 5321
rect 31179 5272 31180 5312
rect 31220 5272 31221 5312
rect 31179 5263 31221 5272
rect 31180 4724 31220 5263
rect 31275 4976 31317 4985
rect 31275 4936 31276 4976
rect 31316 4936 31317 4976
rect 31275 4927 31317 4936
rect 31276 4842 31316 4927
rect 31180 4684 31316 4724
rect 31276 4220 31316 4684
rect 31276 4171 31316 4180
rect 31180 4136 31220 4145
rect 31180 3893 31220 4096
rect 31179 3884 31221 3893
rect 31179 3844 31180 3884
rect 31220 3844 31221 3884
rect 31179 3835 31221 3844
rect 31372 1793 31412 5692
rect 31468 5683 31508 5692
rect 31564 5564 31604 5860
rect 31660 5851 31700 5860
rect 31756 6404 31796 6413
rect 31468 5524 31604 5564
rect 31468 3809 31508 5524
rect 31756 4304 31796 6364
rect 31852 6152 31892 6532
rect 31948 6522 31988 6607
rect 31852 6112 31988 6152
rect 31851 5984 31893 5993
rect 31851 5944 31852 5984
rect 31892 5944 31893 5984
rect 31851 5935 31893 5944
rect 31852 5648 31892 5935
rect 31852 5599 31892 5608
rect 31564 4264 31796 4304
rect 31467 3800 31509 3809
rect 31467 3760 31468 3800
rect 31508 3760 31509 3800
rect 31467 3751 31509 3760
rect 31467 3296 31509 3305
rect 31467 3256 31468 3296
rect 31508 3256 31509 3296
rect 31467 3247 31509 3256
rect 31468 2885 31508 3247
rect 31467 2876 31509 2885
rect 31467 2836 31468 2876
rect 31508 2836 31509 2876
rect 31467 2827 31509 2836
rect 31468 2624 31508 2827
rect 31564 2633 31604 4264
rect 31756 4136 31796 4147
rect 31756 4061 31796 4096
rect 31755 4052 31797 4061
rect 31755 4012 31756 4052
rect 31796 4012 31797 4052
rect 31755 4003 31797 4012
rect 31659 3800 31701 3809
rect 31659 3760 31660 3800
rect 31700 3760 31701 3800
rect 31659 3751 31701 3760
rect 31660 2876 31700 3751
rect 31852 3464 31892 3473
rect 31852 3305 31892 3424
rect 31851 3296 31893 3305
rect 31851 3256 31852 3296
rect 31892 3256 31893 3296
rect 31851 3247 31893 3256
rect 31948 2876 31988 6112
rect 32044 4649 32084 6952
rect 32140 6749 32180 9043
rect 32236 7832 32276 9388
rect 32332 8672 32372 9472
rect 32428 8849 32468 9472
rect 32524 9017 32564 10672
rect 32619 9260 32661 9269
rect 32619 9220 32620 9260
rect 32660 9220 32661 9260
rect 32619 9211 32661 9220
rect 32620 9126 32660 9211
rect 32523 9008 32565 9017
rect 32523 8968 32524 9008
rect 32564 8968 32565 9008
rect 32523 8959 32565 8968
rect 32716 8849 32756 10672
rect 32811 9680 32853 9689
rect 32811 9640 32812 9680
rect 32852 9640 32853 9680
rect 32811 9631 32853 9640
rect 32812 9512 32852 9631
rect 32812 9463 32852 9472
rect 32908 8924 32948 10672
rect 33100 9017 33140 10672
rect 33292 9428 33332 10672
rect 33196 9388 33332 9428
rect 33196 9101 33236 9388
rect 33291 9260 33333 9269
rect 33291 9220 33292 9260
rect 33332 9220 33333 9260
rect 33291 9211 33333 9220
rect 33195 9092 33237 9101
rect 33195 9052 33196 9092
rect 33236 9052 33237 9092
rect 33195 9043 33237 9052
rect 33099 9008 33141 9017
rect 33099 8968 33100 9008
rect 33140 8968 33141 9008
rect 33099 8959 33141 8968
rect 32812 8884 32948 8924
rect 32427 8840 32469 8849
rect 32427 8800 32428 8840
rect 32468 8800 32469 8840
rect 32427 8791 32469 8800
rect 32715 8840 32757 8849
rect 32715 8800 32716 8840
rect 32756 8800 32757 8840
rect 32715 8791 32757 8800
rect 32524 8756 32564 8765
rect 32332 8632 32468 8672
rect 32332 8504 32372 8513
rect 32332 8345 32372 8464
rect 32331 8336 32373 8345
rect 32331 8296 32332 8336
rect 32372 8296 32373 8336
rect 32331 8287 32373 8296
rect 32428 7916 32468 8632
rect 32524 8429 32564 8716
rect 32715 8504 32757 8513
rect 32715 8464 32716 8504
rect 32756 8464 32757 8504
rect 32715 8455 32757 8464
rect 32523 8420 32565 8429
rect 32523 8380 32524 8420
rect 32564 8380 32565 8420
rect 32523 8371 32565 8380
rect 32716 8370 32756 8455
rect 32619 8336 32661 8345
rect 32619 8296 32620 8336
rect 32660 8296 32661 8336
rect 32619 8287 32661 8296
rect 32523 8252 32565 8261
rect 32523 8212 32524 8252
rect 32564 8212 32565 8252
rect 32523 8203 32565 8212
rect 32524 8093 32564 8203
rect 32523 8084 32565 8093
rect 32523 8044 32524 8084
rect 32564 8044 32565 8084
rect 32523 8035 32565 8044
rect 32524 8009 32564 8035
rect 32524 7960 32564 7969
rect 32620 8000 32660 8287
rect 32620 7960 32756 8000
rect 32428 7876 32660 7916
rect 32236 7792 32564 7832
rect 32235 7664 32277 7673
rect 32235 7624 32236 7664
rect 32276 7624 32277 7664
rect 32235 7615 32277 7624
rect 32427 7664 32469 7673
rect 32427 7624 32428 7664
rect 32468 7624 32469 7664
rect 32427 7615 32469 7624
rect 32139 6740 32181 6749
rect 32139 6700 32140 6740
rect 32180 6700 32181 6740
rect 32139 6691 32181 6700
rect 32139 6404 32181 6413
rect 32139 6364 32140 6404
rect 32180 6364 32181 6404
rect 32139 6355 32181 6364
rect 32140 6270 32180 6355
rect 32043 4640 32085 4649
rect 32043 4600 32044 4640
rect 32084 4600 32085 4640
rect 32043 4591 32085 4600
rect 32236 4304 32276 7615
rect 32332 6236 32372 6245
rect 32332 4481 32372 6196
rect 32428 5405 32468 7615
rect 32524 6656 32564 7792
rect 32524 6607 32564 6616
rect 32523 5648 32565 5657
rect 32523 5608 32524 5648
rect 32564 5608 32565 5648
rect 32523 5599 32565 5608
rect 32427 5396 32469 5405
rect 32427 5356 32428 5396
rect 32468 5356 32469 5396
rect 32427 5347 32469 5356
rect 32524 4976 32564 5599
rect 32524 4927 32564 4936
rect 32427 4892 32469 4901
rect 32427 4852 32428 4892
rect 32468 4852 32469 4892
rect 32427 4843 32469 4852
rect 32331 4472 32373 4481
rect 32331 4432 32332 4472
rect 32372 4432 32373 4472
rect 32331 4423 32373 4432
rect 32236 4264 32372 4304
rect 32236 4141 32276 4150
rect 32236 3716 32276 4101
rect 32044 3676 32276 3716
rect 32044 3632 32084 3676
rect 32044 3583 32084 3592
rect 32235 3464 32277 3473
rect 32235 3424 32236 3464
rect 32276 3424 32277 3464
rect 32235 3415 32277 3424
rect 32236 3053 32276 3415
rect 32235 3044 32277 3053
rect 32235 3004 32236 3044
rect 32276 3004 32277 3044
rect 32235 2995 32277 3004
rect 32044 2876 32084 2885
rect 31948 2836 32044 2876
rect 31660 2827 31700 2836
rect 32044 2827 32084 2836
rect 31852 2708 31892 2717
rect 31468 2575 31508 2584
rect 31563 2624 31605 2633
rect 31563 2584 31564 2624
rect 31604 2584 31605 2624
rect 31563 2575 31605 2584
rect 31755 2288 31797 2297
rect 31755 2248 31756 2288
rect 31796 2248 31797 2288
rect 31755 2239 31797 2248
rect 31564 2045 31604 2076
rect 31563 2036 31605 2045
rect 31563 1996 31564 2036
rect 31604 1996 31605 2036
rect 31563 1987 31605 1996
rect 31564 1952 31604 1987
rect 31371 1784 31413 1793
rect 31371 1744 31372 1784
rect 31412 1744 31413 1784
rect 31371 1735 31413 1744
rect 31564 1541 31604 1912
rect 31756 1952 31796 2239
rect 31756 1903 31796 1912
rect 31755 1700 31797 1709
rect 31755 1660 31756 1700
rect 31796 1660 31797 1700
rect 31755 1651 31797 1660
rect 31563 1532 31605 1541
rect 31563 1492 31564 1532
rect 31604 1492 31605 1532
rect 31563 1483 31605 1492
rect 31563 1364 31605 1373
rect 31563 1324 31564 1364
rect 31604 1324 31605 1364
rect 31563 1315 31605 1324
rect 31275 1280 31317 1289
rect 31275 1240 31276 1280
rect 31316 1240 31317 1280
rect 31275 1231 31317 1240
rect 31467 1280 31509 1289
rect 31467 1240 31468 1280
rect 31508 1240 31509 1280
rect 31467 1231 31509 1240
rect 31276 1112 31316 1231
rect 31276 1063 31316 1072
rect 31468 869 31508 1231
rect 31564 1230 31604 1315
rect 31467 860 31509 869
rect 31467 820 31468 860
rect 31508 820 31509 860
rect 31467 811 31509 820
rect 31756 80 31796 1651
rect 31852 1037 31892 2668
rect 32236 2708 32276 2717
rect 32236 1205 32276 2668
rect 32332 1280 32372 4264
rect 32428 4052 32468 4843
rect 32523 4640 32565 4649
rect 32523 4600 32524 4640
rect 32564 4600 32565 4640
rect 32523 4591 32565 4600
rect 32428 4003 32468 4012
rect 32524 1877 32564 4591
rect 32620 3641 32660 7876
rect 32716 6833 32756 7960
rect 32715 6824 32757 6833
rect 32715 6784 32716 6824
rect 32756 6784 32757 6824
rect 32715 6775 32757 6784
rect 32716 6404 32756 6413
rect 32716 5321 32756 6364
rect 32812 6245 32852 8884
rect 32908 8756 32948 8765
rect 32948 8716 33236 8756
rect 32908 8707 32948 8716
rect 33196 8168 33236 8716
rect 33292 8672 33332 9211
rect 33292 8623 33332 8632
rect 33388 8672 33428 8683
rect 33388 8597 33428 8632
rect 33387 8588 33429 8597
rect 33387 8548 33388 8588
rect 33428 8548 33429 8588
rect 33387 8539 33429 8548
rect 33196 8119 33236 8128
rect 33484 8084 33524 10672
rect 39627 10648 39628 10688
rect 39668 10648 39669 10688
rect 39627 10639 39669 10648
rect 35883 10604 35925 10613
rect 35883 10564 35884 10604
rect 35924 10564 35925 10604
rect 35883 10555 35925 10564
rect 34923 10520 34965 10529
rect 34923 10480 34924 10520
rect 34964 10480 34965 10520
rect 34923 10471 34965 10480
rect 34443 9680 34485 9689
rect 34443 9640 34444 9680
rect 34484 9640 34485 9680
rect 34443 9631 34485 9640
rect 34059 9512 34101 9521
rect 34059 9472 34060 9512
rect 34100 9472 34101 9512
rect 34059 9463 34101 9472
rect 34444 9512 34484 9631
rect 34444 9463 34484 9472
rect 34060 9378 34100 9463
rect 34252 9260 34292 9269
rect 34292 9220 34868 9260
rect 34252 9211 34292 9220
rect 33928 9092 34296 9101
rect 33968 9052 34010 9092
rect 34050 9052 34092 9092
rect 34132 9052 34174 9092
rect 34214 9052 34256 9092
rect 33928 9043 34296 9052
rect 34443 9092 34485 9101
rect 34443 9052 34444 9092
rect 34484 9052 34485 9092
rect 34443 9043 34485 9052
rect 33771 8672 33813 8681
rect 33771 8632 33772 8672
rect 33812 8632 33813 8672
rect 33771 8623 33813 8632
rect 33868 8672 33908 8681
rect 33772 8538 33812 8623
rect 33868 8597 33908 8632
rect 34347 8672 34389 8681
rect 34347 8632 34348 8672
rect 34388 8632 34389 8672
rect 34347 8623 34389 8632
rect 33867 8588 33909 8597
rect 33867 8548 33868 8588
rect 33908 8548 33909 8588
rect 33867 8539 33909 8548
rect 33868 8093 33908 8539
rect 34348 8261 34388 8623
rect 34347 8252 34389 8261
rect 34347 8212 34348 8252
rect 34388 8212 34389 8252
rect 34347 8203 34389 8212
rect 34059 8168 34101 8177
rect 34059 8128 34060 8168
rect 34100 8128 34101 8168
rect 34059 8119 34101 8128
rect 33867 8084 33909 8093
rect 33484 8044 33812 8084
rect 33052 7990 33524 8000
rect 33092 7960 33524 7990
rect 33052 7941 33092 7950
rect 33291 7664 33333 7673
rect 33291 7624 33292 7664
rect 33332 7624 33333 7664
rect 33291 7615 33333 7624
rect 33195 7412 33237 7421
rect 33195 7372 33196 7412
rect 33236 7372 33237 7412
rect 33195 7363 33237 7372
rect 32907 6908 32949 6917
rect 32907 6868 32908 6908
rect 32948 6868 32949 6908
rect 32907 6859 32949 6868
rect 32908 6413 32948 6859
rect 33099 6572 33141 6581
rect 33099 6532 33100 6572
rect 33140 6532 33141 6572
rect 33099 6523 33141 6532
rect 33004 6488 33044 6497
rect 32907 6404 32949 6413
rect 32907 6364 32908 6404
rect 32948 6364 32949 6404
rect 32907 6355 32949 6364
rect 32811 6236 32853 6245
rect 32811 6196 32812 6236
rect 32852 6196 32853 6236
rect 32811 6187 32853 6196
rect 32811 5648 32853 5657
rect 32811 5608 32812 5648
rect 32852 5608 32853 5648
rect 32811 5599 32853 5608
rect 32715 5312 32757 5321
rect 32715 5272 32716 5312
rect 32756 5272 32757 5312
rect 32715 5263 32757 5272
rect 32716 4724 32756 4733
rect 32716 4136 32756 4684
rect 32812 4304 32852 5599
rect 32908 4892 32948 6355
rect 33004 5396 33044 6448
rect 33100 6488 33140 6523
rect 33100 6437 33140 6448
rect 33196 5657 33236 7363
rect 33292 7160 33332 7615
rect 33484 7412 33524 7960
rect 33675 7832 33717 7841
rect 33675 7792 33676 7832
rect 33716 7792 33717 7832
rect 33675 7783 33717 7792
rect 33579 7748 33621 7757
rect 33579 7708 33580 7748
rect 33620 7708 33621 7748
rect 33579 7699 33621 7708
rect 33484 7363 33524 7372
rect 33292 7111 33332 7120
rect 33580 6488 33620 7699
rect 33676 7698 33716 7783
rect 33675 7412 33717 7421
rect 33675 7372 33676 7412
rect 33716 7372 33717 7412
rect 33675 7363 33717 7372
rect 33676 7160 33716 7363
rect 33676 7111 33716 7120
rect 33675 6656 33717 6665
rect 33675 6616 33676 6656
rect 33716 6616 33717 6656
rect 33675 6607 33717 6616
rect 33580 6439 33620 6448
rect 33484 6404 33524 6413
rect 33388 6364 33484 6404
rect 33100 5648 33140 5657
rect 33195 5648 33237 5657
rect 33140 5608 33196 5648
rect 33236 5608 33237 5648
rect 33100 5599 33140 5608
rect 33195 5599 33237 5608
rect 33196 5514 33236 5599
rect 33292 5480 33332 5489
rect 33292 5396 33332 5440
rect 33004 5356 33332 5396
rect 33292 4976 33332 4985
rect 33099 4892 33141 4901
rect 32908 4852 33044 4892
rect 32907 4724 32949 4733
rect 32907 4684 32908 4724
rect 32948 4684 32949 4724
rect 32907 4675 32949 4684
rect 32908 4590 32948 4675
rect 32812 4264 32948 4304
rect 32716 4087 32756 4096
rect 32811 4136 32853 4145
rect 32811 4096 32812 4136
rect 32852 4096 32853 4136
rect 32811 4087 32853 4096
rect 32812 4002 32852 4087
rect 32619 3632 32661 3641
rect 32619 3592 32620 3632
rect 32660 3592 32661 3632
rect 32619 3583 32661 3592
rect 32908 3473 32948 4264
rect 32907 3464 32949 3473
rect 32907 3424 32908 3464
rect 32948 3424 32949 3464
rect 32907 3415 32949 3424
rect 32812 2624 32852 2633
rect 32812 2297 32852 2584
rect 32908 2624 32948 2633
rect 33004 2624 33044 4852
rect 33099 4852 33100 4892
rect 33140 4852 33141 4892
rect 33099 4843 33141 4852
rect 33100 4758 33140 4843
rect 33292 4472 33332 4936
rect 33100 4432 33332 4472
rect 33100 3725 33140 4432
rect 33195 4304 33237 4313
rect 33195 4264 33196 4304
rect 33236 4264 33237 4304
rect 33195 4255 33237 4264
rect 33196 4136 33236 4255
rect 33291 4220 33333 4229
rect 33291 4180 33292 4220
rect 33332 4180 33333 4220
rect 33291 4171 33333 4180
rect 33196 3893 33236 4096
rect 33292 4086 33332 4171
rect 33195 3884 33237 3893
rect 33195 3844 33196 3884
rect 33236 3844 33237 3884
rect 33195 3835 33237 3844
rect 33099 3716 33141 3725
rect 33099 3676 33100 3716
rect 33140 3676 33141 3716
rect 33099 3667 33141 3676
rect 33099 3380 33141 3389
rect 33099 3340 33100 3380
rect 33140 3340 33141 3380
rect 33099 3331 33141 3340
rect 32948 2584 33044 2624
rect 32908 2575 32948 2584
rect 33100 2540 33140 3331
rect 33291 2708 33333 2717
rect 33291 2668 33292 2708
rect 33332 2668 33333 2708
rect 33291 2659 33333 2668
rect 33388 2708 33428 6364
rect 33484 6355 33524 6364
rect 33579 6236 33621 6245
rect 33579 6196 33580 6236
rect 33620 6196 33621 6236
rect 33579 6187 33621 6196
rect 33484 5648 33524 5657
rect 33484 5153 33524 5608
rect 33483 5144 33525 5153
rect 33483 5104 33484 5144
rect 33524 5104 33525 5144
rect 33483 5095 33525 5104
rect 33483 3464 33525 3473
rect 33483 3424 33484 3464
rect 33524 3424 33525 3464
rect 33483 3415 33525 3424
rect 33484 3330 33524 3415
rect 33292 2574 33332 2659
rect 33004 2500 33140 2540
rect 32811 2288 32853 2297
rect 32811 2248 32812 2288
rect 32852 2248 32853 2288
rect 32811 2239 32853 2248
rect 33004 1952 33044 2500
rect 33195 2288 33237 2297
rect 33195 2248 33196 2288
rect 33236 2248 33237 2288
rect 33195 2239 33237 2248
rect 33196 2120 33236 2239
rect 33388 2129 33428 2668
rect 33196 2071 33236 2080
rect 33387 2120 33429 2129
rect 33387 2080 33388 2120
rect 33428 2080 33429 2120
rect 33387 2071 33429 2080
rect 33388 1961 33428 2071
rect 33004 1903 33044 1912
rect 33387 1952 33429 1961
rect 33387 1912 33388 1952
rect 33428 1912 33429 1952
rect 33387 1903 33429 1912
rect 32523 1868 32565 1877
rect 32523 1828 32524 1868
rect 32564 1828 32565 1868
rect 32523 1819 32565 1828
rect 32907 1868 32949 1877
rect 32907 1828 32908 1868
rect 32948 1828 32949 1868
rect 32907 1819 32949 1828
rect 32428 1280 32468 1289
rect 32332 1240 32428 1280
rect 32428 1231 32468 1240
rect 32811 1280 32853 1289
rect 32811 1240 32812 1280
rect 32852 1240 32853 1280
rect 32811 1231 32853 1240
rect 32235 1196 32277 1205
rect 32235 1156 32236 1196
rect 32276 1156 32277 1196
rect 32235 1147 32277 1156
rect 32620 1196 32660 1205
rect 31851 1028 31893 1037
rect 31851 988 31852 1028
rect 31892 988 31893 1028
rect 31851 979 31893 988
rect 32620 281 32660 1156
rect 32812 1146 32852 1231
rect 32619 272 32661 281
rect 32619 232 32620 272
rect 32660 232 32661 272
rect 32619 223 32661 232
rect 32908 80 32948 1819
rect 33004 1196 33044 1205
rect 33004 197 33044 1156
rect 33387 1112 33429 1121
rect 33387 1072 33388 1112
rect 33428 1072 33429 1112
rect 33387 1063 33429 1072
rect 33388 978 33428 1063
rect 33580 1037 33620 6187
rect 33676 3977 33716 6607
rect 33772 6329 33812 8044
rect 33867 8044 33868 8084
rect 33908 8044 33909 8084
rect 33867 8035 33909 8044
rect 34060 8000 34100 8119
rect 34060 7951 34100 7960
rect 33867 7916 33909 7925
rect 33867 7876 33868 7916
rect 33908 7876 33909 7916
rect 33867 7867 33909 7876
rect 33868 7782 33908 7867
rect 33928 7580 34296 7589
rect 33968 7540 34010 7580
rect 34050 7540 34092 7580
rect 34132 7540 34174 7580
rect 34214 7540 34256 7580
rect 33928 7531 34296 7540
rect 34060 6488 34100 6497
rect 33771 6320 33813 6329
rect 33771 6280 33772 6320
rect 33812 6280 33813 6320
rect 33771 6271 33813 6280
rect 34060 6236 34100 6448
rect 34444 6320 34484 9043
rect 34731 8756 34773 8765
rect 34731 8716 34732 8756
rect 34772 8716 34773 8756
rect 34731 8707 34773 8716
rect 34732 6656 34772 8707
rect 34828 8686 34868 9220
rect 34828 8637 34868 8646
rect 34924 7664 34964 10471
rect 35168 9848 35536 9857
rect 35208 9808 35250 9848
rect 35290 9808 35332 9848
rect 35372 9808 35414 9848
rect 35454 9808 35496 9848
rect 35168 9799 35536 9808
rect 35691 9764 35733 9773
rect 35691 9724 35692 9764
rect 35732 9724 35733 9764
rect 35691 9715 35733 9724
rect 35692 9512 35732 9715
rect 35692 9437 35732 9472
rect 35691 9428 35733 9437
rect 35691 9388 35692 9428
rect 35732 9388 35733 9428
rect 35691 9379 35733 9388
rect 35884 9017 35924 10555
rect 37611 10520 37653 10529
rect 37611 10480 37612 10520
rect 37652 10480 37653 10520
rect 37611 10471 37653 10480
rect 35979 9680 36021 9689
rect 35979 9640 35980 9680
rect 36020 9640 36021 9680
rect 35979 9631 36021 9640
rect 37323 9680 37365 9689
rect 37323 9640 37324 9680
rect 37364 9640 37365 9680
rect 37323 9631 37365 9640
rect 35595 9008 35637 9017
rect 35595 8968 35596 9008
rect 35636 8968 35637 9008
rect 35595 8959 35637 8968
rect 35883 9008 35925 9017
rect 35883 8968 35884 9008
rect 35924 8968 35925 9008
rect 35883 8959 35925 8968
rect 35403 8756 35445 8765
rect 35403 8716 35404 8756
rect 35444 8716 35445 8756
rect 35403 8707 35445 8716
rect 35404 8622 35444 8707
rect 35212 8513 35252 8598
rect 35020 8504 35060 8513
rect 35020 7925 35060 8464
rect 35211 8504 35253 8513
rect 35211 8464 35212 8504
rect 35252 8464 35253 8504
rect 35211 8455 35253 8464
rect 35168 8336 35536 8345
rect 35208 8296 35250 8336
rect 35290 8296 35332 8336
rect 35372 8296 35414 8336
rect 35454 8296 35496 8336
rect 35168 8287 35536 8296
rect 35596 8168 35636 8959
rect 35788 8672 35828 8681
rect 35404 8128 35636 8168
rect 35692 8168 35732 8177
rect 35788 8168 35828 8632
rect 35884 8672 35924 8959
rect 35884 8623 35924 8632
rect 35732 8128 35828 8168
rect 35307 8000 35349 8009
rect 35307 7960 35308 8000
rect 35348 7960 35349 8000
rect 35307 7951 35349 7960
rect 35019 7916 35061 7925
rect 35019 7876 35020 7916
rect 35060 7876 35061 7916
rect 35019 7867 35061 7876
rect 35019 7748 35061 7757
rect 35019 7708 35020 7748
rect 35060 7708 35061 7748
rect 35019 7699 35061 7708
rect 34828 7624 34964 7664
rect 34828 6665 34868 7624
rect 34923 7496 34965 7505
rect 34923 7456 34924 7496
rect 34964 7456 34965 7496
rect 34923 7447 34965 7456
rect 34924 7169 34964 7447
rect 34923 7160 34965 7169
rect 34923 7120 34924 7160
rect 34964 7120 34965 7160
rect 34923 7111 34965 7120
rect 34924 7026 34964 7111
rect 34732 6607 34772 6616
rect 34827 6656 34869 6665
rect 34827 6616 34828 6656
rect 34868 6616 34869 6656
rect 34827 6607 34869 6616
rect 35020 6488 35060 7699
rect 35308 7421 35348 7951
rect 35307 7412 35349 7421
rect 35307 7372 35308 7412
rect 35348 7372 35349 7412
rect 35307 7363 35349 7372
rect 35404 7412 35444 8128
rect 35692 8119 35732 8128
rect 35883 8000 35925 8009
rect 35980 8000 36020 9631
rect 36076 9512 36116 9521
rect 36076 9353 36116 9472
rect 37324 9512 37364 9631
rect 37324 9463 37364 9472
rect 36075 9344 36117 9353
rect 36075 9304 36076 9344
rect 36116 9304 36117 9344
rect 36075 9295 36117 9304
rect 37227 9344 37269 9353
rect 37227 9304 37228 9344
rect 37268 9304 37269 9344
rect 37227 9295 37269 9304
rect 36076 9101 36116 9295
rect 36075 9092 36117 9101
rect 36075 9052 36076 9092
rect 36116 9052 36117 9092
rect 36075 9043 36117 9052
rect 36844 8765 36884 8796
rect 36843 8756 36885 8765
rect 36843 8716 36844 8756
rect 36884 8716 36885 8756
rect 36843 8707 36885 8716
rect 35883 7960 35884 8000
rect 35924 7960 36020 8000
rect 36268 8672 36308 8681
rect 35883 7951 35925 7960
rect 35884 7866 35924 7951
rect 35499 7748 35541 7757
rect 35499 7708 35500 7748
rect 35540 7708 35541 7748
rect 35499 7699 35541 7708
rect 35500 7614 35540 7699
rect 36268 7673 36308 8632
rect 36364 8672 36404 8683
rect 36364 8597 36404 8632
rect 36844 8672 36884 8707
rect 36363 8588 36405 8597
rect 36363 8548 36364 8588
rect 36404 8548 36405 8588
rect 36363 8539 36405 8548
rect 36267 7664 36309 7673
rect 36267 7624 36268 7664
rect 36308 7624 36309 7664
rect 36267 7615 36309 7624
rect 35404 7363 35444 7372
rect 35596 7244 35636 7253
rect 35787 7244 35829 7253
rect 35636 7204 35732 7244
rect 35596 7195 35636 7204
rect 35168 6824 35536 6833
rect 35208 6784 35250 6824
rect 35290 6784 35332 6824
rect 35372 6784 35414 6824
rect 35454 6784 35496 6824
rect 35168 6775 35536 6784
rect 35211 6656 35253 6665
rect 35211 6616 35212 6656
rect 35252 6616 35253 6656
rect 35211 6607 35253 6616
rect 35116 6488 35156 6497
rect 34588 6446 34628 6455
rect 35020 6448 35116 6488
rect 35116 6439 35156 6448
rect 35212 6488 35252 6607
rect 35692 6572 35732 7204
rect 35787 7204 35788 7244
rect 35828 7204 35829 7244
rect 35787 7195 35829 7204
rect 36364 7244 36404 7253
rect 35788 7110 35828 7195
rect 36267 7076 36309 7085
rect 36267 7036 36268 7076
rect 36308 7036 36309 7076
rect 36267 7027 36309 7036
rect 35883 6992 35925 7001
rect 35883 6952 35884 6992
rect 35924 6952 35925 6992
rect 35883 6943 35925 6952
rect 35980 6992 36020 7001
rect 35692 6532 35828 6572
rect 35596 6488 35636 6497
rect 35212 6439 35252 6448
rect 35500 6448 35596 6488
rect 34588 6404 34628 6406
rect 34588 6364 34964 6404
rect 34444 6280 34868 6320
rect 34060 6196 34676 6236
rect 33928 6068 34296 6077
rect 33968 6028 34010 6068
rect 34050 6028 34092 6068
rect 34132 6028 34174 6068
rect 34214 6028 34256 6068
rect 33928 6019 34296 6028
rect 34539 5648 34581 5657
rect 34539 5608 34540 5648
rect 34580 5608 34581 5648
rect 34539 5599 34581 5608
rect 34540 4976 34580 5599
rect 34540 4927 34580 4936
rect 34347 4724 34389 4733
rect 34347 4684 34348 4724
rect 34388 4684 34389 4724
rect 34347 4675 34389 4684
rect 33928 4556 34296 4565
rect 33968 4516 34010 4556
rect 34050 4516 34092 4556
rect 34132 4516 34174 4556
rect 34214 4516 34256 4556
rect 33928 4507 34296 4516
rect 34348 4220 34388 4675
rect 34443 4556 34485 4565
rect 34443 4516 34444 4556
rect 34484 4516 34485 4556
rect 34443 4507 34485 4516
rect 34300 4180 34388 4220
rect 34300 4178 34340 4180
rect 33772 4136 33812 4147
rect 34300 4129 34340 4138
rect 33772 4061 33812 4096
rect 33771 4052 33813 4061
rect 33771 4012 33772 4052
rect 33812 4012 33813 4052
rect 33771 4003 33813 4012
rect 34444 4052 34484 4507
rect 34444 4003 34484 4012
rect 33675 3968 33717 3977
rect 33675 3928 33676 3968
rect 33716 3928 33717 3968
rect 33675 3919 33717 3928
rect 34539 3884 34581 3893
rect 34539 3844 34540 3884
rect 34580 3844 34581 3884
rect 34539 3835 34581 3844
rect 33675 3632 33717 3641
rect 33675 3592 33676 3632
rect 33716 3592 33717 3632
rect 33675 3583 33717 3592
rect 33676 3498 33716 3583
rect 34252 3464 34292 3473
rect 34292 3424 34388 3464
rect 34252 3415 34292 3424
rect 33868 3380 33908 3389
rect 33772 3340 33868 3380
rect 33675 2120 33717 2129
rect 33675 2080 33676 2120
rect 33716 2080 33717 2120
rect 33675 2071 33717 2080
rect 33676 2036 33716 2071
rect 33676 1985 33716 1996
rect 33772 1709 33812 3340
rect 33868 3331 33908 3340
rect 33928 3044 34296 3053
rect 33968 3004 34010 3044
rect 34050 3004 34092 3044
rect 34132 3004 34174 3044
rect 34214 3004 34256 3044
rect 33928 2995 34296 3004
rect 34348 2885 34388 3424
rect 34347 2876 34389 2885
rect 34347 2836 34348 2876
rect 34388 2836 34389 2876
rect 34347 2827 34389 2836
rect 34251 2792 34293 2801
rect 34251 2752 34252 2792
rect 34292 2752 34293 2792
rect 34251 2743 34293 2752
rect 33867 2708 33909 2717
rect 33867 2668 33868 2708
rect 33908 2668 33909 2708
rect 33867 2659 33909 2668
rect 33868 2624 33908 2659
rect 33868 2573 33908 2584
rect 34060 1952 34100 1961
rect 34252 1952 34292 2743
rect 34396 2633 34436 2642
rect 34436 2593 34484 2624
rect 34396 2584 34484 2593
rect 34444 2129 34484 2584
rect 34540 2456 34580 3835
rect 34636 3221 34676 6196
rect 34731 5984 34773 5993
rect 34731 5944 34732 5984
rect 34772 5944 34773 5984
rect 34731 5935 34773 5944
rect 34732 5657 34772 5935
rect 34731 5648 34773 5657
rect 34731 5608 34732 5648
rect 34772 5608 34773 5648
rect 34731 5599 34773 5608
rect 34732 5514 34772 5599
rect 34732 4733 34772 4818
rect 34731 4724 34773 4733
rect 34731 4684 34732 4724
rect 34772 4684 34773 4724
rect 34731 4675 34773 4684
rect 34828 4556 34868 6280
rect 34924 5900 34964 6364
rect 35500 6329 35540 6448
rect 35596 6439 35636 6448
rect 35692 6446 35732 6455
rect 35692 6329 35732 6406
rect 35499 6320 35541 6329
rect 35499 6280 35500 6320
rect 35540 6280 35541 6320
rect 35499 6271 35541 6280
rect 35691 6320 35733 6329
rect 35691 6280 35692 6320
rect 35732 6280 35733 6320
rect 35691 6271 35733 6280
rect 34924 5851 34964 5860
rect 35212 5732 35252 5741
rect 35212 5489 35252 5692
rect 35595 5648 35637 5657
rect 35595 5608 35596 5648
rect 35636 5608 35637 5648
rect 35595 5599 35637 5608
rect 35404 5489 35444 5574
rect 35596 5514 35636 5599
rect 35211 5480 35253 5489
rect 35211 5440 35212 5480
rect 35252 5440 35253 5480
rect 35211 5431 35253 5440
rect 35403 5480 35445 5489
rect 35403 5440 35404 5480
rect 35444 5440 35445 5480
rect 35403 5431 35445 5440
rect 35168 5312 35536 5321
rect 35208 5272 35250 5312
rect 35290 5272 35332 5312
rect 35372 5272 35414 5312
rect 35454 5272 35496 5312
rect 35168 5263 35536 5272
rect 35500 4976 35540 4985
rect 35116 4892 35156 4901
rect 34923 4808 34965 4817
rect 34923 4768 34924 4808
rect 34964 4768 34965 4808
rect 34923 4759 34965 4768
rect 34924 4674 34964 4759
rect 35116 4565 35156 4852
rect 34732 4516 34868 4556
rect 35115 4556 35157 4565
rect 35115 4516 35116 4556
rect 35156 4516 35157 4556
rect 34635 3212 34677 3221
rect 34635 3172 34636 3212
rect 34676 3172 34677 3212
rect 34635 3163 34677 3172
rect 34636 2717 34676 3163
rect 34635 2708 34677 2717
rect 34635 2668 34636 2708
rect 34676 2668 34677 2708
rect 34635 2659 34677 2668
rect 34540 2407 34580 2416
rect 34443 2120 34485 2129
rect 34443 2080 34444 2120
rect 34484 2080 34485 2120
rect 34443 2071 34485 2080
rect 34252 1912 34676 1952
rect 34060 1793 34100 1912
rect 34059 1784 34101 1793
rect 34059 1744 34060 1784
rect 34100 1744 34101 1784
rect 34059 1735 34101 1744
rect 33771 1700 33813 1709
rect 33771 1660 33772 1700
rect 33812 1660 33813 1700
rect 33771 1651 33813 1660
rect 33928 1532 34296 1541
rect 33968 1492 34010 1532
rect 34050 1492 34092 1532
rect 34132 1492 34174 1532
rect 34214 1492 34256 1532
rect 33928 1483 34296 1492
rect 34636 1112 34676 1912
rect 34636 1063 34676 1072
rect 33579 1028 33621 1037
rect 33579 988 33580 1028
rect 33620 988 33621 1028
rect 33579 979 33621 988
rect 34732 944 34772 4516
rect 35115 4507 35157 4516
rect 35500 4304 35540 4936
rect 35595 4976 35637 4985
rect 35595 4936 35596 4976
rect 35636 4936 35637 4976
rect 35595 4927 35637 4936
rect 35596 4842 35636 4927
rect 35500 4264 35732 4304
rect 35596 4136 35636 4145
rect 35116 3968 35156 3977
rect 35020 3928 35116 3968
rect 34924 2633 34964 2718
rect 34923 2624 34965 2633
rect 34923 2584 34924 2624
rect 34964 2584 34965 2624
rect 34923 2575 34965 2584
rect 34827 2120 34869 2129
rect 34827 2080 34828 2120
rect 34868 2080 34869 2120
rect 34827 2071 34869 2080
rect 34828 1280 34868 2071
rect 34923 1952 34965 1961
rect 35020 1952 35060 3928
rect 35116 3919 35156 3928
rect 35168 3800 35536 3809
rect 35208 3760 35250 3800
rect 35290 3760 35332 3800
rect 35372 3760 35414 3800
rect 35454 3760 35496 3800
rect 35168 3751 35536 3760
rect 35500 3464 35540 3475
rect 35500 3389 35540 3424
rect 35499 3380 35541 3389
rect 35499 3340 35500 3380
rect 35540 3340 35541 3380
rect 35499 3331 35541 3340
rect 35500 2801 35540 3331
rect 35499 2792 35541 2801
rect 35499 2752 35500 2792
rect 35540 2752 35541 2792
rect 35499 2743 35541 2752
rect 35168 2288 35536 2297
rect 35208 2248 35250 2288
rect 35290 2248 35332 2288
rect 35372 2248 35414 2288
rect 35454 2248 35496 2288
rect 35168 2239 35536 2248
rect 34923 1912 34924 1952
rect 34964 1912 35060 1952
rect 34923 1903 34965 1912
rect 34924 1818 34964 1903
rect 34828 1231 34868 1240
rect 35212 1196 35252 1205
rect 35212 953 35252 1156
rect 35596 1112 35636 4096
rect 35692 3632 35732 4264
rect 35788 3809 35828 6532
rect 35884 6329 35924 6943
rect 35883 6320 35925 6329
rect 35883 6280 35884 6320
rect 35924 6280 35925 6320
rect 35883 6271 35925 6280
rect 35787 3800 35829 3809
rect 35787 3760 35788 3800
rect 35828 3760 35829 3800
rect 35787 3751 35829 3760
rect 35692 3583 35732 3592
rect 35884 2120 35924 6271
rect 35980 5069 36020 6952
rect 36171 6992 36213 7001
rect 36171 6952 36172 6992
rect 36212 6952 36213 6992
rect 36171 6943 36213 6952
rect 36172 6858 36212 6943
rect 36172 6488 36212 6497
rect 36268 6488 36308 7027
rect 36364 6665 36404 7204
rect 36556 7160 36596 7169
rect 36844 7160 36884 8632
rect 37131 8000 37173 8009
rect 37131 7960 37132 8000
rect 37172 7960 37173 8000
rect 37131 7951 37173 7960
rect 37132 7673 37172 7951
rect 37131 7664 37173 7673
rect 37131 7624 37132 7664
rect 37172 7624 37173 7664
rect 37131 7615 37173 7624
rect 36363 6656 36405 6665
rect 36363 6616 36364 6656
rect 36404 6616 36405 6656
rect 36363 6607 36405 6616
rect 36212 6448 36308 6488
rect 36172 6439 36212 6448
rect 36268 5657 36308 6448
rect 36267 5648 36309 5657
rect 36267 5608 36268 5648
rect 36308 5608 36309 5648
rect 36267 5599 36309 5608
rect 36556 5573 36596 7120
rect 36748 7120 36884 7160
rect 36652 6474 36692 6483
rect 36652 5909 36692 6434
rect 36651 5900 36693 5909
rect 36651 5860 36652 5900
rect 36692 5860 36693 5900
rect 36651 5851 36693 5860
rect 36555 5564 36597 5573
rect 36555 5524 36556 5564
rect 36596 5524 36597 5564
rect 36555 5515 36597 5524
rect 36363 5480 36405 5489
rect 36363 5440 36364 5480
rect 36404 5440 36405 5480
rect 36363 5431 36405 5440
rect 36171 5144 36213 5153
rect 36171 5104 36172 5144
rect 36212 5104 36213 5144
rect 36171 5095 36213 5104
rect 35979 5060 36021 5069
rect 35979 5020 35980 5060
rect 36020 5020 36021 5060
rect 35979 5011 36021 5020
rect 35979 4892 36021 4901
rect 35979 4852 35980 4892
rect 36020 4852 36021 4892
rect 35979 4843 36021 4852
rect 36076 4892 36116 4901
rect 35980 4758 36020 4843
rect 36076 4397 36116 4852
rect 36075 4388 36117 4397
rect 36075 4348 36076 4388
rect 36116 4348 36117 4388
rect 36075 4339 36117 4348
rect 35980 4136 36020 4145
rect 35980 3296 36020 4096
rect 36075 4136 36117 4145
rect 36075 4096 36076 4136
rect 36116 4096 36117 4136
rect 36075 4087 36117 4096
rect 36076 4002 36116 4087
rect 36172 3464 36212 5095
rect 36364 3968 36404 5431
rect 36556 5153 36596 5515
rect 36555 5144 36597 5153
rect 36555 5104 36556 5144
rect 36596 5104 36597 5144
rect 36555 5095 36597 5104
rect 36556 4976 36596 4985
rect 36596 4936 36692 4976
rect 36556 4927 36596 4936
rect 36555 4640 36597 4649
rect 36555 4600 36556 4640
rect 36596 4600 36597 4640
rect 36555 4591 36597 4600
rect 36459 4388 36501 4397
rect 36459 4348 36460 4388
rect 36500 4348 36501 4388
rect 36459 4339 36501 4348
rect 36460 4220 36500 4339
rect 36460 4171 36500 4180
rect 36556 4220 36596 4591
rect 36556 4171 36596 4180
rect 36652 4061 36692 4936
rect 36651 4052 36693 4061
rect 36651 4012 36652 4052
rect 36692 4012 36693 4052
rect 36651 4003 36693 4012
rect 36364 3928 36500 3968
rect 36172 3415 36212 3424
rect 35980 3256 36404 3296
rect 36364 2876 36404 3256
rect 36364 2827 36404 2836
rect 36171 2792 36213 2801
rect 36171 2752 36172 2792
rect 36212 2752 36213 2792
rect 36171 2743 36213 2752
rect 36172 2624 36212 2743
rect 36172 2575 36212 2584
rect 36076 2120 36116 2129
rect 35884 2080 36076 2120
rect 36076 2071 36116 2080
rect 36267 1280 36309 1289
rect 36267 1240 36268 1280
rect 36308 1240 36309 1280
rect 36267 1231 36309 1240
rect 36268 1146 36308 1231
rect 36363 1196 36405 1205
rect 36363 1156 36364 1196
rect 36404 1156 36405 1196
rect 36363 1147 36405 1156
rect 35596 1063 35636 1072
rect 35020 944 35060 953
rect 34732 904 35020 944
rect 35020 895 35060 904
rect 35211 944 35253 953
rect 35211 904 35212 944
rect 35252 904 35253 944
rect 35211 895 35253 904
rect 35168 776 35536 785
rect 35208 736 35250 776
rect 35290 736 35332 776
rect 35372 736 35414 776
rect 35454 736 35496 776
rect 35168 727 35536 736
rect 35211 608 35253 617
rect 35211 568 35212 608
rect 35252 568 35253 608
rect 35211 559 35253 568
rect 34059 272 34101 281
rect 34059 232 34060 272
rect 34100 232 34101 272
rect 34059 223 34101 232
rect 33003 188 33045 197
rect 33003 148 33004 188
rect 33044 148 33045 188
rect 33003 139 33045 148
rect 34060 80 34100 223
rect 35212 80 35252 559
rect 36364 80 36404 1147
rect 36460 1121 36500 3928
rect 36556 2708 36596 2717
rect 36596 2668 36692 2708
rect 36556 2659 36596 2668
rect 36555 2540 36597 2549
rect 36555 2500 36556 2540
rect 36596 2500 36597 2540
rect 36555 2491 36597 2500
rect 36556 2036 36596 2491
rect 36556 1987 36596 1996
rect 36555 1700 36597 1709
rect 36555 1660 36556 1700
rect 36596 1660 36597 1700
rect 36555 1651 36597 1660
rect 36459 1112 36501 1121
rect 36459 1072 36460 1112
rect 36500 1072 36501 1112
rect 36459 1063 36501 1072
rect 36556 1112 36596 1651
rect 36652 1457 36692 2668
rect 36748 2624 36788 7120
rect 36843 6656 36885 6665
rect 36843 6616 36844 6656
rect 36884 6616 36885 6656
rect 36843 6607 36885 6616
rect 36844 6522 36884 6607
rect 37228 6404 37268 9295
rect 37516 9260 37556 9269
rect 37372 8681 37412 8690
rect 37516 8672 37556 9220
rect 37412 8641 37556 8672
rect 37372 8632 37556 8641
rect 37516 8504 37556 8513
rect 37516 7916 37556 8464
rect 37516 7867 37556 7876
rect 37323 7748 37365 7757
rect 37323 7708 37324 7748
rect 37364 7708 37365 7748
rect 37323 7699 37365 7708
rect 37324 7614 37364 7699
rect 37420 6656 37460 6665
rect 37612 6656 37652 10471
rect 38475 10184 38517 10193
rect 38475 10144 38476 10184
rect 38516 10144 38517 10184
rect 38475 10135 38517 10144
rect 37900 9512 37940 9521
rect 37708 9260 37748 9269
rect 37748 9220 37844 9260
rect 37708 9211 37748 9220
rect 37707 9092 37749 9101
rect 37707 9052 37708 9092
rect 37748 9052 37749 9092
rect 37707 9043 37749 9052
rect 37708 7916 37748 9043
rect 37804 8672 37844 9220
rect 37900 8849 37940 9472
rect 38091 9176 38133 9185
rect 38091 9136 38092 9176
rect 38132 9136 38133 9176
rect 38091 9127 38133 9136
rect 37899 8840 37941 8849
rect 37899 8800 37900 8840
rect 37940 8800 37941 8840
rect 37899 8791 37941 8800
rect 37804 8623 37844 8632
rect 37900 8672 37940 8681
rect 37940 8632 38036 8672
rect 37900 8623 37940 8632
rect 37803 8504 37845 8513
rect 37803 8464 37804 8504
rect 37844 8464 37845 8504
rect 37803 8455 37845 8464
rect 37708 7169 37748 7876
rect 37804 7421 37844 8455
rect 37899 8252 37941 8261
rect 37899 8212 37900 8252
rect 37940 8212 37941 8252
rect 37899 8203 37941 8212
rect 37900 8168 37940 8203
rect 37900 8117 37940 8128
rect 37803 7412 37845 7421
rect 37803 7372 37804 7412
rect 37844 7372 37845 7412
rect 37803 7363 37845 7372
rect 37803 7244 37845 7253
rect 37803 7204 37804 7244
rect 37844 7204 37845 7244
rect 37803 7195 37845 7204
rect 37707 7160 37749 7169
rect 37707 7120 37708 7160
rect 37748 7120 37749 7160
rect 37707 7111 37749 7120
rect 37804 7160 37844 7195
rect 37996 7160 38036 8632
rect 38092 8261 38132 9127
rect 38284 8672 38324 8681
rect 38188 8632 38284 8672
rect 38091 8252 38133 8261
rect 38091 8212 38092 8252
rect 38132 8212 38133 8252
rect 38091 8203 38133 8212
rect 38091 7748 38133 7757
rect 38091 7708 38092 7748
rect 38132 7708 38133 7748
rect 38091 7699 38133 7708
rect 38092 7614 38132 7699
rect 38188 7244 38228 8632
rect 38284 8623 38324 8632
rect 38380 8672 38420 8681
rect 38283 8504 38325 8513
rect 38283 8464 38284 8504
rect 38324 8464 38325 8504
rect 38283 8455 38325 8464
rect 38284 7916 38324 8455
rect 38284 7867 38324 7876
rect 38380 7328 38420 8632
rect 38476 8009 38516 10135
rect 38955 9848 38997 9857
rect 38955 9808 38956 9848
rect 38996 9808 38997 9848
rect 38955 9799 38997 9808
rect 38763 9512 38805 9521
rect 38763 9472 38764 9512
rect 38804 9472 38805 9512
rect 38763 9463 38805 9472
rect 38571 8924 38613 8933
rect 38571 8884 38572 8924
rect 38612 8884 38613 8924
rect 38571 8875 38613 8884
rect 38475 8000 38517 8009
rect 38475 7960 38476 8000
rect 38516 7960 38517 8000
rect 38475 7951 38517 7960
rect 38476 7748 38516 7757
rect 38476 7589 38516 7708
rect 38475 7580 38517 7589
rect 38475 7540 38476 7580
rect 38516 7540 38517 7580
rect 38475 7531 38517 7540
rect 37804 7109 37844 7120
rect 37900 7120 38036 7160
rect 38092 7204 38228 7244
rect 38284 7288 38420 7328
rect 37707 6992 37749 7001
rect 37707 6952 37708 6992
rect 37748 6952 37749 6992
rect 37707 6943 37749 6952
rect 37460 6616 37652 6656
rect 37420 6607 37460 6616
rect 37708 6488 37748 6943
rect 37708 6439 37748 6448
rect 37804 6488 37844 6497
rect 37900 6488 37940 7120
rect 37995 6992 38037 7001
rect 37995 6952 37996 6992
rect 38036 6952 38037 6992
rect 37995 6943 38037 6952
rect 37996 6858 38036 6943
rect 38092 6749 38132 7204
rect 38188 6992 38228 7001
rect 38188 6833 38228 6952
rect 38187 6824 38229 6833
rect 38187 6784 38188 6824
rect 38228 6784 38229 6824
rect 38187 6775 38229 6784
rect 38091 6740 38133 6749
rect 38091 6700 38092 6740
rect 38132 6700 38133 6740
rect 38091 6691 38133 6700
rect 37995 6656 38037 6665
rect 37995 6616 37996 6656
rect 38036 6616 38037 6656
rect 37995 6607 38037 6616
rect 37844 6448 37940 6488
rect 37228 6355 37268 6364
rect 37804 6161 37844 6448
rect 37803 6152 37845 6161
rect 37803 6112 37804 6152
rect 37844 6112 37845 6152
rect 37803 6103 37845 6112
rect 36843 5984 36885 5993
rect 36843 5944 36844 5984
rect 36884 5944 36885 5984
rect 36843 5935 36885 5944
rect 37515 5984 37557 5993
rect 37515 5944 37516 5984
rect 37556 5944 37557 5984
rect 37515 5935 37557 5944
rect 36844 5648 36884 5935
rect 37035 5900 37077 5909
rect 37035 5860 37036 5900
rect 37076 5860 37077 5900
rect 37035 5851 37077 5860
rect 37036 5766 37076 5851
rect 37420 5732 37460 5741
rect 36844 5599 36884 5608
rect 37324 5692 37420 5732
rect 37227 5480 37269 5489
rect 37227 5440 37228 5480
rect 37268 5440 37269 5480
rect 37227 5431 37269 5440
rect 36939 5396 36981 5405
rect 36939 5356 36940 5396
rect 36980 5356 36981 5396
rect 36939 5347 36981 5356
rect 36843 4304 36885 4313
rect 36843 4264 36844 4304
rect 36884 4264 36885 4304
rect 36843 4255 36885 4264
rect 36844 3893 36884 4255
rect 36843 3884 36885 3893
rect 36843 3844 36844 3884
rect 36884 3844 36885 3884
rect 36843 3835 36885 3844
rect 36940 2876 36980 5347
rect 37228 5346 37268 5431
rect 37228 5144 37268 5153
rect 37324 5144 37364 5692
rect 37420 5683 37460 5692
rect 37268 5104 37364 5144
rect 37228 5095 37268 5104
rect 37420 5060 37460 5069
rect 37324 5020 37420 5060
rect 37324 4976 37364 5020
rect 37420 5011 37460 5020
rect 37084 4966 37364 4976
rect 37124 4936 37364 4966
rect 37516 4976 37556 5935
rect 37611 5732 37653 5741
rect 37611 5692 37612 5732
rect 37652 5692 37653 5732
rect 37611 5683 37653 5692
rect 37996 5732 38036 6607
rect 38092 6488 38132 6691
rect 38284 6581 38324 7288
rect 38475 7244 38517 7253
rect 38380 7204 38476 7244
rect 38516 7204 38517 7244
rect 38380 7160 38420 7204
rect 38475 7195 38517 7204
rect 38380 7111 38420 7120
rect 38572 6908 38612 8875
rect 38668 7916 38708 7925
rect 38668 7589 38708 7876
rect 38667 7580 38709 7589
rect 38667 7540 38668 7580
rect 38708 7540 38709 7580
rect 38667 7531 38709 7540
rect 38667 7412 38709 7421
rect 38667 7372 38668 7412
rect 38708 7372 38709 7412
rect 38667 7363 38709 7372
rect 38380 6868 38612 6908
rect 38283 6572 38325 6581
rect 38283 6532 38284 6572
rect 38324 6532 38325 6572
rect 38283 6523 38325 6532
rect 38188 6488 38228 6497
rect 38092 6448 38188 6488
rect 38188 6439 38228 6448
rect 38284 6488 38324 6523
rect 38284 6438 38324 6448
rect 38187 6236 38229 6245
rect 38187 6196 38188 6236
rect 38228 6196 38229 6236
rect 38187 6187 38229 6196
rect 38188 5900 38228 6187
rect 38188 5851 38228 5860
rect 37996 5683 38036 5692
rect 38380 5732 38420 6868
rect 38668 6572 38708 7363
rect 38764 6749 38804 9463
rect 38859 8672 38901 8681
rect 38859 8632 38860 8672
rect 38900 8632 38901 8672
rect 38859 8623 38901 8632
rect 38860 8538 38900 8623
rect 38956 8168 38996 9799
rect 39147 9512 39189 9521
rect 39147 9472 39148 9512
rect 39188 9472 39189 9512
rect 39147 9463 39189 9472
rect 39340 9512 39380 9521
rect 39148 9378 39188 9463
rect 39340 9353 39380 9472
rect 39339 9344 39381 9353
rect 39339 9304 39340 9344
rect 39380 9304 39381 9344
rect 39339 9295 39381 9304
rect 39435 9008 39477 9017
rect 39435 8968 39436 9008
rect 39476 8968 39477 9008
rect 39435 8959 39477 8968
rect 39339 8756 39381 8765
rect 39339 8716 39340 8756
rect 39380 8716 39381 8756
rect 39339 8707 39381 8716
rect 39340 8686 39380 8707
rect 39340 8621 39380 8646
rect 38860 8128 38996 8168
rect 38860 7076 38900 8128
rect 38955 8000 38997 8009
rect 38955 7960 38956 8000
rect 38996 7960 38997 8000
rect 38955 7951 38997 7960
rect 39052 8000 39092 8009
rect 39436 8000 39476 8959
rect 39531 8504 39573 8513
rect 39531 8464 39532 8504
rect 39572 8464 39573 8504
rect 39531 8455 39573 8464
rect 39532 8370 39572 8455
rect 38956 7866 38996 7951
rect 38860 7036 38996 7076
rect 38859 6824 38901 6833
rect 38859 6784 38860 6824
rect 38900 6784 38901 6824
rect 38859 6775 38901 6784
rect 38763 6740 38805 6749
rect 38763 6700 38764 6740
rect 38804 6700 38805 6740
rect 38763 6691 38805 6700
rect 38380 5683 38420 5692
rect 38476 6532 38708 6572
rect 37612 5598 37652 5683
rect 38476 5564 38516 6532
rect 38668 6404 38708 6532
rect 38764 6488 38804 6497
rect 38764 6404 38804 6448
rect 38668 6364 38804 6404
rect 38571 5900 38613 5909
rect 38571 5860 38572 5900
rect 38612 5860 38613 5900
rect 38571 5851 38613 5860
rect 38572 5766 38612 5851
rect 38763 5816 38805 5825
rect 38763 5776 38764 5816
rect 38804 5776 38805 5816
rect 38763 5767 38805 5776
rect 38380 5524 38516 5564
rect 37804 5480 37844 5489
rect 37612 4976 37652 4985
rect 37516 4936 37612 4976
rect 37084 4917 37124 4926
rect 37516 4892 37556 4936
rect 37612 4927 37652 4936
rect 37420 4852 37556 4892
rect 37036 4136 37076 4147
rect 37036 4061 37076 4096
rect 37035 4052 37077 4061
rect 37035 4012 37036 4052
rect 37076 4012 37077 4052
rect 37035 4003 37077 4012
rect 37420 3464 37460 4852
rect 37564 4145 37604 4154
rect 37604 4105 37652 4136
rect 37564 4096 37652 4105
rect 37515 3800 37557 3809
rect 37515 3760 37516 3800
rect 37556 3760 37557 3800
rect 37515 3751 37557 3760
rect 37420 3415 37460 3424
rect 36940 2827 36980 2836
rect 37132 2708 37172 2717
rect 36748 2584 36884 2624
rect 36748 2456 36788 2465
rect 36651 1448 36693 1457
rect 36651 1408 36652 1448
rect 36692 1408 36693 1448
rect 36651 1399 36693 1408
rect 36556 1063 36596 1072
rect 36748 785 36788 2416
rect 36844 1280 36884 2584
rect 36940 1952 36980 1961
rect 36940 1373 36980 1912
rect 37132 1877 37172 2668
rect 37131 1868 37173 1877
rect 37131 1828 37132 1868
rect 37172 1828 37173 1868
rect 37131 1819 37173 1828
rect 36939 1364 36981 1373
rect 36939 1324 36940 1364
rect 36980 1324 36981 1364
rect 36939 1315 36981 1324
rect 36844 1231 36884 1240
rect 36747 776 36789 785
rect 36747 736 36748 776
rect 36788 736 36789 776
rect 36747 727 36789 736
rect 37516 80 37556 3751
rect 37612 3632 37652 4096
rect 37612 3583 37652 3592
rect 37708 3968 37748 3977
rect 37708 3389 37748 3928
rect 37707 3380 37749 3389
rect 37707 3340 37708 3380
rect 37748 3340 37749 3380
rect 37707 3331 37749 3340
rect 37611 3128 37653 3137
rect 37611 3088 37612 3128
rect 37652 3088 37653 3128
rect 37611 3079 37653 3088
rect 37612 2876 37652 3079
rect 37612 2827 37652 2836
rect 37804 2120 37844 5440
rect 37995 4304 38037 4313
rect 37995 4264 37996 4304
rect 38036 4264 38132 4304
rect 37995 4255 38037 4264
rect 38092 4220 38132 4264
rect 38092 4171 38132 4180
rect 38283 4220 38325 4229
rect 38283 4180 38284 4220
rect 38324 4180 38325 4220
rect 38283 4171 38325 4180
rect 38284 4086 38324 4171
rect 37899 3968 37941 3977
rect 37899 3928 37900 3968
rect 37940 3928 37941 3968
rect 37899 3919 37941 3928
rect 37900 3834 37940 3919
rect 38284 3464 38324 3473
rect 38091 3380 38133 3389
rect 38091 3340 38092 3380
rect 38132 3340 38133 3380
rect 38091 3331 38133 3340
rect 38092 3246 38132 3331
rect 37899 3212 37941 3221
rect 37899 3172 37900 3212
rect 37940 3172 37941 3212
rect 37899 3163 37941 3172
rect 37900 3078 37940 3163
rect 38091 3128 38133 3137
rect 38091 3088 38092 3128
rect 38132 3088 38133 3128
rect 38091 3079 38133 3088
rect 37995 2120 38037 2129
rect 37804 2080 37940 2120
rect 37803 1952 37845 1961
rect 37803 1912 37804 1952
rect 37844 1912 37845 1952
rect 37803 1903 37845 1912
rect 37804 1818 37844 1903
rect 37900 113 37940 2080
rect 37995 2080 37996 2120
rect 38036 2080 38037 2120
rect 37995 2071 38037 2080
rect 37996 1112 38036 2071
rect 38092 2045 38132 3079
rect 38284 2633 38324 3424
rect 38380 3221 38420 5524
rect 38764 4145 38804 5767
rect 38860 5648 38900 6775
rect 38956 5909 38996 7036
rect 38955 5900 38997 5909
rect 38955 5860 38956 5900
rect 38996 5860 38997 5900
rect 38955 5851 38997 5860
rect 38860 5599 38900 5608
rect 38956 5648 38996 5657
rect 39052 5648 39092 7960
rect 39340 7960 39436 8000
rect 39147 7328 39189 7337
rect 39147 7288 39148 7328
rect 39188 7288 39189 7328
rect 39147 7279 39189 7288
rect 38996 5608 39092 5648
rect 38956 5599 38996 5608
rect 38955 5480 38997 5489
rect 38955 5440 38956 5480
rect 38996 5440 38997 5480
rect 38955 5431 38997 5440
rect 38860 4976 38900 4985
rect 38860 4229 38900 4936
rect 38859 4220 38901 4229
rect 38859 4180 38860 4220
rect 38900 4180 38901 4220
rect 38859 4171 38901 4180
rect 38763 4136 38805 4145
rect 38763 4096 38764 4136
rect 38804 4096 38805 4136
rect 38763 4087 38805 4096
rect 38476 3968 38516 3977
rect 38379 3212 38421 3221
rect 38379 3172 38380 3212
rect 38420 3172 38421 3212
rect 38379 3163 38421 3172
rect 38283 2624 38325 2633
rect 38283 2584 38284 2624
rect 38324 2584 38325 2624
rect 38283 2575 38325 2584
rect 38091 2036 38133 2045
rect 38091 1996 38092 2036
rect 38132 1996 38133 2036
rect 38091 1987 38133 1996
rect 37996 1063 38036 1072
rect 38476 449 38516 3928
rect 38764 2624 38804 2633
rect 38764 2129 38804 2584
rect 38859 2288 38901 2297
rect 38859 2248 38860 2288
rect 38900 2248 38901 2288
rect 38859 2239 38901 2248
rect 38763 2120 38805 2129
rect 38763 2080 38764 2120
rect 38804 2080 38805 2120
rect 38763 2071 38805 2080
rect 38667 1616 38709 1625
rect 38667 1576 38668 1616
rect 38708 1576 38709 1616
rect 38667 1567 38709 1576
rect 38475 440 38517 449
rect 38475 400 38476 440
rect 38516 400 38517 440
rect 38475 391 38517 400
rect 37899 104 37941 113
rect 30795 55 31124 60
rect 30796 20 31124 55
rect 31736 0 31816 80
rect 32888 0 32968 80
rect 34040 0 34120 80
rect 35192 0 35272 80
rect 36344 0 36424 80
rect 37496 0 37576 80
rect 37899 64 37900 104
rect 37940 64 37941 104
rect 38668 80 38708 1567
rect 38860 1112 38900 2239
rect 38956 2120 38996 5431
rect 39052 4985 39092 5608
rect 39148 5060 39188 7279
rect 39244 6497 39284 6578
rect 39243 6488 39285 6497
rect 39243 6443 39244 6488
rect 39284 6443 39285 6488
rect 39243 6439 39285 6443
rect 39244 6434 39284 6439
rect 39340 5732 39380 7960
rect 39436 7951 39476 7960
rect 39532 8000 39572 8009
rect 39628 8000 39668 10639
rect 40299 9512 40341 9521
rect 40299 9472 40300 9512
rect 40340 9472 40341 9512
rect 40299 9463 40341 9472
rect 40588 9512 40628 9521
rect 39915 8672 39957 8681
rect 39915 8632 39916 8672
rect 39956 8632 39957 8672
rect 39915 8623 39957 8632
rect 39916 8538 39956 8623
rect 39724 8504 39764 8513
rect 39724 8009 39764 8464
rect 39572 7960 39668 8000
rect 39723 8000 39765 8009
rect 39723 7960 39724 8000
rect 39764 7960 39765 8000
rect 39435 7580 39477 7589
rect 39435 7540 39436 7580
rect 39476 7540 39477 7580
rect 39435 7531 39477 7540
rect 39436 6656 39476 7531
rect 39436 6607 39476 6616
rect 39148 5020 39284 5060
rect 39051 4976 39093 4985
rect 39051 4936 39052 4976
rect 39092 4936 39093 4976
rect 39051 4927 39093 4936
rect 39052 4640 39092 4927
rect 39147 4892 39189 4901
rect 39147 4852 39148 4892
rect 39188 4852 39189 4892
rect 39147 4843 39189 4852
rect 39148 4758 39188 4843
rect 39244 4733 39284 5020
rect 39340 4976 39380 5692
rect 39436 5732 39476 5741
rect 39532 5732 39572 7960
rect 39723 7951 39765 7960
rect 40012 8000 40052 8009
rect 39915 7580 39957 7589
rect 39915 7540 39916 7580
rect 39956 7540 39957 7580
rect 39915 7531 39957 7540
rect 39628 7160 39668 7169
rect 39628 6245 39668 7120
rect 39819 7160 39861 7169
rect 39819 7120 39820 7160
rect 39860 7120 39861 7160
rect 39819 7111 39861 7120
rect 39820 7026 39860 7111
rect 39723 6488 39765 6497
rect 39723 6448 39724 6488
rect 39764 6448 39765 6488
rect 39723 6439 39765 6448
rect 39627 6236 39669 6245
rect 39627 6196 39628 6236
rect 39668 6196 39669 6236
rect 39627 6187 39669 6196
rect 39476 5692 39572 5732
rect 39436 5683 39476 5692
rect 39532 5060 39572 5692
rect 39628 5237 39668 6187
rect 39627 5228 39669 5237
rect 39627 5188 39628 5228
rect 39668 5188 39669 5228
rect 39627 5179 39669 5188
rect 39532 5020 39668 5060
rect 39340 4936 39476 4976
rect 39339 4808 39381 4817
rect 39339 4768 39340 4808
rect 39380 4768 39381 4808
rect 39339 4759 39381 4768
rect 39243 4724 39285 4733
rect 39243 4684 39244 4724
rect 39284 4684 39285 4724
rect 39243 4675 39285 4684
rect 39340 4674 39380 4759
rect 39052 4600 39188 4640
rect 39052 4136 39092 4145
rect 39052 3641 39092 4096
rect 39148 4136 39188 4600
rect 39436 4220 39476 4936
rect 39532 4934 39572 4943
rect 39532 4733 39572 4894
rect 39531 4724 39573 4733
rect 39531 4684 39532 4724
rect 39572 4684 39573 4724
rect 39531 4675 39573 4684
rect 39628 4313 39668 5020
rect 39627 4304 39669 4313
rect 39627 4264 39628 4304
rect 39668 4264 39669 4304
rect 39627 4255 39669 4264
rect 39532 4220 39572 4229
rect 39436 4180 39532 4220
rect 39532 4171 39572 4180
rect 39628 4220 39668 4255
rect 39628 4170 39668 4180
rect 39148 4087 39188 4096
rect 39147 3968 39189 3977
rect 39147 3928 39148 3968
rect 39188 3928 39189 3968
rect 39147 3919 39189 3928
rect 39051 3632 39093 3641
rect 39051 3592 39052 3632
rect 39092 3592 39093 3632
rect 39051 3583 39093 3592
rect 38956 2071 38996 2080
rect 39148 1112 39188 3919
rect 39724 3632 39764 6439
rect 39820 6404 39860 6413
rect 39916 6404 39956 7531
rect 40012 6824 40052 7960
rect 40012 6784 40148 6824
rect 40011 6572 40053 6581
rect 40011 6532 40012 6572
rect 40052 6532 40053 6572
rect 40011 6523 40053 6532
rect 39860 6364 39956 6404
rect 39820 6355 39860 6364
rect 40012 6320 40052 6523
rect 40012 6271 40052 6280
rect 40011 5900 40053 5909
rect 40011 5860 40012 5900
rect 40052 5860 40053 5900
rect 40011 5851 40053 5860
rect 39916 5648 39956 5657
rect 39916 5489 39956 5608
rect 39915 5480 39957 5489
rect 39915 5440 39916 5480
rect 39956 5440 39957 5480
rect 39915 5431 39957 5440
rect 39916 3641 39956 3726
rect 39724 3583 39764 3592
rect 39915 3632 39957 3641
rect 39915 3592 39916 3632
rect 39956 3592 39957 3632
rect 39915 3583 39957 3592
rect 39531 3548 39573 3557
rect 39531 3508 39532 3548
rect 39572 3508 39573 3548
rect 39531 3499 39573 3508
rect 39532 3464 39572 3499
rect 40012 3464 40052 5851
rect 40108 4397 40148 6784
rect 40203 6320 40245 6329
rect 40203 6280 40204 6320
rect 40244 6280 40245 6320
rect 40203 6271 40245 6280
rect 40204 6186 40244 6271
rect 40300 4817 40340 9463
rect 40588 8681 40628 9472
rect 40971 9428 41013 9437
rect 40971 9388 40972 9428
rect 41012 9388 41013 9428
rect 40971 9379 41013 9388
rect 40972 9294 41012 9379
rect 41356 9344 41396 9353
rect 41396 9304 41492 9344
rect 41356 9295 41396 9304
rect 40780 9260 40820 9269
rect 40780 8765 40820 9220
rect 41164 9260 41204 9269
rect 41204 9220 41300 9260
rect 41164 9211 41204 9220
rect 40779 8756 40821 8765
rect 40779 8716 40780 8756
rect 40820 8716 40821 8756
rect 40779 8707 40821 8716
rect 40587 8672 40629 8681
rect 40587 8632 40588 8672
rect 40628 8632 40629 8672
rect 40587 8623 40629 8632
rect 41164 8672 41204 8681
rect 40683 8420 40725 8429
rect 40683 8380 40684 8420
rect 40724 8380 40725 8420
rect 40683 8371 40725 8380
rect 40684 8168 40724 8371
rect 40684 8119 40724 8128
rect 40492 7986 40532 7995
rect 40492 7421 40532 7946
rect 40876 7916 40916 7925
rect 40876 7505 40916 7876
rect 41068 7748 41108 7757
rect 41068 7505 41108 7708
rect 41164 7589 41204 8632
rect 41260 8513 41300 9220
rect 41356 8756 41396 8765
rect 41259 8504 41301 8513
rect 41259 8464 41260 8504
rect 41300 8464 41301 8504
rect 41259 8455 41301 8464
rect 41356 8177 41396 8716
rect 41355 8168 41397 8177
rect 41355 8128 41356 8168
rect 41396 8128 41397 8168
rect 41355 8119 41397 8128
rect 41452 8000 41492 9304
rect 42507 8840 42549 8849
rect 42507 8800 42508 8840
rect 42548 8800 42549 8840
rect 42507 8791 42549 8800
rect 41548 8504 41588 8513
rect 41548 8177 41588 8464
rect 41547 8168 41589 8177
rect 41547 8128 41548 8168
rect 41588 8128 41589 8168
rect 41547 8119 41589 8128
rect 41356 7960 41492 8000
rect 41259 7916 41301 7925
rect 41259 7876 41260 7916
rect 41300 7876 41301 7916
rect 41259 7867 41301 7876
rect 41260 7782 41300 7867
rect 41163 7580 41205 7589
rect 41163 7540 41164 7580
rect 41204 7540 41205 7580
rect 41163 7531 41205 7540
rect 40875 7496 40917 7505
rect 40875 7456 40876 7496
rect 40916 7456 40917 7496
rect 40875 7447 40917 7456
rect 41067 7496 41109 7505
rect 41067 7456 41068 7496
rect 41108 7456 41109 7496
rect 41067 7447 41109 7456
rect 40491 7412 40533 7421
rect 40491 7372 40492 7412
rect 40532 7372 40533 7412
rect 40491 7363 40533 7372
rect 41259 7412 41301 7421
rect 41259 7372 41260 7412
rect 41300 7372 41301 7412
rect 41259 7363 41301 7372
rect 41260 7278 41300 7363
rect 40971 7160 41013 7169
rect 41068 7160 41108 7169
rect 40971 7120 40972 7160
rect 41012 7120 41068 7160
rect 40971 7111 41013 7120
rect 41068 7111 41108 7120
rect 41067 6824 41109 6833
rect 41067 6784 41068 6824
rect 41108 6784 41109 6824
rect 41067 6775 41109 6784
rect 41068 6656 41108 6775
rect 41068 6607 41108 6616
rect 40396 6404 40436 6413
rect 40876 6404 40916 6413
rect 40436 6364 40532 6404
rect 40396 6355 40436 6364
rect 40396 5653 40436 5662
rect 40396 5153 40436 5613
rect 40492 5564 40532 6364
rect 40876 6245 40916 6364
rect 41259 6404 41301 6413
rect 41259 6364 41260 6404
rect 41300 6364 41301 6404
rect 41259 6355 41301 6364
rect 41260 6270 41300 6355
rect 40875 6236 40917 6245
rect 40875 6196 40876 6236
rect 40916 6196 40917 6236
rect 40875 6187 40917 6196
rect 41067 6152 41109 6161
rect 41067 6112 41068 6152
rect 41108 6112 41109 6152
rect 41067 6103 41109 6112
rect 41068 5900 41108 6103
rect 41356 5909 41396 7960
rect 41451 7832 41493 7841
rect 41451 7792 41452 7832
rect 41492 7792 41493 7832
rect 41451 7783 41493 7792
rect 41452 7698 41492 7783
rect 41451 7328 41493 7337
rect 41451 7288 41452 7328
rect 41492 7288 41493 7328
rect 41451 7279 41493 7288
rect 41452 7244 41492 7279
rect 41452 7193 41492 7204
rect 41643 7160 41685 7169
rect 41643 7120 41644 7160
rect 41684 7120 41685 7160
rect 41643 7111 41685 7120
rect 41644 6992 41684 7111
rect 41644 6943 41684 6952
rect 42508 6581 42548 8791
rect 42507 6572 42549 6581
rect 42507 6532 42508 6572
rect 42548 6532 42549 6572
rect 42507 6523 42549 6532
rect 41451 6488 41493 6497
rect 41451 6448 41452 6488
rect 41492 6448 41493 6488
rect 41451 6439 41493 6448
rect 41452 6320 41492 6439
rect 41452 6271 41492 6280
rect 41068 5851 41108 5860
rect 41355 5900 41397 5909
rect 41355 5860 41356 5900
rect 41396 5860 41397 5900
rect 41355 5851 41397 5860
rect 41451 5816 41493 5825
rect 41451 5776 41452 5816
rect 41492 5776 41493 5816
rect 41451 5767 41493 5776
rect 40876 5732 40916 5741
rect 40588 5564 40628 5573
rect 40492 5524 40588 5564
rect 40588 5515 40628 5524
rect 40395 5144 40437 5153
rect 40876 5144 40916 5692
rect 41260 5732 41300 5741
rect 40972 5153 41012 5238
rect 40395 5104 40396 5144
rect 40436 5104 40437 5144
rect 40395 5095 40437 5104
rect 40684 5104 40916 5144
rect 40971 5144 41013 5153
rect 40971 5104 40972 5144
rect 41012 5104 41013 5144
rect 40299 4808 40341 4817
rect 40299 4768 40300 4808
rect 40340 4768 40341 4808
rect 40299 4759 40341 4768
rect 40107 4388 40149 4397
rect 40107 4348 40108 4388
rect 40148 4348 40149 4388
rect 40107 4339 40149 4348
rect 40108 4136 40148 4339
rect 40588 4141 40628 4150
rect 40148 4096 40244 4136
rect 40108 4087 40148 4096
rect 40107 3548 40149 3557
rect 40107 3508 40108 3548
rect 40148 3508 40149 3548
rect 40107 3499 40149 3508
rect 39532 3413 39572 3424
rect 39916 3424 40052 3464
rect 40108 3464 40148 3499
rect 39628 2624 39668 2633
rect 39916 2624 39956 3424
rect 40108 3413 40148 3424
rect 40204 3296 40244 4096
rect 39668 2584 39956 2624
rect 40012 3256 40244 3296
rect 40299 3296 40341 3305
rect 40299 3256 40300 3296
rect 40340 3256 40341 3296
rect 40012 2624 40052 3256
rect 40299 3247 40341 3256
rect 39628 2575 39668 2584
rect 40012 2575 40052 2584
rect 40204 2624 40244 2633
rect 40300 2624 40340 3247
rect 40588 2801 40628 4101
rect 40684 3725 40724 5104
rect 40971 5095 41013 5104
rect 40779 4976 40821 4985
rect 40779 4936 40780 4976
rect 40820 4936 40821 4976
rect 40779 4927 40821 4936
rect 40780 4842 40820 4927
rect 41260 4901 41300 5692
rect 41452 5682 41492 5767
rect 41355 5480 41397 5489
rect 41355 5440 41356 5480
rect 41396 5440 41397 5480
rect 41355 5431 41397 5440
rect 41164 4892 41204 4901
rect 40876 4852 41164 4892
rect 40779 4052 40821 4061
rect 40779 4012 40780 4052
rect 40820 4012 40821 4052
rect 40779 4003 40821 4012
rect 40780 3918 40820 4003
rect 40683 3716 40725 3725
rect 40683 3676 40684 3716
rect 40724 3676 40725 3716
rect 40683 3667 40725 3676
rect 40587 2792 40629 2801
rect 40587 2752 40588 2792
rect 40628 2752 40629 2792
rect 40587 2743 40629 2752
rect 40244 2584 40340 2624
rect 40204 2575 40244 2584
rect 40876 2465 40916 4852
rect 41164 4843 41204 4852
rect 41259 4892 41301 4901
rect 41259 4852 41260 4892
rect 41300 4852 41301 4892
rect 41259 4843 41301 4852
rect 41356 4808 41396 5431
rect 41451 5144 41493 5153
rect 41451 5104 41452 5144
rect 41492 5104 41493 5144
rect 41451 5095 41493 5104
rect 41356 4759 41396 4768
rect 41067 4724 41109 4733
rect 41067 4684 41068 4724
rect 41108 4684 41109 4724
rect 41067 4675 41109 4684
rect 40972 4220 41012 4229
rect 40972 3137 41012 4180
rect 40971 3128 41013 3137
rect 40971 3088 40972 3128
rect 41012 3088 41013 3128
rect 40971 3079 41013 3088
rect 41068 2633 41108 4675
rect 41452 4388 41492 5095
rect 41740 4892 41780 4901
rect 41547 4724 41589 4733
rect 41547 4684 41548 4724
rect 41588 4684 41589 4724
rect 41547 4675 41589 4684
rect 41548 4590 41588 4675
rect 41548 4388 41588 4397
rect 41452 4348 41548 4388
rect 41548 4339 41588 4348
rect 41355 4220 41397 4229
rect 41355 4180 41356 4220
rect 41396 4180 41397 4220
rect 41355 4171 41397 4180
rect 41356 4086 41396 4171
rect 41740 4061 41780 4852
rect 41739 4052 41781 4061
rect 41739 4012 41740 4052
rect 41780 4012 41781 4052
rect 41739 4003 41781 4012
rect 41164 3968 41204 3977
rect 41067 2624 41109 2633
rect 41067 2584 41068 2624
rect 41108 2584 41109 2624
rect 41067 2575 41109 2584
rect 40875 2456 40917 2465
rect 40875 2416 40876 2456
rect 40916 2416 40917 2456
rect 40875 2407 40917 2416
rect 39723 2372 39765 2381
rect 39723 2332 39724 2372
rect 39764 2332 39765 2372
rect 39723 2323 39765 2332
rect 39243 1952 39285 1961
rect 39243 1912 39244 1952
rect 39284 1912 39285 1952
rect 39243 1903 39285 1912
rect 39244 1818 39284 1903
rect 39531 1700 39573 1709
rect 39531 1660 39532 1700
rect 39572 1660 39573 1700
rect 39531 1651 39573 1660
rect 39532 1566 39572 1651
rect 39627 1196 39669 1205
rect 39627 1156 39628 1196
rect 39668 1156 39669 1196
rect 39627 1147 39669 1156
rect 39244 1112 39284 1121
rect 39148 1072 39244 1112
rect 38860 1063 38900 1072
rect 39244 1063 39284 1072
rect 39628 1062 39668 1147
rect 39435 1028 39477 1037
rect 39435 988 39436 1028
rect 39476 988 39477 1028
rect 39435 979 39477 988
rect 39436 944 39476 979
rect 39436 893 39476 904
rect 39724 524 39764 2323
rect 40780 1952 40820 1961
rect 40587 1784 40629 1793
rect 40587 1744 40588 1784
rect 40628 1744 40629 1784
rect 40587 1735 40629 1744
rect 40203 1364 40245 1373
rect 40203 1324 40204 1364
rect 40244 1324 40245 1364
rect 40203 1315 40245 1324
rect 40204 1280 40244 1315
rect 40204 1229 40244 1240
rect 40588 1280 40628 1735
rect 40780 1289 40820 1912
rect 41164 1793 41204 3928
rect 41451 3548 41493 3557
rect 41451 3508 41452 3548
rect 41492 3508 41493 3548
rect 41451 3499 41493 3508
rect 41355 3464 41397 3473
rect 41355 3424 41356 3464
rect 41396 3424 41397 3464
rect 41355 3415 41397 3424
rect 41356 3330 41396 3415
rect 41259 3296 41301 3305
rect 41259 3256 41260 3296
rect 41300 3256 41301 3296
rect 41259 3247 41301 3256
rect 41260 2297 41300 3247
rect 41355 2960 41397 2969
rect 41355 2920 41356 2960
rect 41396 2920 41397 2960
rect 41355 2911 41397 2920
rect 41259 2288 41301 2297
rect 41259 2248 41260 2288
rect 41300 2248 41301 2288
rect 41259 2239 41301 2248
rect 41259 2120 41301 2129
rect 41259 2080 41260 2120
rect 41300 2080 41301 2120
rect 41259 2071 41301 2080
rect 41260 1986 41300 2071
rect 41163 1784 41205 1793
rect 41163 1744 41164 1784
rect 41204 1744 41205 1784
rect 41163 1735 41205 1744
rect 40588 1231 40628 1240
rect 40779 1280 40821 1289
rect 40779 1240 40780 1280
rect 40820 1240 40821 1280
rect 40779 1231 40821 1240
rect 40012 1196 40052 1205
rect 39820 944 39860 953
rect 39820 701 39860 904
rect 39819 692 39861 701
rect 39819 652 39820 692
rect 39860 652 39861 692
rect 39819 643 39861 652
rect 39724 484 39860 524
rect 39820 80 39860 484
rect 40012 281 40052 1156
rect 41164 1196 41204 1205
rect 40971 944 41013 953
rect 40971 904 40972 944
rect 41012 904 41013 944
rect 40971 895 41013 904
rect 40972 810 41012 895
rect 41164 617 41204 1156
rect 41356 1196 41396 2911
rect 41452 2624 41492 3499
rect 41547 3296 41589 3305
rect 41547 3256 41548 3296
rect 41588 3256 41589 3296
rect 41547 3247 41589 3256
rect 41548 3162 41588 3247
rect 41643 2792 41685 2801
rect 41643 2752 41644 2792
rect 41684 2752 41685 2792
rect 41643 2743 41685 2752
rect 41644 2658 41684 2743
rect 41452 2575 41492 2584
rect 41547 2624 41589 2633
rect 41547 2584 41548 2624
rect 41588 2584 41589 2624
rect 41547 2575 41589 2584
rect 41548 1364 41588 2575
rect 41548 1315 41588 1324
rect 41356 1147 41396 1156
rect 41163 608 41205 617
rect 41163 568 41164 608
rect 41204 568 41205 608
rect 41163 559 41205 568
rect 40011 272 40053 281
rect 40011 232 40012 272
rect 40052 232 40053 272
rect 40011 223 40053 232
rect 37899 55 37941 64
rect 38648 0 38728 80
rect 39800 0 39880 80
<< via2 >>
rect 1708 10480 1748 10520
rect 1612 10144 1652 10184
rect 1612 8884 1652 8924
rect 4684 9808 4724 9848
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 2956 9472 2996 9512
rect 3244 9472 3284 9512
rect 3436 9304 3476 9344
rect 2092 8716 2132 8756
rect 2860 8716 2900 8756
rect 1708 8380 1748 8420
rect 1324 8128 1364 8168
rect 1900 8128 1940 8168
rect 1804 7960 1844 8000
rect 1708 7540 1748 7580
rect 1132 6448 1172 6488
rect 1420 6952 1460 6992
rect 1804 7372 1844 7412
rect 1324 5944 1364 5984
rect 1132 5524 1172 5564
rect 1324 5440 1364 5480
rect 1324 5188 1364 5228
rect 1132 4432 1172 4472
rect 1324 4096 1364 4136
rect 1420 3592 1460 3632
rect 1324 3424 1364 3464
rect 1324 2752 1364 2792
rect 1132 2500 1172 2540
rect 1516 3340 1556 3380
rect 1516 1996 1556 2036
rect 2572 8632 2612 8672
rect 3052 8632 3092 8672
rect 3148 8212 3188 8252
rect 3052 7708 3092 7748
rect 2956 7288 2996 7328
rect 2476 7036 2516 7076
rect 1804 5944 1844 5984
rect 2956 6448 2996 6488
rect 2668 6280 2708 6320
rect 3148 7288 3188 7328
rect 3148 7120 3188 7160
rect 2860 5692 2900 5732
rect 2284 5356 2324 5396
rect 2668 4936 2708 4976
rect 2764 4852 2804 4892
rect 2956 5020 2996 5060
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 4684 8968 4724 9008
rect 4972 9472 5012 9512
rect 4876 9136 4916 9176
rect 3820 8800 3860 8840
rect 4780 8800 4820 8840
rect 3340 8128 3380 8168
rect 4012 8716 4052 8756
rect 3916 8548 3956 8588
rect 4396 8637 4436 8672
rect 4396 8632 4436 8637
rect 5932 9472 5972 9512
rect 5068 8632 5108 8672
rect 3820 8128 3860 8168
rect 3820 7960 3860 8000
rect 4300 7960 4340 8000
rect 4588 7960 4628 8000
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 4780 8044 4820 8084
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 4588 7540 4628 7580
rect 3820 7288 3860 7328
rect 4204 7288 4244 7328
rect 3532 7120 3572 7160
rect 3436 6868 3476 6908
rect 3340 6364 3380 6404
rect 4204 7120 4244 7160
rect 3820 7036 3860 7076
rect 3628 6448 3668 6488
rect 3820 6364 3860 6404
rect 3724 6196 3764 6236
rect 4012 6448 4052 6488
rect 5356 6952 5396 6992
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 5164 6616 5204 6656
rect 4876 6364 4916 6404
rect 6124 9304 6164 9344
rect 5932 8800 5972 8840
rect 6220 8800 6260 8840
rect 6412 8632 6452 8672
rect 6220 8464 6260 8504
rect 5836 8128 5876 8168
rect 6028 8128 6068 8168
rect 5740 7624 5780 7664
rect 5548 7456 5588 7496
rect 5452 6448 5492 6488
rect 6124 7960 6164 8000
rect 6316 7960 6356 8000
rect 6028 7624 6068 7664
rect 6124 7540 6164 7580
rect 5836 7120 5876 7160
rect 5932 6616 5972 6656
rect 5164 6364 5204 6404
rect 4204 6280 4244 6320
rect 4492 6280 4532 6320
rect 5068 6280 5108 6320
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 3148 5776 3188 5816
rect 3436 5776 3476 5816
rect 2956 4852 2996 4892
rect 3340 5608 3380 5648
rect 4300 6196 4340 6236
rect 3628 5440 3668 5480
rect 4108 5440 4148 5480
rect 4972 6196 5012 6236
rect 4972 5692 5012 5732
rect 3532 5272 3572 5312
rect 3436 5104 3476 5144
rect 3724 5272 3764 5312
rect 3724 5020 3764 5060
rect 3244 4936 3284 4976
rect 2764 3844 2804 3884
rect 2764 3592 2804 3632
rect 1804 3088 1844 3128
rect 2284 3088 2324 3128
rect 1708 2080 1748 2120
rect 1612 1324 1652 1364
rect 1420 904 1460 944
rect 1996 2836 2036 2876
rect 1804 1996 1844 2036
rect 1900 1912 1940 1952
rect 1900 1408 1940 1448
rect 2668 3424 2708 3464
rect 2572 2584 2612 2624
rect 2764 3172 2804 3212
rect 2956 3424 2996 3464
rect 2956 3088 2996 3128
rect 2860 2920 2900 2960
rect 2764 2584 2804 2624
rect 2668 1744 2708 1784
rect 3148 4096 3188 4136
rect 3436 4684 3476 4724
rect 4012 4684 4052 4724
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 3148 3844 3188 3884
rect 3148 2920 3188 2960
rect 3532 3928 3572 3968
rect 3244 2500 3284 2540
rect 3436 2584 3476 2624
rect 2956 2164 2996 2204
rect 3340 2164 3380 2204
rect 3244 2080 3284 2120
rect 3148 1912 3188 1952
rect 3628 3424 3668 3464
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 3916 2836 3956 2876
rect 3820 2752 3860 2792
rect 3628 2248 3668 2288
rect 3532 2164 3572 2204
rect 3724 1744 3764 1784
rect 3628 1660 3668 1700
rect 4012 1660 4052 1700
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 4300 5104 4340 5144
rect 4492 4971 4532 4976
rect 4492 4936 4532 4971
rect 4876 5608 4916 5648
rect 5452 6280 5492 6320
rect 5356 5608 5396 5648
rect 4972 5440 5012 5480
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 5068 5020 5108 5060
rect 5260 5020 5300 5060
rect 4204 4348 4244 4388
rect 4684 4348 4724 4388
rect 4588 4264 4628 4304
rect 4396 3508 4436 3548
rect 4492 3424 4532 3464
rect 4780 3928 4820 3968
rect 4684 3844 4724 3884
rect 4300 3340 4340 3380
rect 4300 2836 4340 2876
rect 4300 2668 4340 2708
rect 5356 3844 5396 3884
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 4972 3256 5012 3296
rect 4876 3172 4916 3212
rect 5548 3424 5588 3464
rect 5452 3256 5492 3296
rect 6220 6784 6260 6824
rect 6700 9472 6740 9512
rect 6604 9220 6644 9260
rect 6796 8800 6836 8840
rect 6508 8464 6548 8504
rect 6892 8632 6932 8672
rect 6892 8128 6932 8168
rect 6700 7960 6740 8000
rect 6700 7456 6740 7496
rect 6604 7036 6644 7076
rect 6412 6868 6452 6908
rect 6796 6868 6836 6908
rect 6220 6448 6260 6488
rect 6508 6532 6548 6572
rect 6988 7540 7028 7580
rect 7276 8800 7316 8840
rect 7468 8800 7508 8840
rect 7180 8548 7220 8588
rect 7276 8128 7316 8168
rect 7084 6868 7124 6908
rect 6892 6448 6932 6488
rect 6316 6112 6356 6152
rect 6220 4684 6260 4724
rect 6412 5272 6452 5312
rect 6412 4432 6452 4472
rect 6604 5020 6644 5060
rect 6604 4684 6644 4724
rect 6892 6028 6932 6068
rect 6796 5524 6836 5564
rect 6892 5188 6932 5228
rect 6796 5104 6836 5144
rect 6796 4936 6836 4976
rect 6988 4936 7028 4976
rect 7276 7876 7316 7916
rect 7276 7708 7316 7748
rect 7372 7624 7412 7664
rect 7276 7540 7316 7580
rect 7564 7708 7604 7748
rect 7756 7876 7796 7916
rect 7276 5020 7316 5060
rect 7180 4936 7220 4976
rect 7276 4852 7316 4892
rect 6700 4600 6740 4640
rect 6028 3508 6068 3548
rect 5740 3340 5780 3380
rect 5740 3172 5780 3212
rect 5068 2920 5108 2960
rect 4972 2584 5012 2624
rect 5356 2584 5396 2624
rect 4780 2500 4820 2540
rect 5356 2416 5396 2456
rect 4780 2248 4820 2288
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 4780 1996 4820 2036
rect 2764 1156 2804 1196
rect 4108 1240 4148 1280
rect 3148 1156 3188 1196
rect 3820 1072 3860 1112
rect 4588 1912 4628 1952
rect 5260 1156 5300 1196
rect 4300 1072 4340 1112
rect 5068 1072 5108 1112
rect 4204 820 4244 860
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 5548 2920 5588 2960
rect 5644 2752 5684 2792
rect 5548 2332 5588 2372
rect 5452 2080 5492 2120
rect 5452 1408 5492 1448
rect 6028 2920 6068 2960
rect 6220 3256 6260 3296
rect 6604 3424 6644 3464
rect 6892 4516 6932 4556
rect 6988 4012 7028 4052
rect 7180 4012 7220 4052
rect 6796 3928 6836 3968
rect 7084 3844 7124 3884
rect 6604 3256 6644 3296
rect 6508 3172 6548 3212
rect 5932 2584 5972 2624
rect 6316 2668 6356 2708
rect 6124 2332 6164 2372
rect 6028 2080 6068 2120
rect 6124 1912 6164 1952
rect 6412 1912 6452 1952
rect 6220 1744 6260 1784
rect 5740 1660 5780 1700
rect 5644 1156 5684 1196
rect 5452 1072 5492 1112
rect 6028 1576 6068 1616
rect 5836 1072 5876 1112
rect 6124 1492 6164 1532
rect 5452 736 5492 776
rect 6316 1660 6356 1700
rect 6700 2332 6740 2372
rect 6988 3172 7028 3212
rect 7180 3592 7220 3632
rect 6604 1660 6644 1700
rect 7372 4516 7412 4556
rect 7564 6616 7604 6656
rect 7660 6112 7700 6152
rect 8140 8800 8180 8840
rect 8140 8632 8180 8672
rect 8428 9220 8468 9260
rect 8332 8637 8372 8672
rect 8332 8632 8372 8637
rect 8332 8464 8372 8504
rect 8812 9472 8852 9512
rect 8524 8632 8564 8672
rect 8428 8128 8468 8168
rect 8236 7540 8276 7580
rect 8140 7372 8180 7412
rect 8044 7120 8084 7160
rect 7852 6616 7892 6656
rect 7564 5020 7604 5060
rect 7756 5020 7796 5060
rect 8140 6616 8180 6656
rect 8236 6532 8276 6572
rect 8140 6448 8180 6488
rect 8812 8716 8852 8756
rect 10252 9976 10292 10016
rect 9100 9556 9140 9596
rect 9484 9472 9524 9512
rect 10156 9472 10196 9512
rect 9100 9052 9140 9092
rect 9388 9052 9428 9092
rect 9100 8632 9140 8672
rect 9196 8128 9236 8168
rect 8812 7624 8852 7664
rect 8812 7036 8852 7076
rect 8812 6448 8852 6488
rect 8428 6280 8468 6320
rect 8236 5524 8276 5564
rect 8044 5272 8084 5312
rect 7948 5188 7988 5228
rect 7468 4012 7508 4052
rect 7372 3844 7412 3884
rect 7084 2500 7124 2540
rect 7372 3340 7412 3380
rect 7372 2500 7412 2540
rect 7276 2332 7316 2372
rect 7564 3928 7604 3968
rect 7564 3424 7604 3464
rect 8332 5188 8372 5228
rect 8524 5524 8564 5564
rect 8812 5440 8852 5480
rect 8524 5020 8564 5060
rect 8812 4971 8852 4976
rect 8812 4936 8852 4971
rect 8044 4684 8084 4724
rect 8428 4432 8468 4472
rect 8140 4180 8180 4220
rect 8332 4096 8372 4136
rect 8524 4264 8564 4304
rect 7948 3592 7988 3632
rect 8428 3760 8468 3800
rect 7660 2752 7700 2792
rect 7852 2584 7892 2624
rect 7852 2416 7892 2456
rect 7564 2164 7604 2204
rect 6988 1828 7028 1868
rect 6796 1660 6836 1700
rect 6892 1156 6932 1196
rect 8044 3424 8084 3464
rect 8332 3088 8372 3128
rect 7948 2248 7988 2288
rect 7756 1744 7796 1784
rect 7660 1660 7700 1700
rect 7180 1072 7220 1112
rect 8812 4348 8852 4388
rect 9100 7960 9140 8000
rect 9196 7708 9236 7748
rect 9004 5524 9044 5564
rect 9004 5020 9044 5060
rect 9580 9388 9620 9428
rect 9676 9304 9716 9344
rect 9580 8968 9620 9008
rect 9868 8800 9908 8840
rect 9964 8296 10004 8336
rect 9676 7876 9716 7916
rect 10348 9220 10388 9260
rect 10540 9976 10580 10016
rect 10252 8800 10292 8840
rect 10732 8968 10772 9008
rect 10540 8464 10580 8504
rect 10444 8128 10484 8168
rect 10924 9388 10964 9428
rect 11404 9808 11444 9848
rect 11212 9304 11252 9344
rect 11212 9052 11252 9092
rect 11020 8716 11060 8756
rect 10636 8044 10676 8084
rect 10252 7372 10292 7412
rect 9484 7120 9524 7160
rect 9388 6784 9428 6824
rect 9676 6952 9716 6992
rect 9580 5692 9620 5732
rect 9772 6448 9812 6488
rect 9484 4600 9524 4640
rect 9388 4516 9428 4556
rect 9772 4936 9812 4976
rect 10732 7708 10772 7748
rect 10636 7204 10676 7244
rect 10924 8044 10964 8084
rect 10924 7624 10964 7664
rect 10636 6952 10676 6992
rect 10060 6280 10100 6320
rect 9964 5860 10004 5900
rect 9998 5692 10038 5732
rect 10156 5440 10196 5480
rect 10060 5188 10100 5228
rect 10732 6448 10772 6488
rect 10828 6280 10868 6320
rect 10540 6112 10580 6152
rect 11116 7792 11156 7832
rect 11020 6616 11060 6656
rect 11308 7708 11348 7748
rect 11404 6532 11444 6572
rect 11116 6280 11156 6320
rect 11020 5944 11060 5984
rect 10540 5860 10580 5900
rect 10540 5692 10580 5732
rect 10156 4936 10196 4976
rect 9388 4264 9428 4304
rect 9100 4180 9140 4220
rect 8812 3760 8852 3800
rect 8716 3592 8756 3632
rect 8908 3592 8948 3632
rect 9388 3508 9428 3548
rect 9100 3424 9140 3464
rect 8716 3088 8756 3128
rect 8140 2416 8180 2456
rect 8332 2164 8372 2204
rect 8524 2164 8564 2204
rect 8140 1828 8180 1868
rect 8524 1744 8564 1784
rect 8140 1408 8180 1448
rect 8044 1240 8084 1280
rect 7852 1072 7892 1112
rect 9100 2668 9140 2708
rect 9292 3172 9332 3212
rect 9292 2920 9332 2960
rect 9676 4180 9716 4220
rect 9580 4096 9620 4136
rect 9772 4012 9812 4052
rect 9580 3844 9620 3884
rect 9484 2836 9524 2876
rect 9388 2584 9428 2624
rect 9196 2416 9236 2456
rect 9292 2332 9332 2372
rect 9484 2332 9524 2372
rect 9868 3676 9908 3716
rect 9676 3256 9716 3296
rect 9772 3172 9812 3212
rect 9676 3088 9716 3128
rect 9772 2332 9812 2372
rect 9580 1240 9620 1280
rect 9772 1072 9812 1112
rect 7564 904 7604 944
rect 6124 400 6164 440
rect 6412 148 6452 188
rect 8716 820 8756 860
rect 8620 652 8660 692
rect 9388 736 9428 776
rect 10444 4768 10484 4808
rect 10348 4600 10388 4640
rect 10252 4348 10292 4388
rect 10348 4264 10388 4304
rect 9964 3088 10004 3128
rect 10924 5776 10964 5816
rect 10828 5692 10868 5732
rect 10636 5188 10676 5228
rect 10732 5020 10772 5060
rect 10636 4936 10676 4976
rect 10732 4432 10772 4472
rect 10156 3928 10196 3968
rect 10348 3760 10388 3800
rect 10252 3508 10292 3548
rect 10252 2752 10292 2792
rect 10156 2668 10196 2708
rect 10060 2416 10100 2456
rect 10060 1996 10100 2036
rect 10348 2584 10388 2624
rect 10348 1240 10388 1280
rect 10540 3844 10580 3884
rect 10732 3928 10772 3968
rect 10636 3592 10676 3632
rect 10924 3508 10964 3548
rect 10828 3424 10868 3464
rect 10636 3172 10676 3212
rect 10636 2836 10676 2876
rect 10828 3004 10868 3044
rect 10732 2752 10772 2792
rect 10924 2500 10964 2540
rect 10924 2080 10964 2120
rect 10732 1240 10772 1280
rect 11308 5272 11348 5312
rect 11884 10312 11924 10352
rect 11788 8968 11828 9008
rect 11596 8464 11636 8504
rect 12268 10564 12308 10604
rect 12172 10312 12212 10352
rect 12172 10144 12212 10184
rect 11980 8716 12020 8756
rect 11788 7456 11828 7496
rect 11596 6700 11636 6740
rect 11692 5692 11732 5732
rect 11596 5188 11636 5228
rect 11212 3088 11252 3128
rect 11596 3676 11636 3716
rect 11500 3424 11540 3464
rect 11404 3340 11444 3380
rect 11308 2752 11348 2792
rect 11212 2416 11252 2456
rect 11596 2080 11636 2120
rect 11404 1912 11444 1952
rect 10444 820 10484 860
rect 11212 1240 11252 1280
rect 12172 8380 12212 8420
rect 12076 7540 12116 7580
rect 11980 6280 12020 6320
rect 11788 5188 11828 5228
rect 12556 10144 12596 10184
rect 13036 9472 13076 9512
rect 12460 9304 12500 9344
rect 12364 8968 12404 9008
rect 12268 6280 12308 6320
rect 12748 9052 12788 9092
rect 12844 7960 12884 8000
rect 12652 7540 12692 7580
rect 12844 7204 12884 7244
rect 12748 6868 12788 6908
rect 12460 6616 12500 6656
rect 12652 6448 12692 6488
rect 12364 6196 12404 6236
rect 12652 6028 12692 6068
rect 12076 5188 12116 5228
rect 11980 4600 12020 4640
rect 11980 4180 12020 4220
rect 12172 4180 12212 4220
rect 11788 4096 11828 4136
rect 11884 3928 11924 3968
rect 12268 3928 12308 3968
rect 12460 4516 12500 4556
rect 12364 3760 12404 3800
rect 12076 3424 12116 3464
rect 12940 5524 12980 5564
rect 12844 4600 12884 4640
rect 12748 4180 12788 4220
rect 12556 4096 12596 4136
rect 12940 4012 12980 4052
rect 13228 9556 13268 9596
rect 13228 9388 13268 9428
rect 13900 9892 13940 9932
rect 14092 9472 14132 9512
rect 13804 8884 13844 8924
rect 13516 8800 13556 8840
rect 13708 8800 13748 8840
rect 14668 10564 14708 10604
rect 14956 10564 14996 10604
rect 14860 9724 14900 9764
rect 14284 8800 14324 8840
rect 13612 7708 13652 7748
rect 13420 7036 13460 7076
rect 13420 6868 13460 6908
rect 13324 6616 13364 6656
rect 13324 4936 13364 4976
rect 13228 4180 13268 4220
rect 13036 3592 13076 3632
rect 12556 3424 12596 3464
rect 11884 2920 11924 2960
rect 11980 2416 12020 2456
rect 11788 2080 11828 2120
rect 11884 1996 11924 2036
rect 11788 1828 11828 1868
rect 11500 1156 11540 1196
rect 10924 736 10964 776
rect 11692 1072 11732 1112
rect 12268 2584 12308 2624
rect 12268 1912 12308 1952
rect 12940 2584 12980 2624
rect 12652 2332 12692 2372
rect 12556 1996 12596 2036
rect 12748 2164 12788 2204
rect 12460 1828 12500 1868
rect 12172 1156 12212 1196
rect 12172 904 12212 944
rect 12652 1408 12692 1448
rect 12460 1240 12500 1280
rect 12748 1240 12788 1280
rect 12364 1072 12404 1112
rect 12556 1072 12596 1112
rect 12844 1072 12884 1112
rect 13036 1912 13076 1952
rect 13420 3928 13460 3968
rect 13324 2752 13364 2792
rect 12652 820 12692 860
rect 12268 232 12308 272
rect 13900 8548 13940 8588
rect 13996 8296 14036 8336
rect 14668 8296 14708 8336
rect 14188 7708 14228 7748
rect 14380 7456 14420 7496
rect 13804 7288 13844 7328
rect 13900 7120 13940 7160
rect 14956 9388 14996 9428
rect 15244 10144 15284 10184
rect 15244 9976 15284 10016
rect 15148 9640 15188 9680
rect 15340 9388 15380 9428
rect 15244 9052 15284 9092
rect 15052 8800 15092 8840
rect 15148 8632 15188 8672
rect 13900 6952 13940 6992
rect 14284 6448 14324 6488
rect 13900 6280 13940 6320
rect 13996 5776 14036 5816
rect 14284 5608 14324 5648
rect 14476 5440 14516 5480
rect 13996 5356 14036 5396
rect 13612 5020 13652 5060
rect 14092 5020 14132 5060
rect 13996 4348 14036 4388
rect 13804 3928 13844 3968
rect 13804 3508 13844 3548
rect 14284 4180 14324 4220
rect 14188 3592 14228 3632
rect 14380 3340 14420 3380
rect 14284 3088 14324 3128
rect 14284 2668 14324 2708
rect 13804 1156 13844 1196
rect 13996 1072 14036 1112
rect 14860 4768 14900 4808
rect 14764 4348 14804 4388
rect 14668 4264 14708 4304
rect 15052 7204 15092 7244
rect 15244 8296 15284 8336
rect 15148 6616 15188 6656
rect 15820 10480 15860 10520
rect 15916 10060 15956 10100
rect 15436 8800 15476 8840
rect 15820 8800 15860 8840
rect 15532 8128 15572 8168
rect 15724 8548 15764 8588
rect 15628 8044 15668 8084
rect 15436 7960 15476 8000
rect 15724 7456 15764 7496
rect 15532 7204 15572 7244
rect 15340 7036 15380 7076
rect 15532 6952 15572 6992
rect 15340 6616 15380 6656
rect 15244 6280 15284 6320
rect 15148 5020 15188 5060
rect 16492 9808 16532 9848
rect 16396 9640 16436 9680
rect 16300 9556 16340 9596
rect 16876 10312 16916 10352
rect 16588 9472 16628 9512
rect 16300 9304 16340 9344
rect 16492 9052 16532 9092
rect 15916 6700 15956 6740
rect 15628 5272 15668 5312
rect 15244 4852 15284 4892
rect 15148 3508 15188 3548
rect 14764 3424 14804 3464
rect 14668 3172 14708 3212
rect 14764 2920 14804 2960
rect 14572 1828 14612 1868
rect 14572 1492 14612 1532
rect 15532 3760 15572 3800
rect 15532 3256 15572 3296
rect 15820 5020 15860 5060
rect 15916 3928 15956 3968
rect 16588 6364 16628 6404
rect 16492 5776 16532 5816
rect 16492 5608 16532 5648
rect 16492 5356 16532 5396
rect 16012 3760 16052 3800
rect 16300 3928 16340 3968
rect 16780 9388 16820 9428
rect 17068 9640 17108 9680
rect 16780 9052 16820 9092
rect 16972 9052 17012 9092
rect 16876 8632 16916 8672
rect 16972 8464 17012 8504
rect 16780 6700 16820 6740
rect 17260 9808 17300 9848
rect 17164 8800 17204 8840
rect 17164 7960 17204 8000
rect 17164 6952 17204 6992
rect 17068 6448 17108 6488
rect 16780 6028 16820 6068
rect 17068 5776 17108 5816
rect 16780 5020 16820 5060
rect 17068 4768 17108 4808
rect 16780 4684 16820 4724
rect 16972 4684 17012 4724
rect 16492 4348 16532 4388
rect 16684 4348 16724 4388
rect 17356 9472 17396 9512
rect 17452 8548 17492 8588
rect 17644 9640 17684 9680
rect 17644 9388 17684 9428
rect 17548 7960 17588 8000
rect 18124 10480 18164 10520
rect 18028 9808 18068 9848
rect 17932 9556 17972 9596
rect 18508 9808 18548 9848
rect 17836 9220 17876 9260
rect 17740 8884 17780 8924
rect 17836 8380 17876 8420
rect 18316 8464 18356 8504
rect 17836 7540 17876 7580
rect 17452 7456 17492 7496
rect 17740 7372 17780 7412
rect 17644 7120 17684 7160
rect 17356 6784 17396 6824
rect 17260 6280 17300 6320
rect 17452 6448 17492 6488
rect 17644 6952 17684 6992
rect 18412 8380 18452 8420
rect 17836 6784 17876 6824
rect 16972 4432 17012 4472
rect 17356 4936 17396 4976
rect 17548 6280 17588 6320
rect 17740 5860 17780 5900
rect 17548 5020 17588 5060
rect 16972 4180 17012 4220
rect 16012 3508 16052 3548
rect 16972 3424 17012 3464
rect 15340 2248 15380 2288
rect 15244 904 15284 944
rect 16684 2836 16724 2876
rect 16684 2668 16724 2708
rect 16204 2584 16244 2624
rect 16588 2584 16628 2624
rect 15820 2080 15860 2120
rect 16300 2500 16340 2540
rect 16780 1996 16820 2036
rect 15916 1912 15956 1952
rect 16204 1828 16244 1868
rect 15916 1492 15956 1532
rect 15820 1156 15860 1196
rect 16780 1240 16820 1280
rect 15820 736 15860 776
rect 17260 3928 17300 3968
rect 17164 2836 17204 2876
rect 17548 4852 17588 4892
rect 18316 7120 18356 7160
rect 18124 6028 18164 6068
rect 18892 9220 18932 9260
rect 19372 10396 19412 10436
rect 19276 9388 19316 9428
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 18892 8800 18932 8840
rect 18700 8212 18740 8252
rect 18988 8464 19028 8504
rect 19180 7960 19220 8000
rect 19180 7708 19220 7748
rect 18508 7624 18548 7664
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 19180 7372 19220 7412
rect 18604 7204 18644 7244
rect 19180 6784 19220 6824
rect 18604 6616 18644 6656
rect 18988 6364 19028 6404
rect 18604 6196 18644 6236
rect 18412 5944 18452 5984
rect 18124 5524 18164 5564
rect 17548 3424 17588 3464
rect 18028 5020 18068 5060
rect 17836 4852 17876 4892
rect 18316 4852 18356 4892
rect 18028 4768 18068 4808
rect 18220 3424 18260 3464
rect 17836 2416 17876 2456
rect 17452 2332 17492 2372
rect 18508 4936 18548 4976
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 19180 5692 19220 5732
rect 19180 5356 19220 5396
rect 19180 4936 19220 4976
rect 18796 4852 18836 4892
rect 19468 9640 19508 9680
rect 19468 9472 19508 9512
rect 19372 8800 19412 8840
rect 19660 8800 19700 8840
rect 19372 8296 19412 8336
rect 19372 7876 19412 7916
rect 20236 10648 20276 10688
rect 20044 9976 20084 10016
rect 20236 9976 20276 10016
rect 20620 10060 20660 10100
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 20332 9640 20372 9680
rect 20140 8716 20180 8756
rect 20812 9808 20852 9848
rect 21292 9892 21332 9932
rect 21196 9640 21236 9680
rect 20716 9472 20756 9512
rect 20428 8464 20468 8504
rect 19948 8296 19988 8336
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 19756 8044 19796 8084
rect 19564 7960 19604 8000
rect 19468 7792 19508 7832
rect 19564 7540 19604 7580
rect 19468 7204 19508 7244
rect 19372 7120 19412 7160
rect 19564 6364 19604 6404
rect 19468 5944 19508 5984
rect 19372 5860 19412 5900
rect 19948 7792 19988 7832
rect 19852 7036 19892 7076
rect 19756 6364 19796 6404
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 19372 4516 19412 4556
rect 18412 4096 18452 4136
rect 18412 3424 18452 3464
rect 18604 3760 18644 3800
rect 18508 3004 18548 3044
rect 18892 3844 18932 3884
rect 18700 3508 18740 3548
rect 19180 3676 19220 3716
rect 19084 3592 19124 3632
rect 18892 3424 18932 3464
rect 19276 3508 19316 3548
rect 19180 3172 19220 3212
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 17836 1912 17876 1952
rect 19756 5524 19796 5564
rect 19756 5188 19796 5228
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 20620 8800 20660 8840
rect 20908 9220 20948 9260
rect 20908 8464 20948 8504
rect 20812 7708 20852 7748
rect 20716 7540 20756 7580
rect 20620 6532 20660 6572
rect 20524 5860 20564 5900
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 20428 5104 20468 5144
rect 20236 4768 20276 4808
rect 19852 4180 19892 4220
rect 20332 4180 20372 4220
rect 19660 3844 19700 3884
rect 20812 5440 20852 5480
rect 20812 5104 20852 5144
rect 21292 8800 21332 8840
rect 21004 7120 21044 7160
rect 21676 10060 21716 10100
rect 21580 9976 21620 10016
rect 21484 9808 21524 9848
rect 21196 5692 21236 5732
rect 21004 5440 21044 5480
rect 20428 4012 20468 4052
rect 19948 3760 19988 3800
rect 19660 3508 19700 3548
rect 19468 3172 19508 3212
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 19852 3592 19892 3632
rect 20044 3424 20084 3464
rect 19756 2752 19796 2792
rect 20428 2500 20468 2540
rect 19276 2332 19316 2372
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 19564 1912 19604 1952
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 18700 1324 18740 1364
rect 19084 1324 19124 1364
rect 17452 1156 17492 1196
rect 17932 1156 17972 1196
rect 18892 1156 18932 1196
rect 17644 1072 17684 1112
rect 17164 820 17204 860
rect 21004 3760 21044 3800
rect 21100 3508 21140 3548
rect 21100 3004 21140 3044
rect 21004 2668 21044 2708
rect 20908 2332 20948 2372
rect 21388 5356 21428 5396
rect 21292 4684 21332 4724
rect 21484 4096 21524 4136
rect 21292 3088 21332 3128
rect 21676 9640 21716 9680
rect 21964 10060 22004 10100
rect 22348 10564 22388 10604
rect 22156 9808 22196 9848
rect 22348 9808 22388 9848
rect 22156 9640 22196 9680
rect 21772 9220 21812 9260
rect 21676 9052 21716 9092
rect 21868 8884 21908 8924
rect 21868 8632 21908 8672
rect 21868 8296 21908 8336
rect 22444 8716 22484 8756
rect 22348 8548 22388 8588
rect 22252 8296 22292 8336
rect 22060 7960 22100 8000
rect 22060 7708 22100 7748
rect 21868 7624 21908 7664
rect 21676 7288 21716 7328
rect 21676 4348 21716 4388
rect 21964 4180 22004 4220
rect 21868 3844 21908 3884
rect 21676 3760 21716 3800
rect 21580 3172 21620 3212
rect 21868 2584 21908 2624
rect 22924 9892 22964 9932
rect 22540 7624 22580 7664
rect 22828 8800 22868 8840
rect 22828 8632 22868 8672
rect 23308 9472 23348 9512
rect 22924 8464 22964 8504
rect 22828 8380 22868 8420
rect 23212 8800 23252 8840
rect 23692 10312 23732 10352
rect 23500 8800 23540 8840
rect 23212 8464 23252 8504
rect 22348 7288 22388 7328
rect 22156 7120 22196 7160
rect 22252 6784 22292 6824
rect 22636 7120 22676 7160
rect 22636 6784 22676 6824
rect 22540 5944 22580 5984
rect 23212 8128 23252 8168
rect 23020 8044 23060 8084
rect 24364 9976 24404 10016
rect 24268 9892 24308 9932
rect 24172 8800 24212 8840
rect 23980 8044 24020 8084
rect 24076 7960 24116 8000
rect 23884 7624 23924 7664
rect 23788 7540 23828 7580
rect 22924 7036 22964 7076
rect 23212 6700 23252 6740
rect 22636 5440 22676 5480
rect 22540 5356 22580 5396
rect 22732 4852 22772 4892
rect 22348 4768 22388 4808
rect 22924 5104 22964 5144
rect 22828 4516 22868 4556
rect 23308 6364 23348 6404
rect 23500 5104 23540 5144
rect 23212 4264 23252 4304
rect 22444 3844 22484 3884
rect 24076 5104 24116 5144
rect 23692 4852 23732 4892
rect 22540 3592 22580 3632
rect 22444 3256 22484 3296
rect 21388 2332 21428 2372
rect 20524 1324 20564 1364
rect 20908 1324 20948 1364
rect 21196 1912 21236 1952
rect 21004 1156 21044 1196
rect 19084 904 19124 944
rect 21100 1072 21140 1112
rect 21196 988 21236 1028
rect 21388 988 21428 1028
rect 21292 904 21332 944
rect 19948 820 19988 860
rect 19468 484 19508 524
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 19948 64 19988 104
rect 20236 64 20276 104
rect 23404 3172 23444 3212
rect 22636 2584 22676 2624
rect 23308 2584 23348 2624
rect 24364 9220 24404 9260
rect 24748 9892 24788 9932
rect 24652 9556 24692 9596
rect 24556 9304 24596 9344
rect 24460 9052 24500 9092
rect 24364 8968 24404 9008
rect 24556 8968 24596 9008
rect 24364 8800 24404 8840
rect 24556 8800 24596 8840
rect 24460 7540 24500 7580
rect 25036 10564 25076 10604
rect 25420 10648 25460 10688
rect 24940 10480 24980 10520
rect 25228 10480 25268 10520
rect 25420 9472 25460 9512
rect 25420 9220 25460 9260
rect 24844 8800 24884 8840
rect 25324 8380 25364 8420
rect 24940 8128 24980 8168
rect 24844 7708 24884 7748
rect 24556 7372 24596 7412
rect 24748 7372 24788 7412
rect 24364 5608 24404 5648
rect 24268 4936 24308 4976
rect 24748 7120 24788 7160
rect 24652 6784 24692 6824
rect 24556 6112 24596 6152
rect 24460 5104 24500 5144
rect 25804 9052 25844 9092
rect 25324 7624 25364 7664
rect 24940 6784 24980 6824
rect 25036 6616 25076 6656
rect 24748 6364 24788 6404
rect 24844 6196 24884 6236
rect 24652 4936 24692 4976
rect 24076 4180 24116 4220
rect 24076 4012 24116 4052
rect 23884 3760 23924 3800
rect 24460 4684 24500 4724
rect 24268 4264 24308 4304
rect 24172 3508 24212 3548
rect 23692 3004 23732 3044
rect 23884 3004 23924 3044
rect 24076 3004 24116 3044
rect 23788 2668 23828 2708
rect 23500 2332 23540 2372
rect 22348 988 22388 1028
rect 22828 1912 22868 1952
rect 24076 1912 24116 1952
rect 23020 1828 23060 1868
rect 23500 1828 23540 1868
rect 24364 2752 24404 2792
rect 24556 4264 24596 4304
rect 24556 3172 24596 3212
rect 24556 2752 24596 2792
rect 25132 6112 25172 6152
rect 24940 5440 24980 5480
rect 24844 4684 24884 4724
rect 24748 3844 24788 3884
rect 25708 8212 25748 8252
rect 26572 9976 26612 10016
rect 26380 9892 26420 9932
rect 27148 10396 27188 10436
rect 27052 9724 27092 9764
rect 26572 9304 26612 9344
rect 25612 6616 25652 6656
rect 25996 7624 26036 7664
rect 26284 8884 26324 8924
rect 26476 8800 26516 8840
rect 26572 8548 26612 8588
rect 26380 8296 26420 8336
rect 26188 7624 26228 7664
rect 26092 6364 26132 6404
rect 25996 5608 26036 5648
rect 26092 5356 26132 5396
rect 25516 5020 25556 5060
rect 25900 4936 25940 4976
rect 25036 4012 25076 4052
rect 25612 3844 25652 3884
rect 24748 3676 24788 3716
rect 24940 3508 24980 3548
rect 25036 3340 25076 3380
rect 25516 3424 25556 3464
rect 25228 3340 25268 3380
rect 24940 3256 24980 3296
rect 24940 3004 24980 3044
rect 24652 2668 24692 2708
rect 24268 1912 24308 1952
rect 24172 1492 24212 1532
rect 23020 1408 23060 1448
rect 22828 1324 22868 1364
rect 24460 1576 24500 1616
rect 24748 2080 24788 2120
rect 24748 1744 24788 1784
rect 25132 3088 25172 3128
rect 25324 3256 25364 3296
rect 25516 2920 25556 2960
rect 26092 2836 26132 2876
rect 26092 1996 26132 2036
rect 25708 1828 25748 1868
rect 25900 1576 25940 1616
rect 25228 1492 25268 1532
rect 25900 1240 25940 1280
rect 26092 1240 26132 1280
rect 26284 4516 26324 4556
rect 26284 3928 26324 3968
rect 26956 9136 26996 9176
rect 26956 8632 26996 8672
rect 27244 9388 27284 9428
rect 27532 9640 27572 9680
rect 27628 9388 27668 9428
rect 27340 8212 27380 8252
rect 27052 7120 27092 7160
rect 26764 6868 26804 6908
rect 26668 6448 26708 6488
rect 26572 5692 26612 5732
rect 26572 4936 26612 4976
rect 27148 6700 27188 6740
rect 27148 6448 27188 6488
rect 27148 4936 27188 4976
rect 27340 7540 27380 7580
rect 27916 10060 27956 10100
rect 28012 8716 28052 8756
rect 28300 8716 28340 8756
rect 27916 8296 27956 8336
rect 27820 7960 27860 8000
rect 28396 8632 28436 8672
rect 28684 8716 28724 8756
rect 28972 9052 29012 9092
rect 28876 8632 28916 8672
rect 28780 8464 28820 8504
rect 28588 8296 28628 8336
rect 28492 8212 28532 8252
rect 28396 7995 28436 8000
rect 28396 7960 28436 7995
rect 28300 7792 28340 7832
rect 28108 7624 28148 7664
rect 27724 7540 27764 7580
rect 28204 7540 28244 7580
rect 27916 6952 27956 6992
rect 27916 6448 27956 6488
rect 27628 6280 27668 6320
rect 27436 5692 27476 5732
rect 27340 5608 27380 5648
rect 27052 4180 27092 4220
rect 27244 4180 27284 4220
rect 27148 3844 27188 3884
rect 26572 3424 26612 3464
rect 26764 3424 26804 3464
rect 26476 3340 26516 3380
rect 27052 3004 27092 3044
rect 26668 2836 26708 2876
rect 27052 2668 27092 2708
rect 26284 2080 26324 2120
rect 26476 1996 26516 2036
rect 27244 2164 27284 2204
rect 26668 1912 26708 1952
rect 26284 1324 26324 1364
rect 26188 1156 26228 1196
rect 26092 1072 26132 1112
rect 26284 1072 26324 1112
rect 25996 988 26036 1028
rect 22444 820 22484 860
rect 24844 820 24884 860
rect 23692 232 23732 272
rect 24844 148 24884 188
rect 27148 904 27188 944
rect 27436 5524 27476 5564
rect 27916 5692 27956 5732
rect 28012 5440 28052 5480
rect 27628 5272 27668 5312
rect 27916 5272 27956 5312
rect 27436 5104 27476 5144
rect 27916 4936 27956 4976
rect 27628 4684 27668 4724
rect 27724 4600 27764 4640
rect 27532 4432 27572 4472
rect 27436 4096 27476 4136
rect 27628 4264 27668 4304
rect 27628 4096 27668 4136
rect 27820 4264 27860 4304
rect 28300 7372 28340 7412
rect 28588 8044 28628 8084
rect 28588 7708 28628 7748
rect 28588 6868 28628 6908
rect 28780 8128 28820 8168
rect 28780 7960 28820 8000
rect 28780 7624 28820 7664
rect 28684 6700 28724 6740
rect 28588 6616 28628 6656
rect 28300 6364 28340 6404
rect 28204 4852 28244 4892
rect 28492 6448 28532 6488
rect 28396 4264 28436 4304
rect 27436 3844 27476 3884
rect 27436 3424 27476 3464
rect 27724 2836 27764 2876
rect 28396 3928 28436 3968
rect 28204 3676 28244 3716
rect 28396 3424 28436 3464
rect 28300 3340 28340 3380
rect 28012 2836 28052 2876
rect 28108 2668 28148 2708
rect 28588 6196 28628 6236
rect 28588 4348 28628 4388
rect 28588 3676 28628 3716
rect 28876 6616 28916 6656
rect 29164 9724 29204 9764
rect 29260 9388 29300 9428
rect 29356 9304 29396 9344
rect 29164 9220 29204 9260
rect 29068 8800 29108 8840
rect 29452 9052 29492 9092
rect 29740 9388 29780 9428
rect 29452 7708 29492 7748
rect 29068 7204 29108 7244
rect 28876 6448 28916 6488
rect 28780 4684 28820 4724
rect 28780 3928 28820 3968
rect 28684 1912 28724 1952
rect 28972 3928 29012 3968
rect 28972 3424 29012 3464
rect 29644 8464 29684 8504
rect 29356 6700 29396 6740
rect 29164 5524 29204 5564
rect 29260 4768 29300 4808
rect 29164 4348 29204 4388
rect 29356 3172 29396 3212
rect 29548 6784 29588 6824
rect 29548 5608 29588 5648
rect 29836 8884 29876 8924
rect 30124 9556 30164 9596
rect 30412 9640 30452 9680
rect 29836 8716 29876 8756
rect 29836 8380 29876 8420
rect 30028 7960 30068 8000
rect 30316 8548 30356 8588
rect 30892 9640 30932 9680
rect 30796 9556 30836 9596
rect 30604 9388 30644 9428
rect 30796 9220 30836 9260
rect 30508 8884 30548 8924
rect 30700 8800 30740 8840
rect 30604 8464 30644 8504
rect 29836 7204 29876 7244
rect 30220 7120 30260 7160
rect 29932 6868 29972 6908
rect 29740 6280 29780 6320
rect 30124 6784 30164 6824
rect 30028 5776 30068 5816
rect 30604 7708 30644 7748
rect 30220 6280 30260 6320
rect 30124 5356 30164 5396
rect 30220 5272 30260 5312
rect 29644 4852 29684 4892
rect 30988 8884 31028 8924
rect 30988 8632 31028 8672
rect 30988 7960 31028 8000
rect 30988 7204 31028 7244
rect 31180 9388 31220 9428
rect 31180 7960 31220 8000
rect 30796 6280 30836 6320
rect 31180 6280 31220 6320
rect 30412 4852 30452 4892
rect 29740 4768 29780 4808
rect 30316 4768 30356 4808
rect 29356 2752 29396 2792
rect 28972 2332 29012 2372
rect 29260 2584 29300 2624
rect 29164 2080 29204 2120
rect 29548 2584 29588 2624
rect 30700 5188 30740 5228
rect 30892 5020 30932 5060
rect 30796 4600 30836 4640
rect 30028 3760 30068 3800
rect 29932 3508 29972 3548
rect 29836 3340 29876 3380
rect 29932 3004 29972 3044
rect 29932 2584 29972 2624
rect 29644 2248 29684 2288
rect 29548 1576 29588 1616
rect 29356 1492 29396 1532
rect 27820 1240 27860 1280
rect 28876 1240 28916 1280
rect 28300 1156 28340 1196
rect 27340 820 27380 860
rect 28108 820 28148 860
rect 30700 3760 30740 3800
rect 30316 3424 30356 3464
rect 30604 3424 30644 3464
rect 30220 3340 30260 3380
rect 30220 3004 30260 3044
rect 29932 1996 29972 2036
rect 29836 1324 29876 1364
rect 29740 820 29780 860
rect 30124 2080 30164 2120
rect 31372 9136 31412 9176
rect 31852 9556 31892 9596
rect 32332 9640 32372 9680
rect 31852 8884 31892 8924
rect 31564 8632 31604 8672
rect 31372 8548 31412 8588
rect 31660 8380 31700 8420
rect 31564 8212 31604 8252
rect 31372 7456 31412 7496
rect 31468 7372 31508 7412
rect 31468 7204 31508 7244
rect 31660 6700 31700 6740
rect 31564 6616 31604 6656
rect 32044 9220 32084 9260
rect 32140 9052 32180 9092
rect 32044 8464 32084 8504
rect 31948 8128 31988 8168
rect 31948 7960 31988 8000
rect 32044 7708 32084 7748
rect 31852 7624 31892 7664
rect 31948 7456 31988 7496
rect 31852 7372 31892 7412
rect 32044 7372 32084 7412
rect 31948 6616 31988 6656
rect 31084 5356 31124 5396
rect 30988 2332 31028 2372
rect 30988 1072 31028 1112
rect 30220 820 30260 860
rect 30892 820 30932 860
rect 29452 64 29492 104
rect 30028 64 30068 104
rect 30604 64 30644 104
rect 30796 64 30836 104
rect 31180 5272 31220 5312
rect 31276 4936 31316 4976
rect 31180 3844 31220 3884
rect 31852 5944 31892 5984
rect 31468 3760 31508 3800
rect 31468 3256 31508 3296
rect 31468 2836 31508 2876
rect 31756 4012 31796 4052
rect 31660 3760 31700 3800
rect 31852 3256 31892 3296
rect 32620 9220 32660 9260
rect 32524 8968 32564 9008
rect 32812 9640 32852 9680
rect 33292 9220 33332 9260
rect 33196 9052 33236 9092
rect 33100 8968 33140 9008
rect 32428 8800 32468 8840
rect 32716 8800 32756 8840
rect 32332 8296 32372 8336
rect 32716 8464 32756 8504
rect 32524 8380 32564 8420
rect 32620 8296 32660 8336
rect 32524 8212 32564 8252
rect 32524 8044 32564 8084
rect 32236 7624 32276 7664
rect 32428 7624 32468 7664
rect 32140 6700 32180 6740
rect 32140 6364 32180 6404
rect 32044 4600 32084 4640
rect 32524 5608 32564 5648
rect 32428 5356 32468 5396
rect 32428 4852 32468 4892
rect 32332 4432 32372 4472
rect 32236 3424 32276 3464
rect 32236 3004 32276 3044
rect 31564 2584 31604 2624
rect 31756 2248 31796 2288
rect 31564 1996 31604 2036
rect 31372 1744 31412 1784
rect 31756 1660 31796 1700
rect 31564 1492 31604 1532
rect 31564 1324 31604 1364
rect 31276 1240 31316 1280
rect 31468 1240 31508 1280
rect 31468 820 31508 860
rect 32524 4600 32564 4640
rect 32716 6784 32756 6824
rect 33388 8548 33428 8588
rect 39628 10648 39668 10688
rect 35884 10564 35924 10604
rect 34924 10480 34964 10520
rect 34444 9640 34484 9680
rect 34060 9472 34100 9512
rect 33928 9052 33968 9092
rect 34010 9052 34050 9092
rect 34092 9052 34132 9092
rect 34174 9052 34214 9092
rect 34256 9052 34296 9092
rect 34444 9052 34484 9092
rect 33772 8632 33812 8672
rect 34348 8632 34388 8672
rect 33868 8548 33908 8588
rect 34348 8212 34388 8252
rect 34060 8128 34100 8168
rect 33292 7624 33332 7664
rect 33196 7372 33236 7412
rect 32908 6868 32948 6908
rect 33100 6532 33140 6572
rect 32908 6364 32948 6404
rect 32812 6196 32852 6236
rect 32812 5608 32852 5648
rect 32716 5272 32756 5312
rect 33676 7792 33716 7832
rect 33580 7708 33620 7748
rect 33676 7372 33716 7412
rect 33676 6616 33716 6656
rect 33196 5608 33236 5648
rect 32908 4684 32948 4724
rect 32812 4096 32852 4136
rect 32620 3592 32660 3632
rect 32908 3424 32948 3464
rect 33100 4852 33140 4892
rect 33196 4264 33236 4304
rect 33292 4180 33332 4220
rect 33196 3844 33236 3884
rect 33100 3676 33140 3716
rect 33100 3340 33140 3380
rect 33292 2668 33332 2708
rect 33580 6196 33620 6236
rect 33484 5104 33524 5144
rect 33484 3424 33524 3464
rect 32812 2248 32852 2288
rect 33196 2248 33236 2288
rect 33388 2080 33428 2120
rect 33388 1912 33428 1952
rect 32524 1828 32564 1868
rect 32908 1828 32948 1868
rect 32812 1240 32852 1280
rect 32236 1156 32276 1196
rect 31852 988 31892 1028
rect 32620 232 32660 272
rect 33388 1072 33428 1112
rect 33868 8044 33908 8084
rect 33868 7876 33908 7916
rect 33928 7540 33968 7580
rect 34010 7540 34050 7580
rect 34092 7540 34132 7580
rect 34174 7540 34214 7580
rect 34256 7540 34296 7580
rect 33772 6280 33812 6320
rect 34732 8716 34772 8756
rect 35168 9808 35208 9848
rect 35250 9808 35290 9848
rect 35332 9808 35372 9848
rect 35414 9808 35454 9848
rect 35496 9808 35536 9848
rect 35692 9724 35732 9764
rect 35692 9388 35732 9428
rect 37612 10480 37652 10520
rect 35980 9640 36020 9680
rect 37324 9640 37364 9680
rect 35596 8968 35636 9008
rect 35884 8968 35924 9008
rect 35404 8716 35444 8756
rect 35212 8464 35252 8504
rect 35168 8296 35208 8336
rect 35250 8296 35290 8336
rect 35332 8296 35372 8336
rect 35414 8296 35454 8336
rect 35496 8296 35536 8336
rect 35308 7960 35348 8000
rect 35020 7876 35060 7916
rect 35020 7708 35060 7748
rect 34924 7456 34964 7496
rect 34924 7120 34964 7160
rect 34828 6616 34868 6656
rect 35308 7372 35348 7412
rect 36076 9304 36116 9344
rect 37228 9304 37268 9344
rect 36076 9052 36116 9092
rect 36844 8716 36884 8756
rect 35884 7960 35924 8000
rect 35500 7708 35540 7748
rect 36364 8548 36404 8588
rect 36268 7624 36308 7664
rect 35168 6784 35208 6824
rect 35250 6784 35290 6824
rect 35332 6784 35372 6824
rect 35414 6784 35454 6824
rect 35496 6784 35536 6824
rect 35212 6616 35252 6656
rect 35788 7204 35828 7244
rect 36268 7036 36308 7076
rect 35884 6952 35924 6992
rect 33928 6028 33968 6068
rect 34010 6028 34050 6068
rect 34092 6028 34132 6068
rect 34174 6028 34214 6068
rect 34256 6028 34296 6068
rect 34540 5608 34580 5648
rect 34348 4684 34388 4724
rect 33928 4516 33968 4556
rect 34010 4516 34050 4556
rect 34092 4516 34132 4556
rect 34174 4516 34214 4556
rect 34256 4516 34296 4556
rect 34444 4516 34484 4556
rect 33772 4012 33812 4052
rect 33676 3928 33716 3968
rect 34540 3844 34580 3884
rect 33676 3592 33716 3632
rect 33676 2080 33716 2120
rect 33928 3004 33968 3044
rect 34010 3004 34050 3044
rect 34092 3004 34132 3044
rect 34174 3004 34214 3044
rect 34256 3004 34296 3044
rect 34348 2836 34388 2876
rect 34252 2752 34292 2792
rect 33868 2668 33908 2708
rect 34732 5944 34772 5984
rect 34732 5608 34772 5648
rect 34732 4684 34772 4724
rect 35500 6280 35540 6320
rect 35692 6280 35732 6320
rect 35596 5608 35636 5648
rect 35212 5440 35252 5480
rect 35404 5440 35444 5480
rect 35168 5272 35208 5312
rect 35250 5272 35290 5312
rect 35332 5272 35372 5312
rect 35414 5272 35454 5312
rect 35496 5272 35536 5312
rect 34924 4768 34964 4808
rect 35116 4516 35156 4556
rect 34636 3172 34676 3212
rect 34636 2668 34676 2708
rect 34444 2080 34484 2120
rect 34060 1744 34100 1784
rect 33772 1660 33812 1700
rect 33928 1492 33968 1532
rect 34010 1492 34050 1532
rect 34092 1492 34132 1532
rect 34174 1492 34214 1532
rect 34256 1492 34296 1532
rect 33580 988 33620 1028
rect 35596 4936 35636 4976
rect 34924 2584 34964 2624
rect 34828 2080 34868 2120
rect 35168 3760 35208 3800
rect 35250 3760 35290 3800
rect 35332 3760 35372 3800
rect 35414 3760 35454 3800
rect 35496 3760 35536 3800
rect 35500 3340 35540 3380
rect 35500 2752 35540 2792
rect 35168 2248 35208 2288
rect 35250 2248 35290 2288
rect 35332 2248 35372 2288
rect 35414 2248 35454 2288
rect 35496 2248 35536 2288
rect 34924 1912 34964 1952
rect 35884 6280 35924 6320
rect 35788 3760 35828 3800
rect 36172 6952 36212 6992
rect 37132 7960 37172 8000
rect 37132 7624 37172 7664
rect 36364 6616 36404 6656
rect 36268 5608 36308 5648
rect 36652 5860 36692 5900
rect 36556 5524 36596 5564
rect 36364 5440 36404 5480
rect 36172 5104 36212 5144
rect 35980 5020 36020 5060
rect 35980 4852 36020 4892
rect 36076 4348 36116 4388
rect 36076 4096 36116 4136
rect 36556 5104 36596 5144
rect 36556 4600 36596 4640
rect 36460 4348 36500 4388
rect 36652 4012 36692 4052
rect 36172 2752 36212 2792
rect 36268 1240 36308 1280
rect 36364 1156 36404 1196
rect 35212 904 35252 944
rect 35168 736 35208 776
rect 35250 736 35290 776
rect 35332 736 35372 776
rect 35414 736 35454 776
rect 35496 736 35536 776
rect 35212 568 35252 608
rect 34060 232 34100 272
rect 33004 148 33044 188
rect 36556 2500 36596 2540
rect 36556 1660 36596 1700
rect 36460 1072 36500 1112
rect 36844 6616 36884 6656
rect 37324 7708 37364 7748
rect 38476 10144 38516 10184
rect 37708 9052 37748 9092
rect 38092 9136 38132 9176
rect 37900 8800 37940 8840
rect 37804 8464 37844 8504
rect 37900 8212 37940 8252
rect 37804 7372 37844 7412
rect 37804 7204 37844 7244
rect 37708 7120 37748 7160
rect 38092 8212 38132 8252
rect 38092 7708 38132 7748
rect 38284 8464 38324 8504
rect 38956 9808 38996 9848
rect 38764 9472 38804 9512
rect 38572 8884 38612 8924
rect 38476 7960 38516 8000
rect 38476 7540 38516 7580
rect 37708 6952 37748 6992
rect 37996 6952 38036 6992
rect 38188 6784 38228 6824
rect 38092 6700 38132 6740
rect 37996 6616 38036 6656
rect 37804 6112 37844 6152
rect 36844 5944 36884 5984
rect 37516 5944 37556 5984
rect 37036 5860 37076 5900
rect 37228 5440 37268 5480
rect 36940 5356 36980 5396
rect 36844 4264 36884 4304
rect 36844 3844 36884 3884
rect 37612 5692 37652 5732
rect 38476 7204 38516 7244
rect 38668 7540 38708 7580
rect 38668 7372 38708 7412
rect 38284 6532 38324 6572
rect 38188 6196 38228 6236
rect 38860 8632 38900 8672
rect 39148 9472 39188 9512
rect 39340 9304 39380 9344
rect 39436 8968 39476 9008
rect 39340 8716 39380 8756
rect 38956 7960 38996 8000
rect 39532 8464 39572 8504
rect 38860 6784 38900 6824
rect 38764 6700 38804 6740
rect 38572 5860 38612 5900
rect 38764 5776 38804 5816
rect 37036 4012 37076 4052
rect 37516 3760 37556 3800
rect 36652 1408 36692 1448
rect 37132 1828 37172 1868
rect 36940 1324 36980 1364
rect 36748 736 36788 776
rect 37708 3340 37748 3380
rect 37612 3088 37652 3128
rect 37996 4264 38036 4304
rect 38284 4180 38324 4220
rect 37900 3928 37940 3968
rect 38092 3340 38132 3380
rect 37900 3172 37940 3212
rect 38092 3088 38132 3128
rect 37804 1912 37844 1952
rect 37996 2080 38036 2120
rect 38956 5860 38996 5900
rect 39148 7288 39188 7328
rect 38956 5440 38996 5480
rect 38860 4180 38900 4220
rect 38764 4096 38804 4136
rect 38380 3172 38420 3212
rect 38284 2584 38324 2624
rect 38092 1996 38132 2036
rect 38860 2248 38900 2288
rect 38764 2080 38804 2120
rect 38668 1576 38708 1616
rect 38476 400 38516 440
rect 37900 64 37940 104
rect 39244 6483 39284 6488
rect 39244 6448 39284 6483
rect 40300 9472 40340 9512
rect 39916 8632 39956 8672
rect 39724 7960 39764 8000
rect 39436 7540 39476 7580
rect 39052 4936 39092 4976
rect 39148 4852 39188 4892
rect 39916 7540 39956 7580
rect 39820 7120 39860 7160
rect 39724 6448 39764 6488
rect 39628 6196 39668 6236
rect 39628 5188 39668 5228
rect 39340 4768 39380 4808
rect 39244 4684 39284 4724
rect 39532 4684 39572 4724
rect 39628 4264 39668 4304
rect 39148 3928 39188 3968
rect 39052 3592 39092 3632
rect 40012 6532 40052 6572
rect 40012 5860 40052 5900
rect 39916 5440 39956 5480
rect 39916 3592 39956 3632
rect 39532 3508 39572 3548
rect 40204 6280 40244 6320
rect 40972 9388 41012 9428
rect 40780 8716 40820 8756
rect 40588 8632 40628 8672
rect 40684 8380 40724 8420
rect 41260 8464 41300 8504
rect 41356 8128 41396 8168
rect 42508 8800 42548 8840
rect 41548 8128 41588 8168
rect 41260 7876 41300 7916
rect 41164 7540 41204 7580
rect 40876 7456 40916 7496
rect 41068 7456 41108 7496
rect 40492 7372 40532 7412
rect 41260 7372 41300 7412
rect 40972 7120 41012 7160
rect 41068 6784 41108 6824
rect 41260 6364 41300 6404
rect 40876 6196 40916 6236
rect 41068 6112 41108 6152
rect 41452 7792 41492 7832
rect 41452 7288 41492 7328
rect 41644 7120 41684 7160
rect 42508 6532 42548 6572
rect 41452 6448 41492 6488
rect 41356 5860 41396 5900
rect 41452 5776 41492 5816
rect 40396 5104 40436 5144
rect 40972 5104 41012 5144
rect 40300 4768 40340 4808
rect 40108 4348 40148 4388
rect 40108 3508 40148 3548
rect 40300 3256 40340 3296
rect 40780 4936 40820 4976
rect 41356 5440 41396 5480
rect 40780 4012 40820 4052
rect 40684 3676 40724 3716
rect 40588 2752 40628 2792
rect 41260 4852 41300 4892
rect 41452 5104 41492 5144
rect 41068 4684 41108 4724
rect 40972 3088 41012 3128
rect 41548 4684 41588 4724
rect 41356 4180 41396 4220
rect 41740 4012 41780 4052
rect 41068 2584 41108 2624
rect 40876 2416 40916 2456
rect 39724 2332 39764 2372
rect 39244 1912 39284 1952
rect 39532 1660 39572 1700
rect 39628 1156 39668 1196
rect 39436 988 39476 1028
rect 40588 1744 40628 1784
rect 40204 1324 40244 1364
rect 41452 3508 41492 3548
rect 41356 3424 41396 3464
rect 41260 3256 41300 3296
rect 41356 2920 41396 2960
rect 41260 2248 41300 2288
rect 41260 2080 41300 2120
rect 41164 1744 41204 1784
rect 40780 1240 40820 1280
rect 39820 652 39860 692
rect 40972 904 41012 944
rect 41548 3256 41588 3296
rect 41644 2752 41684 2792
rect 41548 2584 41588 2624
rect 41164 568 41204 608
rect 40012 232 40052 272
<< metal3 >>
rect 12268 10648 20236 10688
rect 20276 10648 20285 10688
rect 25411 10648 25420 10688
rect 25460 10648 39628 10688
rect 39668 10648 39677 10688
rect 12268 10604 12308 10648
rect 14659 10604 14717 10605
rect 12259 10564 12268 10604
rect 12308 10564 12317 10604
rect 14574 10564 14668 10604
rect 14708 10564 14717 10604
rect 14947 10564 14956 10604
rect 14996 10564 22348 10604
rect 22388 10564 22397 10604
rect 25027 10564 25036 10604
rect 25076 10564 35884 10604
rect 35924 10564 35933 10604
rect 14659 10563 14717 10564
rect 0 10520 80 10540
rect 15811 10520 15869 10521
rect 42928 10520 43008 10540
rect 0 10480 1708 10520
rect 1748 10480 1757 10520
rect 15726 10480 15820 10520
rect 15860 10480 15869 10520
rect 18115 10480 18124 10520
rect 18164 10480 24940 10520
rect 24980 10480 24989 10520
rect 25219 10480 25228 10520
rect 25268 10480 34924 10520
rect 34964 10480 34973 10520
rect 37603 10480 37612 10520
rect 37652 10480 43008 10520
rect 0 10460 80 10480
rect 15811 10479 15869 10480
rect 42928 10460 43008 10480
rect 19363 10396 19372 10436
rect 19412 10396 27148 10436
rect 27188 10396 27197 10436
rect 11875 10312 11884 10352
rect 11924 10312 12172 10352
rect 12212 10312 12221 10352
rect 16867 10312 16876 10352
rect 16916 10312 23692 10352
rect 23732 10312 23741 10352
rect 0 10184 80 10204
rect 15235 10184 15293 10185
rect 42928 10184 43008 10204
rect 0 10144 1612 10184
rect 1652 10144 1661 10184
rect 12163 10144 12172 10184
rect 12212 10144 12556 10184
rect 12596 10144 12605 10184
rect 15150 10144 15244 10184
rect 15284 10144 15293 10184
rect 38467 10144 38476 10184
rect 38516 10144 43008 10184
rect 0 10124 80 10144
rect 15235 10143 15293 10144
rect 42928 10124 43008 10144
rect 28291 10100 28349 10101
rect 15907 10060 15916 10100
rect 15956 10060 20620 10100
rect 20660 10060 20669 10100
rect 21667 10060 21676 10100
rect 21716 10060 21964 10100
rect 22004 10060 22013 10100
rect 27907 10060 27916 10100
rect 27956 10060 28300 10100
rect 28340 10060 28349 10100
rect 28291 10059 28349 10060
rect 21187 10016 21245 10017
rect 21571 10016 21629 10017
rect 10243 9976 10252 10016
rect 10292 9976 10540 10016
rect 10580 9976 10589 10016
rect 15235 9976 15244 10016
rect 15284 9976 20044 10016
rect 20084 9976 20093 10016
rect 20227 9976 20236 10016
rect 20276 9976 21196 10016
rect 21236 9976 21245 10016
rect 21486 9976 21580 10016
rect 21620 9976 21629 10016
rect 24355 9976 24364 10016
rect 24404 9976 26572 10016
rect 26612 9976 26621 10016
rect 21187 9975 21245 9976
rect 21571 9975 21629 9976
rect 17059 9932 17117 9933
rect 26275 9932 26333 9933
rect 13891 9892 13900 9932
rect 13940 9892 17068 9932
rect 17108 9892 17117 9932
rect 21283 9892 21292 9932
rect 21332 9892 22924 9932
rect 22964 9892 22973 9932
rect 24259 9892 24268 9932
rect 24308 9892 24748 9932
rect 24788 9892 24797 9932
rect 26275 9892 26284 9932
rect 26324 9892 26380 9932
rect 26420 9892 26429 9932
rect 17059 9891 17117 9892
rect 26275 9891 26333 9892
rect 0 9848 80 9868
rect 18499 9848 18557 9849
rect 20803 9848 20861 9849
rect 26947 9848 27005 9849
rect 42928 9848 43008 9868
rect 0 9808 4684 9848
rect 4724 9808 4733 9848
rect 4919 9808 4928 9848
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 5296 9808 5305 9848
rect 11320 9808 11404 9848
rect 11444 9808 11453 9848
rect 16483 9808 16492 9848
rect 16532 9808 17260 9848
rect 17300 9808 18028 9848
rect 18068 9808 18077 9848
rect 18414 9808 18508 9848
rect 18548 9808 18557 9848
rect 20039 9808 20048 9848
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20416 9808 20425 9848
rect 20718 9808 20812 9848
rect 20852 9808 20861 9848
rect 21475 9808 21484 9848
rect 21524 9808 22156 9848
rect 22196 9808 22205 9848
rect 22339 9808 22348 9848
rect 22388 9808 26956 9848
rect 26996 9808 27005 9848
rect 35159 9808 35168 9848
rect 35208 9808 35250 9848
rect 35290 9808 35332 9848
rect 35372 9808 35414 9848
rect 35454 9808 35496 9848
rect 35536 9808 35545 9848
rect 38947 9808 38956 9848
rect 38996 9808 43008 9848
rect 0 9788 80 9808
rect 11320 9764 11360 9808
rect 18499 9807 18557 9808
rect 20803 9807 20861 9808
rect 26947 9807 27005 9808
rect 42928 9788 43008 9808
rect 10156 9724 11360 9764
rect 14851 9724 14860 9764
rect 14900 9724 27052 9764
rect 27092 9724 27101 9764
rect 29155 9724 29164 9764
rect 29204 9724 35692 9764
rect 35732 9724 35741 9764
rect 1900 9556 9100 9596
rect 9140 9556 9149 9596
rect 0 9512 80 9532
rect 1900 9512 1940 9556
rect 10156 9512 10196 9724
rect 21091 9680 21149 9681
rect 32419 9680 32477 9681
rect 11020 9640 15148 9680
rect 15188 9640 16340 9680
rect 16387 9640 16396 9680
rect 16436 9640 17068 9680
rect 17108 9640 17117 9680
rect 17635 9640 17644 9680
rect 17684 9640 19412 9680
rect 19459 9640 19468 9680
rect 19508 9640 20332 9680
rect 20372 9640 20381 9680
rect 21091 9640 21100 9680
rect 21140 9640 21196 9680
rect 21236 9640 21245 9680
rect 21667 9640 21676 9680
rect 21716 9640 22156 9680
rect 22196 9640 27532 9680
rect 27572 9640 27581 9680
rect 30403 9640 30412 9680
rect 30452 9640 30892 9680
rect 30932 9640 30941 9680
rect 32323 9640 32332 9680
rect 32372 9640 32428 9680
rect 32468 9640 32477 9680
rect 32803 9640 32812 9680
rect 32852 9640 34444 9680
rect 34484 9640 35980 9680
rect 36020 9640 37324 9680
rect 37364 9640 37373 9680
rect 0 9472 1940 9512
rect 2947 9472 2956 9512
rect 2996 9472 3244 9512
rect 3284 9472 4972 9512
rect 5012 9472 5021 9512
rect 5923 9472 5932 9512
rect 5972 9472 6700 9512
rect 6740 9472 6749 9512
rect 8803 9472 8812 9512
rect 8852 9472 9484 9512
rect 9524 9472 9533 9512
rect 10147 9472 10156 9512
rect 10196 9472 10205 9512
rect 0 9452 80 9472
rect 9571 9388 9580 9428
rect 9620 9388 10924 9428
rect 10964 9388 10973 9428
rect 11020 9344 11060 9640
rect 16300 9596 16340 9640
rect 17923 9596 17981 9597
rect 13219 9556 13228 9596
rect 13268 9556 13277 9596
rect 16291 9556 16300 9596
rect 16340 9556 16349 9596
rect 17838 9556 17932 9596
rect 17972 9556 17981 9596
rect 13228 9512 13268 9556
rect 17923 9555 17981 9556
rect 15619 9512 15677 9513
rect 16579 9512 16637 9513
rect 19267 9512 19325 9513
rect 13027 9472 13036 9512
rect 13076 9472 13268 9512
rect 14083 9472 14092 9512
rect 14132 9472 15628 9512
rect 15668 9472 15677 9512
rect 16494 9472 16588 9512
rect 16628 9472 16637 9512
rect 17347 9472 17356 9512
rect 17396 9472 19276 9512
rect 19316 9472 19325 9512
rect 19372 9512 19412 9640
rect 21091 9639 21149 9640
rect 32419 9639 32477 9640
rect 24643 9556 24652 9596
rect 24692 9556 30124 9596
rect 30164 9556 30173 9596
rect 30787 9556 30796 9596
rect 30836 9556 31852 9596
rect 31892 9556 31901 9596
rect 19459 9512 19517 9513
rect 42928 9512 43008 9532
rect 19372 9472 19468 9512
rect 19508 9472 19602 9512
rect 20707 9472 20716 9512
rect 20756 9472 23308 9512
rect 23348 9472 23357 9512
rect 25411 9472 25420 9512
rect 25460 9472 34060 9512
rect 34100 9472 38764 9512
rect 38804 9472 39148 9512
rect 39188 9472 39197 9512
rect 40291 9472 40300 9512
rect 40340 9472 43008 9512
rect 15619 9471 15677 9472
rect 16579 9471 16637 9472
rect 19267 9471 19325 9472
rect 19459 9471 19517 9472
rect 42928 9452 43008 9472
rect 13219 9428 13277 9429
rect 21667 9428 21725 9429
rect 40963 9428 41021 9429
rect 13134 9388 13228 9428
rect 13268 9388 13277 9428
rect 14947 9388 14956 9428
rect 14996 9388 15340 9428
rect 15380 9388 15389 9428
rect 16204 9388 16780 9428
rect 16820 9388 17644 9428
rect 17684 9388 17693 9428
rect 19267 9388 19276 9428
rect 19316 9388 21676 9428
rect 21716 9388 21725 9428
rect 13219 9387 13277 9388
rect 16204 9344 16244 9388
rect 21667 9387 21725 9388
rect 26440 9388 27092 9428
rect 27235 9388 27244 9428
rect 27284 9388 27628 9428
rect 27668 9388 27677 9428
rect 29251 9388 29260 9428
rect 29300 9388 29740 9428
rect 29780 9388 29789 9428
rect 30595 9388 30604 9428
rect 30644 9388 31180 9428
rect 31220 9388 31229 9428
rect 35683 9388 35692 9428
rect 35732 9388 37268 9428
rect 40878 9388 40972 9428
rect 41012 9388 41021 9428
rect 3427 9304 3436 9344
rect 3476 9304 6124 9344
rect 6164 9304 6173 9344
rect 9667 9304 9676 9344
rect 9716 9304 11060 9344
rect 11203 9304 11212 9344
rect 11252 9304 12460 9344
rect 12500 9304 16244 9344
rect 16291 9304 16300 9344
rect 16340 9304 24556 9344
rect 24596 9304 24605 9344
rect 20707 9260 20765 9261
rect 6595 9220 6604 9260
rect 6644 9220 8428 9260
rect 8468 9220 8477 9260
rect 10339 9220 10348 9260
rect 10388 9220 17836 9260
rect 17876 9220 17885 9260
rect 18883 9220 18892 9260
rect 18932 9220 20716 9260
rect 20756 9220 20765 9260
rect 20899 9220 20908 9260
rect 20948 9220 21772 9260
rect 21812 9220 21821 9260
rect 24355 9220 24364 9260
rect 24404 9220 25420 9260
rect 25460 9220 25469 9260
rect 20707 9219 20765 9220
rect 0 9176 80 9196
rect 26440 9176 26480 9388
rect 26659 9344 26717 9345
rect 26563 9304 26572 9344
rect 26612 9304 26668 9344
rect 26708 9304 26717 9344
rect 27052 9344 27092 9388
rect 37228 9344 37268 9388
rect 40963 9387 41021 9388
rect 27052 9304 29356 9344
rect 29396 9304 36076 9344
rect 36116 9304 36125 9344
rect 37219 9304 37228 9344
rect 37268 9304 39340 9344
rect 39380 9304 39389 9344
rect 26659 9303 26717 9304
rect 26947 9260 27005 9261
rect 27715 9260 27773 9261
rect 26947 9220 26956 9260
rect 26996 9220 27007 9260
rect 27715 9220 27724 9260
rect 27764 9220 29164 9260
rect 29204 9220 29213 9260
rect 30787 9220 30796 9260
rect 30836 9220 32044 9260
rect 32084 9220 32093 9260
rect 32611 9220 32620 9260
rect 32660 9220 33292 9260
rect 33332 9220 33341 9260
rect 26947 9219 27005 9220
rect 27715 9219 27773 9220
rect 26956 9176 26996 9219
rect 42928 9176 43008 9196
rect 0 9136 4876 9176
rect 4916 9136 26480 9176
rect 26947 9136 26956 9176
rect 26996 9136 27005 9176
rect 31363 9136 31372 9176
rect 31412 9136 34484 9176
rect 38083 9136 38092 9176
rect 38132 9136 43008 9176
rect 0 9116 80 9136
rect 16963 9092 17021 9093
rect 21571 9092 21629 9093
rect 26467 9092 26525 9093
rect 34444 9092 34484 9136
rect 42928 9116 43008 9136
rect 3679 9052 3688 9092
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 4056 9052 4065 9092
rect 9091 9052 9100 9092
rect 9140 9052 9388 9092
rect 9428 9052 11212 9092
rect 11252 9052 11261 9092
rect 12739 9052 12748 9092
rect 12788 9052 15244 9092
rect 15284 9052 15293 9092
rect 16483 9052 16492 9092
rect 16532 9052 16780 9092
rect 16820 9052 16829 9092
rect 16878 9052 16972 9092
rect 17012 9052 17021 9092
rect 18799 9052 18808 9092
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 19176 9052 19185 9092
rect 21571 9052 21580 9092
rect 21620 9052 21676 9092
rect 21716 9052 21725 9092
rect 24451 9052 24460 9092
rect 24500 9052 24509 9092
rect 25795 9052 25804 9092
rect 25844 9052 26476 9092
rect 26516 9052 26525 9092
rect 28963 9052 28972 9092
rect 29012 9052 29452 9092
rect 29492 9052 29501 9092
rect 32131 9052 32140 9092
rect 32180 9052 33196 9092
rect 33236 9052 33245 9092
rect 33919 9052 33928 9092
rect 33968 9052 34010 9092
rect 34050 9052 34092 9092
rect 34132 9052 34174 9092
rect 34214 9052 34256 9092
rect 34296 9052 34305 9092
rect 34435 9052 34444 9092
rect 34484 9052 34493 9092
rect 36067 9052 36076 9092
rect 36116 9052 37708 9092
rect 37748 9052 37757 9092
rect 16963 9051 17021 9052
rect 21571 9051 21629 9052
rect 4675 8968 4684 9008
rect 4724 8968 9580 9008
rect 9620 8968 9629 9008
rect 10723 8968 10732 9008
rect 10772 8968 11788 9008
rect 11828 8968 11837 9008
rect 12355 8968 12364 9008
rect 12404 8968 24364 9008
rect 24404 8968 24413 9008
rect 12364 8924 12404 8968
rect 24460 8924 24500 9052
rect 26467 9051 26525 9052
rect 32515 9008 32573 9009
rect 24547 8968 24556 9008
rect 24596 8968 32084 9008
rect 32430 8968 32524 9008
rect 32564 8968 32573 9008
rect 33091 8968 33100 9008
rect 33140 8968 35596 9008
rect 35636 8968 35645 9008
rect 35875 8968 35884 9008
rect 35924 8968 39436 9008
rect 39476 8968 39485 9008
rect 32044 8924 32084 8968
rect 32515 8967 32573 8968
rect 1603 8884 1612 8924
rect 1652 8884 12404 8924
rect 13795 8884 13804 8924
rect 13844 8884 17740 8924
rect 17780 8884 17789 8924
rect 21859 8884 21868 8924
rect 21908 8884 24500 8924
rect 26275 8884 26284 8924
rect 26324 8884 29836 8924
rect 29876 8884 29885 8924
rect 30499 8884 30508 8924
rect 30548 8884 30988 8924
rect 31028 8884 31037 8924
rect 31843 8884 31852 8924
rect 31892 8884 31901 8924
rect 32044 8884 38572 8924
rect 38612 8884 38621 8924
rect 0 8840 80 8860
rect 5923 8840 5981 8841
rect 13507 8840 13565 8841
rect 0 8800 3820 8840
rect 3860 8800 3869 8840
rect 4771 8800 4780 8840
rect 4820 8800 4829 8840
rect 5838 8800 5932 8840
rect 5972 8800 5981 8840
rect 6211 8800 6220 8840
rect 6260 8800 6796 8840
rect 6836 8800 7276 8840
rect 7316 8800 7325 8840
rect 7459 8800 7468 8840
rect 7508 8800 8140 8840
rect 8180 8800 8189 8840
rect 9859 8800 9868 8840
rect 9908 8800 10252 8840
rect 10292 8800 10301 8840
rect 13422 8800 13516 8840
rect 13556 8800 13565 8840
rect 0 8780 80 8800
rect 4780 8756 4820 8800
rect 5923 8799 5981 8800
rect 13507 8799 13565 8800
rect 13699 8840 13757 8841
rect 14275 8840 14333 8841
rect 15043 8840 15101 8841
rect 15523 8840 15581 8841
rect 21283 8840 21341 8841
rect 24364 8840 24404 8884
rect 31852 8840 31892 8884
rect 13699 8800 13708 8840
rect 13748 8800 13842 8840
rect 14190 8800 14284 8840
rect 14324 8800 14333 8840
rect 14958 8800 15052 8840
rect 15092 8800 15101 8840
rect 15427 8800 15436 8840
rect 15476 8800 15532 8840
rect 15572 8800 15581 8840
rect 15811 8800 15820 8840
rect 15860 8800 17164 8840
rect 17204 8800 17213 8840
rect 18883 8800 18892 8840
rect 18932 8800 19372 8840
rect 19412 8800 19421 8840
rect 19651 8800 19660 8840
rect 19700 8800 20620 8840
rect 20660 8800 20669 8840
rect 21198 8800 21292 8840
rect 21332 8800 21341 8840
rect 13699 8799 13757 8800
rect 14275 8799 14333 8800
rect 15043 8799 15101 8800
rect 15523 8799 15581 8800
rect 21283 8799 21341 8800
rect 22348 8800 22828 8840
rect 22868 8800 23212 8840
rect 23252 8800 23261 8840
rect 23491 8800 23500 8840
rect 23540 8800 24172 8840
rect 24212 8800 24221 8840
rect 24355 8800 24364 8840
rect 24404 8800 24413 8840
rect 24547 8800 24556 8840
rect 24596 8800 24844 8840
rect 24884 8800 24893 8840
rect 24940 8800 26476 8840
rect 26516 8800 29068 8840
rect 29108 8800 29117 8840
rect 30691 8800 30700 8840
rect 30740 8800 31892 8840
rect 31939 8840 31997 8841
rect 32611 8840 32669 8841
rect 35299 8840 35357 8841
rect 37891 8840 37949 8841
rect 42928 8840 43008 8860
rect 31939 8800 31948 8840
rect 31988 8800 32428 8840
rect 32468 8800 32477 8840
rect 32611 8800 32620 8840
rect 32660 8800 32716 8840
rect 32756 8800 32765 8840
rect 32812 8800 35308 8840
rect 35348 8800 35357 8840
rect 37806 8800 37900 8840
rect 37940 8800 37949 8840
rect 42499 8800 42508 8840
rect 42548 8800 43008 8840
rect 11011 8756 11069 8757
rect 20899 8756 20957 8757
rect 22348 8756 22388 8800
rect 24940 8756 24980 8800
rect 2083 8716 2092 8756
rect 2132 8716 2860 8756
rect 2900 8716 2909 8756
rect 4003 8716 4012 8756
rect 4052 8716 4820 8756
rect 8428 8716 8812 8756
rect 8852 8716 8861 8756
rect 10926 8716 11020 8756
rect 11060 8716 11069 8756
rect 11971 8716 11980 8756
rect 12020 8716 20140 8756
rect 20180 8716 20189 8756
rect 20899 8716 20908 8756
rect 20948 8716 22388 8756
rect 22435 8716 22444 8756
rect 22484 8716 24980 8756
rect 26440 8716 26516 8800
rect 31939 8799 31997 8800
rect 32611 8799 32669 8800
rect 26659 8756 26717 8757
rect 32812 8756 32852 8800
rect 35299 8799 35357 8800
rect 37891 8799 37949 8800
rect 37900 8756 37940 8799
rect 42928 8780 43008 8800
rect 26659 8716 26668 8756
rect 26708 8716 28012 8756
rect 28052 8716 28061 8756
rect 28291 8716 28300 8756
rect 28340 8716 28684 8756
rect 28724 8716 28733 8756
rect 29827 8716 29836 8756
rect 29876 8716 32852 8756
rect 34723 8716 34732 8756
rect 34772 8716 35404 8756
rect 35444 8716 35453 8756
rect 35500 8716 36844 8756
rect 36884 8716 36893 8756
rect 37900 8716 39284 8756
rect 39331 8716 39340 8756
rect 39380 8716 40780 8756
rect 40820 8716 40829 8756
rect 2563 8632 2572 8672
rect 2612 8632 3052 8672
rect 3092 8632 4396 8672
rect 4436 8632 5068 8672
rect 5108 8632 5117 8672
rect 6403 8632 6412 8672
rect 6452 8632 6892 8672
rect 6932 8632 6941 8672
rect 8131 8632 8140 8672
rect 8180 8632 8332 8672
rect 8372 8632 8381 8672
rect 4195 8588 4253 8589
rect 8428 8588 8468 8716
rect 11011 8715 11069 8716
rect 20899 8715 20957 8716
rect 26659 8715 26717 8716
rect 26431 8672 26489 8673
rect 8515 8632 8524 8672
rect 8564 8632 9100 8672
rect 9140 8632 9149 8672
rect 15139 8632 15148 8672
rect 15188 8632 16724 8672
rect 16867 8632 16876 8672
rect 16916 8632 21868 8672
rect 21908 8632 21917 8672
rect 22819 8632 22828 8672
rect 22868 8632 26440 8672
rect 26480 8632 26489 8672
rect 16684 8588 16724 8632
rect 26431 8631 26489 8632
rect 26563 8672 26621 8673
rect 28387 8672 28445 8673
rect 35500 8672 35540 8716
rect 39244 8672 39284 8716
rect 40771 8672 40829 8673
rect 26563 8632 26572 8672
rect 26612 8632 26956 8672
rect 26996 8632 27005 8672
rect 28302 8632 28396 8672
rect 28436 8632 28445 8672
rect 28867 8632 28876 8672
rect 28916 8632 30988 8672
rect 31028 8632 31037 8672
rect 31555 8632 31564 8672
rect 31604 8632 33772 8672
rect 33812 8632 33821 8672
rect 34339 8632 34348 8672
rect 34388 8632 35540 8672
rect 36364 8632 38860 8672
rect 38900 8632 38909 8672
rect 39244 8632 39916 8672
rect 39956 8632 40588 8672
rect 40628 8632 40780 8672
rect 40820 8632 40829 8672
rect 26563 8631 26621 8632
rect 28387 8631 28445 8632
rect 30115 8588 30173 8589
rect 30307 8588 30365 8589
rect 3907 8548 3916 8588
rect 3956 8548 4204 8588
rect 4244 8548 7180 8588
rect 7220 8548 7229 8588
rect 8332 8548 8468 8588
rect 13891 8548 13900 8588
rect 13940 8548 15724 8588
rect 15764 8548 15773 8588
rect 16684 8548 17452 8588
rect 17492 8548 22348 8588
rect 22388 8548 26572 8588
rect 26612 8548 30124 8588
rect 30164 8548 30173 8588
rect 30222 8548 30316 8588
rect 30356 8548 30365 8588
rect 4195 8547 4253 8548
rect 0 8504 80 8524
rect 4579 8504 4637 8505
rect 8332 8504 8372 8548
rect 30115 8547 30173 8548
rect 30307 8547 30365 8548
rect 16387 8504 16445 8505
rect 21475 8504 21533 8505
rect 30988 8504 31028 8632
rect 36364 8588 36404 8632
rect 31363 8548 31372 8588
rect 31412 8548 33388 8588
rect 33428 8548 33437 8588
rect 33859 8548 33868 8588
rect 33908 8548 36364 8588
rect 36404 8548 36413 8588
rect 32227 8504 32285 8505
rect 34339 8504 34397 8505
rect 37900 8504 37940 8632
rect 40771 8631 40829 8632
rect 42928 8504 43008 8524
rect 0 8464 4588 8504
rect 4628 8464 4637 8504
rect 6211 8464 6220 8504
rect 6260 8464 6508 8504
rect 6548 8464 8332 8504
rect 8372 8464 8381 8504
rect 10531 8464 10540 8504
rect 10580 8464 11540 8504
rect 11587 8464 11596 8504
rect 11636 8464 16396 8504
rect 16436 8464 16445 8504
rect 16963 8464 16972 8504
rect 17012 8464 18316 8504
rect 18356 8464 18988 8504
rect 19028 8464 19037 8504
rect 20419 8464 20428 8504
rect 20468 8464 20908 8504
rect 20948 8464 20957 8504
rect 21475 8464 21484 8504
rect 21524 8464 22924 8504
rect 22964 8464 22973 8504
rect 23203 8464 23212 8504
rect 23252 8464 28780 8504
rect 28820 8464 28829 8504
rect 29635 8464 29644 8504
rect 29684 8464 30604 8504
rect 30644 8464 30653 8504
rect 30988 8464 32044 8504
rect 32084 8464 32093 8504
rect 32227 8464 32236 8504
rect 32276 8464 32716 8504
rect 32756 8464 32765 8504
rect 34339 8464 34348 8504
rect 34388 8464 35212 8504
rect 35252 8464 35261 8504
rect 37795 8464 37804 8504
rect 37844 8464 37940 8504
rect 38275 8464 38284 8504
rect 38324 8464 39532 8504
rect 39572 8464 39581 8504
rect 41251 8464 41260 8504
rect 41300 8464 43008 8504
rect 0 8444 80 8464
rect 4579 8463 4637 8464
rect 11395 8420 11453 8421
rect 1699 8380 1708 8420
rect 1748 8380 11404 8420
rect 11444 8380 11453 8420
rect 11500 8420 11540 8464
rect 16387 8463 16445 8464
rect 21475 8463 21533 8464
rect 32227 8463 32285 8464
rect 34339 8463 34397 8464
rect 42928 8444 43008 8464
rect 31651 8420 31709 8421
rect 11500 8380 12172 8420
rect 12212 8380 12221 8420
rect 17827 8380 17836 8420
rect 17876 8380 18412 8420
rect 18452 8380 18461 8420
rect 18508 8380 22828 8420
rect 22868 8380 22877 8420
rect 25315 8380 25324 8420
rect 25364 8380 29836 8420
rect 29876 8380 29885 8420
rect 31566 8380 31660 8420
rect 31700 8380 31709 8420
rect 32515 8380 32524 8420
rect 32564 8380 40684 8420
rect 40724 8380 40733 8420
rect 11395 8379 11453 8380
rect 18508 8336 18548 8380
rect 31651 8379 31709 8380
rect 26275 8336 26333 8337
rect 4919 8296 4928 8336
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 5296 8296 5305 8336
rect 9955 8296 9964 8336
rect 10004 8296 13996 8336
rect 14036 8296 14045 8336
rect 14659 8296 14668 8336
rect 14708 8296 15244 8336
rect 15284 8296 18548 8336
rect 19363 8296 19372 8336
rect 19412 8296 19948 8336
rect 19988 8296 19997 8336
rect 20039 8296 20048 8336
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20416 8296 20425 8336
rect 21859 8296 21868 8336
rect 21908 8296 22252 8336
rect 22292 8296 22301 8336
rect 26275 8296 26284 8336
rect 26324 8296 26380 8336
rect 26420 8296 26429 8336
rect 27907 8296 27916 8336
rect 27956 8296 28588 8336
rect 28628 8296 28637 8336
rect 32323 8296 32332 8336
rect 32372 8296 32620 8336
rect 32660 8296 32669 8336
rect 35159 8296 35168 8336
rect 35208 8296 35250 8336
rect 35290 8296 35332 8336
rect 35372 8296 35414 8336
rect 35454 8296 35496 8336
rect 35536 8296 35545 8336
rect 26275 8295 26333 8296
rect 11395 8252 11453 8253
rect 15427 8252 15485 8253
rect 3139 8212 3148 8252
rect 3188 8212 5876 8252
rect 0 8168 80 8188
rect 1603 8168 1661 8169
rect 5836 8168 5876 8212
rect 11395 8212 11404 8252
rect 11444 8212 15436 8252
rect 15476 8212 15485 8252
rect 18691 8212 18700 8252
rect 18740 8212 25708 8252
rect 25748 8212 25757 8252
rect 27331 8212 27340 8252
rect 27380 8212 28492 8252
rect 28532 8212 31564 8252
rect 31604 8212 31613 8252
rect 32515 8212 32524 8252
rect 32564 8212 34348 8252
rect 34388 8212 34397 8252
rect 37891 8212 37900 8252
rect 37940 8212 38092 8252
rect 38132 8212 38141 8252
rect 11395 8211 11453 8212
rect 15427 8211 15485 8212
rect 13795 8168 13853 8169
rect 32707 8168 32765 8169
rect 42928 8168 43008 8188
rect 0 8128 1324 8168
rect 1364 8128 1612 8168
rect 1652 8128 1661 8168
rect 1891 8128 1900 8168
rect 1940 8128 3340 8168
rect 3380 8128 3389 8168
rect 3811 8128 3820 8168
rect 3860 8128 4820 8168
rect 5827 8128 5836 8168
rect 5876 8128 6028 8168
rect 6068 8128 6077 8168
rect 6883 8128 6892 8168
rect 6932 8128 7276 8168
rect 7316 8128 7325 8168
rect 8419 8128 8428 8168
rect 8468 8128 9196 8168
rect 9236 8128 9245 8168
rect 10435 8128 10444 8168
rect 10484 8128 13804 8168
rect 13844 8128 13853 8168
rect 15523 8128 15532 8168
rect 15572 8128 23212 8168
rect 23252 8128 23261 8168
rect 24931 8128 24940 8168
rect 24980 8128 28724 8168
rect 28771 8128 28780 8168
rect 28820 8128 31948 8168
rect 31988 8128 31997 8168
rect 32707 8128 32716 8168
rect 32756 8128 34060 8168
rect 34100 8128 41356 8168
rect 41396 8128 41405 8168
rect 41539 8128 41548 8168
rect 41588 8128 43008 8168
rect 0 8108 80 8128
rect 1603 8127 1661 8128
rect 3340 8084 3380 8128
rect 4780 8084 4820 8128
rect 13795 8127 13853 8128
rect 23011 8084 23069 8085
rect 28579 8084 28637 8085
rect 3340 8044 4340 8084
rect 4771 8044 4780 8084
rect 4820 8044 10636 8084
rect 10676 8044 10685 8084
rect 10915 8044 10924 8084
rect 10964 8044 12884 8084
rect 15619 8044 15628 8084
rect 15668 8044 19756 8084
rect 19796 8044 19805 8084
rect 22926 8044 23020 8084
rect 23060 8044 23069 8084
rect 4300 8000 4340 8044
rect 12844 8000 12884 8044
rect 23011 8043 23069 8044
rect 23884 8044 23980 8084
rect 24020 8044 24029 8084
rect 28494 8044 28588 8084
rect 28628 8044 28637 8084
rect 28684 8084 28724 8128
rect 32707 8127 32765 8128
rect 42928 8108 43008 8128
rect 28684 8044 32524 8084
rect 32564 8044 32573 8084
rect 33859 8044 33868 8084
rect 33908 8044 33917 8084
rect 15427 8000 15485 8001
rect 19555 8000 19613 8001
rect 22051 8000 22109 8001
rect 1795 7960 1804 8000
rect 1844 7960 3820 8000
rect 3860 7960 3869 8000
rect 4291 7960 4300 8000
rect 4340 7960 4349 8000
rect 4579 7960 4588 8000
rect 4628 7960 4637 8000
rect 6115 7960 6124 8000
rect 6164 7960 6316 8000
rect 6356 7960 6700 8000
rect 6740 7960 9100 8000
rect 9140 7960 9149 8000
rect 12835 7960 12844 8000
rect 12884 7960 12893 8000
rect 15342 7960 15436 8000
rect 15476 7960 15485 8000
rect 17155 7960 17164 8000
rect 17204 7960 17548 8000
rect 17588 7960 19180 8000
rect 19220 7960 19229 8000
rect 19470 7960 19564 8000
rect 19604 7960 19613 8000
rect 21966 7960 22060 8000
rect 22100 7960 22109 8000
rect 0 7832 80 7852
rect 1699 7832 1757 7833
rect 0 7792 1708 7832
rect 1748 7792 1757 7832
rect 4588 7832 4628 7960
rect 15427 7959 15485 7960
rect 19555 7959 19613 7960
rect 22051 7959 22109 7960
rect 7555 7916 7613 7917
rect 7267 7876 7276 7916
rect 7316 7876 7564 7916
rect 7604 7876 7613 7916
rect 7555 7875 7613 7876
rect 7747 7916 7805 7917
rect 16387 7916 16445 7917
rect 23884 7916 23924 8044
rect 28579 8043 28637 8044
rect 24067 8000 24125 8001
rect 28771 8000 28829 8001
rect 30019 8000 30077 8001
rect 33868 8000 33908 8044
rect 37123 8000 37181 8001
rect 23982 7960 24076 8000
rect 24116 7960 24125 8000
rect 27811 7960 27820 8000
rect 27860 7960 28396 8000
rect 28436 7960 28445 8000
rect 28686 7960 28780 8000
rect 28820 7960 28829 8000
rect 29934 7960 30028 8000
rect 30068 7960 30988 8000
rect 31028 7960 31180 8000
rect 31220 7960 31229 8000
rect 31939 7960 31948 8000
rect 31988 7960 33908 8000
rect 35299 7960 35308 8000
rect 35348 7960 35884 8000
rect 35924 7960 35933 8000
rect 37038 7960 37132 8000
rect 37172 7960 37181 8000
rect 24067 7959 24125 7960
rect 28771 7959 28829 7960
rect 30019 7959 30077 7960
rect 37123 7959 37181 7960
rect 38179 8000 38237 8001
rect 38179 7960 38188 8000
rect 38228 7960 38476 8000
rect 38516 7960 38525 8000
rect 38947 7960 38956 8000
rect 38996 7960 39724 8000
rect 39764 7960 39773 8000
rect 38179 7959 38237 7960
rect 28867 7916 28925 7917
rect 7747 7876 7756 7916
rect 7796 7876 7890 7916
rect 9667 7876 9676 7916
rect 9716 7876 16396 7916
rect 16436 7876 16445 7916
rect 19363 7876 19372 7916
rect 19412 7876 23924 7916
rect 23980 7876 28876 7916
rect 28916 7876 28925 7916
rect 33859 7876 33868 7916
rect 33908 7876 35020 7916
rect 35060 7876 35069 7916
rect 37780 7876 41260 7916
rect 41300 7876 41309 7916
rect 7747 7875 7805 7876
rect 16387 7875 16445 7876
rect 23875 7832 23933 7833
rect 4588 7792 11116 7832
rect 11156 7792 11165 7832
rect 19459 7792 19468 7832
rect 19508 7792 19948 7832
rect 19988 7792 23884 7832
rect 23924 7792 23933 7832
rect 0 7772 80 7792
rect 1699 7791 1757 7792
rect 23875 7791 23933 7792
rect 17635 7748 17693 7749
rect 21475 7748 21533 7749
rect 23980 7748 24020 7876
rect 28867 7875 28925 7876
rect 33667 7832 33725 7833
rect 37780 7832 37820 7876
rect 42928 7832 43008 7852
rect 24076 7792 28300 7832
rect 28340 7792 33236 7832
rect 33582 7792 33676 7832
rect 33716 7792 33725 7832
rect 24076 7749 24116 7792
rect 3043 7708 3052 7748
rect 3092 7708 7276 7748
rect 7316 7708 7325 7748
rect 7555 7708 7564 7748
rect 7604 7708 9196 7748
rect 9236 7708 9245 7748
rect 10723 7708 10732 7748
rect 10772 7708 11308 7748
rect 11348 7708 13612 7748
rect 13652 7708 14188 7748
rect 14228 7708 17644 7748
rect 17684 7708 17693 7748
rect 19171 7708 19180 7748
rect 19220 7708 20812 7748
rect 20852 7708 20861 7748
rect 21475 7708 21484 7748
rect 21524 7708 22060 7748
rect 22100 7708 24020 7748
rect 24067 7748 24125 7749
rect 28867 7748 28925 7749
rect 33196 7748 33236 7792
rect 33667 7791 33725 7792
rect 33772 7792 37820 7832
rect 41443 7792 41452 7832
rect 41492 7792 43008 7832
rect 33772 7748 33812 7792
rect 42928 7772 43008 7792
rect 37315 7748 37373 7749
rect 38083 7748 38141 7749
rect 24067 7708 24076 7748
rect 24116 7708 24125 7748
rect 24835 7708 24844 7748
rect 24884 7708 28588 7748
rect 28628 7708 28637 7748
rect 28867 7708 28876 7748
rect 28916 7708 29452 7748
rect 29492 7708 29501 7748
rect 30595 7708 30604 7748
rect 30644 7708 32044 7748
rect 32084 7708 32093 7748
rect 33196 7708 33580 7748
rect 33620 7708 33629 7748
rect 33676 7708 33812 7748
rect 35011 7708 35020 7748
rect 35060 7708 35500 7748
rect 35540 7708 35549 7748
rect 37230 7708 37324 7748
rect 37364 7708 37373 7748
rect 37998 7708 38092 7748
rect 38132 7708 38141 7748
rect 17635 7707 17693 7708
rect 21475 7707 21533 7708
rect 24067 7707 24125 7708
rect 28867 7707 28925 7708
rect 7459 7664 7517 7665
rect 32419 7664 32477 7665
rect 33283 7664 33341 7665
rect 33676 7664 33716 7708
rect 37315 7707 37373 7708
rect 38083 7707 38141 7708
rect 5731 7624 5740 7664
rect 5780 7624 6028 7664
rect 6068 7624 6077 7664
rect 7363 7624 7372 7664
rect 7412 7624 7468 7664
rect 7508 7624 8812 7664
rect 8852 7624 8861 7664
rect 10915 7624 10924 7664
rect 10964 7624 18508 7664
rect 18548 7624 21868 7664
rect 21908 7624 22540 7664
rect 22580 7624 22589 7664
rect 23875 7624 23884 7664
rect 23924 7624 25324 7664
rect 25364 7624 25373 7664
rect 25987 7624 25996 7664
rect 26036 7624 26188 7664
rect 26228 7624 26237 7664
rect 28099 7624 28108 7664
rect 28148 7624 28780 7664
rect 28820 7624 31700 7664
rect 31843 7624 31852 7664
rect 31892 7624 32236 7664
rect 32276 7624 32285 7664
rect 32419 7624 32428 7664
rect 32468 7624 32562 7664
rect 33198 7624 33292 7664
rect 33332 7624 33716 7664
rect 33772 7624 36268 7664
rect 36308 7624 36317 7664
rect 37123 7624 37132 7664
rect 37172 7624 39956 7664
rect 7459 7623 7517 7624
rect 1699 7580 1757 7581
rect 4579 7580 4637 7581
rect 10924 7580 10964 7624
rect 31660 7580 31700 7624
rect 32419 7623 32477 7624
rect 33283 7623 33341 7624
rect 33772 7580 33812 7624
rect 35299 7580 35357 7581
rect 39916 7580 39956 7624
rect 1614 7540 1708 7580
rect 1748 7540 1757 7580
rect 3679 7540 3688 7580
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 4056 7540 4065 7580
rect 4494 7540 4588 7580
rect 4628 7540 4637 7580
rect 6115 7540 6124 7580
rect 6164 7540 6988 7580
rect 7028 7540 7276 7580
rect 7316 7540 8236 7580
rect 8276 7540 8285 7580
rect 8800 7540 10964 7580
rect 12067 7540 12076 7580
rect 12116 7540 12652 7580
rect 12692 7540 12701 7580
rect 14380 7540 17836 7580
rect 17876 7540 17885 7580
rect 18799 7540 18808 7580
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 19176 7540 19185 7580
rect 19555 7540 19564 7580
rect 19604 7540 20716 7580
rect 20756 7540 20765 7580
rect 23779 7540 23788 7580
rect 23828 7540 24460 7580
rect 24500 7540 27340 7580
rect 27380 7540 27389 7580
rect 27715 7540 27724 7580
rect 27764 7540 28204 7580
rect 28244 7540 28253 7580
rect 31660 7540 33812 7580
rect 33919 7540 33928 7580
rect 33968 7540 34010 7580
rect 34050 7540 34092 7580
rect 34132 7540 34174 7580
rect 34214 7540 34256 7580
rect 34296 7540 34305 7580
rect 35299 7540 35308 7580
rect 35348 7540 38476 7580
rect 38516 7540 38525 7580
rect 38659 7540 38668 7580
rect 38708 7540 39436 7580
rect 39476 7540 39485 7580
rect 39907 7540 39916 7580
rect 39956 7540 41164 7580
rect 41204 7540 41213 7580
rect 1699 7539 1757 7540
rect 4579 7539 4637 7540
rect 0 7496 80 7516
rect 8800 7496 8840 7540
rect 14380 7496 14420 7540
rect 35299 7539 35357 7540
rect 26563 7496 26621 7497
rect 31939 7496 31997 7497
rect 42928 7496 43008 7516
rect 0 7456 1844 7496
rect 5539 7456 5548 7496
rect 5588 7456 6700 7496
rect 6740 7456 8840 7496
rect 11779 7456 11788 7496
rect 11828 7456 14380 7496
rect 14420 7456 14429 7496
rect 15715 7456 15724 7496
rect 15764 7456 17452 7496
rect 17492 7456 17501 7496
rect 20140 7456 26572 7496
rect 26612 7456 26621 7496
rect 31363 7456 31372 7496
rect 31412 7456 31421 7496
rect 31854 7456 31948 7496
rect 31988 7456 31997 7496
rect 34915 7456 34924 7496
rect 34964 7456 40876 7496
rect 40916 7456 40925 7496
rect 41059 7456 41068 7496
rect 41108 7456 43008 7496
rect 0 7436 80 7456
rect 1804 7412 1844 7456
rect 6883 7412 6941 7413
rect 1795 7372 1804 7412
rect 1844 7372 6892 7412
rect 6932 7372 6941 7412
rect 6883 7371 6941 7372
rect 7555 7412 7613 7413
rect 20140 7412 20180 7456
rect 26563 7455 26621 7456
rect 31372 7412 31412 7456
rect 31939 7455 31997 7456
rect 42928 7436 43008 7456
rect 7555 7372 7564 7412
rect 7604 7372 8140 7412
rect 8180 7372 9812 7412
rect 10243 7372 10252 7412
rect 10292 7372 17740 7412
rect 17780 7372 17789 7412
rect 19171 7372 19180 7412
rect 19220 7372 20180 7412
rect 24547 7372 24556 7412
rect 24596 7372 24748 7412
rect 24788 7372 28300 7412
rect 28340 7372 31412 7412
rect 31459 7372 31468 7412
rect 31508 7372 31852 7412
rect 31892 7372 31901 7412
rect 32035 7372 32044 7412
rect 32084 7372 33196 7412
rect 33236 7372 33676 7412
rect 33716 7372 35308 7412
rect 35348 7372 35357 7412
rect 37795 7372 37804 7412
rect 37844 7372 38668 7412
rect 38708 7372 38717 7412
rect 40483 7372 40492 7412
rect 40532 7372 41260 7412
rect 41300 7372 41309 7412
rect 7555 7371 7613 7372
rect 9772 7328 9812 7372
rect 24739 7328 24797 7329
rect 2947 7288 2956 7328
rect 2996 7288 3148 7328
rect 3188 7288 3197 7328
rect 3811 7288 3820 7328
rect 3860 7288 4204 7328
rect 4244 7288 4253 7328
rect 9772 7288 13804 7328
rect 13844 7288 21676 7328
rect 21716 7288 22348 7328
rect 22388 7288 22397 7328
rect 24739 7288 24748 7328
rect 24788 7288 39148 7328
rect 39188 7288 41452 7328
rect 41492 7288 41501 7328
rect 24739 7287 24797 7288
rect 8803 7244 8861 7245
rect 11203 7244 11261 7245
rect 12835 7244 12893 7245
rect 35779 7244 35837 7245
rect 37795 7244 37853 7245
rect 2500 7204 8812 7244
rect 8852 7204 8861 7244
rect 10627 7204 10636 7244
rect 10676 7204 11212 7244
rect 11252 7204 11261 7244
rect 12750 7204 12844 7244
rect 12884 7204 12893 7244
rect 15043 7204 15052 7244
rect 15092 7204 15532 7244
rect 15572 7204 15581 7244
rect 18595 7204 18604 7244
rect 18644 7204 19468 7244
rect 19508 7204 19517 7244
rect 29059 7204 29068 7244
rect 29108 7204 29836 7244
rect 29876 7204 29885 7244
rect 30979 7204 30988 7244
rect 31028 7204 31468 7244
rect 31508 7204 31517 7244
rect 35694 7204 35788 7244
rect 35828 7204 35837 7244
rect 37710 7204 37804 7244
rect 37844 7204 38476 7244
rect 38516 7204 38525 7244
rect 0 7160 80 7180
rect 2500 7160 2540 7204
rect 8803 7203 8861 7204
rect 11203 7203 11261 7204
rect 12835 7203 12893 7204
rect 35779 7203 35837 7204
rect 37795 7203 37853 7204
rect 9475 7160 9533 7161
rect 17155 7160 17213 7161
rect 20995 7160 21053 7161
rect 22627 7160 22685 7161
rect 24739 7160 24797 7161
rect 30211 7160 30269 7161
rect 40771 7160 40829 7161
rect 42928 7160 43008 7180
rect 0 7120 2540 7160
rect 3139 7120 3148 7160
rect 3188 7120 3532 7160
rect 3572 7120 4204 7160
rect 4244 7120 4253 7160
rect 5827 7120 5836 7160
rect 5876 7120 8044 7160
rect 8084 7120 8093 7160
rect 9390 7120 9484 7160
rect 9524 7120 9533 7160
rect 13891 7120 13900 7160
rect 13940 7120 17164 7160
rect 17204 7120 17644 7160
rect 17684 7120 17693 7160
rect 18307 7120 18316 7160
rect 18356 7120 19372 7160
rect 19412 7120 19421 7160
rect 20910 7120 21004 7160
rect 21044 7120 22156 7160
rect 22196 7120 22205 7160
rect 22542 7120 22636 7160
rect 22676 7120 22685 7160
rect 24654 7120 24748 7160
rect 24788 7120 24797 7160
rect 27043 7120 27052 7160
rect 27092 7120 28148 7160
rect 30126 7120 30220 7160
rect 30260 7120 34924 7160
rect 34964 7120 34973 7160
rect 37699 7120 37708 7160
rect 37748 7120 39820 7160
rect 39860 7120 39869 7160
rect 40771 7120 40780 7160
rect 40820 7120 40972 7160
rect 41012 7120 41021 7160
rect 41635 7120 41644 7160
rect 41684 7120 43008 7160
rect 0 7100 80 7120
rect 9475 7119 9533 7120
rect 17155 7119 17213 7120
rect 20995 7119 21053 7120
rect 22627 7119 22685 7120
rect 24739 7119 24797 7120
rect 6595 7076 6653 7077
rect 28108 7076 28148 7120
rect 30211 7119 30269 7120
rect 40771 7119 40829 7120
rect 42928 7100 43008 7120
rect 2467 7036 2476 7076
rect 2516 7036 3820 7076
rect 3860 7036 3869 7076
rect 6510 7036 6604 7076
rect 6644 7036 6653 7076
rect 8803 7036 8812 7076
rect 8852 7036 13420 7076
rect 13460 7036 13469 7076
rect 15331 7036 15340 7076
rect 15380 7036 19852 7076
rect 19892 7036 19901 7076
rect 22915 7036 22924 7076
rect 22964 7036 28052 7076
rect 28108 7036 36268 7076
rect 36308 7036 36317 7076
rect 6595 7035 6653 7036
rect 21091 6992 21149 6993
rect 28012 6992 28052 7036
rect 30115 6992 30173 6993
rect 36163 6992 36221 6993
rect 1411 6952 1420 6992
rect 1460 6952 5356 6992
rect 5396 6952 5405 6992
rect 9667 6952 9676 6992
rect 9716 6952 10636 6992
rect 10676 6952 10685 6992
rect 11212 6952 13900 6992
rect 13940 6952 13949 6992
rect 15523 6952 15532 6992
rect 15572 6952 17164 6992
rect 17204 6952 17213 6992
rect 17635 6952 17644 6992
rect 17684 6952 21100 6992
rect 21140 6952 27916 6992
rect 27956 6952 27965 6992
rect 28012 6952 29972 6992
rect 3331 6908 3389 6909
rect 6403 6908 6461 6909
rect 11212 6908 11252 6952
rect 21091 6951 21149 6952
rect 20803 6908 20861 6909
rect 29932 6908 29972 6952
rect 30115 6952 30124 6992
rect 30164 6952 35884 6992
rect 35924 6952 35933 6992
rect 36078 6952 36172 6992
rect 36212 6952 36221 6992
rect 37699 6952 37708 6992
rect 37748 6952 37996 6992
rect 38036 6952 38045 6992
rect 30115 6951 30173 6952
rect 36163 6951 36221 6952
rect 3331 6868 3340 6908
rect 3380 6868 3436 6908
rect 3476 6868 3485 6908
rect 6318 6868 6412 6908
rect 6452 6868 6461 6908
rect 6787 6868 6796 6908
rect 6836 6868 7084 6908
rect 7124 6868 11252 6908
rect 11320 6868 12748 6908
rect 12788 6868 12797 6908
rect 13411 6868 13420 6908
rect 13460 6868 20812 6908
rect 20852 6868 26764 6908
rect 26804 6868 26813 6908
rect 28579 6868 28588 6908
rect 28628 6868 29876 6908
rect 29923 6868 29932 6908
rect 29972 6868 29981 6908
rect 30028 6868 32908 6908
rect 32948 6868 32957 6908
rect 3331 6867 3389 6868
rect 6403 6867 6461 6868
rect 0 6824 80 6844
rect 11320 6824 11360 6868
rect 17356 6824 17396 6868
rect 20803 6867 20861 6868
rect 26467 6824 26525 6825
rect 29836 6824 29876 6868
rect 30028 6824 30068 6868
rect 42928 6824 43008 6844
rect 0 6784 2540 6824
rect 4919 6784 4928 6824
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 5296 6784 5305 6824
rect 6211 6784 6220 6824
rect 6260 6784 9388 6824
rect 9428 6784 11360 6824
rect 17347 6784 17356 6824
rect 17396 6784 17436 6824
rect 17827 6784 17836 6824
rect 17876 6784 19180 6824
rect 19220 6784 19229 6824
rect 20039 6784 20048 6824
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20416 6784 20425 6824
rect 22243 6784 22252 6824
rect 22292 6784 22636 6824
rect 22676 6784 22685 6824
rect 24643 6784 24652 6824
rect 24692 6784 24940 6824
rect 24980 6784 24989 6824
rect 26467 6784 26476 6824
rect 26516 6784 29548 6824
rect 29588 6784 29597 6824
rect 29836 6784 30068 6824
rect 30115 6784 30124 6824
rect 30164 6784 32716 6824
rect 32756 6784 32765 6824
rect 35159 6784 35168 6824
rect 35208 6784 35250 6824
rect 35290 6784 35332 6824
rect 35372 6784 35414 6824
rect 35454 6784 35496 6824
rect 35536 6784 35545 6824
rect 38179 6784 38188 6824
rect 38228 6784 38860 6824
rect 38900 6784 38909 6824
rect 41059 6784 41068 6824
rect 41108 6784 43008 6824
rect 0 6764 80 6784
rect 2500 6572 2540 6784
rect 26467 6783 26525 6784
rect 42928 6764 43008 6784
rect 5164 6700 11596 6740
rect 11636 6700 11645 6740
rect 12364 6700 15916 6740
rect 15956 6700 16780 6740
rect 16820 6700 16829 6740
rect 23203 6700 23212 6740
rect 23252 6700 27148 6740
rect 27188 6700 27197 6740
rect 28675 6700 28684 6740
rect 28724 6700 29356 6740
rect 29396 6700 29405 6740
rect 31651 6700 31660 6740
rect 31700 6700 32140 6740
rect 32180 6700 32189 6740
rect 35212 6700 38092 6740
rect 38132 6700 38141 6740
rect 38284 6700 38764 6740
rect 38804 6700 38813 6740
rect 5164 6656 5204 6700
rect 5923 6656 5981 6657
rect 12364 6656 12404 6700
rect 31555 6656 31613 6657
rect 35212 6656 35252 6700
rect 38284 6656 38324 6700
rect 5155 6616 5164 6656
rect 5204 6616 5213 6656
rect 5838 6616 5932 6656
rect 5972 6616 5981 6656
rect 7555 6616 7564 6656
rect 7604 6616 7852 6656
rect 7892 6616 8140 6656
rect 8180 6616 8189 6656
rect 11011 6616 11020 6656
rect 11060 6616 12404 6656
rect 12451 6616 12460 6656
rect 12500 6616 13324 6656
rect 13364 6616 13373 6656
rect 15139 6616 15148 6656
rect 15188 6616 15340 6656
rect 15380 6616 15389 6656
rect 18595 6616 18604 6656
rect 18644 6616 25036 6656
rect 25076 6616 25085 6656
rect 25603 6616 25612 6656
rect 25652 6616 25661 6656
rect 28579 6616 28588 6656
rect 28628 6616 28876 6656
rect 28916 6616 28925 6656
rect 31470 6616 31564 6656
rect 31604 6616 31613 6656
rect 31939 6616 31948 6656
rect 31988 6616 33676 6656
rect 33716 6616 33725 6656
rect 34819 6616 34828 6656
rect 34868 6616 35212 6656
rect 35252 6616 35261 6656
rect 36355 6616 36364 6656
rect 36404 6616 36844 6656
rect 36884 6616 36893 6656
rect 37987 6616 37996 6656
rect 38036 6616 38324 6656
rect 5923 6615 5981 6616
rect 25612 6572 25652 6616
rect 31555 6615 31613 6616
rect 2500 6532 5204 6572
rect 6499 6532 6508 6572
rect 6548 6532 8236 6572
rect 8276 6532 8285 6572
rect 11395 6532 11404 6572
rect 11444 6532 20620 6572
rect 20660 6532 20669 6572
rect 25612 6532 33100 6572
rect 33140 6532 38284 6572
rect 38324 6532 38333 6572
rect 40003 6532 40012 6572
rect 40052 6532 42508 6572
rect 42548 6532 42557 6572
rect 0 6488 80 6508
rect 4195 6488 4253 6489
rect 0 6448 1132 6488
rect 1172 6448 1181 6488
rect 2947 6448 2956 6488
rect 2996 6448 3628 6488
rect 3668 6448 3677 6488
rect 4003 6448 4012 6488
rect 4052 6448 4204 6488
rect 4244 6448 4253 6488
rect 0 6428 80 6448
rect 4195 6447 4253 6448
rect 3427 6404 3485 6405
rect 4099 6404 4157 6405
rect 5164 6404 5204 6532
rect 6211 6488 6269 6489
rect 8803 6488 8861 6489
rect 17635 6488 17693 6489
rect 42928 6488 43008 6508
rect 5443 6448 5452 6488
rect 5492 6448 6220 6488
rect 6260 6448 6269 6488
rect 6883 6448 6892 6488
rect 6932 6448 8140 6488
rect 8180 6448 8189 6488
rect 8718 6448 8812 6488
rect 8852 6448 8861 6488
rect 9763 6448 9772 6488
rect 9812 6448 10732 6488
rect 10772 6448 10781 6488
rect 12643 6448 12652 6488
rect 12692 6448 14284 6488
rect 14324 6448 14333 6488
rect 17059 6448 17068 6488
rect 17108 6448 17452 6488
rect 17492 6448 17644 6488
rect 17684 6448 17693 6488
rect 6211 6447 6269 6448
rect 8803 6447 8861 6448
rect 17635 6447 17693 6448
rect 17740 6448 26668 6488
rect 26708 6448 26717 6488
rect 27139 6448 27148 6488
rect 27188 6448 27916 6488
rect 27956 6448 27965 6488
rect 28483 6448 28492 6488
rect 28532 6448 28876 6488
rect 28916 6448 28925 6488
rect 35212 6448 36116 6488
rect 39235 6448 39244 6488
rect 39284 6448 39724 6488
rect 39764 6448 39773 6488
rect 41443 6448 41452 6488
rect 41492 6448 43008 6488
rect 15427 6404 15485 6405
rect 17740 6404 17780 6448
rect 28291 6404 28349 6405
rect 32131 6404 32189 6405
rect 35212 6404 35252 6448
rect 3331 6364 3340 6404
rect 3380 6364 3436 6404
rect 3476 6364 3485 6404
rect 3811 6364 3820 6404
rect 3860 6364 4108 6404
rect 4148 6364 4157 6404
rect 3427 6363 3485 6364
rect 4099 6363 4157 6364
rect 4204 6364 4876 6404
rect 4916 6364 4925 6404
rect 5155 6364 5164 6404
rect 5204 6364 15436 6404
rect 15476 6364 15485 6404
rect 16579 6364 16588 6404
rect 16628 6364 17780 6404
rect 18979 6364 18988 6404
rect 19028 6364 19564 6404
rect 19604 6364 19756 6404
rect 19796 6364 19805 6404
rect 20140 6364 23308 6404
rect 23348 6364 23357 6404
rect 24739 6364 24748 6404
rect 24788 6364 26092 6404
rect 26132 6364 26141 6404
rect 28206 6364 28300 6404
rect 28340 6364 28349 6404
rect 32046 6364 32140 6404
rect 32180 6364 32189 6404
rect 32899 6364 32908 6404
rect 32948 6364 35252 6404
rect 4204 6320 4244 6364
rect 15427 6363 15485 6364
rect 9859 6320 9917 6321
rect 17548 6320 17588 6364
rect 19267 6320 19325 6321
rect 20140 6320 20180 6364
rect 28291 6363 28349 6364
rect 32131 6363 32189 6364
rect 2659 6280 2668 6320
rect 2708 6280 4204 6320
rect 4244 6280 4253 6320
rect 4483 6280 4492 6320
rect 4532 6280 5068 6320
rect 5108 6280 5117 6320
rect 5443 6280 5452 6320
rect 5492 6280 8428 6320
rect 8468 6280 8477 6320
rect 9859 6280 9868 6320
rect 9908 6280 10060 6320
rect 10100 6280 10109 6320
rect 10819 6280 10828 6320
rect 10868 6280 11116 6320
rect 11156 6280 11165 6320
rect 11971 6280 11980 6320
rect 12020 6280 12268 6320
rect 12308 6280 13900 6320
rect 13940 6280 15244 6320
rect 15284 6280 17260 6320
rect 17300 6280 17309 6320
rect 17539 6280 17548 6320
rect 17588 6280 17628 6320
rect 19267 6280 19276 6320
rect 19316 6280 20180 6320
rect 21475 6320 21533 6321
rect 35299 6320 35357 6321
rect 36076 6320 36116 6448
rect 42928 6428 43008 6448
rect 38947 6404 39005 6405
rect 38947 6364 38956 6404
rect 38996 6364 41260 6404
rect 41300 6364 41309 6404
rect 38947 6363 39005 6364
rect 40195 6320 40253 6321
rect 21475 6280 21484 6320
rect 21524 6280 27628 6320
rect 27668 6280 27677 6320
rect 29731 6280 29740 6320
rect 29780 6280 30220 6320
rect 30260 6280 30796 6320
rect 30836 6280 30845 6320
rect 31171 6280 31180 6320
rect 31220 6280 33772 6320
rect 33812 6280 33821 6320
rect 35299 6280 35308 6320
rect 35348 6280 35500 6320
rect 35540 6280 35549 6320
rect 35683 6280 35692 6320
rect 35732 6280 35884 6320
rect 35924 6280 35933 6320
rect 36076 6280 37652 6320
rect 40110 6280 40204 6320
rect 40244 6280 40253 6320
rect 9859 6279 9917 6280
rect 19267 6279 19325 6280
rect 21475 6279 21533 6280
rect 35299 6279 35357 6280
rect 3715 6196 3724 6236
rect 3764 6196 4300 6236
rect 4340 6196 4349 6236
rect 4963 6196 4972 6236
rect 5012 6196 12364 6236
rect 12404 6196 18604 6236
rect 18644 6196 18653 6236
rect 24835 6196 24844 6236
rect 24884 6196 28588 6236
rect 28628 6196 28637 6236
rect 32803 6196 32812 6236
rect 32852 6196 33580 6236
rect 33620 6196 33629 6236
rect 0 6152 80 6172
rect 5347 6152 5405 6153
rect 6403 6152 6461 6153
rect 7651 6152 7709 6153
rect 21379 6152 21437 6153
rect 37612 6152 37652 6280
rect 40195 6279 40253 6280
rect 38179 6236 38237 6237
rect 38094 6196 38188 6236
rect 38228 6196 38237 6236
rect 39619 6196 39628 6236
rect 39668 6196 40876 6236
rect 40916 6196 40925 6236
rect 38179 6195 38237 6196
rect 42928 6152 43008 6172
rect 0 6112 5356 6152
rect 5396 6112 5405 6152
rect 6307 6112 6316 6152
rect 6356 6112 6412 6152
rect 6452 6112 6461 6152
rect 7566 6112 7660 6152
rect 7700 6112 7709 6152
rect 10531 6112 10540 6152
rect 10580 6112 21388 6152
rect 21428 6112 21437 6152
rect 24547 6112 24556 6152
rect 24596 6112 25132 6152
rect 25172 6112 25181 6152
rect 37612 6112 37804 6152
rect 37844 6112 37853 6152
rect 41059 6112 41068 6152
rect 41108 6112 43008 6152
rect 0 6092 80 6112
rect 5347 6111 5405 6112
rect 6403 6111 6461 6112
rect 7651 6111 7709 6112
rect 21379 6111 21437 6112
rect 42928 6092 43008 6112
rect 3679 6028 3688 6068
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 4056 6028 4065 6068
rect 6883 6028 6892 6068
rect 6932 6028 12652 6068
rect 12692 6028 12701 6068
rect 16771 6028 16780 6068
rect 16820 6028 18124 6068
rect 18164 6028 18173 6068
rect 18799 6028 18808 6068
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 19176 6028 19185 6068
rect 33919 6028 33928 6068
rect 33968 6028 34010 6068
rect 34050 6028 34092 6068
rect 34132 6028 34174 6068
rect 34214 6028 34256 6068
rect 34296 6028 34305 6068
rect 24739 5984 24797 5985
rect 1315 5944 1324 5984
rect 1364 5944 1804 5984
rect 1844 5944 1853 5984
rect 3148 5944 11020 5984
rect 11060 5944 11069 5984
rect 18403 5944 18412 5984
rect 18452 5944 19468 5984
rect 19508 5944 19517 5984
rect 22531 5944 22540 5984
rect 22580 5944 24748 5984
rect 24788 5944 31852 5984
rect 31892 5944 31901 5984
rect 34723 5944 34732 5984
rect 34772 5944 36844 5984
rect 36884 5944 37516 5984
rect 37556 5944 37565 5984
rect 0 5816 80 5836
rect 3148 5816 3188 5944
rect 24739 5943 24797 5944
rect 9955 5860 9964 5900
rect 10004 5860 10013 5900
rect 10531 5860 10540 5900
rect 10580 5860 10964 5900
rect 17731 5860 17740 5900
rect 17780 5860 19372 5900
rect 19412 5860 20524 5900
rect 20564 5860 20573 5900
rect 36643 5860 36652 5900
rect 36692 5860 37036 5900
rect 37076 5860 37085 5900
rect 38563 5860 38572 5900
rect 38612 5860 38956 5900
rect 38996 5860 39005 5900
rect 40003 5860 40012 5900
rect 40052 5860 41356 5900
rect 41396 5860 41405 5900
rect 3619 5816 3677 5817
rect 0 5776 3148 5816
rect 3188 5776 3197 5816
rect 3427 5776 3436 5816
rect 3476 5776 3628 5816
rect 3668 5776 3677 5816
rect 9964 5816 10004 5860
rect 10924 5816 10964 5860
rect 19267 5816 19325 5817
rect 42928 5816 43008 5836
rect 9964 5776 10580 5816
rect 10915 5776 10924 5816
rect 10964 5776 10973 5816
rect 13987 5776 13996 5816
rect 14036 5776 16052 5816
rect 16483 5776 16492 5816
rect 16532 5776 17068 5816
rect 17108 5776 17117 5816
rect 19267 5776 19276 5816
rect 19316 5776 29000 5816
rect 30019 5776 30028 5816
rect 30068 5776 38764 5816
rect 38804 5776 38813 5816
rect 41443 5776 41452 5816
rect 41492 5776 43008 5816
rect 0 5756 80 5776
rect 3619 5775 3677 5776
rect 10540 5732 10580 5776
rect 15907 5732 15965 5733
rect 2851 5692 2860 5732
rect 2900 5692 4972 5732
rect 5012 5692 5021 5732
rect 9571 5692 9580 5732
rect 9620 5692 9998 5732
rect 10038 5692 10047 5732
rect 10531 5692 10540 5732
rect 10580 5692 10828 5732
rect 10868 5692 10877 5732
rect 11683 5692 11692 5732
rect 11732 5692 15916 5732
rect 15956 5692 15965 5732
rect 16012 5732 16052 5776
rect 19267 5775 19325 5776
rect 19555 5732 19613 5733
rect 21187 5732 21245 5733
rect 26659 5732 26717 5733
rect 28960 5732 29000 5776
rect 42928 5756 43008 5776
rect 16012 5692 19180 5732
rect 19220 5692 19229 5732
rect 19555 5692 19564 5732
rect 19604 5692 20180 5732
rect 21102 5692 21196 5732
rect 21236 5692 21245 5732
rect 26563 5692 26572 5732
rect 26612 5692 26668 5732
rect 26708 5692 27436 5732
rect 27476 5692 27916 5732
rect 27956 5692 27965 5732
rect 28960 5692 37612 5732
rect 37652 5692 37661 5732
rect 15907 5691 15965 5692
rect 19555 5691 19613 5692
rect 3331 5648 3389 5649
rect 20140 5648 20180 5692
rect 21187 5691 21245 5692
rect 26659 5691 26717 5692
rect 24355 5648 24413 5649
rect 27916 5648 27956 5692
rect 30019 5648 30077 5649
rect 35587 5648 35645 5649
rect 3246 5608 3340 5648
rect 3380 5608 3389 5648
rect 4867 5608 4876 5648
rect 4916 5608 5356 5648
rect 5396 5608 5405 5648
rect 14275 5608 14284 5648
rect 14324 5608 16492 5648
rect 16532 5608 16541 5648
rect 20140 5608 24364 5648
rect 24404 5608 24413 5648
rect 25987 5608 25996 5648
rect 26036 5608 27340 5648
rect 27380 5608 27389 5648
rect 27916 5608 29548 5648
rect 29588 5608 30028 5648
rect 30068 5608 30077 5648
rect 32515 5608 32524 5648
rect 32564 5608 32812 5648
rect 32852 5608 33196 5648
rect 33236 5608 34540 5648
rect 34580 5608 34732 5648
rect 34772 5608 34781 5648
rect 35502 5608 35596 5648
rect 35636 5608 35645 5648
rect 36259 5608 36268 5648
rect 36308 5608 38996 5648
rect 3331 5607 3389 5608
rect 24355 5607 24413 5608
rect 30019 5607 30077 5608
rect 35587 5607 35645 5608
rect 18115 5564 18173 5565
rect 1123 5524 1132 5564
rect 1172 5524 6796 5564
rect 6836 5524 6845 5564
rect 8227 5524 8236 5564
rect 8276 5524 8524 5564
rect 8564 5524 8573 5564
rect 8995 5524 9004 5564
rect 9044 5524 11360 5564
rect 12931 5524 12940 5564
rect 12980 5524 18068 5564
rect 0 5480 80 5500
rect 3619 5480 3677 5481
rect 11320 5480 11360 5524
rect 0 5440 1324 5480
rect 1364 5440 1373 5480
rect 3534 5440 3628 5480
rect 3668 5440 3677 5480
rect 4099 5440 4108 5480
rect 4148 5440 4972 5480
rect 5012 5440 5021 5480
rect 8803 5440 8812 5480
rect 8852 5440 10156 5480
rect 10196 5440 10205 5480
rect 11320 5440 14476 5480
rect 14516 5440 14525 5480
rect 0 5420 80 5440
rect 3619 5439 3677 5440
rect 17827 5396 17885 5397
rect 2275 5356 2284 5396
rect 2324 5356 13996 5396
rect 14036 5356 14045 5396
rect 16483 5356 16492 5396
rect 16532 5356 17836 5396
rect 17876 5356 17885 5396
rect 17827 5355 17885 5356
rect 18028 5312 18068 5524
rect 18115 5524 18124 5564
rect 18164 5524 18258 5564
rect 19747 5524 19756 5564
rect 19796 5524 27436 5564
rect 27476 5524 27485 5564
rect 27532 5524 29164 5564
rect 29204 5524 36556 5564
rect 36596 5524 36605 5564
rect 18115 5523 18173 5524
rect 27532 5480 27572 5524
rect 37219 5480 37277 5481
rect 38956 5480 38996 5608
rect 42928 5480 43008 5500
rect 20803 5440 20812 5480
rect 20852 5440 21004 5480
rect 21044 5440 22636 5480
rect 22676 5440 22685 5480
rect 24931 5440 24940 5480
rect 24980 5440 27572 5480
rect 28003 5440 28012 5480
rect 28052 5440 35212 5480
rect 35252 5440 35261 5480
rect 35395 5440 35404 5480
rect 35444 5440 36364 5480
rect 36404 5440 36413 5480
rect 37134 5440 37228 5480
rect 37268 5440 37277 5480
rect 38947 5440 38956 5480
rect 38996 5440 39916 5480
rect 39956 5440 39965 5480
rect 41347 5440 41356 5480
rect 41396 5440 43008 5480
rect 37219 5439 37277 5440
rect 42928 5420 43008 5440
rect 23875 5396 23933 5397
rect 26467 5396 26525 5397
rect 19171 5356 19180 5396
rect 19220 5356 21388 5396
rect 21428 5356 22540 5396
rect 22580 5356 22589 5396
rect 23875 5356 23884 5396
rect 23924 5356 26092 5396
rect 26132 5356 26141 5396
rect 26467 5356 26476 5396
rect 26516 5356 30124 5396
rect 30164 5356 30173 5396
rect 31075 5356 31084 5396
rect 31124 5356 31316 5396
rect 32419 5356 32428 5396
rect 32468 5356 36940 5396
rect 36980 5356 36989 5396
rect 23875 5355 23933 5356
rect 3523 5272 3532 5312
rect 3572 5272 3724 5312
rect 3764 5272 3773 5312
rect 4919 5272 4928 5312
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 5296 5272 5305 5312
rect 6403 5272 6412 5312
rect 6452 5272 8044 5312
rect 8084 5272 8093 5312
rect 11299 5272 11308 5312
rect 11348 5272 15628 5312
rect 15668 5272 15677 5312
rect 18028 5272 19892 5312
rect 20039 5272 20048 5312
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20416 5272 20425 5312
rect 12451 5228 12509 5229
rect 19852 5228 19892 5272
rect 26092 5228 26132 5356
rect 26467 5355 26525 5356
rect 31276 5312 31316 5356
rect 27619 5272 27628 5312
rect 27668 5272 27916 5312
rect 27956 5272 27965 5312
rect 30211 5272 30220 5312
rect 30260 5272 31180 5312
rect 31220 5272 31229 5312
rect 31276 5272 32716 5312
rect 32756 5272 32765 5312
rect 35159 5272 35168 5312
rect 35208 5272 35250 5312
rect 35290 5272 35332 5312
rect 35372 5272 35414 5312
rect 35454 5272 35496 5312
rect 35536 5272 35545 5312
rect 1315 5188 1324 5228
rect 1364 5188 6892 5228
rect 6932 5188 6941 5228
rect 7939 5188 7948 5228
rect 7988 5188 8332 5228
rect 8372 5188 8381 5228
rect 10051 5188 10060 5228
rect 10100 5188 10636 5228
rect 10676 5188 10685 5228
rect 11587 5188 11596 5228
rect 11636 5188 11788 5228
rect 11828 5188 11837 5228
rect 12067 5188 12076 5228
rect 12116 5188 12125 5228
rect 12451 5188 12460 5228
rect 12500 5188 19756 5228
rect 19796 5188 19805 5228
rect 19852 5188 25652 5228
rect 26092 5188 30700 5228
rect 30740 5188 39628 5228
rect 39668 5188 39677 5228
rect 0 5144 80 5164
rect 1315 5144 1373 5145
rect 4099 5144 4157 5145
rect 12076 5144 12116 5188
rect 12451 5187 12509 5188
rect 0 5104 1324 5144
rect 1364 5104 1373 5144
rect 3427 5104 3436 5144
rect 3476 5104 3485 5144
rect 4099 5104 4108 5144
rect 4148 5104 4300 5144
rect 4340 5104 4349 5144
rect 6787 5104 6796 5144
rect 6836 5104 11360 5144
rect 12076 5104 20180 5144
rect 20419 5104 20428 5144
rect 20468 5104 20812 5144
rect 20852 5104 20861 5144
rect 22915 5104 22924 5144
rect 22964 5104 23500 5144
rect 23540 5104 23549 5144
rect 24067 5104 24076 5144
rect 24116 5104 24460 5144
rect 24500 5104 24509 5144
rect 0 5084 80 5104
rect 1315 5103 1373 5104
rect 3436 5060 3476 5104
rect 4099 5103 4157 5104
rect 5347 5060 5405 5061
rect 11320 5060 11360 5104
rect 12547 5060 12605 5061
rect 20140 5060 20180 5104
rect 25612 5060 25652 5188
rect 42928 5144 43008 5164
rect 27427 5104 27436 5144
rect 27476 5104 33484 5144
rect 33524 5104 33533 5144
rect 36163 5104 36172 5144
rect 36212 5104 36556 5144
rect 36596 5104 36605 5144
rect 40387 5104 40396 5144
rect 40436 5104 40972 5144
rect 41012 5104 41021 5144
rect 41443 5104 41452 5144
rect 41492 5104 43008 5144
rect 42928 5084 43008 5104
rect 27715 5060 27773 5061
rect 30883 5060 30941 5061
rect 40291 5060 40349 5061
rect 2947 5020 2956 5060
rect 2996 5020 3476 5060
rect 3715 5020 3724 5060
rect 3764 5020 5068 5060
rect 5108 5020 5117 5060
rect 5251 5020 5260 5060
rect 5300 5020 5356 5060
rect 5396 5020 5405 5060
rect 6595 5020 6604 5060
rect 6644 5020 7276 5060
rect 7316 5020 7325 5060
rect 7555 5020 7564 5060
rect 7604 5020 7756 5060
rect 7796 5020 7805 5060
rect 8515 5020 8524 5060
rect 8564 5020 8852 5060
rect 8995 5020 9004 5060
rect 9044 5020 10732 5060
rect 10772 5020 10781 5060
rect 11320 5020 12556 5060
rect 12596 5020 12605 5060
rect 13603 5020 13612 5060
rect 13652 5020 14092 5060
rect 14132 5020 14141 5060
rect 15139 5020 15148 5060
rect 15188 5020 15820 5060
rect 15860 5020 15869 5060
rect 16771 5020 16780 5060
rect 16820 5020 16829 5060
rect 17539 5020 17548 5060
rect 17588 5020 18028 5060
rect 18068 5020 18077 5060
rect 20140 5020 25516 5060
rect 25556 5020 25565 5060
rect 25612 5020 27724 5060
rect 27764 5020 27773 5060
rect 30798 5020 30892 5060
rect 30932 5020 30941 5060
rect 35971 5020 35980 5060
rect 36020 5020 40300 5060
rect 40340 5020 40349 5060
rect 5347 5019 5405 5020
rect 7171 4976 7229 4977
rect 8812 4976 8852 5020
rect 12547 5019 12605 5020
rect 10627 4976 10685 4977
rect 16780 4976 16820 5020
rect 27715 5019 27773 5020
rect 30883 5019 30941 5020
rect 40291 5019 40349 5020
rect 19363 4976 19421 4977
rect 27139 4976 27197 4977
rect 28003 4976 28061 4977
rect 31267 4976 31325 4977
rect 40771 4976 40829 4977
rect 2659 4936 2668 4976
rect 2708 4936 3244 4976
rect 3284 4936 4492 4976
rect 4532 4936 6796 4976
rect 6836 4936 6845 4976
rect 6979 4936 6988 4976
rect 7028 4936 7037 4976
rect 7171 4936 7180 4976
rect 7220 4936 7314 4976
rect 8803 4936 8812 4976
rect 8852 4936 9772 4976
rect 9812 4936 10156 4976
rect 10196 4936 10205 4976
rect 10542 4936 10636 4976
rect 10676 4936 10685 4976
rect 13315 4936 13324 4976
rect 13364 4936 16820 4976
rect 17347 4936 17356 4976
rect 17396 4936 18508 4976
rect 18548 4936 18557 4976
rect 19171 4936 19180 4976
rect 19220 4936 19372 4976
rect 19412 4936 19421 4976
rect 24259 4936 24268 4976
rect 24308 4936 24652 4976
rect 24692 4936 24701 4976
rect 25891 4936 25900 4976
rect 25940 4936 26572 4976
rect 26612 4936 26621 4976
rect 27054 4936 27148 4976
rect 27188 4936 27197 4976
rect 27907 4936 27916 4976
rect 27956 4936 28012 4976
rect 28052 4936 28061 4976
rect 31182 4936 31276 4976
rect 31316 4936 31325 4976
rect 6988 4892 7028 4936
rect 7171 4935 7229 4936
rect 10627 4935 10685 4936
rect 19363 4935 19421 4936
rect 8803 4892 8861 4893
rect 9475 4892 9533 4893
rect 17827 4892 17885 4893
rect 25900 4892 25940 4936
rect 27139 4935 27197 4936
rect 28003 4935 28061 4936
rect 31267 4935 31325 4936
rect 32332 4936 35596 4976
rect 35636 4936 39052 4976
rect 39092 4936 39101 4976
rect 40686 4936 40780 4976
rect 40820 4936 40829 4976
rect 32332 4892 32372 4936
rect 40771 4935 40829 4936
rect 37891 4892 37949 4893
rect 41251 4892 41309 4893
rect 2755 4852 2764 4892
rect 2804 4852 2956 4892
rect 2996 4852 7028 4892
rect 7267 4852 7276 4892
rect 7316 4852 8812 4892
rect 8852 4852 9484 4892
rect 9524 4852 9533 4892
rect 15235 4852 15244 4892
rect 15284 4852 17548 4892
rect 17588 4852 17597 4892
rect 17742 4852 17836 4892
rect 17876 4852 17885 4892
rect 18307 4852 18316 4892
rect 18356 4852 18796 4892
rect 18836 4852 18845 4892
rect 22723 4852 22732 4892
rect 22772 4852 23692 4892
rect 23732 4852 25940 4892
rect 28195 4852 28204 4892
rect 28244 4852 29396 4892
rect 29635 4852 29644 4892
rect 29684 4852 30412 4892
rect 30452 4852 32372 4892
rect 32419 4852 32428 4892
rect 32468 4852 33100 4892
rect 33140 4852 33149 4892
rect 33196 4852 35980 4892
rect 36020 4852 36029 4892
rect 37891 4852 37900 4892
rect 37940 4852 39148 4892
rect 39188 4852 39197 4892
rect 41166 4852 41260 4892
rect 41300 4852 41309 4892
rect 8803 4851 8861 4852
rect 9475 4851 9533 4852
rect 17827 4851 17885 4852
rect 0 4808 80 4828
rect 19939 4808 19997 4809
rect 29356 4808 29396 4852
rect 33196 4808 33236 4852
rect 37891 4851 37949 4852
rect 41251 4851 41309 4852
rect 34915 4808 34973 4809
rect 42928 4808 43008 4828
rect 0 4768 10444 4808
rect 10484 4768 10493 4808
rect 14851 4768 14860 4808
rect 14900 4768 17068 4808
rect 17108 4768 18028 4808
rect 18068 4768 18077 4808
rect 19939 4768 19948 4808
rect 19988 4768 20236 4808
rect 20276 4768 20285 4808
rect 22339 4768 22348 4808
rect 22388 4768 29260 4808
rect 29300 4768 29309 4808
rect 29356 4768 29740 4808
rect 29780 4768 30316 4808
rect 30356 4768 33236 4808
rect 34830 4768 34924 4808
rect 34964 4768 34973 4808
rect 39331 4768 39340 4808
rect 39380 4768 40300 4808
rect 40340 4768 40349 4808
rect 41068 4768 43008 4808
rect 0 4748 80 4768
rect 19939 4767 19997 4768
rect 34915 4767 34973 4768
rect 3427 4724 3485 4725
rect 4195 4724 4253 4725
rect 7171 4724 7229 4725
rect 9859 4724 9917 4725
rect 27619 4724 27677 4725
rect 32899 4724 32957 4725
rect 41068 4724 41108 4768
rect 42928 4748 43008 4768
rect 41539 4724 41597 4725
rect 3342 4684 3436 4724
rect 3476 4684 3485 4724
rect 4003 4684 4012 4724
rect 4052 4684 4204 4724
rect 4244 4684 4253 4724
rect 6211 4684 6220 4724
rect 6260 4684 6604 4724
rect 6644 4684 7180 4724
rect 7220 4684 7229 4724
rect 8035 4684 8044 4724
rect 8084 4684 9868 4724
rect 9908 4684 9917 4724
rect 16771 4684 16780 4724
rect 16820 4684 16972 4724
rect 17012 4684 17021 4724
rect 20140 4684 21292 4724
rect 21332 4684 21341 4724
rect 24451 4684 24460 4724
rect 24500 4684 24844 4724
rect 24884 4684 24893 4724
rect 27534 4684 27628 4724
rect 27668 4684 27677 4724
rect 3427 4683 3485 4684
rect 4195 4683 4253 4684
rect 7171 4683 7229 4684
rect 9859 4683 9917 4684
rect 6691 4600 6700 4640
rect 6740 4600 9484 4640
rect 9524 4600 10348 4640
rect 10388 4600 10397 4640
rect 11971 4600 11980 4640
rect 12020 4600 12844 4640
rect 12884 4600 19412 4640
rect 4195 4556 4253 4557
rect 19372 4556 19412 4600
rect 20140 4556 20180 4684
rect 27619 4683 27677 4684
rect 27724 4684 28780 4724
rect 28820 4684 32756 4724
rect 32814 4684 32908 4724
rect 32948 4684 32957 4724
rect 34339 4684 34348 4724
rect 34388 4684 34732 4724
rect 34772 4684 34781 4724
rect 39235 4684 39244 4724
rect 39284 4684 39532 4724
rect 39572 4684 39581 4724
rect 41059 4684 41068 4724
rect 41108 4684 41117 4724
rect 41454 4684 41548 4724
rect 41588 4684 41597 4724
rect 27724 4640 27764 4684
rect 32716 4640 32756 4684
rect 32899 4683 32957 4684
rect 41539 4683 41597 4684
rect 27715 4600 27724 4640
rect 27764 4600 27773 4640
rect 28960 4600 30796 4640
rect 30836 4600 30845 4640
rect 32035 4600 32044 4640
rect 32084 4600 32524 4640
rect 32564 4600 32573 4640
rect 32716 4600 36556 4640
rect 36596 4600 36605 4640
rect 28960 4556 29000 4600
rect 3679 4516 3688 4556
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 4056 4516 4065 4556
rect 4195 4516 4204 4556
rect 4244 4516 6836 4556
rect 6883 4516 6892 4556
rect 6932 4516 7372 4556
rect 7412 4516 7421 4556
rect 9379 4516 9388 4556
rect 9428 4516 12460 4556
rect 12500 4516 16916 4556
rect 18799 4516 18808 4556
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 19176 4516 19185 4556
rect 19363 4516 19372 4556
rect 19412 4516 20180 4556
rect 21196 4516 22828 4556
rect 22868 4516 22877 4556
rect 26275 4516 26284 4556
rect 26324 4516 29000 4556
rect 33919 4516 33928 4556
rect 33968 4516 34010 4556
rect 34050 4516 34092 4556
rect 34132 4516 34174 4556
rect 34214 4516 34256 4556
rect 34296 4516 34305 4556
rect 34435 4516 34444 4556
rect 34484 4516 35116 4556
rect 35156 4516 35165 4556
rect 4195 4515 4253 4516
rect 0 4472 80 4492
rect 6796 4472 6836 4516
rect 0 4432 1132 4472
rect 1172 4432 1181 4472
rect 4684 4432 6412 4472
rect 6452 4432 6461 4472
rect 6796 4432 8428 4472
rect 8468 4432 10732 4472
rect 10772 4432 10781 4472
rect 0 4412 80 4432
rect 4684 4388 4724 4432
rect 16876 4388 16916 4516
rect 21196 4472 21236 4516
rect 16963 4432 16972 4472
rect 17012 4432 21236 4472
rect 22051 4472 22109 4473
rect 42928 4472 43008 4492
rect 22051 4432 22060 4472
rect 22100 4432 27532 4472
rect 27572 4432 27581 4472
rect 32323 4432 32332 4472
rect 32372 4432 43008 4472
rect 22051 4431 22109 4432
rect 42928 4412 43008 4432
rect 21091 4388 21149 4389
rect 4195 4348 4204 4388
rect 4244 4348 4684 4388
rect 4724 4348 4733 4388
rect 8803 4348 8812 4388
rect 8852 4348 10252 4388
rect 10292 4348 10301 4388
rect 13987 4348 13996 4388
rect 14036 4348 14764 4388
rect 14804 4348 14813 4388
rect 16483 4348 16492 4388
rect 16532 4348 16684 4388
rect 16724 4348 16733 4388
rect 16876 4348 21100 4388
rect 21140 4348 21149 4388
rect 21091 4347 21149 4348
rect 21379 4388 21437 4389
rect 27139 4388 27197 4389
rect 21379 4348 21388 4388
rect 21428 4348 21676 4388
rect 21716 4348 27148 4388
rect 27188 4348 27197 4388
rect 28579 4348 28588 4388
rect 28628 4348 29164 4388
rect 29204 4348 29213 4388
rect 35260 4348 36076 4388
rect 36116 4348 36460 4388
rect 36500 4348 40108 4388
rect 40148 4348 40157 4388
rect 21379 4347 21437 4348
rect 27139 4347 27197 4348
rect 35260 4304 35300 4348
rect 4579 4264 4588 4304
rect 4628 4264 8524 4304
rect 8564 4264 9388 4304
rect 9428 4264 9437 4304
rect 10339 4264 10348 4304
rect 10388 4264 14668 4304
rect 14708 4264 23212 4304
rect 23252 4264 23261 4304
rect 24259 4264 24268 4304
rect 24308 4264 24556 4304
rect 24596 4264 24605 4304
rect 27052 4264 27628 4304
rect 27668 4264 27677 4304
rect 27811 4264 27820 4304
rect 27860 4264 28396 4304
rect 28436 4264 28445 4304
rect 33187 4264 33196 4304
rect 33236 4264 35300 4304
rect 36835 4264 36844 4304
rect 36884 4264 37996 4304
rect 38036 4264 38045 4304
rect 38668 4264 39628 4304
rect 39668 4264 39677 4304
rect 7171 4220 7229 4221
rect 12547 4220 12605 4221
rect 21091 4220 21149 4221
rect 21283 4220 21341 4221
rect 27052 4220 27092 4264
rect 33475 4220 33533 4221
rect 76 4180 212 4220
rect 76 4156 116 4180
rect 0 4096 116 4156
rect 0 4076 80 4096
rect 172 3968 212 4180
rect 7171 4180 7180 4220
rect 7220 4180 8140 4220
rect 8180 4180 9100 4220
rect 9140 4180 9676 4220
rect 9716 4180 9725 4220
rect 9772 4180 11980 4220
rect 12020 4180 12029 4220
rect 12163 4180 12172 4220
rect 12212 4180 12556 4220
rect 12596 4180 12605 4220
rect 12739 4180 12748 4220
rect 12788 4180 13228 4220
rect 13268 4180 14284 4220
rect 14324 4180 16972 4220
rect 17012 4180 17021 4220
rect 19843 4180 19852 4220
rect 19892 4180 20332 4220
rect 20372 4180 20381 4220
rect 21091 4180 21100 4220
rect 21140 4180 21292 4220
rect 21332 4180 21964 4220
rect 22004 4180 22013 4220
rect 24067 4180 24076 4220
rect 24116 4180 27052 4220
rect 27092 4180 27101 4220
rect 27235 4180 27244 4220
rect 27284 4180 33292 4220
rect 33332 4180 33341 4220
rect 33475 4180 33484 4220
rect 33524 4180 38284 4220
rect 38324 4180 38333 4220
rect 7171 4179 7229 4180
rect 1315 4136 1373 4137
rect 9772 4136 9812 4180
rect 12547 4179 12605 4180
rect 21091 4179 21149 4180
rect 21283 4179 21341 4180
rect 33475 4179 33533 4180
rect 1230 4096 1324 4136
rect 1364 4096 1373 4136
rect 3139 4096 3148 4136
rect 3188 4096 8332 4136
rect 8372 4096 8381 4136
rect 9571 4096 9580 4136
rect 9620 4096 9812 4136
rect 9859 4136 9917 4137
rect 13795 4136 13853 4137
rect 38668 4136 38708 4264
rect 38851 4220 38909 4221
rect 38766 4180 38860 4220
rect 38900 4180 41356 4220
rect 41396 4180 41405 4220
rect 38851 4179 38909 4180
rect 42928 4136 43008 4156
rect 9859 4096 9868 4136
rect 9908 4096 11788 4136
rect 11828 4096 11837 4136
rect 12547 4096 12556 4136
rect 12596 4096 13804 4136
rect 13844 4096 13853 4136
rect 18403 4096 18412 4136
rect 18452 4096 21484 4136
rect 21524 4096 21533 4136
rect 21580 4096 27436 4136
rect 27476 4096 27485 4136
rect 27619 4096 27628 4136
rect 27668 4096 32812 4136
rect 32852 4096 32861 4136
rect 36067 4096 36076 4136
rect 36116 4096 38708 4136
rect 38755 4096 38764 4136
rect 38804 4096 43008 4136
rect 1315 4095 1373 4096
rect 9859 4095 9917 4096
rect 13795 4095 13853 4096
rect 7171 4052 7229 4053
rect 7459 4052 7517 4053
rect 20035 4052 20093 4053
rect 21580 4052 21620 4096
rect 42928 4076 43008 4096
rect 6979 4012 6988 4052
rect 7028 4012 7180 4052
rect 7220 4012 7229 4052
rect 7374 4012 7468 4052
rect 7508 4012 9772 4052
rect 9812 4012 9821 4052
rect 10348 4012 12940 4052
rect 12980 4012 20044 4052
rect 20084 4012 20093 4052
rect 20419 4012 20428 4052
rect 20468 4012 21620 4052
rect 24067 4012 24076 4052
rect 24116 4012 25036 4052
rect 25076 4012 25085 4052
rect 26380 4012 31756 4052
rect 31796 4012 33772 4052
rect 33812 4012 36652 4052
rect 36692 4012 37036 4052
rect 37076 4012 39188 4052
rect 40771 4012 40780 4052
rect 40820 4012 41740 4052
rect 41780 4012 41789 4052
rect 7171 4011 7229 4012
rect 7459 4011 7517 4012
rect 7843 3968 7901 3969
rect 172 3928 3532 3968
rect 3572 3928 3581 3968
rect 4771 3928 4780 3968
rect 4820 3928 6796 3968
rect 6836 3928 6845 3968
rect 7555 3928 7564 3968
rect 7604 3928 7852 3968
rect 7892 3928 10156 3968
rect 10196 3928 10205 3968
rect 7843 3927 7901 3928
rect 2755 3844 2764 3884
rect 2804 3844 3148 3884
rect 3188 3844 3197 3884
rect 4675 3844 4684 3884
rect 4724 3844 5356 3884
rect 5396 3844 5405 3884
rect 7075 3844 7084 3884
rect 7124 3844 7372 3884
rect 7412 3844 9580 3884
rect 9620 3844 9629 3884
rect 0 3800 80 3820
rect 8803 3800 8861 3801
rect 10348 3800 10388 4012
rect 20035 4011 20093 4012
rect 20131 3968 20189 3969
rect 10723 3928 10732 3968
rect 10772 3928 11884 3968
rect 11924 3928 11933 3968
rect 12259 3928 12268 3968
rect 12308 3928 13420 3968
rect 13460 3928 13804 3968
rect 13844 3928 13853 3968
rect 15907 3928 15916 3968
rect 15956 3928 16300 3968
rect 16340 3928 16349 3968
rect 17251 3928 17260 3968
rect 17300 3928 20140 3968
rect 20180 3928 20189 3968
rect 20131 3927 20189 3928
rect 20323 3968 20381 3969
rect 20323 3928 20332 3968
rect 20372 3928 26284 3968
rect 26324 3928 26333 3968
rect 20323 3927 20381 3928
rect 10531 3844 10540 3884
rect 10580 3844 18892 3884
rect 18932 3844 18941 3884
rect 19651 3844 19660 3884
rect 19700 3844 19709 3884
rect 21484 3844 21812 3884
rect 21859 3844 21868 3884
rect 21908 3844 22444 3884
rect 22484 3844 24748 3884
rect 24788 3844 25612 3884
rect 25652 3844 25661 3884
rect 19660 3800 19700 3844
rect 21484 3800 21524 3844
rect 21667 3800 21725 3801
rect 0 3760 4820 3800
rect 4919 3760 4928 3800
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 5296 3760 5305 3800
rect 5356 3760 8428 3800
rect 8468 3760 8477 3800
rect 8718 3760 8812 3800
rect 8852 3760 8861 3800
rect 10339 3760 10348 3800
rect 10388 3760 10397 3800
rect 12355 3760 12364 3800
rect 12404 3760 12413 3800
rect 15523 3760 15532 3800
rect 15572 3760 16012 3800
rect 16052 3760 18604 3800
rect 18644 3760 18653 3800
rect 19180 3760 19700 3800
rect 19939 3760 19948 3800
rect 19988 3760 19997 3800
rect 20039 3760 20048 3800
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20416 3760 20425 3800
rect 20995 3760 21004 3800
rect 21044 3760 21524 3800
rect 21582 3760 21676 3800
rect 21716 3760 21725 3800
rect 21772 3800 21812 3844
rect 26380 3800 26420 4012
rect 28387 3968 28445 3969
rect 37603 3968 37661 3969
rect 28302 3928 28396 3968
rect 28436 3928 28445 3968
rect 28771 3928 28780 3968
rect 28820 3928 28972 3968
rect 29012 3928 29021 3968
rect 33667 3928 33676 3968
rect 33716 3928 37612 3968
rect 37652 3928 37661 3968
rect 28387 3927 28445 3928
rect 37603 3927 37661 3928
rect 37795 3968 37853 3969
rect 39148 3968 39188 4012
rect 37795 3928 37804 3968
rect 37844 3928 37900 3968
rect 37940 3928 37949 3968
rect 39139 3928 39148 3968
rect 39188 3928 39197 3968
rect 37795 3927 37853 3928
rect 27139 3884 27197 3885
rect 27054 3844 27148 3884
rect 27188 3844 27197 3884
rect 27427 3844 27436 3884
rect 27476 3844 31180 3884
rect 31220 3844 33196 3884
rect 33236 3844 33245 3884
rect 34531 3844 34540 3884
rect 34580 3844 36844 3884
rect 36884 3844 36893 3884
rect 27139 3843 27197 3844
rect 37699 3800 37757 3801
rect 42928 3800 43008 3820
rect 21772 3760 23884 3800
rect 23924 3760 23933 3800
rect 24556 3760 26420 3800
rect 30019 3760 30028 3800
rect 30068 3760 30700 3800
rect 30740 3760 30749 3800
rect 31459 3760 31468 3800
rect 31508 3760 31660 3800
rect 31700 3760 31709 3800
rect 35159 3760 35168 3800
rect 35208 3760 35250 3800
rect 35290 3760 35332 3800
rect 35372 3760 35414 3800
rect 35454 3760 35496 3800
rect 35536 3760 35545 3800
rect 35779 3760 35788 3800
rect 35828 3760 37516 3800
rect 37556 3760 37565 3800
rect 37699 3760 37708 3800
rect 37748 3760 43008 3800
rect 0 3740 80 3760
rect 4780 3716 4820 3760
rect 5356 3716 5396 3760
rect 8803 3759 8861 3760
rect 12364 3716 12404 3760
rect 19180 3716 19220 3760
rect 19948 3716 19988 3760
rect 21667 3759 21725 3760
rect 24556 3716 24596 3760
rect 37699 3759 37757 3760
rect 42928 3740 43008 3760
rect 4780 3676 5396 3716
rect 9859 3676 9868 3716
rect 9908 3676 11596 3716
rect 11636 3676 11645 3716
rect 12364 3676 19180 3716
rect 19220 3676 19229 3716
rect 19948 3676 24596 3716
rect 24739 3716 24797 3717
rect 24739 3676 24748 3716
rect 24788 3676 24882 3716
rect 28195 3676 28204 3716
rect 28244 3676 28588 3716
rect 28628 3676 28637 3716
rect 28960 3676 33100 3716
rect 33140 3676 40684 3716
rect 40724 3676 40733 3716
rect 12364 3632 12404 3676
rect 24739 3675 24797 3676
rect 21187 3632 21245 3633
rect 28960 3632 29000 3676
rect 1411 3592 1420 3632
rect 1460 3592 2764 3632
rect 2804 3592 2813 3632
rect 7171 3592 7180 3632
rect 7220 3592 7948 3632
rect 7988 3592 8716 3632
rect 8756 3592 8765 3632
rect 8899 3592 8908 3632
rect 8948 3592 10636 3632
rect 10676 3592 10685 3632
rect 10732 3592 12404 3632
rect 13027 3592 13036 3632
rect 13076 3592 14188 3632
rect 14228 3592 14237 3632
rect 19075 3592 19084 3632
rect 19124 3592 19852 3632
rect 19892 3592 19901 3632
rect 21187 3592 21196 3632
rect 21236 3592 22540 3632
rect 22580 3592 29000 3632
rect 32611 3592 32620 3632
rect 32660 3592 33676 3632
rect 33716 3592 33725 3632
rect 39043 3592 39052 3632
rect 39092 3592 39916 3632
rect 39956 3592 39965 3632
rect 10732 3548 10772 3592
rect 21187 3591 21245 3592
rect 40771 3548 40829 3549
rect 4387 3508 4396 3548
rect 4436 3508 6028 3548
rect 6068 3508 6077 3548
rect 6412 3508 9388 3548
rect 9428 3508 9437 3548
rect 10243 3508 10252 3548
rect 10292 3508 10772 3548
rect 10915 3508 10924 3548
rect 10964 3508 11360 3548
rect 13795 3508 13804 3548
rect 13844 3508 15148 3548
rect 15188 3508 16012 3548
rect 16052 3508 16061 3548
rect 18691 3508 18700 3548
rect 18740 3508 19276 3548
rect 19316 3508 19660 3548
rect 19700 3508 21100 3548
rect 21140 3508 21149 3548
rect 24163 3508 24172 3548
rect 24212 3508 24940 3548
rect 24980 3508 24989 3548
rect 29923 3508 29932 3548
rect 29972 3508 33524 3548
rect 39523 3508 39532 3548
rect 39572 3508 40108 3548
rect 40148 3508 40780 3548
rect 40820 3508 41452 3548
rect 41492 3508 41501 3548
rect 0 3464 80 3484
rect 1315 3464 1373 3465
rect 2947 3464 3005 3465
rect 6412 3464 6452 3508
rect 11320 3464 11360 3508
rect 12547 3464 12605 3465
rect 16291 3464 16349 3465
rect 18403 3464 18461 3465
rect 33484 3464 33524 3508
rect 40771 3507 40829 3508
rect 41635 3464 41693 3465
rect 42928 3464 43008 3484
rect 0 3424 1172 3464
rect 1230 3424 1324 3464
rect 1364 3424 1373 3464
rect 2659 3424 2668 3464
rect 2708 3424 2956 3464
rect 2996 3424 3005 3464
rect 3619 3424 3628 3464
rect 3668 3424 4492 3464
rect 4532 3424 5548 3464
rect 5588 3424 6452 3464
rect 6595 3424 6604 3464
rect 6644 3424 6653 3464
rect 7555 3424 7564 3464
rect 7604 3424 8044 3464
rect 8084 3424 8093 3464
rect 9091 3424 9100 3464
rect 9140 3424 10828 3464
rect 10868 3424 10877 3464
rect 11320 3424 11500 3464
rect 11540 3424 11549 3464
rect 12067 3424 12076 3464
rect 12116 3424 12125 3464
rect 12462 3424 12556 3464
rect 12596 3424 12605 3464
rect 14755 3424 14764 3464
rect 14804 3424 16300 3464
rect 16340 3424 16349 3464
rect 16963 3424 16972 3464
rect 17012 3424 17548 3464
rect 17588 3424 17597 3464
rect 18211 3424 18220 3464
rect 18260 3424 18412 3464
rect 18452 3424 18461 3464
rect 18883 3424 18892 3464
rect 18932 3424 20044 3464
rect 20084 3424 25516 3464
rect 25556 3424 25565 3464
rect 26563 3424 26572 3464
rect 26612 3424 26764 3464
rect 26804 3424 27436 3464
rect 27476 3424 28396 3464
rect 28436 3424 28972 3464
rect 29012 3424 30316 3464
rect 30356 3424 30604 3464
rect 30644 3424 30653 3464
rect 32227 3424 32236 3464
rect 32276 3424 32908 3464
rect 32948 3424 32957 3464
rect 33475 3424 33484 3464
rect 33524 3424 41356 3464
rect 41396 3424 41405 3464
rect 41635 3424 41644 3464
rect 41684 3424 43008 3464
rect 0 3404 80 3424
rect 1132 3380 1172 3424
rect 1315 3423 1373 3424
rect 2947 3423 3005 3424
rect 6604 3380 6644 3424
rect 12076 3380 12116 3424
rect 12547 3423 12605 3424
rect 16291 3423 16349 3424
rect 18403 3423 18461 3424
rect 25219 3380 25277 3381
rect 32908 3380 32948 3424
rect 41635 3423 41693 3424
rect 42928 3404 43008 3424
rect 1132 3340 1516 3380
rect 1556 3340 1565 3380
rect 4291 3340 4300 3380
rect 4340 3340 5740 3380
rect 5780 3340 5789 3380
rect 6604 3340 7372 3380
rect 7412 3340 11348 3380
rect 11395 3340 11404 3380
rect 11444 3340 12116 3380
rect 14371 3340 14380 3380
rect 14420 3340 25036 3380
rect 25076 3340 25085 3380
rect 25219 3340 25228 3380
rect 25268 3340 25362 3380
rect 26467 3340 26476 3380
rect 26516 3340 28300 3380
rect 28340 3340 28349 3380
rect 29827 3340 29836 3380
rect 29876 3340 30220 3380
rect 30260 3340 30269 3380
rect 32908 3340 33100 3380
rect 33140 3340 35500 3380
rect 35540 3340 35549 3380
rect 37699 3340 37708 3380
rect 37748 3340 38092 3380
rect 38132 3340 38141 3380
rect 9676 3296 9716 3340
rect 11308 3296 11348 3340
rect 25219 3339 25277 3340
rect 16387 3296 16445 3297
rect 24931 3296 24989 3297
rect 26371 3296 26429 3297
rect 4963 3256 4972 3296
rect 5012 3256 5452 3296
rect 5492 3256 6220 3296
rect 6260 3256 6604 3296
rect 6644 3256 6653 3296
rect 9667 3256 9676 3296
rect 9716 3256 9725 3296
rect 11308 3256 15532 3296
rect 15572 3256 15581 3296
rect 16387 3256 16396 3296
rect 16436 3256 22444 3296
rect 22484 3256 22493 3296
rect 24846 3256 24940 3296
rect 24980 3256 24989 3296
rect 25315 3256 25324 3296
rect 25364 3256 26380 3296
rect 26420 3256 26429 3296
rect 31459 3256 31468 3296
rect 31508 3256 31852 3296
rect 31892 3256 40300 3296
rect 40340 3256 40349 3296
rect 41251 3256 41260 3296
rect 41300 3256 41548 3296
rect 41588 3256 41597 3296
rect 16387 3255 16445 3256
rect 24931 3255 24989 3256
rect 26371 3255 26429 3256
rect 6115 3212 6173 3213
rect 9859 3212 9917 3213
rect 24547 3212 24605 3213
rect 2755 3172 2764 3212
rect 2804 3172 4876 3212
rect 4916 3172 4925 3212
rect 5731 3172 5740 3212
rect 5780 3172 6124 3212
rect 6164 3172 6173 3212
rect 6499 3172 6508 3212
rect 6548 3172 6988 3212
rect 7028 3172 9292 3212
rect 9332 3172 9341 3212
rect 9763 3172 9772 3212
rect 9812 3172 9868 3212
rect 9908 3172 9917 3212
rect 10627 3172 10636 3212
rect 10676 3172 14668 3212
rect 14708 3172 14717 3212
rect 19171 3172 19180 3212
rect 19220 3172 19468 3212
rect 19508 3172 19517 3212
rect 20140 3172 21580 3212
rect 21620 3172 23404 3212
rect 23444 3172 23453 3212
rect 24462 3172 24556 3212
rect 24596 3172 24605 3212
rect 6115 3171 6173 3172
rect 9859 3171 9917 3172
rect 0 3128 80 3148
rect 20140 3128 20180 3172
rect 24547 3171 24605 3172
rect 26563 3212 26621 3213
rect 28195 3212 28253 3213
rect 37891 3212 37949 3213
rect 26563 3172 26572 3212
rect 26612 3172 28204 3212
rect 28244 3172 28253 3212
rect 29347 3172 29356 3212
rect 29396 3172 34636 3212
rect 34676 3172 34685 3212
rect 37806 3172 37900 3212
rect 37940 3172 37949 3212
rect 26563 3171 26621 3172
rect 28195 3171 28253 3172
rect 37891 3171 37949 3172
rect 37996 3172 38380 3212
rect 38420 3172 38429 3212
rect 37996 3128 38036 3172
rect 41731 3128 41789 3129
rect 42928 3128 43008 3148
rect 0 3088 1804 3128
rect 1844 3088 2284 3128
rect 2324 3088 2333 3128
rect 2947 3088 2956 3128
rect 2996 3088 8332 3128
rect 8372 3088 8381 3128
rect 8707 3088 8716 3128
rect 8756 3088 9676 3128
rect 9716 3088 9725 3128
rect 9955 3088 9964 3128
rect 10004 3088 11212 3128
rect 11252 3088 11261 3128
rect 14275 3088 14284 3128
rect 14324 3088 20180 3128
rect 21283 3088 21292 3128
rect 21332 3088 25132 3128
rect 25172 3088 37612 3128
rect 37652 3088 38036 3128
rect 38083 3088 38092 3128
rect 38132 3088 40972 3128
rect 41012 3088 41021 3128
rect 41731 3088 41740 3128
rect 41780 3088 43008 3128
rect 0 3068 80 3088
rect 9964 3044 10004 3088
rect 41731 3087 41789 3088
rect 42928 3068 43008 3088
rect 3679 3004 3688 3044
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 4056 3004 4065 3044
rect 5548 3004 10004 3044
rect 10819 3004 10828 3044
rect 10868 3004 18508 3044
rect 18548 3004 18557 3044
rect 18799 3004 18808 3044
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 19176 3004 19185 3044
rect 21091 3004 21100 3044
rect 21140 3004 23692 3044
rect 23732 3004 23741 3044
rect 23875 3004 23884 3044
rect 23924 3004 24076 3044
rect 24116 3004 24940 3044
rect 24980 3004 24989 3044
rect 27043 3004 27052 3044
rect 27092 3004 29932 3044
rect 29972 3004 29981 3044
rect 30211 3004 30220 3044
rect 30260 3004 32236 3044
rect 32276 3004 32285 3044
rect 33919 3004 33928 3044
rect 33968 3004 34010 3044
rect 34050 3004 34092 3044
rect 34132 3004 34174 3044
rect 34214 3004 34256 3044
rect 34296 3004 34305 3044
rect 4195 2960 4253 2961
rect 5548 2960 5588 3004
rect 5923 2960 5981 2961
rect 20899 2960 20957 2961
rect 2851 2920 2860 2960
rect 2900 2920 3148 2960
rect 3188 2920 3197 2960
rect 3820 2920 4204 2960
rect 4244 2920 5068 2960
rect 5108 2920 5117 2960
rect 5539 2920 5548 2960
rect 5588 2920 5597 2960
rect 5923 2920 5932 2960
rect 5972 2920 6028 2960
rect 6068 2920 6077 2960
rect 9283 2920 9292 2960
rect 9332 2920 11360 2960
rect 11875 2920 11884 2960
rect 11924 2920 14764 2960
rect 14804 2920 20908 2960
rect 20948 2920 20957 2960
rect 25507 2920 25516 2960
rect 25556 2920 34388 2960
rect 3820 2876 3860 2920
rect 4195 2919 4253 2920
rect 5923 2919 5981 2920
rect 5827 2876 5885 2877
rect 6595 2876 6653 2877
rect 11320 2876 11360 2920
rect 20899 2919 20957 2920
rect 17155 2876 17213 2877
rect 28195 2876 28253 2877
rect 28963 2876 29021 2877
rect 34348 2876 34388 2920
rect 37780 2920 41356 2960
rect 41396 2920 41405 2960
rect 37780 2876 37820 2920
rect 1987 2836 1996 2876
rect 2036 2836 3860 2876
rect 3907 2836 3916 2876
rect 3956 2836 4300 2876
rect 4340 2836 4349 2876
rect 5827 2836 5836 2876
rect 5876 2836 6604 2876
rect 6644 2836 9484 2876
rect 9524 2836 10636 2876
rect 10676 2836 10685 2876
rect 11320 2836 16684 2876
rect 16724 2836 16733 2876
rect 17070 2836 17164 2876
rect 17204 2836 17213 2876
rect 26083 2836 26092 2876
rect 26132 2836 26668 2876
rect 26708 2836 26717 2876
rect 27715 2836 27724 2876
rect 27764 2836 28012 2876
rect 28052 2836 28061 2876
rect 28195 2836 28204 2876
rect 28244 2836 28916 2876
rect 5827 2835 5885 2836
rect 6595 2835 6653 2836
rect 17155 2835 17213 2836
rect 28195 2835 28253 2836
rect 0 2792 80 2812
rect 5635 2792 5693 2793
rect 0 2752 1324 2792
rect 1364 2752 1373 2792
rect 3811 2752 3820 2792
rect 3860 2752 5644 2792
rect 5684 2752 5693 2792
rect 0 2732 80 2752
rect 5635 2751 5693 2752
rect 6019 2792 6077 2793
rect 7651 2792 7709 2793
rect 11299 2792 11357 2793
rect 28876 2792 28916 2836
rect 28963 2836 28972 2876
rect 29012 2836 31468 2876
rect 31508 2836 31517 2876
rect 34339 2836 34348 2876
rect 34388 2836 37820 2876
rect 28963 2835 29021 2836
rect 42499 2792 42557 2793
rect 42928 2792 43008 2812
rect 6019 2752 6028 2792
rect 6068 2752 7660 2792
rect 7700 2752 10196 2792
rect 10243 2752 10252 2792
rect 10292 2752 10732 2792
rect 10772 2752 10781 2792
rect 11214 2752 11308 2792
rect 11348 2752 11357 2792
rect 13315 2752 13324 2792
rect 13364 2752 19756 2792
rect 19796 2752 19805 2792
rect 24355 2752 24364 2792
rect 24404 2752 24556 2792
rect 24596 2752 28820 2792
rect 28876 2752 29356 2792
rect 29396 2752 29405 2792
rect 34243 2752 34252 2792
rect 34292 2752 35500 2792
rect 35540 2752 36172 2792
rect 36212 2752 36221 2792
rect 40579 2752 40588 2792
rect 40628 2752 41644 2792
rect 41684 2752 41693 2792
rect 42499 2752 42508 2792
rect 42548 2752 43008 2792
rect 6019 2751 6077 2752
rect 7651 2751 7709 2752
rect 10156 2708 10196 2752
rect 11299 2751 11357 2752
rect 25123 2708 25181 2709
rect 28291 2708 28349 2709
rect 28675 2708 28733 2709
rect 4291 2668 4300 2708
rect 4340 2668 6316 2708
rect 6356 2668 9100 2708
rect 9140 2668 9149 2708
rect 10147 2668 10156 2708
rect 10196 2668 10205 2708
rect 10828 2668 14284 2708
rect 14324 2668 14333 2708
rect 16675 2668 16684 2708
rect 16724 2668 21004 2708
rect 21044 2668 21053 2708
rect 23779 2668 23788 2708
rect 23828 2668 24652 2708
rect 24692 2668 24701 2708
rect 25123 2668 25132 2708
rect 25172 2668 27052 2708
rect 27092 2668 27101 2708
rect 28099 2668 28108 2708
rect 28148 2668 28300 2708
rect 28340 2668 28684 2708
rect 28724 2668 28733 2708
rect 10828 2624 10868 2668
rect 25123 2667 25181 2668
rect 28291 2667 28349 2668
rect 28675 2667 28733 2668
rect 26371 2624 26429 2625
rect 28780 2624 28820 2752
rect 42499 2751 42557 2752
rect 42928 2732 43008 2752
rect 28867 2708 28925 2709
rect 36547 2708 36605 2709
rect 28867 2668 28876 2708
rect 28916 2668 33292 2708
rect 33332 2668 33341 2708
rect 33859 2668 33868 2708
rect 33908 2668 34636 2708
rect 34676 2668 36556 2708
rect 36596 2668 36605 2708
rect 28867 2667 28925 2668
rect 36547 2667 36605 2668
rect 28963 2624 29021 2625
rect 2563 2584 2572 2624
rect 2612 2584 2764 2624
rect 2804 2584 2813 2624
rect 3427 2584 3436 2624
rect 3476 2584 4972 2624
rect 5012 2584 5356 2624
rect 5396 2584 5405 2624
rect 5923 2584 5932 2624
rect 5972 2584 7852 2624
rect 7892 2584 7901 2624
rect 9379 2584 9388 2624
rect 9428 2584 10348 2624
rect 10388 2584 10868 2624
rect 11020 2584 11360 2624
rect 2563 2540 2621 2541
rect 3427 2540 3485 2541
rect 11020 2540 11060 2584
rect 1123 2500 1132 2540
rect 1172 2500 2572 2540
rect 2612 2500 2621 2540
rect 3204 2500 3244 2540
rect 3284 2500 3293 2540
rect 3427 2500 3436 2540
rect 3476 2500 4780 2540
rect 4820 2500 5492 2540
rect 7075 2500 7084 2540
rect 7124 2500 7372 2540
rect 7412 2500 7421 2540
rect 7660 2500 7988 2540
rect 10915 2500 10924 2540
rect 10964 2500 11060 2540
rect 11320 2540 11360 2584
rect 11404 2584 12268 2624
rect 12308 2584 12940 2624
rect 12980 2584 12989 2624
rect 16195 2584 16204 2624
rect 16244 2584 16588 2624
rect 16628 2584 16637 2624
rect 20428 2584 21868 2624
rect 21908 2584 21917 2624
rect 22627 2584 22636 2624
rect 22676 2584 23308 2624
rect 23348 2584 23357 2624
rect 26371 2584 26380 2624
rect 26420 2584 28724 2624
rect 28780 2584 28972 2624
rect 29012 2584 29021 2624
rect 11404 2540 11444 2584
rect 16291 2540 16349 2541
rect 20428 2540 20468 2584
rect 26371 2583 26429 2584
rect 28684 2540 28724 2584
rect 28963 2583 29021 2584
rect 29068 2584 29260 2624
rect 29300 2584 29309 2624
rect 29539 2584 29548 2624
rect 29588 2584 29932 2624
rect 29972 2584 31564 2624
rect 31604 2584 34924 2624
rect 34964 2584 38284 2624
rect 38324 2584 38333 2624
rect 41059 2584 41068 2624
rect 41108 2584 41548 2624
rect 41588 2584 41597 2624
rect 29068 2540 29108 2584
rect 36547 2540 36605 2541
rect 11320 2500 11444 2540
rect 16206 2500 16300 2540
rect 16340 2500 16349 2540
rect 20419 2500 20428 2540
rect 20468 2500 20477 2540
rect 28684 2500 29108 2540
rect 36462 2500 36556 2540
rect 36596 2500 36605 2540
rect 2563 2499 2621 2500
rect 0 2456 80 2476
rect 3244 2456 3284 2500
rect 3427 2499 3485 2500
rect 5452 2456 5492 2500
rect 6019 2456 6077 2457
rect 7660 2456 7700 2500
rect 7843 2456 7901 2457
rect 0 2416 2540 2456
rect 3244 2416 5356 2456
rect 5396 2416 5405 2456
rect 5452 2416 6028 2456
rect 6068 2416 6077 2456
rect 0 2396 80 2416
rect 2500 2372 2540 2416
rect 6019 2415 6077 2416
rect 6124 2416 7700 2456
rect 7758 2416 7852 2456
rect 7892 2416 7901 2456
rect 7948 2456 7988 2500
rect 16291 2499 16349 2500
rect 36547 2499 36605 2500
rect 42499 2456 42557 2457
rect 42928 2456 43008 2476
rect 7948 2416 8140 2456
rect 8180 2416 8189 2456
rect 9187 2416 9196 2456
rect 9236 2416 10060 2456
rect 10100 2416 10109 2456
rect 11203 2416 11212 2456
rect 11252 2416 11980 2456
rect 12020 2416 12029 2456
rect 17827 2416 17836 2456
rect 17876 2416 40876 2456
rect 40916 2416 40925 2456
rect 42499 2416 42508 2456
rect 42548 2416 43008 2456
rect 5923 2372 5981 2373
rect 6124 2372 6164 2416
rect 7843 2415 7901 2416
rect 42499 2415 42557 2416
rect 42928 2396 43008 2416
rect 2500 2332 5548 2372
rect 5588 2332 5597 2372
rect 5923 2332 5932 2372
rect 5972 2332 6124 2372
rect 6164 2332 6173 2372
rect 6691 2332 6700 2372
rect 6740 2332 7276 2372
rect 7316 2332 9292 2372
rect 9332 2332 9341 2372
rect 9475 2332 9484 2372
rect 9524 2332 9772 2372
rect 9812 2332 9821 2372
rect 12643 2332 12652 2372
rect 12692 2332 17452 2372
rect 17492 2332 18836 2372
rect 19267 2332 19276 2372
rect 19316 2332 20908 2372
rect 20948 2332 20957 2372
rect 21379 2332 21388 2372
rect 21428 2332 23500 2372
rect 23540 2332 23549 2372
rect 23920 2332 28972 2372
rect 29012 2332 30932 2372
rect 30979 2332 30988 2372
rect 31028 2332 39724 2372
rect 39764 2332 39773 2372
rect 5923 2331 5981 2332
rect 11299 2288 11357 2289
rect 3619 2248 3628 2288
rect 3668 2248 4780 2288
rect 4820 2248 4829 2288
rect 4919 2248 4928 2288
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 5296 2248 5305 2288
rect 5740 2248 7948 2288
rect 7988 2248 7997 2288
rect 11299 2248 11308 2288
rect 11348 2248 15340 2288
rect 15380 2248 15389 2288
rect 5740 2204 5780 2248
rect 11299 2247 11357 2248
rect 18796 2204 18836 2332
rect 23920 2288 23960 2332
rect 20039 2248 20048 2288
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20416 2248 20425 2288
rect 20524 2248 23960 2288
rect 24547 2288 24605 2289
rect 30892 2288 30932 2332
rect 24547 2248 24556 2288
rect 24596 2248 29644 2288
rect 29684 2248 29693 2288
rect 30892 2248 31756 2288
rect 31796 2248 31805 2288
rect 32803 2248 32812 2288
rect 32852 2248 33196 2288
rect 33236 2248 33245 2288
rect 35159 2248 35168 2288
rect 35208 2248 35250 2288
rect 35290 2248 35332 2288
rect 35372 2248 35414 2288
rect 35454 2248 35496 2288
rect 35536 2248 35545 2288
rect 38851 2248 38860 2288
rect 38900 2248 41260 2288
rect 41300 2248 41309 2288
rect 20524 2204 20564 2248
rect 24547 2247 24605 2248
rect 2500 2164 2956 2204
rect 2996 2164 3340 2204
rect 3380 2164 3389 2204
rect 3523 2164 3532 2204
rect 3572 2164 5780 2204
rect 7555 2164 7564 2204
rect 7604 2164 8332 2204
rect 8372 2164 8381 2204
rect 8515 2164 8524 2204
rect 8564 2164 12748 2204
rect 12788 2164 12797 2204
rect 18796 2164 20564 2204
rect 27235 2164 27244 2204
rect 27284 2164 41600 2204
rect 0 2120 80 2140
rect 451 2120 509 2121
rect 2500 2120 2540 2164
rect 6115 2120 6173 2121
rect 41560 2120 41600 2164
rect 42928 2120 43008 2140
rect 0 2080 460 2120
rect 500 2080 509 2120
rect 1699 2080 1708 2120
rect 1748 2080 2540 2120
rect 3235 2080 3244 2120
rect 3284 2080 5452 2120
rect 5492 2080 5501 2120
rect 6019 2080 6028 2120
rect 6068 2080 6124 2120
rect 6164 2080 6173 2120
rect 10915 2080 10924 2120
rect 10964 2080 11596 2120
rect 11636 2080 11645 2120
rect 11779 2080 11788 2120
rect 11828 2080 11837 2120
rect 15811 2080 15820 2120
rect 15860 2080 24748 2120
rect 24788 2080 24797 2120
rect 25132 2080 26284 2120
rect 26324 2080 26333 2120
rect 29155 2080 29164 2120
rect 29204 2080 30124 2120
rect 30164 2080 30173 2120
rect 33379 2080 33388 2120
rect 33428 2080 33676 2120
rect 33716 2080 33725 2120
rect 34435 2080 34444 2120
rect 34484 2080 34828 2120
rect 34868 2080 34877 2120
rect 37987 2080 37996 2120
rect 38036 2080 38764 2120
rect 38804 2080 41260 2120
rect 41300 2080 41309 2120
rect 41560 2080 43008 2120
rect 0 2060 80 2080
rect 451 2079 509 2080
rect 6115 2079 6173 2080
rect 11788 2036 11828 2080
rect 25132 2036 25172 2080
rect 42928 2060 43008 2080
rect 29923 2036 29981 2037
rect 1507 1996 1516 2036
rect 1556 1996 1804 2036
rect 1844 1996 1853 2036
rect 4771 1996 4780 2036
rect 4820 1996 8180 2036
rect 10051 1996 10060 2036
rect 10100 1996 11828 2036
rect 11875 1996 11884 2036
rect 11924 1996 12556 2036
rect 12596 1996 12605 2036
rect 16771 1996 16780 2036
rect 16820 1996 25172 2036
rect 26083 1996 26092 2036
rect 26132 1996 26476 2036
rect 26516 1996 26525 2036
rect 29838 1996 29932 2036
rect 29972 1996 29981 2036
rect 31555 1996 31564 2036
rect 31604 1996 38092 2036
rect 38132 1996 38141 2036
rect 1891 1952 1949 1953
rect 1806 1912 1900 1952
rect 1940 1912 1949 1952
rect 3139 1912 3148 1952
rect 3188 1912 4588 1952
rect 4628 1912 4637 1952
rect 6115 1912 6124 1952
rect 6164 1912 6412 1952
rect 6452 1912 6461 1952
rect 1891 1911 1949 1912
rect 8140 1868 8180 1996
rect 11788 1952 11828 1996
rect 29923 1995 29981 1996
rect 19267 1952 19325 1953
rect 22819 1952 22877 1953
rect 39235 1952 39293 1953
rect 11395 1912 11404 1952
rect 11444 1912 11453 1952
rect 11788 1912 12268 1952
rect 12308 1912 13036 1952
rect 13076 1912 13085 1952
rect 15907 1912 15916 1952
rect 15956 1912 17836 1952
rect 17876 1912 19276 1952
rect 19316 1912 19325 1952
rect 19555 1912 19564 1952
rect 19604 1912 21196 1952
rect 21236 1912 21245 1952
rect 22734 1912 22828 1952
rect 22868 1912 22877 1952
rect 11404 1868 11444 1912
rect 19267 1911 19325 1912
rect 21196 1868 21236 1912
rect 22819 1911 22877 1912
rect 23920 1912 24076 1952
rect 24116 1912 24268 1952
rect 24308 1912 26668 1952
rect 26708 1912 26717 1952
rect 28675 1912 28684 1952
rect 28724 1912 33388 1952
rect 33428 1912 33437 1952
rect 34915 1912 34924 1952
rect 34964 1912 37804 1952
rect 37844 1912 37853 1952
rect 39150 1912 39244 1952
rect 39284 1912 39293 1952
rect 23920 1868 23960 1912
rect 28684 1868 28724 1912
rect 39235 1911 39293 1912
rect 3724 1828 6988 1868
rect 7028 1828 7037 1868
rect 8131 1828 8140 1868
rect 8180 1828 8189 1868
rect 11404 1828 11788 1868
rect 11828 1828 11837 1868
rect 12451 1828 12460 1868
rect 12500 1828 14572 1868
rect 14612 1828 14621 1868
rect 15100 1828 16204 1868
rect 16244 1828 16253 1868
rect 21196 1828 23020 1868
rect 23060 1828 23069 1868
rect 23491 1828 23500 1868
rect 23540 1828 23960 1868
rect 25699 1828 25708 1868
rect 25748 1828 28724 1868
rect 28780 1828 32524 1868
rect 32564 1828 32573 1868
rect 32899 1828 32908 1868
rect 32948 1828 37132 1868
rect 37172 1828 37181 1868
rect 0 1784 80 1804
rect 3724 1784 3764 1828
rect 6211 1784 6269 1785
rect 0 1744 2668 1784
rect 2708 1744 2717 1784
rect 3715 1744 3724 1784
rect 3764 1744 3773 1784
rect 6126 1744 6220 1784
rect 6260 1744 6269 1784
rect 7747 1744 7756 1784
rect 7796 1744 8524 1784
rect 8564 1744 8573 1784
rect 0 1724 80 1744
rect 6211 1743 6269 1744
rect 15100 1700 15140 1828
rect 28780 1784 28820 1828
rect 42928 1784 43008 1804
rect 24739 1744 24748 1784
rect 24788 1744 28820 1784
rect 31363 1744 31372 1784
rect 31412 1744 34004 1784
rect 34051 1744 34060 1784
rect 34100 1744 40588 1784
rect 40628 1744 40637 1784
rect 41155 1744 41164 1784
rect 41204 1744 43008 1784
rect 3619 1660 3628 1700
rect 3668 1660 4012 1700
rect 4052 1660 5740 1700
rect 5780 1660 5789 1700
rect 6307 1660 6316 1700
rect 6356 1660 6604 1700
rect 6644 1660 6796 1700
rect 6836 1660 6845 1700
rect 7651 1660 7660 1700
rect 7700 1660 7709 1700
rect 7756 1660 15140 1700
rect 31747 1660 31756 1700
rect 31796 1660 33772 1700
rect 33812 1660 33821 1700
rect 7660 1616 7700 1660
rect 6019 1576 6028 1616
rect 6068 1576 7700 1616
rect 7756 1532 7796 1660
rect 33964 1616 34004 1744
rect 42928 1724 43008 1744
rect 36547 1660 36556 1700
rect 36596 1660 39532 1700
rect 39572 1660 39581 1700
rect 11320 1576 24460 1616
rect 24500 1576 24509 1616
rect 25891 1576 25900 1616
rect 25940 1576 29548 1616
rect 29588 1576 29597 1616
rect 33964 1576 38668 1616
rect 38708 1576 38717 1616
rect 11320 1532 11360 1576
rect 3679 1492 3688 1532
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 4056 1492 4065 1532
rect 6115 1492 6124 1532
rect 6164 1492 7796 1532
rect 7852 1492 11360 1532
rect 14563 1492 14572 1532
rect 14612 1492 15916 1532
rect 15956 1492 15965 1532
rect 18799 1492 18808 1532
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 19176 1492 19185 1532
rect 19276 1492 24172 1532
rect 24212 1492 24221 1532
rect 25219 1492 25228 1532
rect 25268 1492 29356 1532
rect 29396 1492 31564 1532
rect 31604 1492 31613 1532
rect 33919 1492 33928 1532
rect 33968 1492 34010 1532
rect 34050 1492 34092 1532
rect 34132 1492 34174 1532
rect 34214 1492 34256 1532
rect 34296 1492 34305 1532
rect 0 1448 80 1468
rect 7852 1448 7892 1492
rect 19276 1448 19316 1492
rect 40291 1448 40349 1449
rect 42928 1448 43008 1468
rect 0 1408 1900 1448
rect 1940 1408 1949 1448
rect 5443 1408 5452 1448
rect 5492 1408 7892 1448
rect 8131 1408 8140 1448
rect 8180 1408 12652 1448
rect 12692 1408 12701 1448
rect 15100 1408 19316 1448
rect 23011 1408 23020 1448
rect 23060 1408 36652 1448
rect 36692 1408 36701 1448
rect 40291 1408 40300 1448
rect 40340 1408 43008 1448
rect 0 1388 80 1408
rect 15100 1364 15140 1408
rect 40291 1407 40349 1408
rect 42928 1388 43008 1408
rect 1603 1324 1612 1364
rect 1652 1324 15140 1364
rect 16588 1324 16916 1364
rect 18691 1324 18700 1364
rect 18740 1324 19084 1364
rect 19124 1324 19133 1364
rect 20515 1324 20524 1364
rect 20564 1324 20908 1364
rect 20948 1324 20957 1364
rect 22819 1324 22828 1364
rect 22868 1324 26284 1364
rect 26324 1324 26333 1364
rect 29827 1324 29836 1364
rect 29876 1324 31564 1364
rect 31604 1324 31613 1364
rect 36931 1324 36940 1364
rect 36980 1324 40204 1364
rect 40244 1324 40253 1364
rect 16588 1280 16628 1324
rect 16771 1280 16829 1281
rect 4099 1240 4108 1280
rect 4148 1240 8044 1280
rect 8084 1240 8093 1280
rect 9571 1240 9580 1280
rect 9620 1240 10348 1280
rect 10388 1240 10732 1280
rect 10772 1240 10781 1280
rect 11203 1240 11212 1280
rect 11252 1240 12460 1280
rect 12500 1240 12509 1280
rect 12739 1240 12748 1280
rect 12788 1240 16628 1280
rect 16686 1240 16780 1280
rect 16820 1240 16829 1280
rect 16876 1280 16916 1324
rect 16876 1240 25900 1280
rect 25940 1240 25949 1280
rect 26083 1240 26092 1280
rect 26132 1240 27820 1280
rect 27860 1240 27869 1280
rect 28867 1240 28876 1280
rect 28916 1240 31276 1280
rect 31316 1240 31325 1280
rect 31459 1240 31468 1280
rect 31508 1240 32812 1280
rect 32852 1240 32861 1280
rect 36259 1240 36268 1280
rect 36308 1240 40780 1280
rect 40820 1240 40829 1280
rect 16771 1239 16829 1240
rect 13795 1196 13853 1197
rect 2755 1156 2764 1196
rect 2804 1156 3148 1196
rect 3188 1156 4340 1196
rect 5251 1156 5260 1196
rect 5300 1156 5644 1196
rect 5684 1156 6892 1196
rect 6932 1156 7892 1196
rect 11491 1156 11500 1196
rect 11540 1156 12172 1196
rect 12212 1156 12221 1196
rect 13710 1156 13804 1196
rect 13844 1156 13853 1196
rect 15811 1156 15820 1196
rect 15860 1156 17452 1196
rect 17492 1156 17932 1196
rect 17972 1156 18892 1196
rect 18932 1156 21004 1196
rect 21044 1156 26188 1196
rect 26228 1156 26237 1196
rect 28291 1156 28300 1196
rect 28340 1156 32236 1196
rect 32276 1156 32285 1196
rect 36355 1156 36364 1196
rect 36404 1156 39628 1196
rect 39668 1156 39677 1196
rect 0 1112 80 1132
rect 4099 1112 4157 1113
rect 4300 1112 4340 1156
rect 7852 1112 7892 1156
rect 13795 1155 13853 1156
rect 9763 1112 9821 1113
rect 13987 1112 14045 1113
rect 30979 1112 31037 1113
rect 0 1072 1844 1112
rect 3811 1072 3820 1112
rect 3860 1072 4108 1112
rect 4148 1072 4157 1112
rect 4291 1072 4300 1112
rect 4340 1072 5068 1112
rect 5108 1072 5452 1112
rect 5492 1072 5501 1112
rect 5827 1072 5836 1112
rect 5876 1072 7180 1112
rect 7220 1072 7229 1112
rect 7843 1072 7852 1112
rect 7892 1072 7901 1112
rect 9678 1072 9772 1112
rect 9812 1072 9821 1112
rect 11683 1072 11692 1112
rect 11732 1072 12364 1112
rect 12404 1072 12413 1112
rect 12547 1072 12556 1112
rect 12596 1072 12844 1112
rect 12884 1072 12893 1112
rect 13902 1072 13996 1112
rect 14036 1072 14045 1112
rect 17635 1072 17644 1112
rect 17684 1072 21100 1112
rect 21140 1072 26092 1112
rect 26132 1072 26141 1112
rect 26275 1072 26284 1112
rect 26324 1072 30988 1112
rect 31028 1072 31037 1112
rect 0 1052 80 1072
rect 1804 1028 1844 1072
rect 4099 1071 4157 1072
rect 9763 1071 9821 1072
rect 13987 1071 14045 1072
rect 17644 1028 17684 1072
rect 30979 1071 31037 1072
rect 31555 1112 31613 1113
rect 32131 1112 32189 1113
rect 42928 1112 43008 1132
rect 31555 1072 31564 1112
rect 31604 1072 32140 1112
rect 32180 1072 33388 1112
rect 33428 1072 33437 1112
rect 36451 1072 36460 1112
rect 36500 1072 43008 1112
rect 31555 1071 31613 1072
rect 32131 1071 32189 1072
rect 42928 1052 43008 1072
rect 1804 988 17684 1028
rect 21187 988 21196 1028
rect 21236 988 21388 1028
rect 21428 988 22348 1028
rect 22388 988 22397 1028
rect 25987 988 25996 1028
rect 26036 988 31852 1028
rect 31892 988 31901 1028
rect 33571 988 33580 1028
rect 33620 988 39436 1028
rect 39476 988 39485 1028
rect 40963 944 41021 945
rect 1411 904 1420 944
rect 1460 904 4148 944
rect 7555 904 7564 944
rect 7604 904 12172 944
rect 12212 904 12221 944
rect 15235 904 15244 944
rect 15284 904 19084 944
rect 19124 904 21292 944
rect 21332 904 21341 944
rect 27139 904 27148 944
rect 27188 904 35212 944
rect 35252 904 35261 944
rect 40878 904 40972 944
rect 41012 904 41021 944
rect 0 776 80 796
rect 0 736 2540 776
rect 0 716 80 736
rect 2500 524 2540 736
rect 4108 692 4148 904
rect 40963 903 41021 904
rect 4195 820 4204 860
rect 4244 820 8716 860
rect 8756 820 8765 860
rect 10435 820 10444 860
rect 10484 820 12652 860
rect 12692 820 12701 860
rect 17155 820 17164 860
rect 17204 820 19948 860
rect 19988 820 22444 860
rect 22484 820 24844 860
rect 24884 820 27340 860
rect 27380 820 28108 860
rect 28148 820 29740 860
rect 29780 820 30220 860
rect 30260 820 30269 860
rect 30883 820 30892 860
rect 30932 820 31468 860
rect 31508 820 31517 860
rect 42928 776 43008 796
rect 4919 736 4928 776
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 5296 736 5305 776
rect 5443 736 5452 776
rect 5492 736 9388 776
rect 9428 736 10924 776
rect 10964 736 15820 776
rect 15860 736 15869 776
rect 20039 736 20048 776
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20416 736 20425 776
rect 35159 736 35168 776
rect 35208 736 35250 776
rect 35290 736 35332 776
rect 35372 736 35414 776
rect 35454 736 35496 776
rect 35536 736 35545 776
rect 36739 736 36748 776
rect 36788 736 43008 776
rect 42928 716 43008 736
rect 19459 692 19517 693
rect 27811 692 27869 693
rect 4108 652 8620 692
rect 8660 652 8669 692
rect 19459 652 19468 692
rect 19508 652 27820 692
rect 27860 652 27869 692
rect 19459 651 19517 652
rect 27811 651 27869 652
rect 32515 692 32573 693
rect 32515 652 32524 692
rect 32564 652 39820 692
rect 39860 652 39869 692
rect 32515 651 32573 652
rect 35203 568 35212 608
rect 35252 568 41164 608
rect 41204 568 41213 608
rect 2500 484 19468 524
rect 19508 484 19517 524
rect 0 440 80 460
rect 42928 440 43008 460
rect 0 400 6124 440
rect 6164 400 6173 440
rect 38467 400 38476 440
rect 38516 400 43008 440
rect 0 380 80 400
rect 42928 380 43008 400
rect 2500 232 12268 272
rect 12308 232 12317 272
rect 23683 232 23692 272
rect 23732 232 32620 272
rect 32660 232 32669 272
rect 34051 232 34060 272
rect 34100 232 40012 272
rect 40052 232 40061 272
rect 0 104 80 124
rect 2500 104 2540 232
rect 19939 188 19997 189
rect 6403 148 6412 188
rect 6452 148 19948 188
rect 19988 148 19997 188
rect 24835 148 24844 188
rect 24884 148 33004 188
rect 33044 148 33053 188
rect 19939 147 19997 148
rect 42928 104 43008 124
rect 0 64 2540 104
rect 19939 64 19948 104
rect 19988 64 20236 104
rect 20276 64 20285 104
rect 29443 64 29452 104
rect 29492 64 30028 104
rect 30068 64 30077 104
rect 30595 64 30604 104
rect 30644 64 30796 104
rect 30836 64 30845 104
rect 37891 64 37900 104
rect 37940 64 43008 104
rect 0 44 80 64
rect 42928 44 43008 64
<< via3 >>
rect 14668 10564 14708 10604
rect 15820 10480 15860 10520
rect 15244 10144 15284 10184
rect 28300 10060 28340 10100
rect 21196 9976 21236 10016
rect 21580 9976 21620 10016
rect 17068 9892 17108 9932
rect 26284 9892 26324 9932
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 18508 9808 18548 9848
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 20812 9808 20852 9848
rect 26956 9808 26996 9848
rect 35168 9808 35208 9848
rect 35250 9808 35290 9848
rect 35332 9808 35372 9848
rect 35414 9808 35454 9848
rect 35496 9808 35536 9848
rect 21100 9640 21140 9680
rect 32428 9640 32468 9680
rect 17932 9556 17972 9596
rect 15628 9472 15668 9512
rect 16588 9472 16628 9512
rect 19276 9472 19316 9512
rect 19468 9472 19508 9512
rect 13228 9388 13268 9428
rect 21676 9388 21716 9428
rect 40972 9388 41012 9428
rect 20716 9220 20756 9260
rect 26668 9304 26708 9344
rect 26956 9220 26996 9260
rect 27724 9220 27764 9260
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 16972 9052 17012 9092
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 21580 9052 21620 9092
rect 26476 9052 26516 9092
rect 33928 9052 33968 9092
rect 34010 9052 34050 9092
rect 34092 9052 34132 9092
rect 34174 9052 34214 9092
rect 34256 9052 34296 9092
rect 32524 8968 32564 9008
rect 5932 8800 5972 8840
rect 13516 8800 13556 8840
rect 13708 8800 13748 8840
rect 14284 8800 14324 8840
rect 15052 8800 15092 8840
rect 15532 8800 15572 8840
rect 21292 8800 21332 8840
rect 31948 8800 31988 8840
rect 32620 8800 32660 8840
rect 35308 8800 35348 8840
rect 37900 8800 37940 8840
rect 11020 8716 11060 8756
rect 20908 8716 20948 8756
rect 26668 8716 26708 8756
rect 26440 8632 26480 8672
rect 26572 8632 26612 8672
rect 28396 8632 28436 8672
rect 40780 8632 40820 8672
rect 4204 8548 4244 8588
rect 30124 8548 30164 8588
rect 30316 8548 30356 8588
rect 4588 8464 4628 8504
rect 16396 8464 16436 8504
rect 21484 8464 21524 8504
rect 32236 8464 32276 8504
rect 34348 8464 34388 8504
rect 11404 8380 11444 8420
rect 31660 8380 31700 8420
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 26284 8296 26324 8336
rect 35168 8296 35208 8336
rect 35250 8296 35290 8336
rect 35332 8296 35372 8336
rect 35414 8296 35454 8336
rect 35496 8296 35536 8336
rect 11404 8212 11444 8252
rect 15436 8212 15476 8252
rect 1612 8128 1652 8168
rect 13804 8128 13844 8168
rect 32716 8128 32756 8168
rect 23020 8044 23060 8084
rect 28588 8044 28628 8084
rect 15436 7960 15476 8000
rect 19564 7960 19604 8000
rect 22060 7960 22100 8000
rect 1708 7792 1748 7832
rect 7564 7876 7604 7916
rect 24076 7960 24116 8000
rect 28780 7960 28820 8000
rect 30028 7960 30068 8000
rect 37132 7960 37172 8000
rect 38188 7960 38228 8000
rect 7756 7876 7796 7916
rect 16396 7876 16436 7916
rect 28876 7876 28916 7916
rect 23884 7792 23924 7832
rect 33676 7792 33716 7832
rect 17644 7708 17684 7748
rect 21484 7708 21524 7748
rect 24076 7708 24116 7748
rect 28876 7708 28916 7748
rect 37324 7708 37364 7748
rect 38092 7708 38132 7748
rect 7468 7624 7508 7664
rect 32428 7624 32468 7664
rect 33292 7624 33332 7664
rect 1708 7540 1748 7580
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 4588 7540 4628 7580
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 33928 7540 33968 7580
rect 34010 7540 34050 7580
rect 34092 7540 34132 7580
rect 34174 7540 34214 7580
rect 34256 7540 34296 7580
rect 35308 7540 35348 7580
rect 26572 7456 26612 7496
rect 31948 7456 31988 7496
rect 6892 7372 6932 7412
rect 7564 7372 7604 7412
rect 24748 7288 24788 7328
rect 8812 7204 8852 7244
rect 11212 7204 11252 7244
rect 12844 7204 12884 7244
rect 35788 7204 35828 7244
rect 37804 7204 37844 7244
rect 9484 7120 9524 7160
rect 17164 7120 17204 7160
rect 21004 7120 21044 7160
rect 22636 7120 22676 7160
rect 24748 7120 24788 7160
rect 30220 7120 30260 7160
rect 40780 7120 40820 7160
rect 6604 7036 6644 7076
rect 21100 6952 21140 6992
rect 30124 6952 30164 6992
rect 36172 6952 36212 6992
rect 3340 6868 3380 6908
rect 6412 6868 6452 6908
rect 20812 6868 20852 6908
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 26476 6784 26516 6824
rect 35168 6784 35208 6824
rect 35250 6784 35290 6824
rect 35332 6784 35372 6824
rect 35414 6784 35454 6824
rect 35496 6784 35536 6824
rect 5932 6616 5972 6656
rect 31564 6616 31604 6656
rect 4204 6448 4244 6488
rect 6220 6448 6260 6488
rect 8812 6448 8852 6488
rect 17644 6448 17684 6488
rect 3436 6364 3476 6404
rect 4108 6364 4148 6404
rect 15436 6364 15476 6404
rect 28300 6364 28340 6404
rect 32140 6364 32180 6404
rect 9868 6280 9908 6320
rect 19276 6280 19316 6320
rect 38956 6364 38996 6404
rect 21484 6280 21524 6320
rect 35308 6280 35348 6320
rect 40204 6280 40244 6320
rect 38188 6196 38228 6236
rect 5356 6112 5396 6152
rect 6412 6112 6452 6152
rect 7660 6112 7700 6152
rect 21388 6112 21428 6152
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 33928 6028 33968 6068
rect 34010 6028 34050 6068
rect 34092 6028 34132 6068
rect 34174 6028 34214 6068
rect 34256 6028 34296 6068
rect 24748 5944 24788 5984
rect 3628 5776 3668 5816
rect 19276 5776 19316 5816
rect 15916 5692 15956 5732
rect 19564 5692 19604 5732
rect 21196 5692 21236 5732
rect 26668 5692 26708 5732
rect 3340 5608 3380 5648
rect 24364 5608 24404 5648
rect 30028 5608 30068 5648
rect 35596 5608 35636 5648
rect 3628 5440 3668 5480
rect 17836 5356 17876 5396
rect 18124 5524 18164 5564
rect 37228 5440 37268 5480
rect 23884 5356 23924 5396
rect 26476 5356 26516 5396
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 35168 5272 35208 5312
rect 35250 5272 35290 5312
rect 35332 5272 35372 5312
rect 35414 5272 35454 5312
rect 35496 5272 35536 5312
rect 12460 5188 12500 5228
rect 1324 5104 1364 5144
rect 4108 5104 4148 5144
rect 5356 5020 5396 5060
rect 12556 5020 12596 5060
rect 27724 5020 27764 5060
rect 30892 5020 30932 5060
rect 40300 5020 40340 5060
rect 7180 4936 7220 4976
rect 10636 4936 10676 4976
rect 19372 4936 19412 4976
rect 27148 4936 27188 4976
rect 28012 4936 28052 4976
rect 31276 4936 31316 4976
rect 40780 4936 40820 4976
rect 8812 4852 8852 4892
rect 9484 4852 9524 4892
rect 17836 4852 17876 4892
rect 37900 4852 37940 4892
rect 41260 4852 41300 4892
rect 19948 4768 19988 4808
rect 34924 4768 34964 4808
rect 3436 4684 3476 4724
rect 4204 4684 4244 4724
rect 7180 4684 7220 4724
rect 9868 4684 9908 4724
rect 27628 4684 27668 4724
rect 32908 4684 32948 4724
rect 41548 4684 41588 4724
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 4204 4516 4244 4556
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 33928 4516 33968 4556
rect 34010 4516 34050 4556
rect 34092 4516 34132 4556
rect 34174 4516 34214 4556
rect 34256 4516 34296 4556
rect 22060 4432 22100 4472
rect 21100 4348 21140 4388
rect 21388 4348 21428 4388
rect 27148 4348 27188 4388
rect 7180 4180 7220 4220
rect 12556 4180 12596 4220
rect 21100 4180 21140 4220
rect 21292 4180 21332 4220
rect 33484 4180 33524 4220
rect 1324 4096 1364 4136
rect 38860 4180 38900 4220
rect 9868 4096 9908 4136
rect 13804 4096 13844 4136
rect 7180 4012 7220 4052
rect 7468 4012 7508 4052
rect 20044 4012 20084 4052
rect 7852 3928 7892 3968
rect 20140 3928 20180 3968
rect 20332 3928 20372 3968
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 8812 3760 8852 3800
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 21676 3760 21716 3800
rect 28396 3928 28436 3968
rect 37612 3928 37652 3968
rect 37804 3928 37844 3968
rect 27148 3844 27188 3884
rect 35168 3760 35208 3800
rect 35250 3760 35290 3800
rect 35332 3760 35372 3800
rect 35414 3760 35454 3800
rect 35496 3760 35536 3800
rect 37708 3760 37748 3800
rect 24748 3676 24788 3716
rect 21196 3592 21236 3632
rect 40780 3508 40820 3548
rect 1324 3424 1364 3464
rect 2956 3424 2996 3464
rect 12556 3424 12596 3464
rect 16300 3424 16340 3464
rect 18412 3424 18452 3464
rect 41644 3424 41684 3464
rect 25228 3340 25268 3380
rect 16396 3256 16436 3296
rect 24940 3256 24980 3296
rect 26380 3256 26420 3296
rect 6124 3172 6164 3212
rect 9868 3172 9908 3212
rect 24556 3172 24596 3212
rect 26572 3172 26612 3212
rect 28204 3172 28244 3212
rect 37900 3172 37940 3212
rect 41740 3088 41780 3128
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 33928 3004 33968 3044
rect 34010 3004 34050 3044
rect 34092 3004 34132 3044
rect 34174 3004 34214 3044
rect 34256 3004 34296 3044
rect 4204 2920 4244 2960
rect 5932 2920 5972 2960
rect 20908 2920 20948 2960
rect 5836 2836 5876 2876
rect 6604 2836 6644 2876
rect 17164 2836 17204 2876
rect 28204 2836 28244 2876
rect 5644 2752 5684 2792
rect 28972 2836 29012 2876
rect 6028 2752 6068 2792
rect 7660 2752 7700 2792
rect 11308 2752 11348 2792
rect 42508 2752 42548 2792
rect 25132 2668 25172 2708
rect 28300 2668 28340 2708
rect 28684 2668 28724 2708
rect 28876 2668 28916 2708
rect 36556 2668 36596 2708
rect 2572 2500 2612 2540
rect 3436 2500 3476 2540
rect 26380 2584 26420 2624
rect 28972 2584 29012 2624
rect 16300 2500 16340 2540
rect 36556 2500 36596 2540
rect 6028 2416 6068 2456
rect 7852 2416 7892 2456
rect 42508 2416 42548 2456
rect 5932 2332 5972 2372
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 11308 2248 11348 2288
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 24556 2248 24596 2288
rect 35168 2248 35208 2288
rect 35250 2248 35290 2288
rect 35332 2248 35372 2288
rect 35414 2248 35454 2288
rect 35496 2248 35536 2288
rect 460 2080 500 2120
rect 6124 2080 6164 2120
rect 29932 1996 29972 2036
rect 1900 1912 1940 1952
rect 19276 1912 19316 1952
rect 22828 1912 22868 1952
rect 39244 1912 39284 1952
rect 6220 1744 6260 1784
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 33928 1492 33968 1532
rect 34010 1492 34050 1532
rect 34092 1492 34132 1532
rect 34174 1492 34214 1532
rect 34256 1492 34296 1532
rect 40300 1408 40340 1448
rect 16780 1240 16820 1280
rect 13804 1156 13844 1196
rect 4108 1072 4148 1112
rect 9772 1072 9812 1112
rect 13996 1072 14036 1112
rect 30988 1072 31028 1112
rect 31564 1072 31604 1112
rect 32140 1072 32180 1112
rect 40972 904 41012 944
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 35168 736 35208 776
rect 35250 736 35290 776
rect 35332 736 35372 776
rect 35414 736 35454 776
rect 35496 736 35536 776
rect 19468 652 19508 692
rect 27820 652 27860 692
rect 32524 652 32564 692
rect 19948 148 19988 188
<< metal4 >>
rect 14668 10604 14708 10613
rect 4928 9848 5296 9857
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 4928 9799 5296 9808
rect 8811 9428 8853 9437
rect 8811 9388 8812 9428
rect 8852 9388 8853 9428
rect 8811 9379 8853 9388
rect 13228 9428 13268 9437
rect 1611 9260 1653 9269
rect 1611 9220 1612 9260
rect 1652 9220 1653 9260
rect 1611 9211 1653 9220
rect 1612 8168 1652 9211
rect 3688 9092 4056 9101
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 3688 9043 4056 9052
rect 1707 8924 1749 8933
rect 1707 8884 1708 8924
rect 1748 8884 1749 8924
rect 1707 8875 1749 8884
rect 1612 8119 1652 8128
rect 1708 7832 1748 8875
rect 5932 8840 5972 8849
rect 1708 7580 1748 7792
rect 4204 8588 4244 8597
rect 1708 7531 1748 7540
rect 3688 7580 4056 7589
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 3688 7531 4056 7540
rect 3340 6908 3380 6917
rect 3340 5657 3380 6868
rect 4204 6488 4244 8548
rect 4588 8504 4628 8513
rect 4588 8009 4628 8464
rect 4928 8336 5296 8345
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 4928 8287 5296 8296
rect 4587 8000 4629 8009
rect 4587 7960 4588 8000
rect 4628 7960 4629 8000
rect 4587 7951 4629 7960
rect 4588 7580 4628 7951
rect 4588 7531 4628 7540
rect 4928 6824 5296 6833
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 4928 6775 5296 6784
rect 5932 6656 5972 8800
rect 7564 7916 7604 7925
rect 7468 7664 7508 7673
rect 6892 7412 6932 7421
rect 6892 7169 6932 7372
rect 6891 7160 6933 7169
rect 6891 7120 6892 7160
rect 6932 7120 6933 7160
rect 6891 7111 6933 7120
rect 6604 7076 6644 7085
rect 5932 6607 5972 6616
rect 6412 6908 6452 6917
rect 3436 6404 3476 6413
rect 3339 5648 3381 5657
rect 3339 5608 3340 5648
rect 3380 5608 3381 5648
rect 3339 5599 3381 5608
rect 3340 5514 3380 5599
rect 1324 5144 1364 5153
rect 1324 4145 1364 5104
rect 3436 4724 3476 6364
rect 4108 6404 4148 6413
rect 3688 6068 4056 6077
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 3688 6019 4056 6028
rect 3628 5816 3668 5825
rect 3628 5480 3668 5776
rect 3628 5431 3668 5440
rect 4108 5144 4148 6364
rect 4108 5095 4148 5104
rect 1323 4136 1365 4145
rect 1323 4096 1324 4136
rect 1364 4096 1365 4136
rect 1323 4087 1365 4096
rect 1324 4002 1364 4087
rect 1323 3548 1365 3557
rect 1323 3508 1324 3548
rect 1364 3508 1365 3548
rect 1323 3499 1365 3508
rect 1324 3464 1364 3499
rect 1324 3413 1364 3424
rect 2956 3464 2996 3475
rect 2956 3389 2996 3424
rect 2955 3380 2997 3389
rect 2955 3340 2956 3380
rect 2996 3340 2997 3380
rect 2955 3331 2997 3340
rect 2572 2540 2612 2549
rect 460 2120 500 2129
rect 460 1877 500 2080
rect 1899 1952 1941 1961
rect 1899 1912 1900 1952
rect 1940 1912 1941 1952
rect 1899 1903 1941 1912
rect 459 1868 501 1877
rect 459 1828 460 1868
rect 500 1828 501 1868
rect 459 1819 501 1828
rect 1900 1818 1940 1903
rect 2572 1121 2612 2500
rect 3436 2540 3476 4684
rect 4204 4724 4244 6448
rect 6220 6488 6260 6497
rect 5356 6152 5396 6161
rect 4928 5312 5296 5321
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 4928 5263 5296 5272
rect 5356 5060 5396 6112
rect 6220 5657 6260 6448
rect 6412 6152 6452 6868
rect 6412 6103 6452 6112
rect 6219 5648 6261 5657
rect 6219 5608 6220 5648
rect 6260 5608 6261 5648
rect 6219 5599 6261 5608
rect 5356 4985 5396 5020
rect 5355 4976 5397 4985
rect 5355 4936 5356 4976
rect 5396 4936 5397 4976
rect 5355 4927 5397 4936
rect 5356 4896 5396 4927
rect 3688 4556 4056 4565
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 3688 4507 4056 4516
rect 4204 4556 4244 4684
rect 3688 3044 4056 3053
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 3688 2995 4056 3004
rect 4204 2960 4244 4516
rect 4928 3800 5296 3809
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 4928 3751 5296 3760
rect 6124 3212 6164 3221
rect 4204 2911 4244 2920
rect 5932 2960 5972 2969
rect 5836 2876 5876 2885
rect 5644 2836 5836 2876
rect 5644 2792 5684 2836
rect 5836 2827 5876 2836
rect 5644 2743 5684 2752
rect 3436 2491 3476 2500
rect 5932 2372 5972 2920
rect 6028 2792 6068 2801
rect 6028 2456 6068 2752
rect 6028 2407 6068 2416
rect 5932 2323 5972 2332
rect 4928 2288 5296 2297
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 4928 2239 5296 2248
rect 6124 2120 6164 3172
rect 6124 2071 6164 2080
rect 4107 1868 4149 1877
rect 4107 1828 4108 1868
rect 4148 1828 4149 1868
rect 4107 1819 4149 1828
rect 3688 1532 4056 1541
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 3688 1483 4056 1492
rect 2571 1112 2613 1121
rect 2571 1072 2572 1112
rect 2612 1072 2613 1112
rect 2571 1063 2613 1072
rect 4108 1112 4148 1819
rect 6220 1784 6260 5599
rect 6604 2876 6644 7036
rect 7180 4976 7220 4985
rect 7180 4724 7220 4936
rect 7180 4220 7220 4684
rect 7180 4052 7220 4180
rect 7180 4003 7220 4012
rect 7468 4052 7508 7624
rect 7564 7412 7604 7876
rect 7564 7363 7604 7372
rect 7756 7916 7796 7925
rect 7468 4003 7508 4012
rect 7660 6152 7700 6161
rect 7756 6152 7796 7876
rect 8812 7244 8852 9379
rect 8812 6488 8852 7204
rect 11020 8756 11060 8765
rect 8812 6439 8852 6448
rect 9484 7160 9524 7169
rect 7700 6112 7796 6152
rect 6604 2827 6644 2836
rect 7660 2792 7700 6112
rect 8812 4892 8852 4901
rect 7660 2743 7700 2752
rect 7852 3968 7892 3977
rect 7852 2456 7892 3928
rect 8812 3800 8852 4852
rect 9484 4892 9524 7120
rect 9484 4843 9524 4852
rect 9868 6320 9908 6329
rect 8812 3751 8852 3760
rect 9868 4724 9908 6280
rect 11020 5909 11060 8716
rect 11404 8420 11444 8429
rect 11404 8252 11444 8380
rect 11404 8203 11444 8212
rect 11212 7244 11252 7253
rect 11019 5900 11061 5909
rect 11019 5860 11020 5900
rect 11060 5860 11061 5900
rect 11019 5851 11061 5860
rect 10635 4976 10677 4985
rect 10635 4936 10636 4976
rect 10676 4936 10677 4976
rect 10635 4927 10677 4936
rect 10636 4733 10676 4927
rect 9868 4136 9908 4684
rect 10635 4724 10677 4733
rect 10635 4684 10636 4724
rect 10676 4684 10677 4724
rect 10635 4675 10677 4684
rect 9868 3212 9908 4096
rect 9868 3163 9908 3172
rect 7852 2407 7892 2416
rect 6220 1735 6260 1744
rect 4108 1063 4148 1072
rect 9771 1112 9813 1121
rect 9771 1072 9772 1112
rect 9812 1072 9813 1112
rect 9771 1063 9813 1072
rect 9772 978 9812 1063
rect 11212 953 11252 7204
rect 12843 7244 12885 7253
rect 12843 7204 12844 7244
rect 12884 7204 12885 7244
rect 12843 7195 12885 7204
rect 12844 7110 12884 7195
rect 12460 5228 12500 5237
rect 12460 3548 12500 5188
rect 12556 5060 12596 5069
rect 12556 4220 12596 5020
rect 12556 3809 12596 4180
rect 12555 3800 12597 3809
rect 12555 3760 12556 3800
rect 12596 3760 12597 3800
rect 12555 3751 12597 3760
rect 12555 3548 12597 3557
rect 12460 3508 12556 3548
rect 12596 3508 12597 3548
rect 12555 3499 12597 3508
rect 12556 3464 12596 3499
rect 12556 3413 12596 3424
rect 11308 2792 11348 2801
rect 11308 2288 11348 2752
rect 11308 2239 11348 2248
rect 11211 944 11253 953
rect 11211 904 11212 944
rect 11252 904 11253 944
rect 11211 895 11253 904
rect 4928 776 5296 785
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 4928 727 5296 736
rect 13228 617 13268 9388
rect 13516 8840 13556 8849
rect 13516 869 13556 8800
rect 13708 8840 13748 8849
rect 13708 1037 13748 8800
rect 14284 8840 14324 8849
rect 13804 8168 13844 8179
rect 13804 8093 13844 8128
rect 13803 8084 13845 8093
rect 13803 8044 13804 8084
rect 13844 8044 13845 8084
rect 13803 8035 13845 8044
rect 14284 5489 14324 8800
rect 14668 5741 14708 10564
rect 15820 10520 15860 10529
rect 15244 10184 15284 10193
rect 15052 8840 15092 8849
rect 15052 5825 15092 8800
rect 15244 7001 15284 10144
rect 15628 9512 15668 9521
rect 15435 9260 15477 9269
rect 15435 9220 15436 9260
rect 15476 9220 15477 9260
rect 15435 9211 15477 9220
rect 15436 8252 15476 9211
rect 15436 8000 15476 8212
rect 15436 7951 15476 7960
rect 15532 8840 15572 8849
rect 15243 6992 15285 7001
rect 15243 6952 15244 6992
rect 15284 6952 15285 6992
rect 15243 6943 15285 6952
rect 15436 6404 15476 6413
rect 15051 5816 15093 5825
rect 15051 5776 15052 5816
rect 15092 5776 15093 5816
rect 15051 5767 15093 5776
rect 14667 5732 14709 5741
rect 14667 5692 14668 5732
rect 14708 5692 14709 5732
rect 14667 5683 14709 5692
rect 14283 5480 14325 5489
rect 14283 5440 14284 5480
rect 14324 5440 14325 5480
rect 14283 5431 14325 5440
rect 15436 5069 15476 6364
rect 15435 5060 15477 5069
rect 15435 5020 15436 5060
rect 15476 5020 15477 5060
rect 15435 5011 15477 5020
rect 13804 4136 13844 4145
rect 13804 1793 13844 4096
rect 15532 2129 15572 8800
rect 15531 2120 15573 2129
rect 15531 2080 15532 2120
rect 15572 2080 15573 2120
rect 15531 2071 15573 2080
rect 15628 2045 15668 9472
rect 15820 7841 15860 10480
rect 28300 10100 28340 10109
rect 21196 10016 21236 10025
rect 17068 9932 17108 9941
rect 16588 9512 16628 9521
rect 16395 8504 16437 8513
rect 16395 8464 16396 8504
rect 16436 8464 16437 8504
rect 16395 8455 16437 8464
rect 16396 8370 16436 8455
rect 16396 7916 16436 7925
rect 15819 7832 15861 7841
rect 15819 7792 15820 7832
rect 15860 7792 15861 7832
rect 15819 7783 15861 7792
rect 15916 5732 15956 5741
rect 15916 3473 15956 5692
rect 16299 3548 16341 3557
rect 16299 3508 16300 3548
rect 16340 3508 16341 3548
rect 16299 3499 16341 3508
rect 15915 3464 15957 3473
rect 15915 3424 15916 3464
rect 15956 3424 15957 3464
rect 15915 3415 15957 3424
rect 16300 3464 16340 3499
rect 16300 2540 16340 3424
rect 16396 3296 16436 7876
rect 16588 4313 16628 9472
rect 16972 9092 17012 9101
rect 16972 7421 17012 9052
rect 16971 7412 17013 7421
rect 16971 7372 16972 7412
rect 17012 7372 17013 7412
rect 16971 7363 17013 7372
rect 16779 6404 16821 6413
rect 16779 6364 16780 6404
rect 16820 6364 16821 6404
rect 16779 6355 16821 6364
rect 16587 4304 16629 4313
rect 16587 4264 16588 4304
rect 16628 4264 16629 4304
rect 16587 4255 16629 4264
rect 16396 3247 16436 3256
rect 16300 2491 16340 2500
rect 15627 2036 15669 2045
rect 15627 1996 15628 2036
rect 15668 1996 15669 2036
rect 15627 1987 15669 1996
rect 13803 1784 13845 1793
rect 13803 1744 13804 1784
rect 13844 1744 13845 1784
rect 13803 1735 13845 1744
rect 16780 1280 16820 6355
rect 17068 3221 17108 9892
rect 18508 9848 18548 9857
rect 17932 9596 17972 9605
rect 17643 7748 17685 7757
rect 17643 7708 17644 7748
rect 17684 7708 17685 7748
rect 17643 7699 17685 7708
rect 17644 7614 17684 7699
rect 17164 7160 17204 7169
rect 17067 3212 17109 3221
rect 17067 3172 17068 3212
rect 17108 3172 17109 3212
rect 17067 3163 17109 3172
rect 17164 2876 17204 7120
rect 17643 7076 17685 7085
rect 17643 7036 17644 7076
rect 17684 7036 17685 7076
rect 17643 7027 17685 7036
rect 17644 6488 17684 7027
rect 17644 6439 17684 6448
rect 17932 6245 17972 9556
rect 17931 6236 17973 6245
rect 17931 6196 17932 6236
rect 17972 6196 17973 6236
rect 17931 6187 17973 6196
rect 18124 5564 18164 5573
rect 17836 5396 17876 5405
rect 17836 4892 17876 5356
rect 18124 4901 18164 5524
rect 17836 4843 17876 4852
rect 18123 4892 18165 4901
rect 18123 4852 18124 4892
rect 18164 4852 18165 4892
rect 18123 4843 18165 4852
rect 18508 3641 18548 9808
rect 20048 9848 20416 9857
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20048 9799 20416 9808
rect 20812 9848 20852 9857
rect 19276 9512 19316 9521
rect 18808 9092 19176 9101
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 18808 9043 19176 9052
rect 18808 7580 19176 7589
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 18808 7531 19176 7540
rect 19276 6320 19316 9472
rect 19468 9512 19508 9521
rect 19468 8177 19508 9472
rect 20716 9260 20756 9269
rect 20048 8336 20416 8345
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20048 8287 20416 8296
rect 19467 8168 19509 8177
rect 19467 8128 19468 8168
rect 19508 8128 19509 8168
rect 19467 8119 19509 8128
rect 19563 8000 19605 8009
rect 19563 7960 19564 8000
rect 19604 7960 19605 8000
rect 19563 7951 19605 7960
rect 19276 6271 19316 6280
rect 18808 6068 19176 6077
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 18808 6019 19176 6028
rect 19276 5816 19316 5825
rect 18808 4556 19176 4565
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 18808 4507 19176 4516
rect 18507 3632 18549 3641
rect 18507 3592 18508 3632
rect 18548 3592 18549 3632
rect 18507 3583 18549 3592
rect 18411 3548 18453 3557
rect 18411 3508 18412 3548
rect 18452 3508 18453 3548
rect 18411 3499 18453 3508
rect 18412 3464 18452 3499
rect 18412 3413 18452 3424
rect 18808 3044 19176 3053
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 18808 2995 19176 3004
rect 17164 2827 17204 2836
rect 19276 1952 19316 5776
rect 19564 5732 19604 7951
rect 20716 7757 20756 9220
rect 20715 7748 20757 7757
rect 20715 7708 20716 7748
rect 20756 7708 20757 7748
rect 20715 7699 20757 7708
rect 20812 6908 20852 9808
rect 21100 9680 21140 9689
rect 21003 9008 21045 9017
rect 21003 8968 21004 9008
rect 21044 8968 21045 9008
rect 21003 8959 21045 8968
rect 20812 6859 20852 6868
rect 20908 8756 20948 8765
rect 20048 6824 20416 6833
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20048 6775 20416 6784
rect 19564 5683 19604 5692
rect 20048 5312 20416 5321
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20048 5263 20416 5272
rect 19276 1903 19316 1912
rect 19372 4976 19412 4985
rect 18808 1532 19176 1541
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 18808 1483 19176 1492
rect 16780 1231 16820 1240
rect 13803 1196 13845 1205
rect 13803 1156 13804 1196
rect 13844 1156 13845 1196
rect 13803 1147 13845 1156
rect 13804 1062 13844 1147
rect 19372 1121 19412 4936
rect 19467 4976 19509 4985
rect 19467 4936 19468 4976
rect 19508 4936 19509 4976
rect 19467 4927 19509 4936
rect 19468 3809 19508 4927
rect 19948 4808 19988 4817
rect 19467 3800 19509 3809
rect 19467 3760 19468 3800
rect 19508 3760 19509 3800
rect 19467 3751 19509 3760
rect 13995 1112 14037 1121
rect 13995 1072 13996 1112
rect 14036 1072 14037 1112
rect 13995 1063 14037 1072
rect 19371 1112 19413 1121
rect 19371 1072 19372 1112
rect 19412 1072 19413 1112
rect 19371 1063 19413 1072
rect 13707 1028 13749 1037
rect 13707 988 13708 1028
rect 13748 988 13749 1028
rect 13707 979 13749 988
rect 13996 978 14036 1063
rect 13515 860 13557 869
rect 13515 820 13516 860
rect 13556 820 13557 860
rect 13515 811 13557 820
rect 13227 608 13269 617
rect 13227 568 13228 608
rect 13268 568 13269 608
rect 13227 559 13269 568
rect 19372 533 19412 1063
rect 19467 860 19509 869
rect 19467 820 19468 860
rect 19508 820 19509 860
rect 19467 811 19509 820
rect 19468 692 19508 811
rect 19468 643 19508 652
rect 19371 524 19413 533
rect 19371 484 19372 524
rect 19412 484 19413 524
rect 19371 475 19413 484
rect 19948 188 19988 4768
rect 20043 4472 20085 4481
rect 20043 4432 20044 4472
rect 20084 4432 20085 4472
rect 20043 4423 20085 4432
rect 20044 4052 20084 4423
rect 20044 4003 20084 4012
rect 20140 3968 20180 3977
rect 20332 3968 20372 3977
rect 20180 3928 20332 3968
rect 20140 3919 20180 3928
rect 20332 3919 20372 3928
rect 20048 3800 20416 3809
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20048 3751 20416 3760
rect 20908 2960 20948 8716
rect 21004 7160 21044 8959
rect 21004 7111 21044 7120
rect 21100 6992 21140 9640
rect 21100 6943 21140 6952
rect 21196 5732 21236 9976
rect 21580 10016 21620 10025
rect 21580 9092 21620 9976
rect 26284 9932 26324 9941
rect 21580 9043 21620 9052
rect 21676 9428 21716 9437
rect 21196 5683 21236 5692
rect 21292 8840 21332 8849
rect 21195 4724 21237 4733
rect 21195 4684 21196 4724
rect 21236 4684 21237 4724
rect 21195 4675 21237 4684
rect 21100 4388 21140 4397
rect 21100 4220 21140 4348
rect 21100 4171 21140 4180
rect 21196 3632 21236 4675
rect 21292 4220 21332 8800
rect 21483 8504 21525 8513
rect 21483 8464 21484 8504
rect 21524 8464 21525 8504
rect 21483 8455 21525 8464
rect 21484 8370 21524 8455
rect 21484 7748 21524 7757
rect 21387 7664 21429 7673
rect 21484 7664 21524 7708
rect 21387 7624 21388 7664
rect 21428 7624 21524 7664
rect 21387 7615 21429 7624
rect 21483 6404 21525 6413
rect 21483 6364 21484 6404
rect 21524 6364 21525 6404
rect 21483 6355 21525 6364
rect 21484 6320 21524 6355
rect 21484 6269 21524 6280
rect 21388 6152 21428 6161
rect 21388 4817 21428 6112
rect 21387 4808 21429 4817
rect 21387 4768 21388 4808
rect 21428 4768 21429 4808
rect 21387 4759 21429 4768
rect 21292 4171 21332 4180
rect 21388 4388 21428 4397
rect 21388 4145 21428 4348
rect 21387 4136 21429 4145
rect 21387 4096 21388 4136
rect 21428 4096 21429 4136
rect 21387 4087 21429 4096
rect 21676 3800 21716 9388
rect 24747 9428 24789 9437
rect 24747 9388 24748 9428
rect 24788 9388 24789 9428
rect 24747 9379 24789 9388
rect 24075 8840 24117 8849
rect 24075 8800 24076 8840
rect 24116 8800 24117 8840
rect 24075 8791 24117 8800
rect 23019 8084 23061 8093
rect 23019 8044 23020 8084
rect 23060 8044 23061 8084
rect 23019 8035 23061 8044
rect 22060 8000 22100 8009
rect 22060 4481 22100 7960
rect 23020 7950 23060 8035
rect 24076 8009 24116 8791
rect 24075 8000 24117 8009
rect 24075 7960 24076 8000
rect 24116 7960 24117 8000
rect 24075 7951 24117 7960
rect 24076 7866 24116 7951
rect 23884 7832 23924 7841
rect 23884 7748 23924 7792
rect 24076 7748 24116 7757
rect 23884 7708 24076 7748
rect 24076 7699 24116 7708
rect 24748 7328 24788 9379
rect 26284 8336 26324 9892
rect 26956 9848 26996 9857
rect 26668 9344 26708 9353
rect 26475 9092 26517 9101
rect 26475 9052 26476 9092
rect 26516 9052 26517 9092
rect 26475 9043 26517 9052
rect 26476 8958 26516 9043
rect 26668 8756 26708 9304
rect 26956 9260 26996 9808
rect 26956 9211 26996 9220
rect 27723 9260 27765 9269
rect 27723 9220 27724 9260
rect 27764 9220 27765 9260
rect 27723 9211 27765 9220
rect 27724 9126 27764 9211
rect 26440 8672 26480 8681
rect 26572 8672 26612 8681
rect 26480 8632 26572 8672
rect 26440 8623 26480 8632
rect 26572 8623 26612 8632
rect 26284 8287 26324 8296
rect 25515 8084 25557 8093
rect 25515 8044 25516 8084
rect 25556 8044 25557 8084
rect 25515 8035 25557 8044
rect 22635 7160 22677 7169
rect 22635 7120 22636 7160
rect 22676 7120 22677 7160
rect 22635 7111 22677 7120
rect 24748 7160 24788 7288
rect 24748 7111 24788 7120
rect 22636 7026 22676 7111
rect 24748 5984 24788 5993
rect 24363 5648 24405 5657
rect 24363 5608 24364 5648
rect 24404 5608 24405 5648
rect 24363 5599 24405 5608
rect 24364 5514 24404 5599
rect 23884 5396 23924 5405
rect 23884 5069 23924 5356
rect 23883 5060 23925 5069
rect 23883 5020 23884 5060
rect 23924 5020 23925 5060
rect 23883 5011 23925 5020
rect 22059 4472 22101 4481
rect 22059 4432 22060 4472
rect 22100 4432 22101 4472
rect 22059 4423 22101 4432
rect 22060 4338 22100 4423
rect 22635 3968 22677 3977
rect 22635 3928 22636 3968
rect 22676 3928 22677 3968
rect 22635 3919 22677 3928
rect 21676 3751 21716 3760
rect 21196 3583 21236 3592
rect 22636 3473 22676 3919
rect 24748 3716 24788 5944
rect 24748 3667 24788 3676
rect 22635 3464 22677 3473
rect 22635 3424 22636 3464
rect 22676 3424 22677 3464
rect 22635 3415 22677 3424
rect 25227 3380 25269 3389
rect 25227 3340 25228 3380
rect 25268 3340 25269 3380
rect 25227 3331 25269 3340
rect 24939 3296 24981 3305
rect 24939 3256 24940 3296
rect 24980 3256 24981 3296
rect 24939 3247 24981 3256
rect 20908 2911 20948 2920
rect 24556 3212 24596 3221
rect 24556 2465 24596 3172
rect 24940 3162 24980 3247
rect 25228 3246 25268 3331
rect 25132 2708 25172 2717
rect 24555 2456 24597 2465
rect 24555 2416 24556 2456
rect 24596 2416 24597 2456
rect 24555 2407 24597 2416
rect 20048 2288 20416 2297
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20048 2239 20416 2248
rect 24556 2288 24596 2297
rect 22827 1952 22869 1961
rect 22827 1912 22828 1952
rect 22868 1912 22869 1952
rect 22827 1903 22869 1912
rect 22828 1818 22868 1903
rect 24556 953 24596 2248
rect 25132 1877 25172 2668
rect 25131 1868 25173 1877
rect 25131 1828 25132 1868
rect 25172 1828 25173 1868
rect 25131 1819 25173 1828
rect 24555 944 24597 953
rect 24555 904 24556 944
rect 24596 904 24597 944
rect 24555 895 24597 904
rect 20048 776 20416 785
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20048 727 20416 736
rect 25516 617 25556 8035
rect 26572 7496 26612 7505
rect 26476 6824 26516 6833
rect 26476 5909 26516 6784
rect 26475 5900 26517 5909
rect 26475 5860 26476 5900
rect 26516 5860 26517 5900
rect 26475 5851 26517 5860
rect 26476 5396 26516 5405
rect 26476 3641 26516 5356
rect 26475 3632 26517 3641
rect 26475 3592 26476 3632
rect 26516 3592 26517 3632
rect 26475 3583 26517 3592
rect 26475 3380 26517 3389
rect 26380 3340 26476 3380
rect 26516 3340 26517 3380
rect 26380 3296 26420 3340
rect 26475 3331 26517 3340
rect 26380 3247 26420 3256
rect 26572 3212 26612 7456
rect 26668 5732 26708 8716
rect 27723 8588 27765 8597
rect 27723 8548 27724 8588
rect 27764 8548 27765 8588
rect 27723 8539 27765 8548
rect 26668 5683 26708 5692
rect 27724 5060 27764 8539
rect 28011 7076 28053 7085
rect 28011 7036 28012 7076
rect 28052 7036 28053 7076
rect 28011 7027 28053 7036
rect 28012 6329 28052 7027
rect 28300 6404 28340 10060
rect 35168 9848 35536 9857
rect 35208 9808 35250 9848
rect 35290 9808 35332 9848
rect 35372 9808 35414 9848
rect 35454 9808 35496 9848
rect 35168 9799 35536 9808
rect 32428 9680 32468 9689
rect 31659 9092 31701 9101
rect 31659 9052 31660 9092
rect 31700 9052 31701 9092
rect 31659 9043 31701 9052
rect 28396 8672 28436 8681
rect 28396 7085 28436 8632
rect 30124 8588 30164 8597
rect 28587 8084 28629 8093
rect 28587 8044 28588 8084
rect 28628 8044 28629 8084
rect 28587 8035 28629 8044
rect 28588 7950 28628 8035
rect 28779 8000 28821 8009
rect 28779 7960 28780 8000
rect 28820 7960 28821 8000
rect 28779 7951 28821 7960
rect 30028 8000 30068 8009
rect 28780 7866 28820 7951
rect 28876 7916 28916 7925
rect 28876 7748 28916 7876
rect 28876 7699 28916 7708
rect 28395 7076 28437 7085
rect 28395 7036 28396 7076
rect 28436 7036 28437 7076
rect 28395 7027 28437 7036
rect 28011 6320 28053 6329
rect 28011 6280 28012 6320
rect 28052 6280 28053 6320
rect 28011 6271 28053 6280
rect 27724 5011 27764 5020
rect 27147 4976 27189 4985
rect 27147 4936 27148 4976
rect 27188 4936 27189 4976
rect 27147 4927 27189 4936
rect 28012 4976 28052 4985
rect 27148 4842 27188 4927
rect 27628 4724 27668 4733
rect 27147 4388 27189 4397
rect 27147 4348 27148 4388
rect 27188 4348 27189 4388
rect 27147 4339 27189 4348
rect 27148 3884 27188 4339
rect 27148 3835 27188 3844
rect 26572 3163 26612 3172
rect 27628 2801 27668 4684
rect 27627 2792 27669 2801
rect 27627 2752 27628 2792
rect 27668 2752 27669 2792
rect 27627 2743 27669 2752
rect 26380 2624 26420 2633
rect 26380 1793 26420 2584
rect 28012 1961 28052 4936
rect 28204 3212 28244 3221
rect 28204 2876 28244 3172
rect 28204 2827 28244 2836
rect 28300 2708 28340 6364
rect 30028 5648 30068 7960
rect 30124 6992 30164 8548
rect 30315 8588 30357 8597
rect 30315 8548 30316 8588
rect 30356 8548 30357 8588
rect 30315 8539 30357 8548
rect 30316 8454 30356 8539
rect 31660 8420 31700 9043
rect 31660 8371 31700 8380
rect 31948 8840 31988 8849
rect 31948 8093 31988 8800
rect 32236 8504 32276 8513
rect 31947 8084 31989 8093
rect 31947 8044 31948 8084
rect 31988 8044 31989 8084
rect 31947 8035 31989 8044
rect 31948 7496 31988 8035
rect 31948 7447 31988 7456
rect 31563 7244 31605 7253
rect 31563 7204 31564 7244
rect 31604 7204 31605 7244
rect 31563 7195 31605 7204
rect 30219 7160 30261 7169
rect 30219 7120 30220 7160
rect 30260 7120 30261 7160
rect 30219 7111 30261 7120
rect 30220 7026 30260 7111
rect 30124 6943 30164 6952
rect 31564 6656 31604 7195
rect 31564 6607 31604 6616
rect 32140 6404 32180 6413
rect 31467 5732 31509 5741
rect 31467 5692 31468 5732
rect 31508 5692 31509 5732
rect 31467 5683 31509 5692
rect 30028 5599 30068 5608
rect 30892 5060 30932 5069
rect 30892 4817 30932 5020
rect 31275 5060 31317 5069
rect 31275 5020 31276 5060
rect 31316 5020 31317 5060
rect 31275 5011 31317 5020
rect 31276 4976 31316 5011
rect 31276 4925 31316 4936
rect 31468 4817 31508 5683
rect 30891 4808 30933 4817
rect 30891 4768 30892 4808
rect 30932 4768 30933 4808
rect 30891 4759 30933 4768
rect 31467 4808 31509 4817
rect 31467 4768 31468 4808
rect 31508 4768 31509 4808
rect 31467 4759 31509 4768
rect 28395 3968 28437 3977
rect 28395 3928 28396 3968
rect 28436 3928 28437 3968
rect 28395 3919 28437 3928
rect 28396 3834 28436 3919
rect 28972 2876 29012 2885
rect 28300 2659 28340 2668
rect 28684 2708 28724 2717
rect 28876 2708 28916 2717
rect 28724 2668 28876 2708
rect 28684 2659 28724 2668
rect 28876 2659 28916 2668
rect 28972 2624 29012 2836
rect 28972 2575 29012 2584
rect 29932 2036 29972 2045
rect 28011 1952 28053 1961
rect 28011 1912 28012 1952
rect 28052 1912 28053 1952
rect 28011 1903 28053 1912
rect 26379 1784 26421 1793
rect 26379 1744 26380 1784
rect 26420 1744 26421 1784
rect 26379 1735 26421 1744
rect 27819 1280 27861 1289
rect 27819 1240 27820 1280
rect 27860 1240 27861 1280
rect 27819 1231 27861 1240
rect 27820 692 27860 1231
rect 29932 1205 29972 1996
rect 29931 1196 29973 1205
rect 29931 1156 29932 1196
rect 29972 1156 29973 1196
rect 29931 1147 29973 1156
rect 30987 1112 31029 1121
rect 30987 1072 30988 1112
rect 31028 1072 31029 1112
rect 30987 1063 31029 1072
rect 31564 1112 31604 1121
rect 30988 978 31028 1063
rect 27820 643 27860 652
rect 25515 608 25557 617
rect 25515 568 25516 608
rect 25556 568 25557 608
rect 25515 559 25557 568
rect 31564 533 31604 1072
rect 32140 1112 32180 6364
rect 32236 5825 32276 8464
rect 32428 7664 32468 9640
rect 40972 9428 41012 9437
rect 33928 9092 34296 9101
rect 33968 9052 34010 9092
rect 34050 9052 34092 9092
rect 34132 9052 34174 9092
rect 34214 9052 34256 9092
rect 33928 9043 34296 9052
rect 32428 7615 32468 7624
rect 32524 9008 32564 9017
rect 32235 5816 32277 5825
rect 32235 5776 32236 5816
rect 32276 5776 32277 5816
rect 32235 5767 32277 5776
rect 32140 1063 32180 1072
rect 32524 692 32564 8968
rect 32715 9008 32757 9017
rect 32715 8968 32716 9008
rect 32756 8968 32757 9008
rect 32715 8959 32757 8968
rect 32620 8840 32660 8849
rect 32620 953 32660 8800
rect 32716 8168 32756 8959
rect 35307 8840 35349 8849
rect 35307 8800 35308 8840
rect 35348 8800 35349 8840
rect 35307 8791 35349 8800
rect 37900 8840 37940 8849
rect 35308 8706 35348 8791
rect 37900 8765 37940 8800
rect 37899 8756 37941 8765
rect 37804 8716 37900 8756
rect 37940 8716 37941 8756
rect 32716 8119 32756 8128
rect 34348 8504 34388 8513
rect 33291 8000 33333 8009
rect 33291 7960 33292 8000
rect 33332 7960 33333 8000
rect 33291 7951 33333 7960
rect 33292 7664 33332 7951
rect 33675 7832 33717 7841
rect 33675 7792 33676 7832
rect 33716 7792 33717 7832
rect 33675 7783 33717 7792
rect 33676 7698 33716 7783
rect 33292 7615 33332 7624
rect 33928 7580 34296 7589
rect 33968 7540 34010 7580
rect 34050 7540 34092 7580
rect 34132 7540 34174 7580
rect 34214 7540 34256 7580
rect 33928 7531 34296 7540
rect 33928 6068 34296 6077
rect 33968 6028 34010 6068
rect 34050 6028 34092 6068
rect 34132 6028 34174 6068
rect 34214 6028 34256 6068
rect 33928 6019 34296 6028
rect 32908 4724 32948 4733
rect 32908 1289 32948 4684
rect 33928 4556 34296 4565
rect 33968 4516 34010 4556
rect 34050 4516 34092 4556
rect 34132 4516 34174 4556
rect 34214 4516 34256 4556
rect 33928 4507 34296 4516
rect 33484 4220 33524 4229
rect 33484 3557 33524 4180
rect 33483 3548 33525 3557
rect 33483 3508 33484 3548
rect 33524 3508 33525 3548
rect 33483 3499 33525 3508
rect 33928 3044 34296 3053
rect 33968 3004 34010 3044
rect 34050 3004 34092 3044
rect 34132 3004 34174 3044
rect 34214 3004 34256 3044
rect 33928 2995 34296 3004
rect 33928 1532 34296 1541
rect 33968 1492 34010 1532
rect 34050 1492 34092 1532
rect 34132 1492 34174 1532
rect 34214 1492 34256 1532
rect 33928 1483 34296 1492
rect 32907 1280 32949 1289
rect 32907 1240 32908 1280
rect 32948 1240 32949 1280
rect 32907 1231 32949 1240
rect 34348 1037 34388 8464
rect 35168 8336 35536 8345
rect 35208 8296 35250 8336
rect 35290 8296 35332 8336
rect 35372 8296 35414 8336
rect 35454 8296 35496 8336
rect 35168 8287 35536 8296
rect 37131 8084 37173 8093
rect 37131 8044 37132 8084
rect 37172 8044 37173 8084
rect 37131 8035 37173 8044
rect 37132 8000 37172 8035
rect 37132 7949 37172 7960
rect 37324 7748 37364 7757
rect 35308 7580 35348 7589
rect 35308 7421 35348 7540
rect 35307 7412 35349 7421
rect 35307 7372 35308 7412
rect 35348 7372 35349 7412
rect 35307 7363 35349 7372
rect 35788 7244 35828 7253
rect 35168 6824 35536 6833
rect 35208 6784 35250 6824
rect 35290 6784 35332 6824
rect 35372 6784 35414 6824
rect 35454 6784 35496 6824
rect 35168 6775 35536 6784
rect 35307 6320 35349 6329
rect 35307 6280 35308 6320
rect 35348 6280 35349 6320
rect 35307 6271 35349 6280
rect 35308 6186 35348 6271
rect 35595 5648 35637 5657
rect 35595 5608 35596 5648
rect 35636 5608 35637 5648
rect 35595 5599 35637 5608
rect 35596 5514 35636 5599
rect 35168 5312 35536 5321
rect 35208 5272 35250 5312
rect 35290 5272 35332 5312
rect 35372 5272 35414 5312
rect 35454 5272 35496 5312
rect 35168 5263 35536 5272
rect 34923 4808 34965 4817
rect 34923 4768 34924 4808
rect 34964 4768 34965 4808
rect 34923 4759 34965 4768
rect 34924 4674 34964 4759
rect 35168 3800 35536 3809
rect 35208 3760 35250 3800
rect 35290 3760 35332 3800
rect 35372 3760 35414 3800
rect 35454 3760 35496 3800
rect 35168 3751 35536 3760
rect 35168 2288 35536 2297
rect 35208 2248 35250 2288
rect 35290 2248 35332 2288
rect 35372 2248 35414 2288
rect 35454 2248 35496 2288
rect 35168 2239 35536 2248
rect 35788 1121 35828 7204
rect 36171 6992 36213 7001
rect 36171 6952 36172 6992
rect 36212 6952 36213 6992
rect 36171 6943 36213 6952
rect 36172 6858 36212 6943
rect 37227 5480 37269 5489
rect 37227 5440 37228 5480
rect 37268 5440 37269 5480
rect 37227 5431 37269 5440
rect 37228 5346 37268 5431
rect 36556 2708 36596 2717
rect 36556 2540 36596 2668
rect 36556 2491 36596 2500
rect 37324 2129 37364 7708
rect 37804 7244 37844 8716
rect 37899 8707 37941 8716
rect 37900 8705 37940 8707
rect 40780 8672 40820 8681
rect 37899 8168 37941 8177
rect 37899 8128 37900 8168
rect 37940 8128 37941 8168
rect 37899 8119 37941 8128
rect 37804 7195 37844 7204
rect 37900 4892 37940 8119
rect 38188 8000 38228 8009
rect 38091 7748 38133 7757
rect 38091 7708 38092 7748
rect 38132 7708 38133 7748
rect 38091 7699 38133 7708
rect 38092 7614 38132 7699
rect 38188 6236 38228 7960
rect 40780 7160 40820 8632
rect 38188 6187 38228 6196
rect 38956 6404 38996 6413
rect 38956 5069 38996 6364
rect 40203 6320 40245 6329
rect 40203 6280 40204 6320
rect 40244 6280 40245 6320
rect 40203 6271 40245 6280
rect 40204 6186 40244 6271
rect 38955 5060 38997 5069
rect 38955 5020 38956 5060
rect 38996 5020 38997 5060
rect 38955 5011 38997 5020
rect 40300 5060 40340 5069
rect 37900 4843 37940 4852
rect 38859 4388 38901 4397
rect 38859 4348 38860 4388
rect 38900 4348 38901 4388
rect 38859 4339 38901 4348
rect 38860 4220 38900 4339
rect 38860 4171 38900 4180
rect 37612 3968 37652 3977
rect 37612 3800 37652 3928
rect 37804 3968 37844 3977
rect 37708 3800 37748 3809
rect 37612 3760 37708 3800
rect 37708 3751 37748 3760
rect 37323 2120 37365 2129
rect 37323 2080 37324 2120
rect 37364 2080 37365 2120
rect 37323 2071 37365 2080
rect 37804 2045 37844 3928
rect 37899 3212 37941 3221
rect 37899 3172 37900 3212
rect 37940 3172 37941 3212
rect 37899 3163 37941 3172
rect 37900 3078 37940 3163
rect 37803 2036 37845 2045
rect 37803 1996 37804 2036
rect 37844 1996 37845 2036
rect 37803 1987 37845 1996
rect 39243 1952 39285 1961
rect 39243 1912 39244 1952
rect 39284 1912 39285 1952
rect 39243 1903 39285 1912
rect 39244 1818 39284 1903
rect 40300 1448 40340 5020
rect 40780 4976 40820 7120
rect 40972 5657 41012 9388
rect 40971 5648 41013 5657
rect 40971 5608 40972 5648
rect 41012 5608 41013 5648
rect 40971 5599 41013 5608
rect 40780 3548 40820 4936
rect 41259 4892 41301 4901
rect 41259 4852 41260 4892
rect 41300 4852 41301 4892
rect 41259 4843 41301 4852
rect 41260 4758 41300 4843
rect 41548 4724 41588 4733
rect 41548 4313 41588 4684
rect 41547 4304 41589 4313
rect 41547 4264 41548 4304
rect 41588 4264 41589 4304
rect 41547 4255 41589 4264
rect 40780 3499 40820 3508
rect 41644 3464 41684 3475
rect 41644 3389 41684 3424
rect 41643 3380 41685 3389
rect 41643 3340 41644 3380
rect 41684 3340 41685 3380
rect 41643 3331 41685 3340
rect 41739 3296 41781 3305
rect 41739 3256 41740 3296
rect 41780 3256 41781 3296
rect 41739 3247 41781 3256
rect 41740 3128 41780 3247
rect 41740 3079 41780 3088
rect 42507 2792 42549 2801
rect 42507 2752 42508 2792
rect 42548 2752 42549 2792
rect 42507 2743 42549 2752
rect 42508 2658 42548 2743
rect 42507 2456 42549 2465
rect 42507 2416 42508 2456
rect 42548 2416 42549 2456
rect 42507 2407 42549 2416
rect 42508 2322 42548 2407
rect 40300 1399 40340 1408
rect 35787 1112 35829 1121
rect 35787 1072 35788 1112
rect 35828 1072 35829 1112
rect 35787 1063 35829 1072
rect 34347 1028 34389 1037
rect 34347 988 34348 1028
rect 34388 988 34389 1028
rect 34347 979 34389 988
rect 32619 944 32661 953
rect 32619 904 32620 944
rect 32660 904 32661 944
rect 32619 895 32661 904
rect 40971 944 41013 953
rect 40971 904 40972 944
rect 41012 904 41013 944
rect 40971 895 41013 904
rect 40972 810 41012 895
rect 35168 776 35536 785
rect 35208 736 35250 776
rect 35290 736 35332 776
rect 35372 736 35414 776
rect 35454 736 35496 776
rect 35168 727 35536 736
rect 32524 643 32564 652
rect 31563 524 31605 533
rect 31563 484 31564 524
rect 31604 484 31605 524
rect 31563 475 31605 484
rect 19948 139 19988 148
<< via4 >>
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 8812 9388 8852 9428
rect 1612 9220 1652 9260
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 1708 8884 1748 8924
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 4588 7960 4628 8000
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 6892 7120 6932 7160
rect 3340 5608 3380 5648
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 1324 4096 1364 4136
rect 1324 3508 1364 3548
rect 2956 3340 2996 3380
rect 1900 1912 1940 1952
rect 460 1828 500 1868
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 6220 5608 6260 5648
rect 5356 4936 5396 4976
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 4108 1828 4148 1868
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 2572 1072 2612 1112
rect 11020 5860 11060 5900
rect 10636 4936 10676 4976
rect 10636 4684 10676 4724
rect 9772 1072 9812 1112
rect 12844 7204 12884 7244
rect 12556 3760 12596 3800
rect 12556 3508 12596 3548
rect 11212 904 11252 944
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 13804 8044 13844 8084
rect 15436 9220 15476 9260
rect 15244 6952 15284 6992
rect 15052 5776 15092 5816
rect 14668 5692 14708 5732
rect 14284 5440 14324 5480
rect 15436 5020 15476 5060
rect 15532 2080 15572 2120
rect 16396 8464 16436 8504
rect 15820 7792 15860 7832
rect 16300 3508 16340 3548
rect 15916 3424 15956 3464
rect 16972 7372 17012 7412
rect 16780 6364 16820 6404
rect 16588 4264 16628 4304
rect 15628 1996 15668 2036
rect 13804 1744 13844 1784
rect 17644 7708 17684 7748
rect 17068 3172 17108 3212
rect 17644 7036 17684 7076
rect 17932 6196 17972 6236
rect 18124 4852 18164 4892
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 19468 8128 19508 8168
rect 19564 7960 19604 8000
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 18508 3592 18548 3632
rect 18412 3508 18452 3548
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 20716 7708 20756 7748
rect 21004 8968 21044 9008
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 13804 1156 13844 1196
rect 19468 4936 19508 4976
rect 19468 3760 19508 3800
rect 13996 1072 14036 1112
rect 19372 1072 19412 1112
rect 13708 988 13748 1028
rect 13516 820 13556 860
rect 13228 568 13268 608
rect 19468 820 19508 860
rect 19372 484 19412 524
rect 20044 4432 20084 4472
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 21196 4684 21236 4724
rect 21484 8464 21524 8504
rect 21388 7624 21428 7664
rect 21484 6364 21524 6404
rect 21388 4768 21428 4808
rect 21388 4096 21428 4136
rect 24748 9388 24788 9428
rect 24076 8800 24116 8840
rect 23020 8044 23060 8084
rect 24076 7960 24116 8000
rect 26476 9052 26516 9092
rect 27724 9220 27764 9260
rect 25516 8044 25556 8084
rect 22636 7120 22676 7160
rect 24364 5608 24404 5648
rect 23884 5020 23924 5060
rect 22060 4432 22100 4472
rect 22636 3928 22676 3968
rect 22636 3424 22676 3464
rect 25228 3340 25268 3380
rect 24940 3256 24980 3296
rect 24556 2416 24596 2456
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 22828 1912 22868 1952
rect 25132 1828 25172 1868
rect 24556 904 24596 944
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 26476 5860 26516 5900
rect 26476 3592 26516 3632
rect 26476 3340 26516 3380
rect 27724 8548 27764 8588
rect 28012 7036 28052 7076
rect 35168 9808 35208 9848
rect 35250 9808 35290 9848
rect 35332 9808 35372 9848
rect 35414 9808 35454 9848
rect 35496 9808 35536 9848
rect 31660 9052 31700 9092
rect 28588 8044 28628 8084
rect 28780 7960 28820 8000
rect 28396 7036 28436 7076
rect 28012 6280 28052 6320
rect 27148 4936 27188 4976
rect 27148 4348 27188 4388
rect 27628 2752 27668 2792
rect 30316 8548 30356 8588
rect 31948 8044 31988 8084
rect 31564 7204 31604 7244
rect 30220 7120 30260 7160
rect 31468 5692 31508 5732
rect 31276 5020 31316 5060
rect 30892 4768 30932 4808
rect 31468 4768 31508 4808
rect 28396 3928 28436 3968
rect 28012 1912 28052 1952
rect 26380 1744 26420 1784
rect 27820 1240 27860 1280
rect 29932 1156 29972 1196
rect 30988 1072 31028 1112
rect 25516 568 25556 608
rect 33928 9052 33968 9092
rect 34010 9052 34050 9092
rect 34092 9052 34132 9092
rect 34174 9052 34214 9092
rect 34256 9052 34296 9092
rect 32236 5776 32276 5816
rect 32716 8968 32756 9008
rect 35308 8800 35348 8840
rect 37900 8716 37940 8756
rect 33292 7960 33332 8000
rect 33676 7792 33716 7832
rect 33928 7540 33968 7580
rect 34010 7540 34050 7580
rect 34092 7540 34132 7580
rect 34174 7540 34214 7580
rect 34256 7540 34296 7580
rect 33928 6028 33968 6068
rect 34010 6028 34050 6068
rect 34092 6028 34132 6068
rect 34174 6028 34214 6068
rect 34256 6028 34296 6068
rect 33928 4516 33968 4556
rect 34010 4516 34050 4556
rect 34092 4516 34132 4556
rect 34174 4516 34214 4556
rect 34256 4516 34296 4556
rect 33484 3508 33524 3548
rect 33928 3004 33968 3044
rect 34010 3004 34050 3044
rect 34092 3004 34132 3044
rect 34174 3004 34214 3044
rect 34256 3004 34296 3044
rect 33928 1492 33968 1532
rect 34010 1492 34050 1532
rect 34092 1492 34132 1532
rect 34174 1492 34214 1532
rect 34256 1492 34296 1532
rect 32908 1240 32948 1280
rect 35168 8296 35208 8336
rect 35250 8296 35290 8336
rect 35332 8296 35372 8336
rect 35414 8296 35454 8336
rect 35496 8296 35536 8336
rect 37132 8044 37172 8084
rect 35308 7372 35348 7412
rect 35168 6784 35208 6824
rect 35250 6784 35290 6824
rect 35332 6784 35372 6824
rect 35414 6784 35454 6824
rect 35496 6784 35536 6824
rect 35308 6280 35348 6320
rect 35596 5608 35636 5648
rect 35168 5272 35208 5312
rect 35250 5272 35290 5312
rect 35332 5272 35372 5312
rect 35414 5272 35454 5312
rect 35496 5272 35536 5312
rect 34924 4768 34964 4808
rect 35168 3760 35208 3800
rect 35250 3760 35290 3800
rect 35332 3760 35372 3800
rect 35414 3760 35454 3800
rect 35496 3760 35536 3800
rect 35168 2248 35208 2288
rect 35250 2248 35290 2288
rect 35332 2248 35372 2288
rect 35414 2248 35454 2288
rect 35496 2248 35536 2288
rect 36172 6952 36212 6992
rect 37228 5440 37268 5480
rect 37900 8128 37940 8168
rect 38092 7708 38132 7748
rect 40204 6280 40244 6320
rect 38956 5020 38996 5060
rect 38860 4348 38900 4388
rect 37324 2080 37364 2120
rect 37900 3172 37940 3212
rect 37804 1996 37844 2036
rect 39244 1912 39284 1952
rect 40972 5608 41012 5648
rect 41260 4852 41300 4892
rect 41548 4264 41588 4304
rect 41644 3340 41684 3380
rect 41740 3256 41780 3296
rect 42508 2752 42548 2792
rect 42508 2416 42548 2456
rect 35788 1072 35828 1112
rect 34348 988 34388 1028
rect 32620 904 32660 944
rect 40972 904 41012 944
rect 35168 736 35208 776
rect 35250 736 35290 776
rect 35332 736 35372 776
rect 35414 736 35454 776
rect 35496 736 35536 776
rect 31564 484 31604 524
<< metal5 >>
rect 4919 9871 5305 9890
rect 4919 9848 4985 9871
rect 5071 9848 5153 9871
rect 5239 9848 5305 9871
rect 4919 9808 4928 9848
rect 4968 9808 4985 9848
rect 5071 9808 5092 9848
rect 5132 9808 5153 9848
rect 5239 9808 5256 9848
rect 5296 9808 5305 9848
rect 4919 9785 4985 9808
rect 5071 9785 5153 9808
rect 5239 9785 5305 9808
rect 4919 9766 5305 9785
rect 20039 9871 20425 9890
rect 20039 9848 20105 9871
rect 20191 9848 20273 9871
rect 20359 9848 20425 9871
rect 20039 9808 20048 9848
rect 20088 9808 20105 9848
rect 20191 9808 20212 9848
rect 20252 9808 20273 9848
rect 20359 9808 20376 9848
rect 20416 9808 20425 9848
rect 20039 9785 20105 9808
rect 20191 9785 20273 9808
rect 20359 9785 20425 9808
rect 20039 9766 20425 9785
rect 35159 9871 35545 9890
rect 35159 9848 35225 9871
rect 35311 9848 35393 9871
rect 35479 9848 35545 9871
rect 35159 9808 35168 9848
rect 35208 9808 35225 9848
rect 35311 9808 35332 9848
rect 35372 9808 35393 9848
rect 35479 9808 35496 9848
rect 35536 9808 35545 9848
rect 35159 9785 35225 9808
rect 35311 9785 35393 9808
rect 35479 9785 35545 9808
rect 35159 9766 35545 9785
rect 8803 9388 8812 9428
rect 8852 9388 24748 9428
rect 24788 9388 24797 9428
rect 1603 9220 1612 9260
rect 1652 9220 11360 9260
rect 15427 9220 15436 9260
rect 15476 9220 27724 9260
rect 27764 9220 27773 9260
rect 3679 9115 4065 9134
rect 3679 9092 3745 9115
rect 3831 9092 3913 9115
rect 3999 9092 4065 9115
rect 3679 9052 3688 9092
rect 3728 9052 3745 9092
rect 3831 9052 3852 9092
rect 3892 9052 3913 9092
rect 3999 9052 4016 9092
rect 4056 9052 4065 9092
rect 3679 9029 3745 9052
rect 3831 9029 3913 9052
rect 3999 9029 4065 9052
rect 3679 9010 4065 9029
rect 11320 8924 11360 9220
rect 18799 9115 19185 9134
rect 18799 9092 18865 9115
rect 18951 9092 19033 9115
rect 19119 9092 19185 9115
rect 33919 9115 34305 9134
rect 33919 9092 33985 9115
rect 34071 9092 34153 9115
rect 34239 9092 34305 9115
rect 18799 9052 18808 9092
rect 18848 9052 18865 9092
rect 18951 9052 18972 9092
rect 19012 9052 19033 9092
rect 19119 9052 19136 9092
rect 19176 9052 19185 9092
rect 26467 9052 26476 9092
rect 26516 9052 31660 9092
rect 31700 9052 31709 9092
rect 33919 9052 33928 9092
rect 33968 9052 33985 9092
rect 34071 9052 34092 9092
rect 34132 9052 34153 9092
rect 34239 9052 34256 9092
rect 34296 9052 34305 9092
rect 18799 9029 18865 9052
rect 18951 9029 19033 9052
rect 19119 9029 19185 9052
rect 18799 9010 19185 9029
rect 33919 9029 33985 9052
rect 34071 9029 34153 9052
rect 34239 9029 34305 9052
rect 33919 9010 34305 9029
rect 20140 8968 21004 9008
rect 21044 8968 32716 9008
rect 32756 8968 32765 9008
rect 20140 8924 20180 8968
rect 1699 8884 1708 8924
rect 1748 8884 2540 8924
rect 11320 8884 20180 8924
rect 2500 8840 2540 8884
rect 2500 8800 24076 8840
rect 24116 8800 24125 8840
rect 35299 8800 35308 8840
rect 35348 8800 35357 8840
rect 35308 8756 35348 8800
rect 35308 8716 37900 8756
rect 37940 8716 37949 8756
rect 27715 8548 27724 8588
rect 27764 8548 30316 8588
rect 30356 8548 30365 8588
rect 16387 8464 16396 8504
rect 16436 8464 21484 8504
rect 21524 8464 21533 8504
rect 4919 8359 5305 8378
rect 4919 8336 4985 8359
rect 5071 8336 5153 8359
rect 5239 8336 5305 8359
rect 4919 8296 4928 8336
rect 4968 8296 4985 8336
rect 5071 8296 5092 8336
rect 5132 8296 5153 8336
rect 5239 8296 5256 8336
rect 5296 8296 5305 8336
rect 4919 8273 4985 8296
rect 5071 8273 5153 8296
rect 5239 8273 5305 8296
rect 4919 8254 5305 8273
rect 20039 8359 20425 8378
rect 20039 8336 20105 8359
rect 20191 8336 20273 8359
rect 20359 8336 20425 8359
rect 20039 8296 20048 8336
rect 20088 8296 20105 8336
rect 20191 8296 20212 8336
rect 20252 8296 20273 8336
rect 20359 8296 20376 8336
rect 20416 8296 20425 8336
rect 20039 8273 20105 8296
rect 20191 8273 20273 8296
rect 20359 8273 20425 8296
rect 20039 8254 20425 8273
rect 35159 8359 35545 8378
rect 35159 8336 35225 8359
rect 35311 8336 35393 8359
rect 35479 8336 35545 8359
rect 35159 8296 35168 8336
rect 35208 8296 35225 8336
rect 35311 8296 35332 8336
rect 35372 8296 35393 8336
rect 35479 8296 35496 8336
rect 35536 8296 35545 8336
rect 35159 8273 35225 8296
rect 35311 8273 35393 8296
rect 35479 8273 35545 8296
rect 35159 8254 35545 8273
rect 19459 8128 19468 8168
rect 19508 8128 37900 8168
rect 37940 8128 37949 8168
rect 13795 8044 13804 8084
rect 13844 8044 23020 8084
rect 23060 8044 23069 8084
rect 25507 8044 25516 8084
rect 25556 8044 28588 8084
rect 28628 8044 28637 8084
rect 31939 8044 31948 8084
rect 31988 8044 37132 8084
rect 37172 8044 37181 8084
rect 4579 7960 4588 8000
rect 4628 7960 19564 8000
rect 19604 7960 19613 8000
rect 24067 7960 24076 8000
rect 24116 7960 28780 8000
rect 28820 7960 33292 8000
rect 33332 7960 33341 8000
rect 15811 7792 15820 7832
rect 15860 7792 33676 7832
rect 33716 7792 33725 7832
rect 17635 7708 17644 7748
rect 17684 7708 20180 7748
rect 20707 7708 20716 7748
rect 20756 7708 38092 7748
rect 38132 7708 38141 7748
rect 20140 7664 20180 7708
rect 20140 7624 21388 7664
rect 21428 7624 21437 7664
rect 3679 7603 4065 7622
rect 3679 7580 3745 7603
rect 3831 7580 3913 7603
rect 3999 7580 4065 7603
rect 3679 7540 3688 7580
rect 3728 7540 3745 7580
rect 3831 7540 3852 7580
rect 3892 7540 3913 7580
rect 3999 7540 4016 7580
rect 4056 7540 4065 7580
rect 3679 7517 3745 7540
rect 3831 7517 3913 7540
rect 3999 7517 4065 7540
rect 3679 7498 4065 7517
rect 18799 7603 19185 7622
rect 18799 7580 18865 7603
rect 18951 7580 19033 7603
rect 19119 7580 19185 7603
rect 18799 7540 18808 7580
rect 18848 7540 18865 7580
rect 18951 7540 18972 7580
rect 19012 7540 19033 7580
rect 19119 7540 19136 7580
rect 19176 7540 19185 7580
rect 18799 7517 18865 7540
rect 18951 7517 19033 7540
rect 19119 7517 19185 7540
rect 18799 7498 19185 7517
rect 33919 7603 34305 7622
rect 33919 7580 33985 7603
rect 34071 7580 34153 7603
rect 34239 7580 34305 7603
rect 33919 7540 33928 7580
rect 33968 7540 33985 7580
rect 34071 7540 34092 7580
rect 34132 7540 34153 7580
rect 34239 7540 34256 7580
rect 34296 7540 34305 7580
rect 33919 7517 33985 7540
rect 34071 7517 34153 7540
rect 34239 7517 34305 7540
rect 33919 7498 34305 7517
rect 16963 7372 16972 7412
rect 17012 7372 35308 7412
rect 35348 7372 35357 7412
rect 12835 7204 12844 7244
rect 12884 7204 31564 7244
rect 31604 7204 31613 7244
rect 6883 7120 6892 7160
rect 6932 7120 22636 7160
rect 22676 7120 30220 7160
rect 30260 7120 30269 7160
rect 17635 7036 17644 7076
rect 17684 7036 28012 7076
rect 28052 7036 28396 7076
rect 28436 7036 28445 7076
rect 15235 6952 15244 6992
rect 15284 6952 36172 6992
rect 36212 6952 36221 6992
rect 4919 6847 5305 6866
rect 4919 6824 4985 6847
rect 5071 6824 5153 6847
rect 5239 6824 5305 6847
rect 4919 6784 4928 6824
rect 4968 6784 4985 6824
rect 5071 6784 5092 6824
rect 5132 6784 5153 6824
rect 5239 6784 5256 6824
rect 5296 6784 5305 6824
rect 4919 6761 4985 6784
rect 5071 6761 5153 6784
rect 5239 6761 5305 6784
rect 4919 6742 5305 6761
rect 20039 6847 20425 6866
rect 20039 6824 20105 6847
rect 20191 6824 20273 6847
rect 20359 6824 20425 6847
rect 20039 6784 20048 6824
rect 20088 6784 20105 6824
rect 20191 6784 20212 6824
rect 20252 6784 20273 6824
rect 20359 6784 20376 6824
rect 20416 6784 20425 6824
rect 20039 6761 20105 6784
rect 20191 6761 20273 6784
rect 20359 6761 20425 6784
rect 20039 6742 20425 6761
rect 35159 6847 35545 6866
rect 35159 6824 35225 6847
rect 35311 6824 35393 6847
rect 35479 6824 35545 6847
rect 35159 6784 35168 6824
rect 35208 6784 35225 6824
rect 35311 6784 35332 6824
rect 35372 6784 35393 6824
rect 35479 6784 35496 6824
rect 35536 6784 35545 6824
rect 35159 6761 35225 6784
rect 35311 6761 35393 6784
rect 35479 6761 35545 6784
rect 35159 6742 35545 6761
rect 16771 6364 16780 6404
rect 16820 6364 21484 6404
rect 21524 6364 21533 6404
rect 28003 6280 28012 6320
rect 28052 6280 35308 6320
rect 35348 6280 35357 6320
rect 37708 6280 40204 6320
rect 40244 6280 40253 6320
rect 37708 6236 37748 6280
rect 17923 6196 17932 6236
rect 17972 6196 37748 6236
rect 3679 6091 4065 6110
rect 3679 6068 3745 6091
rect 3831 6068 3913 6091
rect 3999 6068 4065 6091
rect 3679 6028 3688 6068
rect 3728 6028 3745 6068
rect 3831 6028 3852 6068
rect 3892 6028 3913 6068
rect 3999 6028 4016 6068
rect 4056 6028 4065 6068
rect 3679 6005 3745 6028
rect 3831 6005 3913 6028
rect 3999 6005 4065 6028
rect 3679 5986 4065 6005
rect 18799 6091 19185 6110
rect 18799 6068 18865 6091
rect 18951 6068 19033 6091
rect 19119 6068 19185 6091
rect 18799 6028 18808 6068
rect 18848 6028 18865 6068
rect 18951 6028 18972 6068
rect 19012 6028 19033 6068
rect 19119 6028 19136 6068
rect 19176 6028 19185 6068
rect 18799 6005 18865 6028
rect 18951 6005 19033 6028
rect 19119 6005 19185 6028
rect 18799 5986 19185 6005
rect 33919 6091 34305 6110
rect 33919 6068 33985 6091
rect 34071 6068 34153 6091
rect 34239 6068 34305 6091
rect 33919 6028 33928 6068
rect 33968 6028 33985 6068
rect 34071 6028 34092 6068
rect 34132 6028 34153 6068
rect 34239 6028 34256 6068
rect 34296 6028 34305 6068
rect 33919 6005 33985 6028
rect 34071 6005 34153 6028
rect 34239 6005 34305 6028
rect 33919 5986 34305 6005
rect 11011 5860 11020 5900
rect 11060 5860 26476 5900
rect 26516 5860 26525 5900
rect 15043 5776 15052 5816
rect 15092 5776 32236 5816
rect 32276 5776 32285 5816
rect 14659 5692 14668 5732
rect 14708 5692 31468 5732
rect 31508 5692 31517 5732
rect 3331 5608 3340 5648
rect 3380 5608 6220 5648
rect 6260 5608 6269 5648
rect 24355 5608 24364 5648
rect 24404 5608 35596 5648
rect 35636 5608 40972 5648
rect 41012 5608 41021 5648
rect 14275 5440 14284 5480
rect 14324 5440 37228 5480
rect 37268 5440 37277 5480
rect 4919 5335 5305 5354
rect 4919 5312 4985 5335
rect 5071 5312 5153 5335
rect 5239 5312 5305 5335
rect 4919 5272 4928 5312
rect 4968 5272 4985 5312
rect 5071 5272 5092 5312
rect 5132 5272 5153 5312
rect 5239 5272 5256 5312
rect 5296 5272 5305 5312
rect 4919 5249 4985 5272
rect 5071 5249 5153 5272
rect 5239 5249 5305 5272
rect 4919 5230 5305 5249
rect 20039 5335 20425 5354
rect 20039 5312 20105 5335
rect 20191 5312 20273 5335
rect 20359 5312 20425 5335
rect 20039 5272 20048 5312
rect 20088 5272 20105 5312
rect 20191 5272 20212 5312
rect 20252 5272 20273 5312
rect 20359 5272 20376 5312
rect 20416 5272 20425 5312
rect 20039 5249 20105 5272
rect 20191 5249 20273 5272
rect 20359 5249 20425 5272
rect 20039 5230 20425 5249
rect 35159 5335 35545 5354
rect 35159 5312 35225 5335
rect 35311 5312 35393 5335
rect 35479 5312 35545 5335
rect 35159 5272 35168 5312
rect 35208 5272 35225 5312
rect 35311 5272 35332 5312
rect 35372 5272 35393 5312
rect 35479 5272 35496 5312
rect 35536 5272 35545 5312
rect 35159 5249 35225 5272
rect 35311 5249 35393 5272
rect 35479 5249 35545 5272
rect 35159 5230 35545 5249
rect 15427 5020 15436 5060
rect 15476 5020 23884 5060
rect 23924 5020 23933 5060
rect 28960 5020 31276 5060
rect 31316 5020 38956 5060
rect 38996 5020 39005 5060
rect 28960 4976 29000 5020
rect 5347 4936 5356 4976
rect 5396 4936 10636 4976
rect 10676 4936 10685 4976
rect 19459 4936 19468 4976
rect 19508 4936 27148 4976
rect 27188 4936 29000 4976
rect 18115 4852 18124 4892
rect 18164 4852 41260 4892
rect 41300 4852 41309 4892
rect 21379 4768 21388 4808
rect 21428 4768 30892 4808
rect 30932 4768 30941 4808
rect 31459 4768 31468 4808
rect 31508 4768 34924 4808
rect 34964 4768 34973 4808
rect 10627 4684 10636 4724
rect 10676 4684 21196 4724
rect 21236 4684 21245 4724
rect 3679 4579 4065 4598
rect 3679 4556 3745 4579
rect 3831 4556 3913 4579
rect 3999 4556 4065 4579
rect 3679 4516 3688 4556
rect 3728 4516 3745 4556
rect 3831 4516 3852 4556
rect 3892 4516 3913 4556
rect 3999 4516 4016 4556
rect 4056 4516 4065 4556
rect 3679 4493 3745 4516
rect 3831 4493 3913 4516
rect 3999 4493 4065 4516
rect 3679 4474 4065 4493
rect 18799 4579 19185 4598
rect 18799 4556 18865 4579
rect 18951 4556 19033 4579
rect 19119 4556 19185 4579
rect 18799 4516 18808 4556
rect 18848 4516 18865 4556
rect 18951 4516 18972 4556
rect 19012 4516 19033 4556
rect 19119 4516 19136 4556
rect 19176 4516 19185 4556
rect 18799 4493 18865 4516
rect 18951 4493 19033 4516
rect 19119 4493 19185 4516
rect 18799 4474 19185 4493
rect 33919 4579 34305 4598
rect 33919 4556 33985 4579
rect 34071 4556 34153 4579
rect 34239 4556 34305 4579
rect 33919 4516 33928 4556
rect 33968 4516 33985 4556
rect 34071 4516 34092 4556
rect 34132 4516 34153 4556
rect 34239 4516 34256 4556
rect 34296 4516 34305 4556
rect 33919 4493 33985 4516
rect 34071 4493 34153 4516
rect 34239 4493 34305 4516
rect 33919 4474 34305 4493
rect 20035 4432 20044 4472
rect 20084 4432 22060 4472
rect 22100 4432 22109 4472
rect 27139 4348 27148 4388
rect 27188 4348 38860 4388
rect 38900 4348 38909 4388
rect 16579 4264 16588 4304
rect 16628 4264 41548 4304
rect 41588 4264 41597 4304
rect 1315 4096 1324 4136
rect 1364 4096 21388 4136
rect 21428 4096 21437 4136
rect 22627 3928 22636 3968
rect 22676 3928 28396 3968
rect 28436 3928 28445 3968
rect 4919 3823 5305 3842
rect 4919 3800 4985 3823
rect 5071 3800 5153 3823
rect 5239 3800 5305 3823
rect 20039 3823 20425 3842
rect 20039 3800 20105 3823
rect 20191 3800 20273 3823
rect 20359 3800 20425 3823
rect 4919 3760 4928 3800
rect 4968 3760 4985 3800
rect 5071 3760 5092 3800
rect 5132 3760 5153 3800
rect 5239 3760 5256 3800
rect 5296 3760 5305 3800
rect 12547 3760 12556 3800
rect 12596 3760 19468 3800
rect 19508 3760 19517 3800
rect 20039 3760 20048 3800
rect 20088 3760 20105 3800
rect 20191 3760 20212 3800
rect 20252 3760 20273 3800
rect 20359 3760 20376 3800
rect 20416 3760 20425 3800
rect 4919 3737 4985 3760
rect 5071 3737 5153 3760
rect 5239 3737 5305 3760
rect 4919 3718 5305 3737
rect 20039 3737 20105 3760
rect 20191 3737 20273 3760
rect 20359 3737 20425 3760
rect 20039 3718 20425 3737
rect 35159 3823 35545 3842
rect 35159 3800 35225 3823
rect 35311 3800 35393 3823
rect 35479 3800 35545 3823
rect 35159 3760 35168 3800
rect 35208 3760 35225 3800
rect 35311 3760 35332 3800
rect 35372 3760 35393 3800
rect 35479 3760 35496 3800
rect 35536 3760 35545 3800
rect 35159 3737 35225 3760
rect 35311 3737 35393 3760
rect 35479 3737 35545 3760
rect 35159 3718 35545 3737
rect 18499 3592 18508 3632
rect 18548 3592 26476 3632
rect 26516 3592 26525 3632
rect 1315 3508 1324 3548
rect 1364 3508 12556 3548
rect 12596 3508 12605 3548
rect 16291 3508 16300 3548
rect 16340 3508 18412 3548
rect 18452 3508 33484 3548
rect 33524 3508 33533 3548
rect 15907 3424 15916 3464
rect 15956 3424 22636 3464
rect 22676 3424 22685 3464
rect 2947 3340 2956 3380
rect 2996 3340 25228 3380
rect 25268 3340 25277 3380
rect 26467 3340 26476 3380
rect 26516 3340 41644 3380
rect 41684 3340 41693 3380
rect 24931 3256 24940 3296
rect 24980 3256 41740 3296
rect 41780 3256 41789 3296
rect 17059 3172 17068 3212
rect 17108 3172 37900 3212
rect 37940 3172 37949 3212
rect 3679 3067 4065 3086
rect 3679 3044 3745 3067
rect 3831 3044 3913 3067
rect 3999 3044 4065 3067
rect 3679 3004 3688 3044
rect 3728 3004 3745 3044
rect 3831 3004 3852 3044
rect 3892 3004 3913 3044
rect 3999 3004 4016 3044
rect 4056 3004 4065 3044
rect 3679 2981 3745 3004
rect 3831 2981 3913 3004
rect 3999 2981 4065 3004
rect 3679 2962 4065 2981
rect 18799 3067 19185 3086
rect 18799 3044 18865 3067
rect 18951 3044 19033 3067
rect 19119 3044 19185 3067
rect 18799 3004 18808 3044
rect 18848 3004 18865 3044
rect 18951 3004 18972 3044
rect 19012 3004 19033 3044
rect 19119 3004 19136 3044
rect 19176 3004 19185 3044
rect 18799 2981 18865 3004
rect 18951 2981 19033 3004
rect 19119 2981 19185 3004
rect 18799 2962 19185 2981
rect 33919 3067 34305 3086
rect 33919 3044 33985 3067
rect 34071 3044 34153 3067
rect 34239 3044 34305 3067
rect 33919 3004 33928 3044
rect 33968 3004 33985 3044
rect 34071 3004 34092 3044
rect 34132 3004 34153 3044
rect 34239 3004 34256 3044
rect 34296 3004 34305 3044
rect 33919 2981 33985 3004
rect 34071 2981 34153 3004
rect 34239 2981 34305 3004
rect 33919 2962 34305 2981
rect 27619 2752 27628 2792
rect 27668 2752 42508 2792
rect 42548 2752 42557 2792
rect 24547 2416 24556 2456
rect 24596 2416 42508 2456
rect 42548 2416 42557 2456
rect 4919 2311 5305 2330
rect 4919 2288 4985 2311
rect 5071 2288 5153 2311
rect 5239 2288 5305 2311
rect 4919 2248 4928 2288
rect 4968 2248 4985 2288
rect 5071 2248 5092 2288
rect 5132 2248 5153 2288
rect 5239 2248 5256 2288
rect 5296 2248 5305 2288
rect 4919 2225 4985 2248
rect 5071 2225 5153 2248
rect 5239 2225 5305 2248
rect 4919 2206 5305 2225
rect 20039 2311 20425 2330
rect 20039 2288 20105 2311
rect 20191 2288 20273 2311
rect 20359 2288 20425 2311
rect 20039 2248 20048 2288
rect 20088 2248 20105 2288
rect 20191 2248 20212 2288
rect 20252 2248 20273 2288
rect 20359 2248 20376 2288
rect 20416 2248 20425 2288
rect 20039 2225 20105 2248
rect 20191 2225 20273 2248
rect 20359 2225 20425 2248
rect 20039 2206 20425 2225
rect 35159 2311 35545 2330
rect 35159 2288 35225 2311
rect 35311 2288 35393 2311
rect 35479 2288 35545 2311
rect 35159 2248 35168 2288
rect 35208 2248 35225 2288
rect 35311 2248 35332 2288
rect 35372 2248 35393 2288
rect 35479 2248 35496 2288
rect 35536 2248 35545 2288
rect 35159 2225 35225 2248
rect 35311 2225 35393 2248
rect 35479 2225 35545 2248
rect 35159 2206 35545 2225
rect 15523 2080 15532 2120
rect 15572 2080 37324 2120
rect 37364 2080 37373 2120
rect 15619 1996 15628 2036
rect 15668 1996 37804 2036
rect 37844 1996 37853 2036
rect 1891 1912 1900 1952
rect 1940 1912 22828 1952
rect 22868 1912 22877 1952
rect 28003 1912 28012 1952
rect 28052 1912 39244 1952
rect 39284 1912 39293 1952
rect 451 1828 460 1868
rect 500 1828 4108 1868
rect 4148 1828 25132 1868
rect 25172 1828 25181 1868
rect 13795 1744 13804 1784
rect 13844 1744 26380 1784
rect 26420 1744 26429 1784
rect 3679 1555 4065 1574
rect 3679 1532 3745 1555
rect 3831 1532 3913 1555
rect 3999 1532 4065 1555
rect 3679 1492 3688 1532
rect 3728 1492 3745 1532
rect 3831 1492 3852 1532
rect 3892 1492 3913 1532
rect 3999 1492 4016 1532
rect 4056 1492 4065 1532
rect 3679 1469 3745 1492
rect 3831 1469 3913 1492
rect 3999 1469 4065 1492
rect 3679 1450 4065 1469
rect 18799 1555 19185 1574
rect 18799 1532 18865 1555
rect 18951 1532 19033 1555
rect 19119 1532 19185 1555
rect 18799 1492 18808 1532
rect 18848 1492 18865 1532
rect 18951 1492 18972 1532
rect 19012 1492 19033 1532
rect 19119 1492 19136 1532
rect 19176 1492 19185 1532
rect 18799 1469 18865 1492
rect 18951 1469 19033 1492
rect 19119 1469 19185 1492
rect 18799 1450 19185 1469
rect 33919 1555 34305 1574
rect 33919 1532 33985 1555
rect 34071 1532 34153 1555
rect 34239 1532 34305 1555
rect 33919 1492 33928 1532
rect 33968 1492 33985 1532
rect 34071 1492 34092 1532
rect 34132 1492 34153 1532
rect 34239 1492 34256 1532
rect 34296 1492 34305 1532
rect 33919 1469 33985 1492
rect 34071 1469 34153 1492
rect 34239 1469 34305 1492
rect 33919 1450 34305 1469
rect 27811 1240 27820 1280
rect 27860 1240 32908 1280
rect 32948 1240 32957 1280
rect 13795 1156 13804 1196
rect 13844 1156 29932 1196
rect 29972 1156 29981 1196
rect 2563 1072 2572 1112
rect 2612 1072 9772 1112
rect 9812 1072 13996 1112
rect 14036 1072 19372 1112
rect 19412 1072 19421 1112
rect 30979 1072 30988 1112
rect 31028 1072 35788 1112
rect 35828 1072 35837 1112
rect 13699 988 13708 1028
rect 13748 988 34348 1028
rect 34388 988 34397 1028
rect 11203 904 11212 944
rect 11252 904 24556 944
rect 24596 904 24605 944
rect 32611 904 32620 944
rect 32660 904 40972 944
rect 41012 904 41021 944
rect 13507 820 13516 860
rect 13556 820 19468 860
rect 19508 820 19517 860
rect 4919 799 5305 818
rect 4919 776 4985 799
rect 5071 776 5153 799
rect 5239 776 5305 799
rect 4919 736 4928 776
rect 4968 736 4985 776
rect 5071 736 5092 776
rect 5132 736 5153 776
rect 5239 736 5256 776
rect 5296 736 5305 776
rect 4919 713 4985 736
rect 5071 713 5153 736
rect 5239 713 5305 736
rect 4919 694 5305 713
rect 20039 799 20425 818
rect 20039 776 20105 799
rect 20191 776 20273 799
rect 20359 776 20425 799
rect 20039 736 20048 776
rect 20088 736 20105 776
rect 20191 736 20212 776
rect 20252 736 20273 776
rect 20359 736 20376 776
rect 20416 736 20425 776
rect 20039 713 20105 736
rect 20191 713 20273 736
rect 20359 713 20425 736
rect 20039 694 20425 713
rect 35159 799 35545 818
rect 35159 776 35225 799
rect 35311 776 35393 799
rect 35479 776 35545 799
rect 35159 736 35168 776
rect 35208 736 35225 776
rect 35311 736 35332 776
rect 35372 736 35393 776
rect 35479 736 35496 776
rect 35536 736 35545 776
rect 35159 713 35225 736
rect 35311 713 35393 736
rect 35479 713 35545 736
rect 35159 694 35545 713
rect 13219 568 13228 608
rect 13268 568 25516 608
rect 25556 568 25565 608
rect 19363 484 19372 524
rect 19412 484 31564 524
rect 31604 484 31613 524
<< via5 >>
rect 4985 9848 5071 9871
rect 5153 9848 5239 9871
rect 4985 9808 5010 9848
rect 5010 9808 5050 9848
rect 5050 9808 5071 9848
rect 5153 9808 5174 9848
rect 5174 9808 5214 9848
rect 5214 9808 5239 9848
rect 4985 9785 5071 9808
rect 5153 9785 5239 9808
rect 20105 9848 20191 9871
rect 20273 9848 20359 9871
rect 20105 9808 20130 9848
rect 20130 9808 20170 9848
rect 20170 9808 20191 9848
rect 20273 9808 20294 9848
rect 20294 9808 20334 9848
rect 20334 9808 20359 9848
rect 20105 9785 20191 9808
rect 20273 9785 20359 9808
rect 35225 9848 35311 9871
rect 35393 9848 35479 9871
rect 35225 9808 35250 9848
rect 35250 9808 35290 9848
rect 35290 9808 35311 9848
rect 35393 9808 35414 9848
rect 35414 9808 35454 9848
rect 35454 9808 35479 9848
rect 35225 9785 35311 9808
rect 35393 9785 35479 9808
rect 3745 9092 3831 9115
rect 3913 9092 3999 9115
rect 3745 9052 3770 9092
rect 3770 9052 3810 9092
rect 3810 9052 3831 9092
rect 3913 9052 3934 9092
rect 3934 9052 3974 9092
rect 3974 9052 3999 9092
rect 3745 9029 3831 9052
rect 3913 9029 3999 9052
rect 18865 9092 18951 9115
rect 19033 9092 19119 9115
rect 33985 9092 34071 9115
rect 34153 9092 34239 9115
rect 18865 9052 18890 9092
rect 18890 9052 18930 9092
rect 18930 9052 18951 9092
rect 19033 9052 19054 9092
rect 19054 9052 19094 9092
rect 19094 9052 19119 9092
rect 33985 9052 34010 9092
rect 34010 9052 34050 9092
rect 34050 9052 34071 9092
rect 34153 9052 34174 9092
rect 34174 9052 34214 9092
rect 34214 9052 34239 9092
rect 18865 9029 18951 9052
rect 19033 9029 19119 9052
rect 33985 9029 34071 9052
rect 34153 9029 34239 9052
rect 4985 8336 5071 8359
rect 5153 8336 5239 8359
rect 4985 8296 5010 8336
rect 5010 8296 5050 8336
rect 5050 8296 5071 8336
rect 5153 8296 5174 8336
rect 5174 8296 5214 8336
rect 5214 8296 5239 8336
rect 4985 8273 5071 8296
rect 5153 8273 5239 8296
rect 20105 8336 20191 8359
rect 20273 8336 20359 8359
rect 20105 8296 20130 8336
rect 20130 8296 20170 8336
rect 20170 8296 20191 8336
rect 20273 8296 20294 8336
rect 20294 8296 20334 8336
rect 20334 8296 20359 8336
rect 20105 8273 20191 8296
rect 20273 8273 20359 8296
rect 35225 8336 35311 8359
rect 35393 8336 35479 8359
rect 35225 8296 35250 8336
rect 35250 8296 35290 8336
rect 35290 8296 35311 8336
rect 35393 8296 35414 8336
rect 35414 8296 35454 8336
rect 35454 8296 35479 8336
rect 35225 8273 35311 8296
rect 35393 8273 35479 8296
rect 3745 7580 3831 7603
rect 3913 7580 3999 7603
rect 3745 7540 3770 7580
rect 3770 7540 3810 7580
rect 3810 7540 3831 7580
rect 3913 7540 3934 7580
rect 3934 7540 3974 7580
rect 3974 7540 3999 7580
rect 3745 7517 3831 7540
rect 3913 7517 3999 7540
rect 18865 7580 18951 7603
rect 19033 7580 19119 7603
rect 18865 7540 18890 7580
rect 18890 7540 18930 7580
rect 18930 7540 18951 7580
rect 19033 7540 19054 7580
rect 19054 7540 19094 7580
rect 19094 7540 19119 7580
rect 18865 7517 18951 7540
rect 19033 7517 19119 7540
rect 33985 7580 34071 7603
rect 34153 7580 34239 7603
rect 33985 7540 34010 7580
rect 34010 7540 34050 7580
rect 34050 7540 34071 7580
rect 34153 7540 34174 7580
rect 34174 7540 34214 7580
rect 34214 7540 34239 7580
rect 33985 7517 34071 7540
rect 34153 7517 34239 7540
rect 4985 6824 5071 6847
rect 5153 6824 5239 6847
rect 4985 6784 5010 6824
rect 5010 6784 5050 6824
rect 5050 6784 5071 6824
rect 5153 6784 5174 6824
rect 5174 6784 5214 6824
rect 5214 6784 5239 6824
rect 4985 6761 5071 6784
rect 5153 6761 5239 6784
rect 20105 6824 20191 6847
rect 20273 6824 20359 6847
rect 20105 6784 20130 6824
rect 20130 6784 20170 6824
rect 20170 6784 20191 6824
rect 20273 6784 20294 6824
rect 20294 6784 20334 6824
rect 20334 6784 20359 6824
rect 20105 6761 20191 6784
rect 20273 6761 20359 6784
rect 35225 6824 35311 6847
rect 35393 6824 35479 6847
rect 35225 6784 35250 6824
rect 35250 6784 35290 6824
rect 35290 6784 35311 6824
rect 35393 6784 35414 6824
rect 35414 6784 35454 6824
rect 35454 6784 35479 6824
rect 35225 6761 35311 6784
rect 35393 6761 35479 6784
rect 3745 6068 3831 6091
rect 3913 6068 3999 6091
rect 3745 6028 3770 6068
rect 3770 6028 3810 6068
rect 3810 6028 3831 6068
rect 3913 6028 3934 6068
rect 3934 6028 3974 6068
rect 3974 6028 3999 6068
rect 3745 6005 3831 6028
rect 3913 6005 3999 6028
rect 18865 6068 18951 6091
rect 19033 6068 19119 6091
rect 18865 6028 18890 6068
rect 18890 6028 18930 6068
rect 18930 6028 18951 6068
rect 19033 6028 19054 6068
rect 19054 6028 19094 6068
rect 19094 6028 19119 6068
rect 18865 6005 18951 6028
rect 19033 6005 19119 6028
rect 33985 6068 34071 6091
rect 34153 6068 34239 6091
rect 33985 6028 34010 6068
rect 34010 6028 34050 6068
rect 34050 6028 34071 6068
rect 34153 6028 34174 6068
rect 34174 6028 34214 6068
rect 34214 6028 34239 6068
rect 33985 6005 34071 6028
rect 34153 6005 34239 6028
rect 4985 5312 5071 5335
rect 5153 5312 5239 5335
rect 4985 5272 5010 5312
rect 5010 5272 5050 5312
rect 5050 5272 5071 5312
rect 5153 5272 5174 5312
rect 5174 5272 5214 5312
rect 5214 5272 5239 5312
rect 4985 5249 5071 5272
rect 5153 5249 5239 5272
rect 20105 5312 20191 5335
rect 20273 5312 20359 5335
rect 20105 5272 20130 5312
rect 20130 5272 20170 5312
rect 20170 5272 20191 5312
rect 20273 5272 20294 5312
rect 20294 5272 20334 5312
rect 20334 5272 20359 5312
rect 20105 5249 20191 5272
rect 20273 5249 20359 5272
rect 35225 5312 35311 5335
rect 35393 5312 35479 5335
rect 35225 5272 35250 5312
rect 35250 5272 35290 5312
rect 35290 5272 35311 5312
rect 35393 5272 35414 5312
rect 35414 5272 35454 5312
rect 35454 5272 35479 5312
rect 35225 5249 35311 5272
rect 35393 5249 35479 5272
rect 3745 4556 3831 4579
rect 3913 4556 3999 4579
rect 3745 4516 3770 4556
rect 3770 4516 3810 4556
rect 3810 4516 3831 4556
rect 3913 4516 3934 4556
rect 3934 4516 3974 4556
rect 3974 4516 3999 4556
rect 3745 4493 3831 4516
rect 3913 4493 3999 4516
rect 18865 4556 18951 4579
rect 19033 4556 19119 4579
rect 18865 4516 18890 4556
rect 18890 4516 18930 4556
rect 18930 4516 18951 4556
rect 19033 4516 19054 4556
rect 19054 4516 19094 4556
rect 19094 4516 19119 4556
rect 18865 4493 18951 4516
rect 19033 4493 19119 4516
rect 33985 4556 34071 4579
rect 34153 4556 34239 4579
rect 33985 4516 34010 4556
rect 34010 4516 34050 4556
rect 34050 4516 34071 4556
rect 34153 4516 34174 4556
rect 34174 4516 34214 4556
rect 34214 4516 34239 4556
rect 33985 4493 34071 4516
rect 34153 4493 34239 4516
rect 4985 3800 5071 3823
rect 5153 3800 5239 3823
rect 20105 3800 20191 3823
rect 20273 3800 20359 3823
rect 4985 3760 5010 3800
rect 5010 3760 5050 3800
rect 5050 3760 5071 3800
rect 5153 3760 5174 3800
rect 5174 3760 5214 3800
rect 5214 3760 5239 3800
rect 20105 3760 20130 3800
rect 20130 3760 20170 3800
rect 20170 3760 20191 3800
rect 20273 3760 20294 3800
rect 20294 3760 20334 3800
rect 20334 3760 20359 3800
rect 4985 3737 5071 3760
rect 5153 3737 5239 3760
rect 20105 3737 20191 3760
rect 20273 3737 20359 3760
rect 35225 3800 35311 3823
rect 35393 3800 35479 3823
rect 35225 3760 35250 3800
rect 35250 3760 35290 3800
rect 35290 3760 35311 3800
rect 35393 3760 35414 3800
rect 35414 3760 35454 3800
rect 35454 3760 35479 3800
rect 35225 3737 35311 3760
rect 35393 3737 35479 3760
rect 3745 3044 3831 3067
rect 3913 3044 3999 3067
rect 3745 3004 3770 3044
rect 3770 3004 3810 3044
rect 3810 3004 3831 3044
rect 3913 3004 3934 3044
rect 3934 3004 3974 3044
rect 3974 3004 3999 3044
rect 3745 2981 3831 3004
rect 3913 2981 3999 3004
rect 18865 3044 18951 3067
rect 19033 3044 19119 3067
rect 18865 3004 18890 3044
rect 18890 3004 18930 3044
rect 18930 3004 18951 3044
rect 19033 3004 19054 3044
rect 19054 3004 19094 3044
rect 19094 3004 19119 3044
rect 18865 2981 18951 3004
rect 19033 2981 19119 3004
rect 33985 3044 34071 3067
rect 34153 3044 34239 3067
rect 33985 3004 34010 3044
rect 34010 3004 34050 3044
rect 34050 3004 34071 3044
rect 34153 3004 34174 3044
rect 34174 3004 34214 3044
rect 34214 3004 34239 3044
rect 33985 2981 34071 3004
rect 34153 2981 34239 3004
rect 4985 2288 5071 2311
rect 5153 2288 5239 2311
rect 4985 2248 5010 2288
rect 5010 2248 5050 2288
rect 5050 2248 5071 2288
rect 5153 2248 5174 2288
rect 5174 2248 5214 2288
rect 5214 2248 5239 2288
rect 4985 2225 5071 2248
rect 5153 2225 5239 2248
rect 20105 2288 20191 2311
rect 20273 2288 20359 2311
rect 20105 2248 20130 2288
rect 20130 2248 20170 2288
rect 20170 2248 20191 2288
rect 20273 2248 20294 2288
rect 20294 2248 20334 2288
rect 20334 2248 20359 2288
rect 20105 2225 20191 2248
rect 20273 2225 20359 2248
rect 35225 2288 35311 2311
rect 35393 2288 35479 2311
rect 35225 2248 35250 2288
rect 35250 2248 35290 2288
rect 35290 2248 35311 2288
rect 35393 2248 35414 2288
rect 35414 2248 35454 2288
rect 35454 2248 35479 2288
rect 35225 2225 35311 2248
rect 35393 2225 35479 2248
rect 3745 1532 3831 1555
rect 3913 1532 3999 1555
rect 3745 1492 3770 1532
rect 3770 1492 3810 1532
rect 3810 1492 3831 1532
rect 3913 1492 3934 1532
rect 3934 1492 3974 1532
rect 3974 1492 3999 1532
rect 3745 1469 3831 1492
rect 3913 1469 3999 1492
rect 18865 1532 18951 1555
rect 19033 1532 19119 1555
rect 18865 1492 18890 1532
rect 18890 1492 18930 1532
rect 18930 1492 18951 1532
rect 19033 1492 19054 1532
rect 19054 1492 19094 1532
rect 19094 1492 19119 1532
rect 18865 1469 18951 1492
rect 19033 1469 19119 1492
rect 33985 1532 34071 1555
rect 34153 1532 34239 1555
rect 33985 1492 34010 1532
rect 34010 1492 34050 1532
rect 34050 1492 34071 1532
rect 34153 1492 34174 1532
rect 34174 1492 34214 1532
rect 34214 1492 34239 1532
rect 33985 1469 34071 1492
rect 34153 1469 34239 1492
rect 4985 776 5071 799
rect 5153 776 5239 799
rect 4985 736 5010 776
rect 5010 736 5050 776
rect 5050 736 5071 776
rect 5153 736 5174 776
rect 5174 736 5214 776
rect 5214 736 5239 776
rect 4985 713 5071 736
rect 5153 713 5239 736
rect 20105 776 20191 799
rect 20273 776 20359 799
rect 20105 736 20130 776
rect 20130 736 20170 776
rect 20170 736 20191 776
rect 20273 736 20294 776
rect 20294 736 20334 776
rect 20334 736 20359 776
rect 20105 713 20191 736
rect 20273 713 20359 736
rect 35225 776 35311 799
rect 35393 776 35479 799
rect 35225 736 35250 776
rect 35250 736 35290 776
rect 35290 736 35311 776
rect 35393 736 35414 776
rect 35414 736 35454 776
rect 35454 736 35479 776
rect 35225 713 35311 736
rect 35393 713 35479 736
<< metal6 >>
rect 3652 9115 4092 10752
rect 3652 9029 3745 9115
rect 3831 9029 3913 9115
rect 3999 9029 4092 9115
rect 3652 7603 4092 9029
rect 3652 7517 3745 7603
rect 3831 7517 3913 7603
rect 3999 7517 4092 7603
rect 3652 6091 4092 7517
rect 3652 6005 3745 6091
rect 3831 6005 3913 6091
rect 3999 6005 4092 6091
rect 3652 4579 4092 6005
rect 3652 4493 3745 4579
rect 3831 4493 3913 4579
rect 3999 4493 4092 4579
rect 3652 3067 4092 4493
rect 3652 2981 3745 3067
rect 3831 2981 3913 3067
rect 3999 2981 4092 3067
rect 3652 1555 4092 2981
rect 3652 1469 3745 1555
rect 3831 1469 3913 1555
rect 3999 1469 4092 1555
rect 3652 0 4092 1469
rect 4892 9871 5332 10752
rect 4892 9785 4985 9871
rect 5071 9785 5153 9871
rect 5239 9785 5332 9871
rect 4892 8359 5332 9785
rect 4892 8273 4985 8359
rect 5071 8273 5153 8359
rect 5239 8273 5332 8359
rect 4892 6847 5332 8273
rect 4892 6761 4985 6847
rect 5071 6761 5153 6847
rect 5239 6761 5332 6847
rect 4892 5335 5332 6761
rect 4892 5249 4985 5335
rect 5071 5249 5153 5335
rect 5239 5249 5332 5335
rect 4892 3823 5332 5249
rect 4892 3737 4985 3823
rect 5071 3737 5153 3823
rect 5239 3737 5332 3823
rect 4892 2311 5332 3737
rect 4892 2225 4985 2311
rect 5071 2225 5153 2311
rect 5239 2225 5332 2311
rect 4892 799 5332 2225
rect 4892 713 4985 799
rect 5071 713 5153 799
rect 5239 713 5332 799
rect 4892 0 5332 713
rect 18772 9115 19212 10752
rect 18772 9029 18865 9115
rect 18951 9029 19033 9115
rect 19119 9029 19212 9115
rect 18772 7603 19212 9029
rect 18772 7517 18865 7603
rect 18951 7517 19033 7603
rect 19119 7517 19212 7603
rect 18772 6091 19212 7517
rect 18772 6005 18865 6091
rect 18951 6005 19033 6091
rect 19119 6005 19212 6091
rect 18772 4579 19212 6005
rect 18772 4493 18865 4579
rect 18951 4493 19033 4579
rect 19119 4493 19212 4579
rect 18772 3067 19212 4493
rect 18772 2981 18865 3067
rect 18951 2981 19033 3067
rect 19119 2981 19212 3067
rect 18772 1555 19212 2981
rect 18772 1469 18865 1555
rect 18951 1469 19033 1555
rect 19119 1469 19212 1555
rect 18772 0 19212 1469
rect 20012 9871 20452 10752
rect 20012 9785 20105 9871
rect 20191 9785 20273 9871
rect 20359 9785 20452 9871
rect 20012 8359 20452 9785
rect 20012 8273 20105 8359
rect 20191 8273 20273 8359
rect 20359 8273 20452 8359
rect 20012 6847 20452 8273
rect 20012 6761 20105 6847
rect 20191 6761 20273 6847
rect 20359 6761 20452 6847
rect 20012 5335 20452 6761
rect 20012 5249 20105 5335
rect 20191 5249 20273 5335
rect 20359 5249 20452 5335
rect 20012 3823 20452 5249
rect 20012 3737 20105 3823
rect 20191 3737 20273 3823
rect 20359 3737 20452 3823
rect 20012 2311 20452 3737
rect 20012 2225 20105 2311
rect 20191 2225 20273 2311
rect 20359 2225 20452 2311
rect 20012 799 20452 2225
rect 20012 713 20105 799
rect 20191 713 20273 799
rect 20359 713 20452 799
rect 20012 0 20452 713
rect 33892 9115 34332 10752
rect 33892 9029 33985 9115
rect 34071 9029 34153 9115
rect 34239 9029 34332 9115
rect 33892 7603 34332 9029
rect 33892 7517 33985 7603
rect 34071 7517 34153 7603
rect 34239 7517 34332 7603
rect 33892 6091 34332 7517
rect 33892 6005 33985 6091
rect 34071 6005 34153 6091
rect 34239 6005 34332 6091
rect 33892 4579 34332 6005
rect 33892 4493 33985 4579
rect 34071 4493 34153 4579
rect 34239 4493 34332 4579
rect 33892 3067 34332 4493
rect 33892 2981 33985 3067
rect 34071 2981 34153 3067
rect 34239 2981 34332 3067
rect 33892 1555 34332 2981
rect 33892 1469 33985 1555
rect 34071 1469 34153 1555
rect 34239 1469 34332 1555
rect 33892 0 34332 1469
rect 35132 9871 35572 10752
rect 35132 9785 35225 9871
rect 35311 9785 35393 9871
rect 35479 9785 35572 9871
rect 35132 8359 35572 9785
rect 35132 8273 35225 8359
rect 35311 8273 35393 8359
rect 35479 8273 35572 8359
rect 35132 6847 35572 8273
rect 35132 6761 35225 6847
rect 35311 6761 35393 6847
rect 35479 6761 35572 6847
rect 35132 5335 35572 6761
rect 35132 5249 35225 5335
rect 35311 5249 35393 5335
rect 35479 5249 35572 5335
rect 35132 3823 35572 5249
rect 35132 3737 35225 3823
rect 35311 3737 35393 3823
rect 35479 3737 35572 3823
rect 35132 2311 35572 3737
rect 35132 2225 35225 2311
rect 35311 2225 35393 2311
rect 35479 2225 35572 2311
rect 35132 799 35572 2225
rect 35132 713 35225 799
rect 35311 713 35393 799
rect 35479 713 35572 799
rect 35132 0 35572 713
use sg13g2_inv_1  _083_
timestamp 1676382929
transform -1 0 6432 0 1 2268
box -48 -56 336 834
use sg13g2_inv_1  _084_
timestamp 1676382929
transform 1 0 8736 0 -1 3780
box -48 -56 336 834
use sg13g2_inv_1  _085_
timestamp 1676382929
transform -1 0 10176 0 1 6804
box -48 -56 336 834
use sg13g2_inv_1  _086_
timestamp 1676382929
transform -1 0 12384 0 1 2268
box -48 -56 336 834
use sg13g2_mux4_1  _087_
timestamp 1677257233
transform 1 0 26496 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _088_
timestamp 1677257233
transform 1 0 18720 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _089_
timestamp 1677257233
transform 1 0 27648 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _090_
timestamp 1677257233
transform 1 0 21120 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _091_
timestamp 1677257233
transform 1 0 28992 0 -1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _092_
timestamp 1677257233
transform 1 0 27360 0 1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _093_
timestamp 1677257233
transform 1 0 20544 0 1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _094_
timestamp 1677257233
transform -1 0 21024 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _095_
timestamp 1677257233
transform -1 0 15936 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _096_
timestamp 1677257233
transform -1 0 13056 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _097_
timestamp 1677257233
transform -1 0 5088 0 1 2268
box -48 -56 2064 834
use sg13g2_o21ai_1  _098_
timestamp 1685175443
transform -1 0 1824 0 1 756
box -48 -56 538 834
use sg13g2_nor2_1  _099_
timestamp 1676627187
transform 1 0 1248 0 1 6804
box -48 -56 432 834
use sg13g2_nand2_1  _100_
timestamp 1676557249
transform 1 0 5280 0 -1 6804
box -48 -56 432 834
use sg13g2_nand3_1  _101_
timestamp 1683988354
transform -1 0 8736 0 -1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  _102_
timestamp 1685175443
transform 1 0 2880 0 1 3780
box -48 -56 538 834
use sg13g2_mux4_1  _103_
timestamp 1677257233
transform 1 0 2784 0 -1 5292
box -48 -56 2064 834
use sg13g2_o21ai_1  _104_
timestamp 1685175443
transform 1 0 3168 0 1 5292
box -48 -56 538 834
use sg13g2_nor2_1  _105_
timestamp 1676627187
transform -1 0 7104 0 -1 5292
box -48 -56 432 834
use sg13g2_nand2_1  _106_
timestamp 1676557249
transform -1 0 4896 0 -1 3780
box -48 -56 432 834
use sg13g2_nand3_1  _107_
timestamp 1683988354
transform -1 0 5472 0 1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  _108_
timestamp 1685175443
transform 1 0 4608 0 1 5292
box -48 -56 538 834
use sg13g2_nand2b_1  _109_
timestamp 1676567195
transform -1 0 4320 0 1 6804
box -48 -56 528 834
use sg13g2_mux4_1  _110_
timestamp 1677257233
transform 1 0 2784 0 -1 6804
box -48 -56 2064 834
use sg13g2_o21ai_1  _111_
timestamp 1685175443
transform 1 0 3360 0 1 6804
box -48 -56 538 834
use sg13g2_o21ai_1  _112_
timestamp 1685175443
transform 1 0 3648 0 1 5292
box -48 -56 538 834
use sg13g2_nand2b_1  _113_
timestamp 1676567195
transform 1 0 4128 0 1 5292
box -48 -56 528 834
use sg13g2_o21ai_1  _114_
timestamp 1685175443
transform 1 0 4800 0 -1 6804
box -48 -56 538 834
use sg13g2_nand2b_1  _115_
timestamp 1676567195
transform -1 0 2688 0 1 8316
box -48 -56 528 834
use sg13g2_mux4_1  _116_
timestamp 1677257233
transform 1 0 2688 0 1 8316
box -48 -56 2064 834
use sg13g2_o21ai_1  _117_
timestamp 1685175443
transform -1 0 5280 0 -1 9828
box -48 -56 538 834
use sg13g2_o21ai_1  _118_
timestamp 1685175443
transform -1 0 2208 0 1 8316
box -48 -56 538 834
use sg13g2_nand2b_1  _119_
timestamp 1676567195
transform 1 0 3744 0 -1 8316
box -48 -56 528 834
use sg13g2_o21ai_1  _120_
timestamp 1685175443
transform 1 0 4224 0 -1 8316
box -48 -56 538 834
use sg13g2_nand2_1  _121_
timestamp 1676557249
transform 1 0 9024 0 -1 8316
box -48 -56 432 834
use sg13g2_nand2b_1  _122_
timestamp 1676567195
transform 1 0 7296 0 -1 9828
box -48 -56 528 834
use sg13g2_a21oi_1  _123_
timestamp 1683973020
transform 1 0 7296 0 1 6804
box -48 -56 528 834
use sg13g2_nor2b_1  _124_
timestamp 1685181386
transform 1 0 6624 0 -1 6804
box -54 -56 528 834
use sg13g2_o21ai_1  _125_
timestamp 1685175443
transform 1 0 6144 0 -1 6804
box -48 -56 538 834
use sg13g2_o21ai_1  _126_
timestamp 1685175443
transform 1 0 8064 0 -1 6804
box -48 -56 538 834
use sg13g2_mux2_1  _127_
timestamp 1677247768
transform 1 0 6144 0 1 6804
box -48 -56 1008 834
use sg13g2_or2_1  _128_
timestamp 1684236171
transform 1 0 6048 0 -1 9828
box -48 -56 528 834
use sg13g2_a21oi_1  _129_
timestamp 1683973020
transform -1 0 6144 0 -1 6804
box -48 -56 528 834
use sg13g2_a221oi_1  _130_
timestamp 1685197497
transform 1 0 6528 0 -1 9828
box -48 -56 816 834
use sg13g2_o21ai_1  _131_
timestamp 1685175443
transform 1 0 8064 0 -1 9828
box -48 -56 538 834
use sg13g2_mux4_1  _132_
timestamp 1677257233
transform 1 0 6624 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _133_
timestamp 1677257233
transform 1 0 6528 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux2_1  _134_
timestamp 1677247768
transform 1 0 8640 0 1 8316
box -48 -56 1008 834
use sg13g2_nand2b_1  _135_
timestamp 1676567195
transform 1 0 8640 0 -1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _136_
timestamp 1685175443
transform 1 0 8544 0 -1 8316
box -48 -56 538 834
use sg13g2_mux2_1  _137_
timestamp 1677247768
transform 1 0 9120 0 -1 5292
box -48 -56 1008 834
use sg13g2_mux2_1  _138_
timestamp 1677247768
transform -1 0 9888 0 1 3780
box -48 -56 1008 834
use sg13g2_nand2b_1  _139_
timestamp 1676567195
transform 1 0 8448 0 1 5292
box -48 -56 528 834
use sg13g2_a21oi_1  _140_
timestamp 1683973020
transform 1 0 9408 0 1 6804
box -48 -56 528 834
use sg13g2_mux2_1  _141_
timestamp 1677247768
transform 1 0 7968 0 1 3780
box -48 -56 1008 834
use sg13g2_nand2b_1  _142_
timestamp 1676567195
transform 1 0 10080 0 -1 5292
box -48 -56 528 834
use sg13g2_mux2_1  _143_
timestamp 1677247768
transform 1 0 8928 0 1 5292
box -48 -56 1008 834
use sg13g2_a21oi_1  _144_
timestamp 1683973020
transform 1 0 10368 0 -1 6804
box -48 -56 528 834
use sg13g2_a221oi_1  _145_
timestamp 1685197497
transform -1 0 10656 0 1 5292
box -48 -56 816 834
use sg13g2_mux2_1  _146_
timestamp 1677247768
transform 1 0 7008 0 1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _147_
timestamp 1677247768
transform 1 0 6048 0 1 3780
box -48 -56 1008 834
use sg13g2_mux2_1  _148_
timestamp 1677247768
transform 1 0 7104 0 -1 6804
box -48 -56 1008 834
use sg13g2_mux2_1  _149_
timestamp 1677247768
transform 1 0 6816 0 -1 3780
box -48 -56 1008 834
use sg13g2_mux4_1  _150_
timestamp 1677257233
transform 1 0 7104 0 -1 5292
box -48 -56 2064 834
use sg13g2_a21o_1  _151_
timestamp 1677175127
transform -1 0 11328 0 1 5292
box -48 -56 720 834
use sg13g2_mux4_1  _152_
timestamp 1677257233
transform 1 0 10080 0 1 2268
box -48 -56 2064 834
use sg13g2_mux2_1  _153_
timestamp 1677247768
transform -1 0 12480 0 -1 2268
box -48 -56 1008 834
use sg13g2_nor2b_1  _154_
timestamp 1685181386
transform 1 0 9984 0 1 3780
box -54 -56 528 834
use sg13g2_o21ai_1  _155_
timestamp 1685175443
transform -1 0 13248 0 1 756
box -48 -56 538 834
use sg13g2_o21ai_1  _156_
timestamp 1685175443
transform -1 0 12768 0 1 756
box -48 -56 538 834
use sg13g2_a21oi_1  _157_
timestamp 1683973020
transform -1 0 11808 0 1 756
box -48 -56 528 834
use sg13g2_o21ai_1  _158_
timestamp 1685175443
transform 1 0 11040 0 -1 2268
box -48 -56 538 834
use sg13g2_mux4_1  _159_
timestamp 1677257233
transform 1 0 9024 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _160_
timestamp 1677257233
transform 1 0 9024 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux2_1  _161_
timestamp 1677247768
transform 1 0 11040 0 -1 3780
box -48 -56 1008 834
use sg13g2_nand2b_1  _162_
timestamp 1676567195
transform 1 0 12000 0 -1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  _163_
timestamp 1685175443
transform 1 0 11808 0 1 756
box -48 -56 538 834
use sg13g2_mux2_1  _164_
timestamp 1677247768
transform 1 0 5184 0 1 2268
box -48 -56 1008 834
use sg13g2_or2_1  _165_
timestamp 1684236171
transform 1 0 5376 0 -1 3780
box -48 -56 528 834
use sg13g2_a21oi_1  _166_
timestamp 1683973020
transform 1 0 5856 0 -1 3780
box -48 -56 528 834
use sg13g2_a221oi_1  _167_
timestamp 1685197497
transform 1 0 5664 0 -1 2268
box -48 -56 816 834
use sg13g2_nor2b_1  _168_
timestamp 1685181386
transform 1 0 6336 0 -1 3780
box -54 -56 528 834
use sg13g2_o21ai_1  _169_
timestamp 1685175443
transform 1 0 6144 0 1 756
box -48 -56 538 834
use sg13g2_nand2_1  _170_
timestamp 1676557249
transform -1 0 3456 0 -1 2268
box -48 -56 432 834
use sg13g2_nand2b_1  _171_
timestamp 1676567195
transform 1 0 4896 0 -1 3780
box -48 -56 528 834
use sg13g2_a21oi_1  _172_
timestamp 1683973020
transform -1 0 5952 0 1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  _173_
timestamp 1685175443
transform 1 0 6624 0 1 756
box -48 -56 538 834
use sg13g2_o21ai_1  _174_
timestamp 1685175443
transform -1 0 3936 0 -1 2268
box -48 -56 538 834
use sg13g2_mux4_1  _175_
timestamp 1677257233
transform 1 0 6624 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _176_
timestamp 1677257233
transform 1 0 6432 0 1 2268
box -48 -56 2064 834
use sg13g2_mux2_1  _177_
timestamp 1677247768
transform -1 0 8064 0 1 756
box -48 -56 1008 834
use sg13g2_nand2b_1  _178_
timestamp 1676567195
transform 1 0 5664 0 1 756
box -48 -56 528 834
use sg13g2_o21ai_1  _179_
timestamp 1685175443
transform 1 0 7776 0 -1 3780
box -48 -56 538 834
use sg13g2_mux4_1  _180_
timestamp 1677257233
transform 1 0 18528 0 1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _181_
timestamp 1677257233
transform 1 0 16416 0 1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _182_
timestamp 1677257233
transform 1 0 37632 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _183_
timestamp 1677257233
transform 1 0 16224 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _184_
timestamp 1677257233
transform 1 0 38784 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _185_
timestamp 1677257233
transform 1 0 23808 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _186_
timestamp 1677257233
transform 1 0 23712 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _187_
timestamp 1677257233
transform 1 0 38688 0 1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _188_
timestamp 1677257233
transform 1 0 12192 0 -1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _189_
timestamp 1677257233
transform 1 0 13152 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _190_
timestamp 1677257233
transform 1 0 21216 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _191_
timestamp 1677257233
transform 1 0 14016 0 1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _192_
timestamp 1677257233
transform 1 0 37536 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _193_
timestamp 1677257233
transform 1 0 14016 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _194_
timestamp 1677257233
transform 1 0 38880 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _195_
timestamp 1677257233
transform 1 0 24384 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _196_
timestamp 1677257233
transform 1 0 24384 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _197_
timestamp 1677257233
transform 1 0 14592 0 -1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _198_
timestamp 1677257233
transform 1 0 33120 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _199_
timestamp 1677257233
transform 1 0 21600 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _200_
timestamp 1677257233
transform 1 0 35616 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _201_
timestamp 1677257233
transform 1 0 34944 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _202_
timestamp 1677257233
transform 1 0 31296 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _203_
timestamp 1677257233
transform 1 0 25728 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _204_
timestamp 1677257233
transform 1 0 32544 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _205_
timestamp 1677257233
transform 1 0 17952 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _206_
timestamp 1677257233
transform 1 0 35328 0 -1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _207_
timestamp 1677257233
transform 1 0 32640 0 1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _208_
timestamp 1677257233
transform 1 0 35808 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _209_
timestamp 1677257233
transform 1 0 32832 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _210_
timestamp 1677257233
transform 1 0 30528 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _211_
timestamp 1677257233
transform 1 0 28032 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _212_
timestamp 1677257233
transform 1 0 23136 0 1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _213_
timestamp 1677257233
transform -1 0 18720 0 -1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _214_
timestamp 1677257233
transform 1 0 26688 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _215_
timestamp 1677257233
transform 1 0 18240 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _216_
timestamp 1677257233
transform -1 0 32256 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _217_
timestamp 1677257233
transform 1 0 21024 0 -1 9828
box -48 -56 2064 834
use sg13g2_mux4_1  _218_
timestamp 1677257233
transform 1 0 29664 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _219_
timestamp 1677257233
transform 1 0 27648 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _220_
timestamp 1677257233
transform 1 0 23616 0 -1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _221_
timestamp 1677257233
transform 1 0 15840 0 -1 6804
box -48 -56 2064 834
use sg13g2_dlhq_1  _222_
timestamp 1678805552
transform -1 0 12576 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _223_
timestamp 1678805552
transform 1 0 9408 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _224_
timestamp 1678805552
transform 1 0 12288 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _225_
timestamp 1678805552
transform -1 0 15552 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _226_
timestamp 1678805552
transform 1 0 17760 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _227_
timestamp 1678805552
transform 1 0 18336 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _228_
timestamp 1678805552
transform 1 0 19488 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _229_
timestamp 1678805552
transform 1 0 21024 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _230_
timestamp 1678805552
transform 1 0 26208 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _231_
timestamp 1678805552
transform -1 0 31680 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _232_
timestamp 1678805552
transform -1 0 30144 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _233_
timestamp 1678805552
transform -1 0 31968 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _234_
timestamp 1678805552
transform 1 0 19680 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _235_
timestamp 1678805552
transform 1 0 21312 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _236_
timestamp 1678805552
transform -1 0 29280 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _237_
timestamp 1678805552
transform -1 0 30336 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _238_
timestamp 1678805552
transform 1 0 17376 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _239_
timestamp 1678805552
transform 1 0 19104 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _240_
timestamp 1678805552
transform 1 0 25440 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _241_
timestamp 1678805552
transform 1 0 27072 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _242_
timestamp 1678805552
transform 1 0 14208 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _243_
timestamp 1678805552
transform 1 0 15840 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _244_
timestamp 1678805552
transform 1 0 22464 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _245_
timestamp 1678805552
transform -1 0 27264 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _246_
timestamp 1678805552
transform -1 0 30912 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _247_
timestamp 1678805552
transform 1 0 26016 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _248_
timestamp 1678805552
transform 1 0 30144 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _249_
timestamp 1678805552
transform 1 0 28704 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _250_
timestamp 1678805552
transform 1 0 20928 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _251_
timestamp 1678805552
transform 1 0 19488 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _252_
timestamp 1678805552
transform -1 0 32544 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _253_
timestamp 1678805552
transform 1 0 29280 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _254_
timestamp 1678805552
transform 1 0 17856 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _255_
timestamp 1678805552
transform 1 0 16224 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _256_
timestamp 1678805552
transform 1 0 25344 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _257_
timestamp 1678805552
transform -1 0 29376 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _258_
timestamp 1678805552
transform 1 0 15840 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _259_
timestamp 1678805552
transform -1 0 18336 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _260_
timestamp 1678805552
transform 1 0 21120 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _261_
timestamp 1678805552
transform -1 0 26208 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _262_
timestamp 1678805552
transform -1 0 31104 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _263_
timestamp 1678805552
transform -1 0 29472 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _264_
timestamp 1678805552
transform -1 0 33600 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _265_
timestamp 1678805552
transform -1 0 31584 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _266_
timestamp 1678805552
transform 1 0 33408 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _267_
timestamp 1678805552
transform 1 0 31776 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _268_
timestamp 1678805552
transform 1 0 36096 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _269_
timestamp 1678805552
transform 1 0 34848 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _270_
timestamp 1678805552
transform 1 0 31680 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _271_
timestamp 1678805552
transform 1 0 33312 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _272_
timestamp 1678805552
transform 1 0 34176 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _273_
timestamp 1678805552
transform -1 0 38976 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _274_
timestamp 1678805552
transform 1 0 16416 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _275_
timestamp 1678805552
transform 1 0 18048 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _276_
timestamp 1678805552
transform 1 0 33216 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _277_
timestamp 1678805552
transform 1 0 31200 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _278_
timestamp 1678805552
transform 1 0 26016 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _279_
timestamp 1678805552
transform 1 0 24672 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _280_
timestamp 1678805552
transform -1 0 35040 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _281_
timestamp 1678805552
transform -1 0 33408 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _282_
timestamp 1678805552
transform 1 0 33984 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _283_
timestamp 1678805552
transform 1 0 35520 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _284_
timestamp 1678805552
transform -1 0 37248 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _285_
timestamp 1678805552
transform 1 0 36000 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _286_
timestamp 1678805552
transform 1 0 19392 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _287_
timestamp 1678805552
transform -1 0 24672 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _288_
timestamp 1678805552
transform -1 0 34176 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _289_
timestamp 1678805552
transform -1 0 35808 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _290_
timestamp 1678805552
transform 1 0 12384 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _291_
timestamp 1678805552
transform 1 0 14688 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _292_
timestamp 1678805552
transform 1 0 22944 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _293_
timestamp 1678805552
transform -1 0 28032 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _294_
timestamp 1678805552
transform 1 0 22752 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _295_
timestamp 1678805552
transform 1 0 25152 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _296_
timestamp 1678805552
transform -1 0 41472 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _297_
timestamp 1678805552
transform 1 0 40128 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _298_
timestamp 1678805552
transform 1 0 12480 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _299_
timestamp 1678805552
transform 1 0 13920 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _300_
timestamp 1678805552
transform 1 0 36480 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _301_
timestamp 1678805552
transform 1 0 38208 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _302_
timestamp 1678805552
transform 1 0 12576 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _303_
timestamp 1678805552
transform 1 0 13920 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _304_
timestamp 1678805552
transform 1 0 19968 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _305_
timestamp 1678805552
transform 1 0 21600 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _306_
timestamp 1678805552
transform 1 0 12576 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _307_
timestamp 1678805552
transform 1 0 10944 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _308_
timestamp 1678805552
transform 1 0 10560 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _309_
timestamp 1678805552
transform 1 0 12096 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _310_
timestamp 1678805552
transform -1 0 39744 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _311_
timestamp 1678805552
transform 1 0 39456 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _312_
timestamp 1678805552
transform 1 0 22560 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _313_
timestamp 1678805552
transform 1 0 24000 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _314_
timestamp 1678805552
transform 1 0 22176 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _315_
timestamp 1678805552
transform 1 0 24288 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _316_
timestamp 1678805552
transform -1 0 41280 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _317_
timestamp 1678805552
transform 1 0 39744 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _318_
timestamp 1678805552
transform 1 0 16704 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _319_
timestamp 1678805552
transform 1 0 15072 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _320_
timestamp 1678805552
transform -1 0 39264 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _321_
timestamp 1678805552
transform 1 0 39264 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _322_
timestamp 1678805552
transform 1 0 14496 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _323_
timestamp 1678805552
transform 1 0 16128 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _324_
timestamp 1678805552
transform 1 0 19392 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _325_
timestamp 1678805552
transform 1 0 17568 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _326_
timestamp 1678805552
transform 1 0 1824 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _327_
timestamp 1678805552
transform 1 0 2880 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _328_
timestamp 1678805552
transform 1 0 3744 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _329_
timestamp 1678805552
transform -1 0 5568 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _330_
timestamp 1678805552
transform 1 0 1248 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _331_
timestamp 1678805552
transform 1 0 1440 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _332_
timestamp 1678805552
transform 1 0 1440 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _333_
timestamp 1678805552
transform 1 0 8448 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _334_
timestamp 1678805552
transform 1 0 8064 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _335_
timestamp 1678805552
transform 1 0 9696 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _336_
timestamp 1678805552
transform 1 0 10464 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _337_
timestamp 1678805552
transform 1 0 1248 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _338_
timestamp 1678805552
transform 1 0 1152 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _339_
timestamp 1678805552
transform 1 0 3360 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _340_
timestamp 1678805552
transform 1 0 5088 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _341_
timestamp 1678805552
transform 1 0 6720 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _342_
timestamp 1678805552
transform 1 0 5088 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _343_
timestamp 1678805552
transform 1 0 8736 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _344_
timestamp 1678805552
transform 1 0 1248 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _345_
timestamp 1678805552
transform 1 0 1632 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _346_
timestamp 1678805552
transform 1 0 1152 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _347_
timestamp 1678805552
transform 1 0 4512 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _348_
timestamp 1678805552
transform 1 0 4704 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _349_
timestamp 1678805552
transform 1 0 4704 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _350_
timestamp 1678805552
transform -1 0 9408 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _351_
timestamp 1678805552
transform -1 0 4800 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _352_
timestamp 1678805552
transform 1 0 1536 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _353_
timestamp 1678805552
transform 1 0 1824 0 -1 8316
box -50 -56 1692 834
use sg13g2_dfrbpq_1  _354_
timestamp 1746535128
transform 1 0 33600 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _355_
timestamp 1746535128
transform -1 0 40128 0 1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _356_
timestamp 1746535128
transform 1 0 36480 0 -1 2268
box -48 -56 2640 834
use sg13g2_dfrbpq_1  _357_
timestamp 1746535128
transform -1 0 39360 0 1 756
box -48 -56 2640 834
use sg13g2_tiehi  _358_
timestamp 1680000651
transform -1 0 40512 0 1 756
box -48 -56 432 834
use sg13g2_tiehi  _359_
timestamp 1680000651
transform -1 0 41856 0 -1 3780
box -48 -56 432 834
use sg13g2_tiehi  _360_
timestamp 1680000651
transform -1 0 40896 0 1 756
box -48 -56 432 834
use sg13g2_tiehi  _361_
timestamp 1680000651
transform -1 0 41664 0 -1 9828
box -48 -56 432 834
use sg13g2_tielo  _362_
timestamp 1680000637
transform -1 0 20640 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _363_
timestamp 1676381911
transform 1 0 37536 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _364_
timestamp 1676381911
transform 1 0 38208 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _365_
timestamp 1676381911
transform 1 0 36480 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _366_
timestamp 1676381911
transform 1 0 35136 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _367_
timestamp 1676381911
transform 1 0 35712 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _368_
timestamp 1676381911
transform 1 0 40896 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _369_
timestamp 1676381911
transform 1 0 26976 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _370_
timestamp 1676381911
transform 1 0 24288 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _371_
timestamp 1676381911
transform 1 0 27360 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _372_
timestamp 1676381911
transform 1 0 24672 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _373_
timestamp 1676381911
transform 1 0 25056 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _374_
timestamp 1676381911
transform 1 0 31680 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _375_
timestamp 1676381911
transform 1 0 29760 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _376_
timestamp 1676381911
transform 1 0 32064 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _377_
timestamp 1676381911
transform 1 0 41280 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _378_
timestamp 1676381911
transform 1 0 41280 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _379_
timestamp 1676381911
transform 1 0 41088 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _380_
timestamp 1676381911
transform 1 0 41184 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _381_
timestamp 1676381911
transform 1 0 40800 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _382_
timestamp 1676381911
transform 1 0 41184 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _383_
timestamp 1676381911
transform 1 0 40800 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _384_
timestamp 1676381911
transform 1 0 41376 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _385_
timestamp 1676381911
transform 1 0 40800 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _386_
timestamp 1676381911
transform 1 0 41184 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _387_
timestamp 1676381911
transform 1 0 41280 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _388_
timestamp 1676381911
transform 1 0 40896 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _389_
timestamp 1676381911
transform 1 0 39744 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _390_
timestamp 1676381911
transform 1 0 37632 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _391_
timestamp 1676381911
transform 1 0 39072 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _392_
timestamp 1676381911
transform 1 0 38304 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _393_
timestamp 1676381911
transform 1 0 37920 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _394_
timestamp 1676381911
transform 1 0 37152 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _395_
timestamp 1676381911
transform 1 0 26016 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _396_
timestamp 1676381911
transform 1 0 29760 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _397_
timestamp 1676381911
transform -1 0 30720 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _398_
timestamp 1676381911
transform -1 0 31104 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _399_
timestamp 1676381911
transform 1 0 29376 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _400_
timestamp 1676381911
transform -1 0 32736 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _401_
timestamp 1676381911
transform -1 0 33120 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _402_
timestamp 1676381911
transform -1 0 31968 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _403_
timestamp 1676381911
transform -1 0 35328 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _404_
timestamp 1676381911
transform -1 0 32352 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _405_
timestamp 1676381911
transform 1 0 30144 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _406_
timestamp 1676381911
transform -1 0 32832 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _407_
timestamp 1676381911
transform -1 0 33984 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _408_
timestamp 1676381911
transform -1 0 37248 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _409_
timestamp 1676381911
transform -1 0 40128 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _410_
timestamp 1676381911
transform -1 0 41280 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _411_
timestamp 1676381911
transform -1 0 39744 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _412_
timestamp 1676381911
transform -1 0 35712 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _413_
timestamp 1676381911
transform 1 0 31392 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _414_
timestamp 1676381911
transform 1 0 31008 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _415_
timestamp 1676381911
transform -1 0 9696 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _416_
timestamp 1676381911
transform -1 0 10080 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _417_
timestamp 1676381911
transform -1 0 10464 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _418_
timestamp 1676381911
transform 1 0 9600 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _419_
timestamp 1676381911
transform -1 0 12576 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _420_
timestamp 1676381911
transform 1 0 9984 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _421_
timestamp 1676381911
transform 1 0 10368 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _422_
timestamp 1676381911
transform -1 0 11136 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _423_
timestamp 1676381911
transform -1 0 11520 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _424_
timestamp 1676381911
transform -1 0 11808 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _425_
timestamp 1676381911
transform 1 0 10176 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _426_
timestamp 1676381911
transform -1 0 12192 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _427_
timestamp 1676381911
transform 1 0 10560 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _428_
timestamp 1676381911
transform -1 0 12960 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _429_
timestamp 1676381911
transform 1 0 11520 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _430_
timestamp 1676381911
transform -1 0 12960 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _431_
timestamp 1676381911
transform 1 0 11904 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _432_
timestamp 1676381911
transform -1 0 13344 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _433_
timestamp 1676381911
transform -1 0 13536 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _434_
timestamp 1676381911
transform -1 0 14496 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _435_
timestamp 1676381911
transform -1 0 13920 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _436_
timestamp 1676381911
transform -1 0 33216 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _437_
timestamp 1676381911
transform -1 0 35520 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _438_
timestamp 1676381911
transform -1 0 38208 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _439_
timestamp 1676381911
transform -1 0 38208 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _440_
timestamp 1676381911
transform -1 0 37536 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _441_
timestamp 1676381911
transform -1 0 15072 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _442_
timestamp 1676381911
transform -1 0 35232 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _443_
timestamp 1676381911
transform -1 0 27360 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _444_
timestamp 1676381911
transform -1 0 33024 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _445_
timestamp 1676381911
transform -1 0 36480 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _446_
timestamp 1676381911
transform -1 0 37632 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _447_
timestamp 1676381911
transform -1 0 23520 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _448_
timestamp 1676381911
transform -1 0 33984 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _449_
timestamp 1676381911
transform -1 0 16416 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _450_
timestamp 1676381911
transform -1 0 16704 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _451_
timestamp 1676381911
transform -1 0 17376 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _452_
timestamp 1676381911
transform -1 0 41856 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _453_
timestamp 1676381911
transform 1 0 16224 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _454_
timestamp 1676381911
transform -1 0 38784 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _455_
timestamp 1676381911
transform 1 0 16032 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _456_
timestamp 1676381911
transform -1 0 23616 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _457_
timestamp 1676381911
transform 1 0 15456 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _458_
timestamp 1676381911
transform 1 0 13536 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _459_
timestamp 1676381911
transform -1 0 40512 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _460_
timestamp 1676381911
transform -1 0 25344 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _461_
timestamp 1676381911
transform -1 0 26016 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _462_
timestamp 1676381911
transform -1 0 32640 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _463_
timestamp 1676381911
transform 1 0 18528 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _464_
timestamp 1676381911
transform -1 0 38400 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _465_
timestamp 1676381911
transform 1 0 18720 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _466_
timestamp 1676381911
transform -1 0 21984 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _467_
timestamp 1676381911
transform -1 0 29856 0 1 2268
box -48 -56 432 834
use sg13g2_buf_8  clkbuf_0_UserCLK
timestamp 1676451365
transform 1 0 27744 0 -1 5292
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_0_UserCLK_regs
timestamp 1676451365
transform -1 0 36768 0 1 756
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_1_0__f_UserCLK_regs
timestamp 1676451365
transform -1 0 35808 0 1 3780
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_1_0__f_UserCLK
timestamp 1676451365
transform 1 0 31104 0 1 756
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_1_1__f_UserCLK_regs
timestamp 1676451365
transform 1 0 40608 0 -1 2268
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_regs_0_UserCLK
timestamp 1676451365
transform 1 0 39072 0 -1 2268
box -48 -56 1296 834
use sg13g2_fill_2  FILLER_0_0
timestamp 1677580104
transform 1 0 1152 0 1 756
box -48 -56 240 834
use sg13g2_fill_2  FILLER_0_24
timestamp 1677580104
transform 1 0 3456 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_26
timestamp 1677579658
transform 1 0 3648 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_44
timestamp 1677580104
transform 1 0 5376 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_46
timestamp 1677579658
transform 1 0 5568 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_126
timestamp 1677580104
transform 1 0 13248 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_128
timestamp 1677579658
transform 1 0 13440 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_150
timestamp 1677580104
transform 1 0 15552 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_152
timestamp 1677579658
transform 1 0 15744 0 1 756
box -48 -56 144 834
use sg13g2_fill_1  FILLER_0_170
timestamp 1677579658
transform 1 0 17472 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_188
timestamp 1677580104
transform 1 0 19200 0 1 756
box -48 -56 240 834
use sg13g2_fill_2  FILLER_0_224
timestamp 1677580104
transform 1 0 22656 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_226
timestamp 1677579658
transform 1 0 22848 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_333
timestamp 1677580104
transform 1 0 33120 0 1 756
box -48 -56 240 834
use sg13g2_fill_2  FILLER_0_356
timestamp 1677580104
transform 1 0 35328 0 1 756
box -48 -56 240 834
use sg13g2_fill_2  FILLER_0_422
timestamp 1677580104
transform 1 0 41664 0 1 756
box -48 -56 240 834
use sg13g2_fill_2  FILLER_1_0
timestamp 1677580104
transform 1 0 1152 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_2
timestamp 1677579658
transform 1 0 1344 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_46
timestamp 1677579658
transform 1 0 5568 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_55
timestamp 1677580104
transform 1 0 6432 0 -1 2268
box -48 -56 240 834
use sg13g2_decap_4  FILLER_1_78
timestamp 1679577901
transform 1 0 8640 0 -1 2268
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_118
timestamp 1677579658
transform 1 0 12480 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_136
timestamp 1677580104
transform 1 0 14208 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_138
timestamp 1677579658
transform 1 0 14400 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_190
timestamp 1677579658
transform 1 0 19392 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_335
timestamp 1677580104
transform 1 0 33312 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_337
timestamp 1677579658
transform 1 0 33504 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_365
timestamp 1677580104
transform 1 0 36192 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_367
timestamp 1677579658
transform 1 0 36384 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_408
timestamp 1677580104
transform 1 0 40320 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_410
timestamp 1677579658
transform 1 0 40512 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_0
timestamp 1677580104
transform 1 0 1152 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_2
timestamp 1677579658
transform 1 0 1344 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_41
timestamp 1677579658
transform 1 0 5088 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_180
timestamp 1677579658
transform 1 0 18432 0 1 2268
box -48 -56 144 834
use sg13g2_decap_4  FILLER_2_223
timestamp 1679577901
transform 1 0 22560 0 1 2268
box -48 -56 432 834
use sg13g2_fill_2  FILLER_2_227
timestamp 1677580104
transform 1 0 22944 0 1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_267
timestamp 1677580104
transform 1 0 26784 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_294
timestamp 1677579658
transform 1 0 29376 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_299
timestamp 1677579658
transform 1 0 29856 0 1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_325
timestamp 1677580104
transform 1 0 32352 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_327
timestamp 1677579658
transform 1 0 32544 0 1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_349
timestamp 1677580104
transform 1 0 34656 0 1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_376
timestamp 1677580104
transform 1 0 37248 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_378
timestamp 1677579658
transform 1 0 37440 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_423
timestamp 1677579658
transform 1 0 41760 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_0
timestamp 1677579658
transform 1 0 1152 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_139
timestamp 1677580104
transform 1 0 14496 0 -1 3780
box -48 -56 240 834
use sg13g2_decap_4  FILLER_3_217
timestamp 1679577901
transform 1 0 21984 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_3_221
timestamp 1677579658
transform 1 0 22368 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_239
timestamp 1677580104
transform 1 0 24096 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_342
timestamp 1677580104
transform 1 0 33984 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_361
timestamp 1677580104
transform 1 0 35808 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_363
timestamp 1677579658
transform 1 0 36000 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_381
timestamp 1677579658
transform 1 0 37728 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_0
timestamp 1677579658
transform 1 0 1152 0 1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_50
timestamp 1677579658
transform 1 0 5952 0 1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_91
timestamp 1677579658
transform 1 0 9888 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_131
timestamp 1677580104
transform 1 0 13728 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_133
timestamp 1677579658
transform 1 0 13920 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_155
timestamp 1677580104
transform 1 0 16032 0 1 3780
box -48 -56 240 834
use sg13g2_decap_4  FILLER_4_161
timestamp 1679577901
transform 1 0 16608 0 1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_4_207
timestamp 1677580104
transform 1 0 21024 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_230
timestamp 1679581782
transform 1 0 23232 0 1 3780
box -48 -56 720 834
use sg13g2_decap_4  FILLER_4_237
timestamp 1679577901
transform 1 0 23904 0 1 3780
box -48 -56 432 834
use sg13g2_fill_1  FILLER_4_241
timestamp 1677579658
transform 1 0 24288 0 1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_263
timestamp 1677579658
transform 1 0 26400 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_390
timestamp 1677580104
transform 1 0 38592 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_392
timestamp 1677579658
transform 1 0 38784 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_422
timestamp 1677580104
transform 1 0 41664 0 1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_5_38
timestamp 1677580104
transform 1 0 4800 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_40
timestamp 1677579658
transform 1 0 4992 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_5_136
timestamp 1679577901
transform 1 0 14208 0 -1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_5_161
timestamp 1677579658
transform 1 0 16608 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_204
timestamp 1679581782
transform 1 0 20736 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_2  FILLER_5_211
timestamp 1677580104
transform 1 0 21408 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_272
timestamp 1677579658
transform 1 0 27264 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_311
timestamp 1677580104
transform 1 0 31008 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_355
timestamp 1677579658
transform 1 0 35232 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_394
timestamp 1677579658
transform 1 0 38976 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_0
timestamp 1677579658
transform 1 0 1152 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_18
timestamp 1677580104
transform 1 0 2880 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_20
timestamp 1677579658
transform 1 0 3072 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_75
timestamp 1677579658
transform 1 0 8352 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_106
timestamp 1677579658
transform 1 0 11328 0 1 5292
box -48 -56 144 834
use sg13g2_decap_4  FILLER_6_119
timestamp 1679577901
transform 1 0 12576 0 1 5292
box -48 -56 432 834
use sg13g2_fill_2  FILLER_6_123
timestamp 1677580104
transform 1 0 12960 0 1 5292
box -48 -56 240 834
use sg13g2_decap_4  FILLER_6_150
timestamp 1679577901
transform 1 0 15552 0 1 5292
box -48 -56 432 834
use sg13g2_fill_1  FILLER_6_154
timestamp 1677579658
transform 1 0 15936 0 1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_6_227
timestamp 1679581782
transform 1 0 22944 0 1 5292
box -48 -56 720 834
use sg13g2_decap_8  FILLER_6_234
timestamp 1679581782
transform 1 0 23616 0 1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_258
timestamp 1677579658
transform 1 0 25920 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_310
timestamp 1677579658
transform 1 0 30912 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_353
timestamp 1677579658
transform 1 0 35040 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_412
timestamp 1677579658
transform 1 0 40704 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_421
timestamp 1677580104
transform 1 0 41568 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_423
timestamp 1677579658
transform 1 0 41760 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_77
timestamp 1677580104
transform 1 0 8544 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_101
timestamp 1677579658
transform 1 0 10848 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_174
timestamp 1679581782
transform 1 0 17856 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_181
timestamp 1677580104
transform 1 0 18528 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_8  FILLER_7_204
timestamp 1679581782
transform 1 0 20736 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_211
timestamp 1679581782
transform 1 0 21408 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_7_218
timestamp 1677579658
transform 1 0 22080 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_257
timestamp 1677580104
transform 1 0 25824 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_351
timestamp 1677579658
transform 1 0 34848 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_373
timestamp 1677580104
transform 1 0 36960 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_400
timestamp 1677580104
transform 1 0 39552 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_7_410
timestamp 1677580104
transform 1 0 40512 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_412
timestamp 1677579658
transform 1 0 40704 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_421
timestamp 1677580104
transform 1 0 41568 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_423
timestamp 1677579658
transform 1 0 41760 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_0
timestamp 1677579658
transform 1 0 1152 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_22
timestamp 1677579658
transform 1 0 3264 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_33
timestamp 1677580104
transform 1 0 4320 0 1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_62
timestamp 1677580104
transform 1 0 7104 0 1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_123
timestamp 1677580104
transform 1 0 12960 0 1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_146
timestamp 1677580104
transform 1 0 15168 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_148
timestamp 1677579658
transform 1 0 15360 0 1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_170
timestamp 1679577901
transform 1 0 17472 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_174
timestamp 1677579658
transform 1 0 17856 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_196
timestamp 1679581782
transform 1 0 19968 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_203
timestamp 1677580104
transform 1 0 20640 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_205
timestamp 1677579658
transform 1 0 20832 0 1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_240
timestamp 1679577901
transform 1 0 24192 0 1 6804
box -48 -56 432 834
use sg13g2_fill_1  FILLER_8_244
timestamp 1677579658
transform 1 0 24576 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_262
timestamp 1679581782
transform 1 0 26304 0 1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_8_269
timestamp 1679581782
transform 1 0 26976 0 1 6804
box -48 -56 720 834
use sg13g2_fill_1  FILLER_8_297
timestamp 1677579658
transform 1 0 29664 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_353
timestamp 1677580104
transform 1 0 35040 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_355
timestamp 1677579658
transform 1 0 35232 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_423
timestamp 1677579658
transform 1 0 41760 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_9_0
timestamp 1679581782
transform 1 0 1152 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_24
timestamp 1677580104
transform 1 0 3456 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_26
timestamp 1677579658
transform 1 0 3648 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_54
timestamp 1677580104
transform 1 0 6336 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_124
timestamp 1679581782
transform 1 0 13056 0 -1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_9_131
timestamp 1677580104
transform 1 0 13728 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_9_150
timestamp 1679581782
transform 1 0 15552 0 -1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_9_233
timestamp 1679577901
transform 1 0 23520 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_237
timestamp 1677579658
transform 1 0 23904 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_263
timestamp 1677580104
transform 1 0 26400 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_265
timestamp 1677579658
transform 1 0 26592 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_312
timestamp 1677580104
transform 1 0 31104 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_335
timestamp 1677580104
transform 1 0 33312 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_337
timestamp 1677579658
transform 1 0 33504 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_421
timestamp 1677580104
transform 1 0 41568 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_423
timestamp 1677579658
transform 1 0 41760 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_10_0
timestamp 1679577901
transform 1 0 1152 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_4
timestamp 1677580104
transform 1 0 1536 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_54
timestamp 1677580104
transform 1 0 6336 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_56
timestamp 1677579658
transform 1 0 6528 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_154
timestamp 1677580104
transform 1 0 15936 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_156
timestamp 1677579658
transform 1 0 16128 0 1 8316
box -48 -56 144 834
use sg13g2_decap_8  FILLER_10_203
timestamp 1679581782
transform 1 0 20640 0 1 8316
box -48 -56 720 834
use sg13g2_fill_2  FILLER_10_210
timestamp 1677580104
transform 1 0 21312 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_212
timestamp 1677579658
transform 1 0 21504 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_234
timestamp 1677579658
transform 1 0 23616 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_302
timestamp 1677579658
transform 1 0 30144 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_332
timestamp 1677579658
transform 1 0 33024 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_358
timestamp 1677579658
transform 1 0 35520 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_10_422
timestamp 1677580104
transform 1 0 41664 0 1 8316
box -48 -56 240 834
use sg13g2_decap_4  FILLER_11_0
timestamp 1679577901
transform 1 0 1152 0 -1 9828
box -48 -56 432 834
use sg13g2_decap_8  FILLER_11_43
timestamp 1679581782
transform 1 0 5280 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_50
timestamp 1677579658
transform 1 0 5952 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_69
timestamp 1677580104
transform 1 0 7776 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_71
timestamp 1677579658
transform 1 0 7968 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_77
timestamp 1677579658
transform 1 0 8544 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_83
timestamp 1677580104
transform 1 0 9120 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_8  FILLER_11_97
timestamp 1679581782
transform 1 0 10464 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_104
timestamp 1679581782
transform 1 0 11136 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_111
timestamp 1679581782
transform 1 0 11808 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_1  FILLER_11_118
timestamp 1677579658
transform 1 0 12480 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_127
timestamp 1679581782
transform 1 0 13344 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_134
timestamp 1679581782
transform 1 0 14016 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_179
timestamp 1677580104
transform 1 0 18336 0 -1 9828
box -48 -56 240 834
use sg13g2_decap_4  FILLER_11_185
timestamp 1679577901
transform 1 0 18912 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_11_189
timestamp 1677579658
transform 1 0 19296 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_245
timestamp 1677580104
transform 1 0 24672 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_247
timestamp 1677579658
transform 1 0 24864 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_273
timestamp 1679581782
transform 1 0 27360 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_8  FILLER_11_280
timestamp 1679581782
transform 1 0 28032 0 -1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_11_287
timestamp 1679577901
transform 1 0 28704 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_2  FILLER_11_291
timestamp 1677580104
transform 1 0 29088 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_361
timestamp 1677580104
transform 1 0 35808 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_422
timestamp 1677580104
transform 1 0 41664 0 -1 9828
box -48 -56 240 834
<< labels >>
flabel metal2 s 4088 0 4168 80 0 FreeSans 320 0 0 0 A_I_top
port 0 nsew signal output
flabel metal2 s 2936 0 3016 80 0 FreeSans 320 0 0 0 A_O_top
port 1 nsew signal input
flabel metal2 s 5240 0 5320 80 0 FreeSans 320 0 0 0 A_T_top
port 2 nsew signal output
flabel metal2 s 7544 0 7624 80 0 FreeSans 320 0 0 0 B_I_top
port 3 nsew signal output
flabel metal2 s 6392 0 6472 80 0 FreeSans 320 0 0 0 B_O_top
port 4 nsew signal input
flabel metal2 s 8696 0 8776 80 0 FreeSans 320 0 0 0 B_T_top
port 5 nsew signal output
flabel metal2 s 11000 0 11080 80 0 FreeSans 320 0 0 0 C_I_top
port 6 nsew signal output
flabel metal2 s 9848 0 9928 80 0 FreeSans 320 0 0 0 C_O_top
port 7 nsew signal input
flabel metal2 s 12152 0 12232 80 0 FreeSans 320 0 0 0 C_T_top
port 8 nsew signal output
flabel metal2 s 19448 10672 19528 10752 0 FreeSans 320 0 0 0 Co
port 9 nsew signal output
flabel metal2 s 14456 0 14536 80 0 FreeSans 320 0 0 0 D_I_top
port 10 nsew signal output
flabel metal2 s 13304 0 13384 80 0 FreeSans 320 0 0 0 D_O_top
port 11 nsew signal input
flabel metal2 s 15608 0 15688 80 0 FreeSans 320 0 0 0 D_T_top
port 12 nsew signal output
flabel metal3 s 0 44 80 124 0 FreeSans 320 0 0 0 FrameData[0]
port 13 nsew signal input
flabel metal3 s 0 3404 80 3484 0 FreeSans 320 0 0 0 FrameData[10]
port 14 nsew signal input
flabel metal3 s 0 3740 80 3820 0 FreeSans 320 0 0 0 FrameData[11]
port 15 nsew signal input
flabel metal3 s 0 4076 80 4156 0 FreeSans 320 0 0 0 FrameData[12]
port 16 nsew signal input
flabel metal3 s 0 4412 80 4492 0 FreeSans 320 0 0 0 FrameData[13]
port 17 nsew signal input
flabel metal3 s 0 4748 80 4828 0 FreeSans 320 0 0 0 FrameData[14]
port 18 nsew signal input
flabel metal3 s 0 5084 80 5164 0 FreeSans 320 0 0 0 FrameData[15]
port 19 nsew signal input
flabel metal3 s 0 5420 80 5500 0 FreeSans 320 0 0 0 FrameData[16]
port 20 nsew signal input
flabel metal3 s 0 5756 80 5836 0 FreeSans 320 0 0 0 FrameData[17]
port 21 nsew signal input
flabel metal3 s 0 6092 80 6172 0 FreeSans 320 0 0 0 FrameData[18]
port 22 nsew signal input
flabel metal3 s 0 6428 80 6508 0 FreeSans 320 0 0 0 FrameData[19]
port 23 nsew signal input
flabel metal3 s 0 380 80 460 0 FreeSans 320 0 0 0 FrameData[1]
port 24 nsew signal input
flabel metal3 s 0 6764 80 6844 0 FreeSans 320 0 0 0 FrameData[20]
port 25 nsew signal input
flabel metal3 s 0 7100 80 7180 0 FreeSans 320 0 0 0 FrameData[21]
port 26 nsew signal input
flabel metal3 s 0 7436 80 7516 0 FreeSans 320 0 0 0 FrameData[22]
port 27 nsew signal input
flabel metal3 s 0 7772 80 7852 0 FreeSans 320 0 0 0 FrameData[23]
port 28 nsew signal input
flabel metal3 s 0 8108 80 8188 0 FreeSans 320 0 0 0 FrameData[24]
port 29 nsew signal input
flabel metal3 s 0 8444 80 8524 0 FreeSans 320 0 0 0 FrameData[25]
port 30 nsew signal input
flabel metal3 s 0 8780 80 8860 0 FreeSans 320 0 0 0 FrameData[26]
port 31 nsew signal input
flabel metal3 s 0 9116 80 9196 0 FreeSans 320 0 0 0 FrameData[27]
port 32 nsew signal input
flabel metal3 s 0 9452 80 9532 0 FreeSans 320 0 0 0 FrameData[28]
port 33 nsew signal input
flabel metal3 s 0 9788 80 9868 0 FreeSans 320 0 0 0 FrameData[29]
port 34 nsew signal input
flabel metal3 s 0 716 80 796 0 FreeSans 320 0 0 0 FrameData[2]
port 35 nsew signal input
flabel metal3 s 0 10124 80 10204 0 FreeSans 320 0 0 0 FrameData[30]
port 36 nsew signal input
flabel metal3 s 0 10460 80 10540 0 FreeSans 320 0 0 0 FrameData[31]
port 37 nsew signal input
flabel metal3 s 0 1052 80 1132 0 FreeSans 320 0 0 0 FrameData[3]
port 38 nsew signal input
flabel metal3 s 0 1388 80 1468 0 FreeSans 320 0 0 0 FrameData[4]
port 39 nsew signal input
flabel metal3 s 0 1724 80 1804 0 FreeSans 320 0 0 0 FrameData[5]
port 40 nsew signal input
flabel metal3 s 0 2060 80 2140 0 FreeSans 320 0 0 0 FrameData[6]
port 41 nsew signal input
flabel metal3 s 0 2396 80 2476 0 FreeSans 320 0 0 0 FrameData[7]
port 42 nsew signal input
flabel metal3 s 0 2732 80 2812 0 FreeSans 320 0 0 0 FrameData[8]
port 43 nsew signal input
flabel metal3 s 0 3068 80 3148 0 FreeSans 320 0 0 0 FrameData[9]
port 44 nsew signal input
flabel metal3 s 42928 44 43008 124 0 FreeSans 320 0 0 0 FrameData_O[0]
port 45 nsew signal output
flabel metal3 s 42928 3404 43008 3484 0 FreeSans 320 0 0 0 FrameData_O[10]
port 46 nsew signal output
flabel metal3 s 42928 3740 43008 3820 0 FreeSans 320 0 0 0 FrameData_O[11]
port 47 nsew signal output
flabel metal3 s 42928 4076 43008 4156 0 FreeSans 320 0 0 0 FrameData_O[12]
port 48 nsew signal output
flabel metal3 s 42928 4412 43008 4492 0 FreeSans 320 0 0 0 FrameData_O[13]
port 49 nsew signal output
flabel metal3 s 42928 4748 43008 4828 0 FreeSans 320 0 0 0 FrameData_O[14]
port 50 nsew signal output
flabel metal3 s 42928 5084 43008 5164 0 FreeSans 320 0 0 0 FrameData_O[15]
port 51 nsew signal output
flabel metal3 s 42928 5420 43008 5500 0 FreeSans 320 0 0 0 FrameData_O[16]
port 52 nsew signal output
flabel metal3 s 42928 5756 43008 5836 0 FreeSans 320 0 0 0 FrameData_O[17]
port 53 nsew signal output
flabel metal3 s 42928 6092 43008 6172 0 FreeSans 320 0 0 0 FrameData_O[18]
port 54 nsew signal output
flabel metal3 s 42928 6428 43008 6508 0 FreeSans 320 0 0 0 FrameData_O[19]
port 55 nsew signal output
flabel metal3 s 42928 380 43008 460 0 FreeSans 320 0 0 0 FrameData_O[1]
port 56 nsew signal output
flabel metal3 s 42928 6764 43008 6844 0 FreeSans 320 0 0 0 FrameData_O[20]
port 57 nsew signal output
flabel metal3 s 42928 7100 43008 7180 0 FreeSans 320 0 0 0 FrameData_O[21]
port 58 nsew signal output
flabel metal3 s 42928 7436 43008 7516 0 FreeSans 320 0 0 0 FrameData_O[22]
port 59 nsew signal output
flabel metal3 s 42928 7772 43008 7852 0 FreeSans 320 0 0 0 FrameData_O[23]
port 60 nsew signal output
flabel metal3 s 42928 8108 43008 8188 0 FreeSans 320 0 0 0 FrameData_O[24]
port 61 nsew signal output
flabel metal3 s 42928 8444 43008 8524 0 FreeSans 320 0 0 0 FrameData_O[25]
port 62 nsew signal output
flabel metal3 s 42928 8780 43008 8860 0 FreeSans 320 0 0 0 FrameData_O[26]
port 63 nsew signal output
flabel metal3 s 42928 9116 43008 9196 0 FreeSans 320 0 0 0 FrameData_O[27]
port 64 nsew signal output
flabel metal3 s 42928 9452 43008 9532 0 FreeSans 320 0 0 0 FrameData_O[28]
port 65 nsew signal output
flabel metal3 s 42928 9788 43008 9868 0 FreeSans 320 0 0 0 FrameData_O[29]
port 66 nsew signal output
flabel metal3 s 42928 716 43008 796 0 FreeSans 320 0 0 0 FrameData_O[2]
port 67 nsew signal output
flabel metal3 s 42928 10124 43008 10204 0 FreeSans 320 0 0 0 FrameData_O[30]
port 68 nsew signal output
flabel metal3 s 42928 10460 43008 10540 0 FreeSans 320 0 0 0 FrameData_O[31]
port 69 nsew signal output
flabel metal3 s 42928 1052 43008 1132 0 FreeSans 320 0 0 0 FrameData_O[3]
port 70 nsew signal output
flabel metal3 s 42928 1388 43008 1468 0 FreeSans 320 0 0 0 FrameData_O[4]
port 71 nsew signal output
flabel metal3 s 42928 1724 43008 1804 0 FreeSans 320 0 0 0 FrameData_O[5]
port 72 nsew signal output
flabel metal3 s 42928 2060 43008 2140 0 FreeSans 320 0 0 0 FrameData_O[6]
port 73 nsew signal output
flabel metal3 s 42928 2396 43008 2476 0 FreeSans 320 0 0 0 FrameData_O[7]
port 74 nsew signal output
flabel metal3 s 42928 2732 43008 2812 0 FreeSans 320 0 0 0 FrameData_O[8]
port 75 nsew signal output
flabel metal3 s 42928 3068 43008 3148 0 FreeSans 320 0 0 0 FrameData_O[9]
port 76 nsew signal output
flabel metal2 s 17912 0 17992 80 0 FreeSans 320 0 0 0 FrameStrobe[0]
port 77 nsew signal input
flabel metal2 s 29432 0 29512 80 0 FreeSans 320 0 0 0 FrameStrobe[10]
port 78 nsew signal input
flabel metal2 s 30584 0 30664 80 0 FreeSans 320 0 0 0 FrameStrobe[11]
port 79 nsew signal input
flabel metal2 s 31736 0 31816 80 0 FreeSans 320 0 0 0 FrameStrobe[12]
port 80 nsew signal input
flabel metal2 s 32888 0 32968 80 0 FreeSans 320 0 0 0 FrameStrobe[13]
port 81 nsew signal input
flabel metal2 s 34040 0 34120 80 0 FreeSans 320 0 0 0 FrameStrobe[14]
port 82 nsew signal input
flabel metal2 s 35192 0 35272 80 0 FreeSans 320 0 0 0 FrameStrobe[15]
port 83 nsew signal input
flabel metal2 s 36344 0 36424 80 0 FreeSans 320 0 0 0 FrameStrobe[16]
port 84 nsew signal input
flabel metal2 s 37496 0 37576 80 0 FreeSans 320 0 0 0 FrameStrobe[17]
port 85 nsew signal input
flabel metal2 s 38648 0 38728 80 0 FreeSans 320 0 0 0 FrameStrobe[18]
port 86 nsew signal input
flabel metal2 s 39800 0 39880 80 0 FreeSans 320 0 0 0 FrameStrobe[19]
port 87 nsew signal input
flabel metal2 s 19064 0 19144 80 0 FreeSans 320 0 0 0 FrameStrobe[1]
port 88 nsew signal input
flabel metal2 s 20216 0 20296 80 0 FreeSans 320 0 0 0 FrameStrobe[2]
port 89 nsew signal input
flabel metal2 s 21368 0 21448 80 0 FreeSans 320 0 0 0 FrameStrobe[3]
port 90 nsew signal input
flabel metal2 s 22520 0 22600 80 0 FreeSans 320 0 0 0 FrameStrobe[4]
port 91 nsew signal input
flabel metal2 s 23672 0 23752 80 0 FreeSans 320 0 0 0 FrameStrobe[5]
port 92 nsew signal input
flabel metal2 s 24824 0 24904 80 0 FreeSans 320 0 0 0 FrameStrobe[6]
port 93 nsew signal input
flabel metal2 s 25976 0 26056 80 0 FreeSans 320 0 0 0 FrameStrobe[7]
port 94 nsew signal input
flabel metal2 s 27128 0 27208 80 0 FreeSans 320 0 0 0 FrameStrobe[8]
port 95 nsew signal input
flabel metal2 s 28280 0 28360 80 0 FreeSans 320 0 0 0 FrameStrobe[9]
port 96 nsew signal input
flabel metal2 s 29816 10672 29896 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[0]
port 97 nsew signal output
flabel metal2 s 31736 10672 31816 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[10]
port 98 nsew signal output
flabel metal2 s 31928 10672 32008 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[11]
port 99 nsew signal output
flabel metal2 s 32120 10672 32200 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[12]
port 100 nsew signal output
flabel metal2 s 32312 10672 32392 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[13]
port 101 nsew signal output
flabel metal2 s 32504 10672 32584 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[14]
port 102 nsew signal output
flabel metal2 s 32696 10672 32776 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[15]
port 103 nsew signal output
flabel metal2 s 32888 10672 32968 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[16]
port 104 nsew signal output
flabel metal2 s 33080 10672 33160 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[17]
port 105 nsew signal output
flabel metal2 s 33272 10672 33352 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[18]
port 106 nsew signal output
flabel metal2 s 33464 10672 33544 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[19]
port 107 nsew signal output
flabel metal2 s 30008 10672 30088 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[1]
port 108 nsew signal output
flabel metal2 s 30200 10672 30280 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[2]
port 109 nsew signal output
flabel metal2 s 30392 10672 30472 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[3]
port 110 nsew signal output
flabel metal2 s 30584 10672 30664 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[4]
port 111 nsew signal output
flabel metal2 s 30776 10672 30856 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[5]
port 112 nsew signal output
flabel metal2 s 30968 10672 31048 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[6]
port 113 nsew signal output
flabel metal2 s 31160 10672 31240 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[7]
port 114 nsew signal output
flabel metal2 s 31352 10672 31432 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[8]
port 115 nsew signal output
flabel metal2 s 31544 10672 31624 10752 0 FreeSans 320 0 0 0 FrameStrobe_O[9]
port 116 nsew signal output
flabel metal2 s 9464 10672 9544 10752 0 FreeSans 320 0 0 0 N1BEG[0]
port 117 nsew signal output
flabel metal2 s 9656 10672 9736 10752 0 FreeSans 320 0 0 0 N1BEG[1]
port 118 nsew signal output
flabel metal2 s 9848 10672 9928 10752 0 FreeSans 320 0 0 0 N1BEG[2]
port 119 nsew signal output
flabel metal2 s 10040 10672 10120 10752 0 FreeSans 320 0 0 0 N1BEG[3]
port 120 nsew signal output
flabel metal2 s 10232 10672 10312 10752 0 FreeSans 320 0 0 0 N2BEG[0]
port 121 nsew signal output
flabel metal2 s 10424 10672 10504 10752 0 FreeSans 320 0 0 0 N2BEG[1]
port 122 nsew signal output
flabel metal2 s 10616 10672 10696 10752 0 FreeSans 320 0 0 0 N2BEG[2]
port 123 nsew signal output
flabel metal2 s 10808 10672 10888 10752 0 FreeSans 320 0 0 0 N2BEG[3]
port 124 nsew signal output
flabel metal2 s 11000 10672 11080 10752 0 FreeSans 320 0 0 0 N2BEG[4]
port 125 nsew signal output
flabel metal2 s 11192 10672 11272 10752 0 FreeSans 320 0 0 0 N2BEG[5]
port 126 nsew signal output
flabel metal2 s 11384 10672 11464 10752 0 FreeSans 320 0 0 0 N2BEG[6]
port 127 nsew signal output
flabel metal2 s 11576 10672 11656 10752 0 FreeSans 320 0 0 0 N2BEG[7]
port 128 nsew signal output
flabel metal2 s 11768 10672 11848 10752 0 FreeSans 320 0 0 0 N2BEGb[0]
port 129 nsew signal output
flabel metal2 s 11960 10672 12040 10752 0 FreeSans 320 0 0 0 N2BEGb[1]
port 130 nsew signal output
flabel metal2 s 12152 10672 12232 10752 0 FreeSans 320 0 0 0 N2BEGb[2]
port 131 nsew signal output
flabel metal2 s 12344 10672 12424 10752 0 FreeSans 320 0 0 0 N2BEGb[3]
port 132 nsew signal output
flabel metal2 s 12536 10672 12616 10752 0 FreeSans 320 0 0 0 N2BEGb[4]
port 133 nsew signal output
flabel metal2 s 12728 10672 12808 10752 0 FreeSans 320 0 0 0 N2BEGb[5]
port 134 nsew signal output
flabel metal2 s 12920 10672 13000 10752 0 FreeSans 320 0 0 0 N2BEGb[6]
port 135 nsew signal output
flabel metal2 s 13112 10672 13192 10752 0 FreeSans 320 0 0 0 N2BEGb[7]
port 136 nsew signal output
flabel metal2 s 13304 10672 13384 10752 0 FreeSans 320 0 0 0 N4BEG[0]
port 137 nsew signal output
flabel metal2 s 15224 10672 15304 10752 0 FreeSans 320 0 0 0 N4BEG[10]
port 138 nsew signal output
flabel metal2 s 15416 10672 15496 10752 0 FreeSans 320 0 0 0 N4BEG[11]
port 139 nsew signal output
flabel metal2 s 15608 10672 15688 10752 0 FreeSans 320 0 0 0 N4BEG[12]
port 140 nsew signal output
flabel metal2 s 15800 10672 15880 10752 0 FreeSans 320 0 0 0 N4BEG[13]
port 141 nsew signal output
flabel metal2 s 15992 10672 16072 10752 0 FreeSans 320 0 0 0 N4BEG[14]
port 142 nsew signal output
flabel metal2 s 16184 10672 16264 10752 0 FreeSans 320 0 0 0 N4BEG[15]
port 143 nsew signal output
flabel metal2 s 13496 10672 13576 10752 0 FreeSans 320 0 0 0 N4BEG[1]
port 144 nsew signal output
flabel metal2 s 13688 10672 13768 10752 0 FreeSans 320 0 0 0 N4BEG[2]
port 145 nsew signal output
flabel metal2 s 13880 10672 13960 10752 0 FreeSans 320 0 0 0 N4BEG[3]
port 146 nsew signal output
flabel metal2 s 14072 10672 14152 10752 0 FreeSans 320 0 0 0 N4BEG[4]
port 147 nsew signal output
flabel metal2 s 14264 10672 14344 10752 0 FreeSans 320 0 0 0 N4BEG[5]
port 148 nsew signal output
flabel metal2 s 14456 10672 14536 10752 0 FreeSans 320 0 0 0 N4BEG[6]
port 149 nsew signal output
flabel metal2 s 14648 10672 14728 10752 0 FreeSans 320 0 0 0 N4BEG[7]
port 150 nsew signal output
flabel metal2 s 14840 10672 14920 10752 0 FreeSans 320 0 0 0 N4BEG[8]
port 151 nsew signal output
flabel metal2 s 15032 10672 15112 10752 0 FreeSans 320 0 0 0 N4BEG[9]
port 152 nsew signal output
flabel metal2 s 16376 10672 16456 10752 0 FreeSans 320 0 0 0 NN4BEG[0]
port 153 nsew signal output
flabel metal2 s 18296 10672 18376 10752 0 FreeSans 320 0 0 0 NN4BEG[10]
port 154 nsew signal output
flabel metal2 s 18488 10672 18568 10752 0 FreeSans 320 0 0 0 NN4BEG[11]
port 155 nsew signal output
flabel metal2 s 18680 10672 18760 10752 0 FreeSans 320 0 0 0 NN4BEG[12]
port 156 nsew signal output
flabel metal2 s 18872 10672 18952 10752 0 FreeSans 320 0 0 0 NN4BEG[13]
port 157 nsew signal output
flabel metal2 s 19064 10672 19144 10752 0 FreeSans 320 0 0 0 NN4BEG[14]
port 158 nsew signal output
flabel metal2 s 19256 10672 19336 10752 0 FreeSans 320 0 0 0 NN4BEG[15]
port 159 nsew signal output
flabel metal2 s 16568 10672 16648 10752 0 FreeSans 320 0 0 0 NN4BEG[1]
port 160 nsew signal output
flabel metal2 s 16760 10672 16840 10752 0 FreeSans 320 0 0 0 NN4BEG[2]
port 161 nsew signal output
flabel metal2 s 16952 10672 17032 10752 0 FreeSans 320 0 0 0 NN4BEG[3]
port 162 nsew signal output
flabel metal2 s 17144 10672 17224 10752 0 FreeSans 320 0 0 0 NN4BEG[4]
port 163 nsew signal output
flabel metal2 s 17336 10672 17416 10752 0 FreeSans 320 0 0 0 NN4BEG[5]
port 164 nsew signal output
flabel metal2 s 17528 10672 17608 10752 0 FreeSans 320 0 0 0 NN4BEG[6]
port 165 nsew signal output
flabel metal2 s 17720 10672 17800 10752 0 FreeSans 320 0 0 0 NN4BEG[7]
port 166 nsew signal output
flabel metal2 s 17912 10672 17992 10752 0 FreeSans 320 0 0 0 NN4BEG[8]
port 167 nsew signal output
flabel metal2 s 18104 10672 18184 10752 0 FreeSans 320 0 0 0 NN4BEG[9]
port 168 nsew signal output
flabel metal2 s 19640 10672 19720 10752 0 FreeSans 320 0 0 0 S1END[0]
port 169 nsew signal input
flabel metal2 s 19832 10672 19912 10752 0 FreeSans 320 0 0 0 S1END[1]
port 170 nsew signal input
flabel metal2 s 20024 10672 20104 10752 0 FreeSans 320 0 0 0 S1END[2]
port 171 nsew signal input
flabel metal2 s 20216 10672 20296 10752 0 FreeSans 320 0 0 0 S1END[3]
port 172 nsew signal input
flabel metal2 s 21944 10672 22024 10752 0 FreeSans 320 0 0 0 S2END[0]
port 173 nsew signal input
flabel metal2 s 22136 10672 22216 10752 0 FreeSans 320 0 0 0 S2END[1]
port 174 nsew signal input
flabel metal2 s 22328 10672 22408 10752 0 FreeSans 320 0 0 0 S2END[2]
port 175 nsew signal input
flabel metal2 s 22520 10672 22600 10752 0 FreeSans 320 0 0 0 S2END[3]
port 176 nsew signal input
flabel metal2 s 22712 10672 22792 10752 0 FreeSans 320 0 0 0 S2END[4]
port 177 nsew signal input
flabel metal2 s 22904 10672 22984 10752 0 FreeSans 320 0 0 0 S2END[5]
port 178 nsew signal input
flabel metal2 s 23096 10672 23176 10752 0 FreeSans 320 0 0 0 S2END[6]
port 179 nsew signal input
flabel metal2 s 23288 10672 23368 10752 0 FreeSans 320 0 0 0 S2END[7]
port 180 nsew signal input
flabel metal2 s 20408 10672 20488 10752 0 FreeSans 320 0 0 0 S2MID[0]
port 181 nsew signal input
flabel metal2 s 20600 10672 20680 10752 0 FreeSans 320 0 0 0 S2MID[1]
port 182 nsew signal input
flabel metal2 s 20792 10672 20872 10752 0 FreeSans 320 0 0 0 S2MID[2]
port 183 nsew signal input
flabel metal2 s 20984 10672 21064 10752 0 FreeSans 320 0 0 0 S2MID[3]
port 184 nsew signal input
flabel metal2 s 21176 10672 21256 10752 0 FreeSans 320 0 0 0 S2MID[4]
port 185 nsew signal input
flabel metal2 s 21368 10672 21448 10752 0 FreeSans 320 0 0 0 S2MID[5]
port 186 nsew signal input
flabel metal2 s 21560 10672 21640 10752 0 FreeSans 320 0 0 0 S2MID[6]
port 187 nsew signal input
flabel metal2 s 21752 10672 21832 10752 0 FreeSans 320 0 0 0 S2MID[7]
port 188 nsew signal input
flabel metal2 s 23480 10672 23560 10752 0 FreeSans 320 0 0 0 S4END[0]
port 189 nsew signal input
flabel metal2 s 25400 10672 25480 10752 0 FreeSans 320 0 0 0 S4END[10]
port 190 nsew signal input
flabel metal2 s 25592 10672 25672 10752 0 FreeSans 320 0 0 0 S4END[11]
port 191 nsew signal input
flabel metal2 s 25784 10672 25864 10752 0 FreeSans 320 0 0 0 S4END[12]
port 192 nsew signal input
flabel metal2 s 25976 10672 26056 10752 0 FreeSans 320 0 0 0 S4END[13]
port 193 nsew signal input
flabel metal2 s 26168 10672 26248 10752 0 FreeSans 320 0 0 0 S4END[14]
port 194 nsew signal input
flabel metal2 s 26360 10672 26440 10752 0 FreeSans 320 0 0 0 S4END[15]
port 195 nsew signal input
flabel metal2 s 23672 10672 23752 10752 0 FreeSans 320 0 0 0 S4END[1]
port 196 nsew signal input
flabel metal2 s 23864 10672 23944 10752 0 FreeSans 320 0 0 0 S4END[2]
port 197 nsew signal input
flabel metal2 s 24056 10672 24136 10752 0 FreeSans 320 0 0 0 S4END[3]
port 198 nsew signal input
flabel metal2 s 24248 10672 24328 10752 0 FreeSans 320 0 0 0 S4END[4]
port 199 nsew signal input
flabel metal2 s 24440 10672 24520 10752 0 FreeSans 320 0 0 0 S4END[5]
port 200 nsew signal input
flabel metal2 s 24632 10672 24712 10752 0 FreeSans 320 0 0 0 S4END[6]
port 201 nsew signal input
flabel metal2 s 24824 10672 24904 10752 0 FreeSans 320 0 0 0 S4END[7]
port 202 nsew signal input
flabel metal2 s 25016 10672 25096 10752 0 FreeSans 320 0 0 0 S4END[8]
port 203 nsew signal input
flabel metal2 s 25208 10672 25288 10752 0 FreeSans 320 0 0 0 S4END[9]
port 204 nsew signal input
flabel metal2 s 26552 10672 26632 10752 0 FreeSans 320 0 0 0 SS4END[0]
port 205 nsew signal input
flabel metal2 s 28472 10672 28552 10752 0 FreeSans 320 0 0 0 SS4END[10]
port 206 nsew signal input
flabel metal2 s 28664 10672 28744 10752 0 FreeSans 320 0 0 0 SS4END[11]
port 207 nsew signal input
flabel metal2 s 28856 10672 28936 10752 0 FreeSans 320 0 0 0 SS4END[12]
port 208 nsew signal input
flabel metal2 s 29048 10672 29128 10752 0 FreeSans 320 0 0 0 SS4END[13]
port 209 nsew signal input
flabel metal2 s 29240 10672 29320 10752 0 FreeSans 320 0 0 0 SS4END[14]
port 210 nsew signal input
flabel metal2 s 29432 10672 29512 10752 0 FreeSans 320 0 0 0 SS4END[15]
port 211 nsew signal input
flabel metal2 s 26744 10672 26824 10752 0 FreeSans 320 0 0 0 SS4END[1]
port 212 nsew signal input
flabel metal2 s 26936 10672 27016 10752 0 FreeSans 320 0 0 0 SS4END[2]
port 213 nsew signal input
flabel metal2 s 27128 10672 27208 10752 0 FreeSans 320 0 0 0 SS4END[3]
port 214 nsew signal input
flabel metal2 s 27320 10672 27400 10752 0 FreeSans 320 0 0 0 SS4END[4]
port 215 nsew signal input
flabel metal2 s 27512 10672 27592 10752 0 FreeSans 320 0 0 0 SS4END[5]
port 216 nsew signal input
flabel metal2 s 27704 10672 27784 10752 0 FreeSans 320 0 0 0 SS4END[6]
port 217 nsew signal input
flabel metal2 s 27896 10672 27976 10752 0 FreeSans 320 0 0 0 SS4END[7]
port 218 nsew signal input
flabel metal2 s 28088 10672 28168 10752 0 FreeSans 320 0 0 0 SS4END[8]
port 219 nsew signal input
flabel metal2 s 28280 10672 28360 10752 0 FreeSans 320 0 0 0 SS4END[9]
port 220 nsew signal input
flabel metal2 s 16760 0 16840 80 0 FreeSans 320 0 0 0 UserCLK
port 221 nsew signal input
flabel metal2 s 29624 10672 29704 10752 0 FreeSans 320 0 0 0 UserCLKo
port 222 nsew signal output
flabel metal6 s 4892 0 5332 10752 0 FreeSans 2624 90 0 0 VGND
port 223 nsew ground bidirectional
flabel metal6 s 4892 0 5332 328 0 FreeSans 2624 0 0 0 VGND
port 223 nsew ground bidirectional
flabel metal6 s 4892 10424 5332 10752 0 FreeSans 2624 0 0 0 VGND
port 223 nsew ground bidirectional
flabel metal6 s 20012 0 20452 10752 0 FreeSans 2624 90 0 0 VGND
port 223 nsew ground bidirectional
flabel metal6 s 20012 0 20452 328 0 FreeSans 2624 0 0 0 VGND
port 223 nsew ground bidirectional
flabel metal6 s 20012 10424 20452 10752 0 FreeSans 2624 0 0 0 VGND
port 223 nsew ground bidirectional
flabel metal6 s 35132 0 35572 10752 0 FreeSans 2624 90 0 0 VGND
port 223 nsew ground bidirectional
flabel metal6 s 35132 0 35572 328 0 FreeSans 2624 0 0 0 VGND
port 223 nsew ground bidirectional
flabel metal6 s 35132 10424 35572 10752 0 FreeSans 2624 0 0 0 VGND
port 223 nsew ground bidirectional
flabel metal6 s 3652 0 4092 10752 0 FreeSans 2624 90 0 0 VPWR
port 224 nsew power bidirectional
flabel metal6 s 3652 0 4092 328 0 FreeSans 2624 0 0 0 VPWR
port 224 nsew power bidirectional
flabel metal6 s 3652 10424 4092 10752 0 FreeSans 2624 0 0 0 VPWR
port 224 nsew power bidirectional
flabel metal6 s 18772 0 19212 10752 0 FreeSans 2624 90 0 0 VPWR
port 224 nsew power bidirectional
flabel metal6 s 18772 0 19212 328 0 FreeSans 2624 0 0 0 VPWR
port 224 nsew power bidirectional
flabel metal6 s 18772 10424 19212 10752 0 FreeSans 2624 0 0 0 VPWR
port 224 nsew power bidirectional
flabel metal6 s 33892 0 34332 10752 0 FreeSans 2624 90 0 0 VPWR
port 224 nsew power bidirectional
flabel metal6 s 33892 0 34332 328 0 FreeSans 2624 0 0 0 VPWR
port 224 nsew power bidirectional
flabel metal6 s 33892 10424 34332 10752 0 FreeSans 2624 0 0 0 VPWR
port 224 nsew power bidirectional
rlabel metal1 21504 9828 21504 9828 0 VGND
rlabel metal1 21504 9072 21504 9072 0 VPWR
rlabel metal2 4128 660 4128 660 0 A_I_top
rlabel metal2 33696 2058 33696 2058 0 A_O_top
rlabel metal2 5280 324 5280 324 0 A_T_top
rlabel metal2 7584 492 7584 492 0 B_I_top
rlabel metal2 31200 3990 31200 3990 0 B_O_top
rlabel metal2 8736 450 8736 450 0 B_T_top
rlabel metal2 11040 492 11040 492 0 C_I_top
rlabel metal2 29328 1932 29328 1932 0 C_O_top
rlabel metal2 12192 72 12192 72 0 C_T_top
rlabel metal2 19488 10176 19488 10176 0 Co
rlabel metal2 14496 2760 14496 2760 0 D_I_top
rlabel metal2 39216 1092 39216 1092 0 D_O_top
rlabel metal2 15648 114 15648 114 0 D_T_top
rlabel metal3 18576 1932 18576 1932 0 FrameData[0]
rlabel metal2 1584 2604 1584 2604 0 FrameData[10]
rlabel metal3 16608 1302 16608 1302 0 FrameData[11]
rlabel metal3 78 4116 78 4116 0 FrameData[12]
rlabel metal3 606 4452 606 4452 0 FrameData[13]
rlabel metal2 18912 3654 18912 3654 0 FrameData[14]
rlabel metal3 702 5124 702 5124 0 FrameData[15]
rlabel metal2 1296 4956 1296 4956 0 FrameData[16]
rlabel metal2 18144 5586 18144 5586 0 FrameData[17]
rlabel metal2 33312 4704 33312 4704 0 FrameData[18]
rlabel metal3 606 6468 606 6468 0 FrameData[19]
rlabel metal2 16224 1974 16224 1974 0 FrameData[1]
rlabel metal4 15456 5712 15456 5712 0 FrameData[20]
rlabel metal3 1290 7140 1290 7140 0 FrameData[21]
rlabel metal3 1584 5964 1584 5964 0 FrameData[22]
rlabel metal2 1728 7350 1728 7350 0 FrameData[23]
rlabel metal3 846 8148 846 8148 0 FrameData[24]
rlabel metal4 19584 6846 19584 6846 0 FrameData[25]
rlabel metal2 24768 1932 24768 1932 0 FrameData[26]
rlabel metal2 36096 9408 36096 9408 0 FrameData[27]
rlabel metal3 990 9492 990 9492 0 FrameData[28]
rlabel metal2 15168 9576 15168 9576 0 FrameData[29]
rlabel metal2 19488 798 19488 798 0 FrameData[2]
rlabel metal2 1632 9198 1632 9198 0 FrameData[30]
rlabel metal2 1920 7896 1920 7896 0 FrameData[31]
rlabel metal3 942 1092 942 1092 0 FrameData[3]
rlabel metal2 1920 1512 1920 1512 0 FrameData[4]
rlabel metal2 29376 1302 29376 1302 0 FrameData[5]
rlabel metal3 270 2100 270 2100 0 FrameData[6]
rlabel metal2 31872 3360 31872 3360 0 FrameData[7]
rlabel metal4 1344 3486 1344 3486 0 FrameData[8]
rlabel metal3 1182 3108 1182 3108 0 FrameData[9]
rlabel metal2 37920 1092 37920 1092 0 FrameData_O[0]
rlabel metal4 26448 3360 26448 3360 0 FrameData_O[10]
rlabel metal2 33696 5292 33696 5292 0 FrameData_O[11]
rlabel metal2 30048 6384 30048 6384 0 FrameData_O[12]
rlabel metal2 32352 5334 32352 5334 0 FrameData_O[13]
rlabel metal3 42018 4788 42018 4788 0 FrameData_O[14]
rlabel metal2 41520 4368 41520 4368 0 FrameData_O[15]
rlabel metal2 41376 5124 41376 5124 0 FrameData_O[16]
rlabel metal3 42210 5796 42210 5796 0 FrameData_O[17]
rlabel metal2 41088 6006 41088 6006 0 FrameData_O[18]
rlabel metal3 42210 6468 42210 6468 0 FrameData_O[19]
rlabel metal3 40722 420 40722 420 0 FrameData_O[1]
rlabel metal2 41088 6720 41088 6720 0 FrameData_O[20]
rlabel metal3 42306 7140 42306 7140 0 FrameData_O[21]
rlabel metal3 42018 7476 42018 7476 0 FrameData_O[22]
rlabel metal3 42210 7812 42210 7812 0 FrameData_O[23]
rlabel metal3 42258 8148 42258 8148 0 FrameData_O[24]
rlabel metal3 42114 8484 42114 8484 0 FrameData_O[25]
rlabel metal2 40032 6426 40032 6426 0 FrameData_O[26]
rlabel metal2 37920 8190 37920 8190 0 FrameData_O[27]
rlabel metal3 39840 4788 39840 4788 0 FrameData_O[28]
rlabel metal3 38784 5880 38784 5880 0 FrameData_O[29]
rlabel metal2 36768 1596 36768 1596 0 FrameData_O[2]
rlabel metal2 38208 6048 38208 6048 0 FrameData_O[30]
rlabel metal2 37536 6636 37536 6636 0 FrameData_O[31]
rlabel metal3 39714 1092 39714 1092 0 FrameData_O[3]
rlabel metal3 41634 1428 41634 1428 0 FrameData_O[4]
rlabel metal3 42066 1764 42066 1764 0 FrameData_O[5]
rlabel metal2 27264 2310 27264 2310 0 FrameData_O[6]
rlabel metal3 42738 2436 42738 2436 0 FrameData_O[7]
rlabel metal4 27648 3738 27648 3738 0 FrameData_O[8]
rlabel metal3 42354 3108 42354 3108 0 FrameData_O[9]
rlabel metal2 20736 1050 20736 1050 0 FrameStrobe[0]
rlabel via2 29472 72 29472 72 0 FrameStrobe[10]
rlabel via2 30624 72 30624 72 0 FrameStrobe[11]
rlabel metal2 31776 870 31776 870 0 FrameStrobe[12]
rlabel metal2 32928 954 32928 954 0 FrameStrobe[13]
rlabel metal2 34080 156 34080 156 0 FrameStrobe[14]
rlabel metal2 35232 324 35232 324 0 FrameStrobe[15]
rlabel metal2 36384 618 36384 618 0 FrameStrobe[16]
rlabel metal3 36672 3780 36672 3780 0 FrameStrobe[17]
rlabel metal2 38688 828 38688 828 0 FrameStrobe[18]
rlabel metal2 39840 282 39840 282 0 FrameStrobe[19]
rlabel metal3 22464 2352 22464 2352 0 FrameStrobe[1]
rlabel metal2 17184 966 17184 966 0 FrameStrobe[2]
rlabel metal2 20976 1932 20976 1932 0 FrameStrobe[3]
rlabel metal2 22560 72 22560 72 0 FrameStrobe[4]
rlabel metal2 23712 156 23712 156 0 FrameStrobe[5]
rlabel metal2 33024 672 33024 672 0 FrameStrobe[6]
rlabel metal2 26016 534 26016 534 0 FrameStrobe[7]
rlabel metal2 35232 1050 35232 1050 0 FrameStrobe[8]
rlabel metal2 28320 618 28320 618 0 FrameStrobe[9]
rlabel metal2 29856 9798 29856 9798 0 FrameStrobe_O[0]
rlabel metal2 30528 4368 30528 4368 0 FrameStrobe_O[10]
rlabel metal2 32544 7224 32544 7224 0 FrameStrobe_O[11]
rlabel metal3 33168 3612 33168 3612 0 FrameStrobe_O[12]
rlabel metal2 36960 4116 36960 4116 0 FrameStrobe_O[13]
rlabel metal2 39840 798 39840 798 0 FrameStrobe_O[14]
rlabel metal5 36816 924 36816 924 0 FrameStrobe_O[15]
rlabel metal2 39456 966 39456 966 0 FrameStrobe_O[16]
rlabel metal2 35424 7770 35424 7770 0 FrameStrobe_O[17]
rlabel metal2 31680 6300 31680 6300 0 FrameStrobe_O[18]
rlabel metal2 31248 5460 31248 5460 0 FrameStrobe_O[19]
rlabel metal2 30048 9756 30048 9756 0 FrameStrobe_O[1]
rlabel metal2 30432 8694 30432 8694 0 FrameStrobe_O[2]
rlabel metal2 30816 8568 30816 8568 0 FrameStrobe_O[3]
rlabel metal3 30144 8484 30144 8484 0 FrameStrobe_O[4]
rlabel metal2 32400 1260 32400 1260 0 FrameStrobe_O[5]
rlabel metal3 31200 840 31200 840 0 FrameStrobe_O[6]
rlabel metal2 31680 3318 31680 3318 0 FrameStrobe_O[7]
rlabel metal2 34896 924 34896 924 0 FrameStrobe_O[8]
rlabel metal2 32016 2856 32016 2856 0 FrameStrobe_O[9]
rlabel metal2 36000 2100 36000 2100 0 Inst_A_IO_1_bidirectional_frame_config_pass.Q
rlabel metal2 37632 2982 37632 2982 0 Inst_B_IO_1_bidirectional_frame_config_pass.Q
rlabel metal2 14688 8484 14688 8484 0 Inst_C_IO_1_bidirectional_frame_config_pass.Q
rlabel metal2 36864 7896 36864 7896 0 Inst_D_IO_1_bidirectional_frame_config_pass.Q
rlabel metal2 16128 2100 16128 2100 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit0.Q
rlabel metal2 17904 2100 17904 2100 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit1.Q
rlabel metal2 2976 2982 2976 2982 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit10.Q
rlabel metal3 12672 1932 12672 1932 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit11.Q
rlabel metal3 11856 2604 11856 2604 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit12.Q
rlabel metal2 12480 1176 12480 1176 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit13.Q
rlabel metal3 12096 3402 12096 3402 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit14.Q
rlabel metal2 2976 4914 2976 4914 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit15.Q
rlabel via2 4512 4953 4512 4953 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit16.Q
rlabel metal2 4896 4452 4896 4452 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit17.Q
rlabel metal3 6912 4704 6912 4704 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit18.Q
rlabel metal2 9696 7056 9696 7056 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit19.Q
rlabel metal3 20736 1344 20736 1344 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit2.Q
rlabel metal2 7296 4914 7296 4914 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit20.Q
rlabel metal2 10224 6636 10224 6636 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit21.Q
rlabel metal3 3312 6468 3312 6468 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 4368 7140 4368 7140 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit23.Q
rlabel metal2 3936 5712 3936 5712 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit24.Q
rlabel metal3 7920 7980 7920 7980 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit25.Q
rlabel metal2 6432 6384 6432 6384 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit26.Q
rlabel metal2 8832 8694 8832 8694 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit27.Q
rlabel metal2 8352 9576 8352 9576 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit28.Q
rlabel metal2 2112 8694 2112 8694 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit29.Q
rlabel metal2 19104 1302 19104 1302 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit3.Q
rlabel via2 4416 8654 4416 8654 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit30.Q
rlabel metal2 1920 8400 1920 8400 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit31.Q
rlabel metal2 3408 1932 3408 1932 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit4.Q
rlabel metal2 6144 2142 6144 2142 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit5.Q
rlabel metal2 6912 1134 6912 1134 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit6.Q
rlabel metal3 4896 1680 4896 1680 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit7.Q
rlabel metal2 1488 1092 1488 1092 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit8.Q
rlabel metal2 1728 3696 1728 3696 0 Inst_S_IO4_ConfigMem.Inst_frame0_bit9.Q
rlabel metal2 13920 3612 13920 3612 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit0.Q
rlabel metal2 16224 3990 16224 3990 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit1.Q
rlabel metal2 37728 6720 37728 6720 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit10.Q
rlabel metal2 39744 5040 39744 5040 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit11.Q
rlabel metal2 14160 2100 14160 2100 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit12.Q
rlabel metal2 15456 1512 15456 1512 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit13.Q
rlabel metal2 21504 3696 21504 3696 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit14.Q
rlabel metal2 22992 4179 22992 4179 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit15.Q
rlabel metal2 14112 6678 14112 6678 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit16.Q
rlabel metal3 12912 6636 12912 6636 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit17.Q
rlabel metal2 12384 4998 12384 4998 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit18.Q
rlabel metal2 13632 4410 13632 4410 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit19.Q
rlabel metal2 24528 1344 24528 1344 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit2.Q
rlabel metal2 38880 6216 38880 6216 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit20.Q
rlabel metal3 40704 5124 40704 5124 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit21.Q
rlabel metal2 24096 7602 24096 7602 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit22.Q
rlabel metal2 25536 8400 25536 8400 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit23.Q
rlabel metal2 24000 6510 24000 6510 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit24.Q
rlabel metal2 25824 6167 25824 6167 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit25.Q
rlabel metal3 39360 7980 39360 7980 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit26.Q
rlabel metal3 40896 7392 40896 7392 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit27.Q
rlabel metal2 18144 9240 18144 9240 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit28.Q
rlabel metal2 16416 8946 16416 8946 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit29.Q
rlabel metal2 26112 1971 26112 1971 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit3.Q
rlabel metal2 37824 8946 37824 8946 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit30.Q
rlabel metal2 39360 8701 39360 8701 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit31.Q
rlabel metal3 24432 4284 24432 4284 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit4.Q
rlabel metal3 26400 2856 26400 2856 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit5.Q
rlabel metal3 39504 3612 39504 3612 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit6.Q
rlabel metal3 41136 2772 41136 2772 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit7.Q
rlabel metal2 14016 3864 14016 3864 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit8.Q
rlabel metal2 15744 4795 15744 4795 0 Inst_S_IO4_ConfigMem.Inst_frame1_bit9.Q
rlabel metal3 17952 4956 17952 4956 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit0.Q
rlabel metal2 16800 4158 16800 4158 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit1.Q
rlabel metal2 37632 3864 37632 3864 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit10.Q
rlabel metal2 36384 3066 36384 3066 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit11.Q
rlabel metal2 33216 2184 33216 2184 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit12.Q
rlabel metal2 34848 1680 34848 1680 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit13.Q
rlabel metal2 35712 3948 35712 3948 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit14.Q
rlabel via1 37104 4951 37104 4951 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit15.Q
rlabel metal2 17952 6510 17952 6510 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit16.Q
rlabel metal2 19632 5880 19632 5880 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit17.Q
rlabel metal2 34320 4179 34320 4179 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit18.Q
rlabel metal2 32736 4410 32736 4410 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit19.Q
rlabel metal3 22992 2604 22992 2604 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit2.Q
rlabel metal2 27504 5880 27504 5880 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit20.Q
rlabel metal2 26208 7518 26208 7518 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit21.Q
rlabel metal2 33504 7686 33504 7686 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit22.Q
rlabel metal3 31680 7392 31680 7392 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit23.Q
rlabel metal2 35088 6468 35088 6468 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit24.Q
rlabel metal3 36864 5880 36864 5880 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit25.Q
rlabel metal2 35760 8148 35760 8148 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit26.Q
rlabel via1 37392 8656 37392 8656 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit27.Q
rlabel metal2 21792 8946 21792 8946 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit28.Q
rlabel metal2 23328 8953 23328 8953 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit29.Q
rlabel metal2 24768 1260 24768 1260 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit3.Q
rlabel metal2 33312 8946 33312 8946 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit30.Q
rlabel metal2 34848 8953 34848 8953 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit31.Q
rlabel metal2 29568 1386 29568 1386 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit4.Q
rlabel metal2 27984 1344 27984 1344 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit5.Q
rlabel metal2 32064 3654 32064 3654 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit6.Q
rlabel metal2 30048 3318 30048 3318 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit7.Q
rlabel metal2 34944 6132 34944 6132 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit8.Q
rlabel metal2 33312 5418 33312 5418 0 Inst_S_IO4_ConfigMem.Inst_frame2_bit9.Q
rlabel metal2 19296 2226 19296 2226 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit0.Q
rlabel metal3 19488 3612 19488 3612 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit1.Q
rlabel metal2 27744 6090 27744 6090 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit10.Q
rlabel metal2 29376 6932 29376 6932 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit11.Q
rlabel metal2 18816 4368 18816 4368 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit12.Q
rlabel metal2 20640 5376 20640 5376 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit13.Q
rlabel metal2 26832 3612 26832 3612 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit14.Q
rlabel metal2 28608 3654 28608 3654 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit15.Q
rlabel metal2 16032 6510 16032 6510 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit16.Q
rlabel metal2 17568 6717 17568 6717 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit17.Q
rlabel metal2 23904 3612 23904 3612 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit18.Q
rlabel metal2 25392 4893 25392 4893 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit19.Q
rlabel metal2 20880 2100 20880 2100 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit2.Q
rlabel metal2 29376 6167 29376 6167 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit20.Q
rlabel metal2 27840 6510 27840 6510 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit21.Q
rlabel via1 31440 6463 31440 6463 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit22.Q
rlabel metal2 29856 6762 29856 6762 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit23.Q
rlabel metal2 22608 7392 22608 7392 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit24.Q
rlabel metal2 21024 8820 21024 8820 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit25.Q
rlabel metal2 30528 8785 30528 8785 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit26.Q
rlabel metal2 32064 8946 32064 8946 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit27.Q
rlabel metal2 19392 8232 19392 8232 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit28.Q
rlabel metal2 17760 8190 17760 8190 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit29.Q
rlabel metal2 22560 1680 22560 1680 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit3.Q
rlabel metal2 26976 8988 26976 8988 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit30.Q
rlabel via2 28416 7977 28416 7977 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit31.Q
rlabel metal2 27696 1260 27696 1260 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit4.Q
rlabel metal3 29664 2100 29664 2100 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit5.Q
rlabel metal2 29184 4662 29184 4662 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit6.Q
rlabel metal2 30480 3612 30480 3612 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit7.Q
rlabel metal2 21264 5880 21264 5880 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit8.Q
rlabel metal2 22848 6923 22848 6923 0 Inst_S_IO4_ConfigMem.Inst_frame3_bit9.Q
rlabel metal2 11040 7686 11040 7686 0 Inst_S_IO4_ConfigMem.Inst_frame4_bit28.Q
rlabel metal3 12864 8022 12864 8022 0 Inst_S_IO4_ConfigMem.Inst_frame4_bit29.Q
rlabel metal2 15744 8610 15744 8610 0 Inst_S_IO4_ConfigMem.Inst_frame4_bit30.Q
rlabel metal2 14064 8148 14064 8148 0 Inst_S_IO4_ConfigMem.Inst_frame4_bit31.Q
rlabel metal2 11136 8358 11136 8358 0 Inst_S_IO4_switch_matrix.N1BEG0
rlabel metal2 14016 8400 14016 8400 0 Inst_S_IO4_switch_matrix.N1BEG1
rlabel metal2 17856 8820 17856 8820 0 Inst_S_IO4_switch_matrix.N1BEG2
rlabel metal4 16416 5586 16416 5586 0 Inst_S_IO4_switch_matrix.N1BEG3
rlabel metal5 20112 1764 20112 1764 0 Inst_S_IO4_switch_matrix.N2BEG0
rlabel metal4 30912 4914 30912 4914 0 Inst_S_IO4_switch_matrix.N2BEG1
rlabel metal4 13824 8106 13824 8106 0 Inst_S_IO4_switch_matrix.N2BEG2
rlabel metal2 29568 6888 29568 6888 0 Inst_S_IO4_switch_matrix.N2BEG3
rlabel metal2 11424 7644 11424 7644 0 Inst_S_IO4_switch_matrix.N2BEG4
rlabel metal4 15936 4578 15936 4578 0 Inst_S_IO4_switch_matrix.N2BEG5
rlabel metal2 17760 7014 17760 7014 0 Inst_S_IO4_switch_matrix.N2BEG6
rlabel metal3 12096 5166 12096 5166 0 Inst_S_IO4_switch_matrix.N2BEG7
rlabel metal4 24576 1596 24576 1596 0 Inst_S_IO4_switch_matrix.N2BEGb0
rlabel metal4 31584 6930 31584 6930 0 Inst_S_IO4_switch_matrix.N2BEGb1
rlabel metal3 14016 8484 14016 8484 0 Inst_S_IO4_switch_matrix.N2BEGb2
rlabel metal3 19872 5250 19872 5250 0 Inst_S_IO4_switch_matrix.N2BEGb3
rlabel metal3 16080 8736 16080 8736 0 Inst_S_IO4_switch_matrix.N2BEGb4
rlabel metal5 19392 588 19392 588 0 Inst_S_IO4_switch_matrix.N2BEGb5
rlabel metal3 16800 4998 16800 4998 0 Inst_S_IO4_switch_matrix.N2BEGb6
rlabel metal2 25056 2940 25056 2940 0 Inst_S_IO4_switch_matrix.N2BEGb7
rlabel metal4 29952 1596 29952 1596 0 Inst_S_IO4_switch_matrix.N4BEG0
rlabel metal3 32784 4872 32784 4872 0 Inst_S_IO4_switch_matrix.N4BEG1
rlabel metal3 36624 6636 36624 6636 0 Inst_S_IO4_switch_matrix.N4BEG10
rlabel metal2 37536 8190 37536 8190 0 Inst_S_IO4_switch_matrix.N4BEG11
rlabel metal2 23472 7896 23472 7896 0 Inst_S_IO4_switch_matrix.N4BEG12
rlabel metal3 34464 7896 34464 7896 0 Inst_S_IO4_switch_matrix.N4BEG13
rlabel metal2 16416 5040 16416 5040 0 Inst_S_IO4_switch_matrix.N4BEG14
rlabel metal3 25152 2058 25152 2058 0 Inst_S_IO4_switch_matrix.N4BEG15
rlabel metal2 34752 7686 34752 7686 0 Inst_S_IO4_switch_matrix.N4BEG2
rlabel metal2 37728 3654 37728 3654 0 Inst_S_IO4_switch_matrix.N4BEG3
rlabel metal2 34560 3150 34560 3150 0 Inst_S_IO4_switch_matrix.N4BEG4
rlabel metal2 37296 5124 37296 5124 0 Inst_S_IO4_switch_matrix.N4BEG5
rlabel metal3 15168 9408 15168 9408 0 Inst_S_IO4_switch_matrix.N4BEG6
rlabel metal2 35136 4704 35136 4704 0 Inst_S_IO4_switch_matrix.N4BEG7
rlabel metal3 27456 9408 27456 9408 0 Inst_S_IO4_switch_matrix.N4BEG8
rlabel metal2 33216 8442 33216 8442 0 Inst_S_IO4_switch_matrix.N4BEG9
rlabel metal2 17280 4074 17280 4074 0 Inst_S_IO4_switch_matrix.NN4BEG0
rlabel metal2 41760 4452 41760 4452 0 Inst_S_IO4_switch_matrix.NN4BEG1
rlabel metal2 25776 6636 25776 6636 0 Inst_S_IO4_switch_matrix.NN4BEG10
rlabel metal2 32544 8568 32544 8568 0 Inst_S_IO4_switch_matrix.NN4BEG11
rlabel metal2 18624 9156 18624 9156 0 Inst_S_IO4_switch_matrix.NN4BEG12
rlabel metal2 38304 8190 38304 8190 0 Inst_S_IO4_switch_matrix.NN4BEG13
rlabel metal2 18336 3696 18336 3696 0 Inst_S_IO4_switch_matrix.NN4BEG14
rlabel metal2 20448 2457 20448 2457 0 Inst_S_IO4_switch_matrix.NN4BEG15
rlabel metal2 16320 4074 16320 4074 0 Inst_S_IO4_switch_matrix.NN4BEG2
rlabel metal2 39456 7098 39456 7098 0 Inst_S_IO4_switch_matrix.NN4BEG3
rlabel metal2 16032 2520 16032 2520 0 Inst_S_IO4_switch_matrix.NN4BEG4
rlabel metal2 23520 4452 23520 4452 0 Inst_S_IO4_switch_matrix.NN4BEG5
rlabel metal3 15312 7224 15312 7224 0 Inst_S_IO4_switch_matrix.NN4BEG6
rlabel metal3 13872 5040 13872 5040 0 Inst_S_IO4_switch_matrix.NN4BEG7
rlabel metal2 40464 6384 40464 6384 0 Inst_S_IO4_switch_matrix.NN4BEG8
rlabel metal2 25248 9198 25248 9198 0 Inst_S_IO4_switch_matrix.NN4BEG9
rlabel metal2 9456 9660 9456 9660 0 N1BEG[0]
rlabel metal2 9744 9660 9744 9660 0 N1BEG[1]
rlabel metal2 10032 9660 10032 9660 0 N1BEG[2]
rlabel metal3 10080 8820 10080 8820 0 N1BEG[3]
rlabel metal2 12240 5880 12240 5880 0 N2BEG[0]
rlabel metal2 10320 8484 10320 8484 0 N2BEG[1]
rlabel metal2 10656 9756 10656 9756 0 N2BEG[2]
rlabel metal2 10848 9756 10848 9756 0 N2BEG[3]
rlabel metal2 11184 8820 11184 8820 0 N2BEG[4]
rlabel metal2 11520 7770 11520 7770 0 N2BEG[5]
rlabel metal2 11424 10260 11424 10260 0 N2BEG[6]
rlabel metal2 11904 7014 11904 7014 0 N2BEG[7]
rlabel metal2 11808 9840 11808 9840 0 N2BEGb[0]
rlabel metal2 12672 7476 12672 7476 0 N2BEGb[1]
rlabel metal2 11856 8820 11856 8820 0 N2BEGb[2]
rlabel metal2 12672 9828 12672 9828 0 N2BEGb[3]
rlabel metal2 12192 9492 12192 9492 0 N2BEGb[4]
rlabel metal2 13056 9828 13056 9828 0 N2BEGb[5]
rlabel metal2 13200 5880 13200 5880 0 N2BEGb[6]
rlabel metal3 13632 3612 13632 3612 0 N2BEGb[7]
rlabel metal2 13584 1260 13584 1260 0 N4BEG[0]
rlabel metal2 15264 10428 15264 10428 0 N4BEG[10]
rlabel metal5 26448 2100 26448 2100 0 N4BEG[11]
rlabel metal2 15648 10050 15648 10050 0 N4BEG[12]
rlabel metal2 15840 10596 15840 10596 0 N4BEG[13]
rlabel metal2 16176 5460 16176 5460 0 N4BEG[14]
rlabel metal2 16416 4242 16416 4242 0 N4BEG[15]
rlabel metal4 19488 756 19488 756 0 N4BEG[1]
rlabel metal5 24048 1008 24048 1008 0 N4BEG[2]
rlabel metal2 13920 10302 13920 10302 0 N4BEG[3]
rlabel metal5 26736 2016 26736 2016 0 N4BEG[4]
rlabel metal2 14304 9756 14304 9756 0 N4BEG[5]
rlabel metal2 14640 9660 14640 9660 0 N4BEG[6]
rlabel metal2 14688 10638 14688 10638 0 N4BEG[7]
rlabel metal2 14880 10218 14880 10218 0 N4BEG[8]
rlabel metal2 15072 9756 15072 9756 0 N4BEG[9]
rlabel metal2 17088 4494 17088 4494 0 NN4BEG[0]
rlabel metal2 18336 10134 18336 10134 0 NN4BEG[10]
rlabel metal2 18528 10260 18528 10260 0 NN4BEG[11]
rlabel metal2 18768 9660 18768 9660 0 NN4BEG[12]
rlabel metal2 18912 9966 18912 9966 0 NN4BEG[13]
rlabel metal2 19152 4788 19152 4788 0 NN4BEG[14]
rlabel metal2 19296 10050 19296 10050 0 NN4BEG[15]
rlabel metal2 16608 10092 16608 10092 0 NN4BEG[1]
rlabel metal3 16608 4368 16608 4368 0 NN4BEG[2]
rlabel metal2 16992 9882 16992 9882 0 NN4BEG[3]
rlabel metal2 16320 3066 16320 3066 0 NN4BEG[4]
rlabel metal2 17376 10092 17376 10092 0 NN4BEG[5]
rlabel metal2 15744 7434 15744 7434 0 NN4BEG[6]
rlabel metal2 13776 5880 13776 5880 0 NN4BEG[7]
rlabel metal2 17952 10134 17952 10134 0 NN4BEG[8]
rlabel metal2 18144 10596 18144 10596 0 NN4BEG[9]
rlabel metal2 19680 9756 19680 9756 0 S1END[0]
rlabel metal2 19872 9462 19872 9462 0 S1END[1]
rlabel metal2 15264 9366 15264 9366 0 S1END[2]
rlabel metal2 12288 9282 12288 9282 0 S1END[3]
rlabel metal2 14304 2856 14304 2856 0 S2END[0]
rlabel metal2 18432 4452 18432 4452 0 S2END[1]
rlabel metal2 14688 3360 14688 3360 0 S2END[2]
rlabel metal2 18528 8148 18528 8148 0 S2END[3]
rlabel metal2 12000 2058 12000 2058 0 S2END[4]
rlabel metal2 2496 7854 2496 7854 0 S2END[5]
rlabel metal2 13200 1092 13200 1092 0 S2END[6]
rlabel metal2 14688 4242 14688 4242 0 S2END[7]
rlabel metal2 16704 2730 16704 2730 0 S2MID[0]
rlabel metal2 16128 6888 16128 6888 0 S2MID[1]
rlabel metal2 13440 7014 13440 7014 0 S2MID[2]
rlabel metal2 19296 2646 19296 2646 0 S2MID[3]
rlabel metal2 17664 7056 17664 7056 0 S2MID[4]
rlabel metal2 19392 3654 19392 3654 0 S2MID[5]
rlabel metal2 13824 7266 13824 7266 0 S2MID[6]
rlabel metal2 12960 4452 12960 4452 0 S2MID[7]
rlabel metal2 24144 6468 24144 6468 0 S4END[0]
rlabel via2 25440 10680 25440 10680 0 S4END[10]
rlabel metal2 33120 6510 33120 6510 0 S4END[11]
rlabel metal2 31680 8190 31680 8190 0 S4END[12]
rlabel metal2 26016 9672 26016 9672 0 S4END[13]
rlabel metal2 30816 4368 30816 4368 0 S4END[14]
rlabel metal2 26478 3696 26478 3696 0 S4END[15]
rlabel metal2 16512 8862 16512 8862 0 S4END[1]
rlabel metal2 24480 7014 24480 7014 0 S4END[2]
rlabel metal2 19008 8568 19008 8568 0 S4END[3]
rlabel metal2 33408 8610 33408 8610 0 S4END[4]
rlabel metal2 21792 8232 21792 8232 0 S4END[5]
rlabel metal2 30432 7182 30432 7182 0 S4END[6]
rlabel metal2 32976 2604 32976 2604 0 S4END[7]
rlabel metal2 35904 9618 35904 9618 0 S4END[8]
rlabel metal2 35232 6552 35232 6552 0 S4END[9]
rlabel metal2 25008 1932 25008 1932 0 SS4END[0]
rlabel metal2 36576 4410 36576 4410 0 SS4END[10]
rlabel metal2 19488 8232 19488 8232 0 SS4END[11]
rlabel metal2 32064 8232 32064 8232 0 SS4END[12]
rlabel metal3 26496 8778 26496 8778 0 SS4END[13]
rlabel metal2 30864 6468 30864 6468 0 SS4END[14]
rlabel metal2 28944 6468 28944 6468 0 SS4END[15]
rlabel metal3 17184 6384 17184 6384 0 SS4END[1]
rlabel metal2 27456 8022 27456 8022 0 SS4END[2]
rlabel metal2 18912 8778 18912 8778 0 SS4END[3]
rlabel metal2 31584 8442 31584 8442 0 SS4END[4]
rlabel metal2 21696 9576 21696 9576 0 SS4END[5]
rlabel metal3 29376 4830 29376 4830 0 SS4END[6]
rlabel metal3 28416 2688 28416 2688 0 SS4END[7]
rlabel metal3 31680 7602 31680 7602 0 SS4END[8]
rlabel metal3 17376 6468 17376 6468 0 SS4END[9]
rlabel metal2 16800 660 16800 660 0 UserCLK
rlabel metal2 36576 1386 36576 1386 0 UserCLK_regs
rlabel metal2 29520 2856 29520 2856 0 UserCLKo
rlabel metal2 6144 3780 6144 3780 0 _000_
rlabel metal3 9792 3612 9792 3612 0 _001_
rlabel metal2 10560 5670 10560 5670 0 _002_
rlabel metal2 11520 1134 11520 1134 0 _003_
rlabel metal2 3120 2520 3120 2520 0 _004_
rlabel metal3 4128 798 4128 798 0 _005_
rlabel metal2 5376 6720 5376 6720 0 _006_
rlabel metal2 8640 4116 8640 4116 0 _007_
rlabel metal3 5760 4116 5760 4116 0 _008_
rlabel metal2 4752 5124 4752 5124 0 _009_
rlabel metal2 5232 4116 5232 4116 0 _010_
rlabel metal2 4800 3696 4800 3696 0 _011_
rlabel metal2 4704 3696 4704 3696 0 _012_
rlabel metal2 5328 4368 5328 4368 0 _013_
rlabel metal2 3840 5754 3840 5754 0 _014_
rlabel metal2 4992 6552 4992 6552 0 _015_
rlabel metal2 4320 5922 4320 5922 0 _016_
rlabel metal2 4128 5628 4128 5628 0 _017_
rlabel metal2 5088 6384 5088 6384 0 _018_
rlabel metal2 2160 8484 2160 8484 0 _019_
rlabel metal2 4416 7896 4416 7896 0 _020_
rlabel metal2 4848 9492 4848 9492 0 _021_
rlabel metal2 1824 8232 1824 8232 0 _022_
rlabel metal2 4128 8169 4128 8169 0 _023_
rlabel metal2 7584 7434 7584 7434 0 _024_
rlabel metal2 7680 8400 7680 8400 0 _025_
rlabel metal2 7440 7392 7440 7392 0 _026_
rlabel metal3 7536 6468 7536 6468 0 _027_
rlabel metal2 8256 6510 8256 6510 0 _028_
rlabel metal2 8400 6636 8400 6636 0 _029_
rlabel via1 7106 9492 7106 9492 0 _030_
rlabel metal2 6912 9576 6912 9576 0 _031_
rlabel metal3 6336 9492 6336 9492 0 _032_
rlabel metal2 8640 8190 8640 8190 0 _033_
rlabel metal2 8736 8358 8736 8358 0 _034_
rlabel metal2 8544 8610 8544 8610 0 _035_
rlabel metal3 8832 8148 8832 8148 0 _036_
rlabel metal3 9168 9492 9168 9492 0 _037_
rlabel metal2 8976 9660 8976 9660 0 _038_
rlabel metal2 9840 7140 9840 7140 0 _039_
rlabel metal2 8784 5628 8784 5628 0 _040_
rlabel metal2 10176 5544 10176 5544 0 _041_
rlabel metal2 10018 5677 10018 5677 0 _042_
rlabel metal2 10272 4662 10272 4662 0 _043_
rlabel metal2 10272 5376 10272 5376 0 _044_
rlabel metal3 10272 6468 10272 6468 0 _045_
rlabel metal2 10464 5922 10464 5922 0 _046_
rlabel metal3 10752 5880 10752 5880 0 _047_
rlabel metal2 7872 4620 7872 4620 0 _048_
rlabel metal2 7392 4746 7392 4746 0 _049_
rlabel metal2 8352 5082 8352 5082 0 _050_
rlabel metal2 7728 3192 7728 3192 0 _051_
rlabel metal3 9888 5040 9888 5040 0 _052_
rlabel metal2 11232 2184 11232 2184 0 _053_
rlabel metal2 11424 1386 11424 1386 0 _054_
rlabel metal2 12672 966 12672 966 0 _055_
rlabel metal3 12720 1092 12720 1092 0 _056_
rlabel metal3 12048 1092 12048 1092 0 _057_
rlabel metal2 11904 1176 11904 1176 0 _058_
rlabel metal2 12000 1302 12000 1302 0 _059_
rlabel metal3 11430 3444 11430 3444 0 _060_
rlabel metal2 11616 2772 11616 2772 0 _061_
rlabel metal2 12192 3360 12192 3360 0 _062_
rlabel metal2 12192 3024 12192 3024 0 _063_
rlabel metal2 6288 2436 6288 2436 0 _064_
rlabel metal2 6048 2016 6048 2016 0 _065_
rlabel metal2 5856 2562 5856 2562 0 _066_
rlabel metal2 5952 2352 5952 2352 0 _067_
rlabel metal2 6768 2100 6768 2100 0 _068_
rlabel metal2 6672 924 6672 924 0 _069_
rlabel metal2 3264 2058 3264 2058 0 _070_
rlabel metal2 5520 4116 5520 4116 0 _071_
rlabel metal2 3888 1932 3888 1932 0 _072_
rlabel metal2 7008 1470 7008 1470 0 _073_
rlabel metal2 3552 2142 3552 2142 0 _074_
rlabel metal2 7680 1092 7680 1092 0 _075_
rlabel metal2 7488 1344 7488 1344 0 _076_
rlabel metal3 6528 1092 6528 1092 0 _077_
rlabel metal2 7632 2352 7632 2352 0 _078_
rlabel metal2 40224 1302 40224 1302 0 _079_
rlabel metal3 40080 2268 40080 2268 0 _080_
rlabel metal2 40608 1512 40608 1512 0 _081_
rlabel metal2 41424 9324 41424 9324 0 _082_
rlabel metal2 31296 1176 31296 1176 0 clknet_0_UserCLK
rlabel metal3 38544 1260 38544 1260 0 clknet_0_UserCLK_regs
rlabel metal3 30720 1344 30720 1344 0 clknet_1_0__leaf_UserCLK
rlabel metal3 36384 1932 36384 1932 0 clknet_1_0__leaf_UserCLK_regs
rlabel metal3 40032 2100 40032 2100 0 clknet_1_1__leaf_UserCLK_regs
<< properties >>
string FIXED_BBOX 0 0 43008 10752
<< end >>
