module SW_term (UserCLK,
    UserCLKo,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N2BEG,
    N2BEGb,
    N4BEG,
    S1END,
    S2END,
    S2MID,
    S4END);
 input UserCLK;
 output UserCLKo;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 output [15:0] N4BEG;
 input [3:0] S1END;
 input [7:0] S2END;
 input [7:0] S2MID;
 input [15:0] S4END;


 sg13g2_buf_1 _00_ (.A(FrameData[0]),
    .X(FrameData_O[0]));
 sg13g2_buf_1 _01_ (.A(FrameData[1]),
    .X(FrameData_O[1]));
 sg13g2_buf_1 _02_ (.A(FrameData[2]),
    .X(FrameData_O[2]));
 sg13g2_buf_1 _03_ (.A(FrameData[3]),
    .X(FrameData_O[3]));
 sg13g2_buf_1 _04_ (.A(FrameData[4]),
    .X(FrameData_O[4]));
 sg13g2_buf_1 _05_ (.A(FrameData[5]),
    .X(FrameData_O[5]));
 sg13g2_buf_1 _06_ (.A(FrameData[6]),
    .X(FrameData_O[6]));
 sg13g2_buf_1 _07_ (.A(FrameData[7]),
    .X(FrameData_O[7]));
 sg13g2_buf_1 _08_ (.A(FrameData[8]),
    .X(FrameData_O[8]));
 sg13g2_buf_1 _09_ (.A(FrameData[9]),
    .X(FrameData_O[9]));
 sg13g2_buf_1 _10_ (.A(FrameData[10]),
    .X(FrameData_O[10]));
 sg13g2_buf_1 _11_ (.A(FrameData[11]),
    .X(FrameData_O[11]));
 sg13g2_buf_1 _12_ (.A(FrameData[12]),
    .X(FrameData_O[12]));
 sg13g2_buf_1 _13_ (.A(FrameData[13]),
    .X(FrameData_O[13]));
 sg13g2_buf_1 _14_ (.A(FrameData[14]),
    .X(FrameData_O[14]));
 sg13g2_buf_1 _15_ (.A(FrameData[15]),
    .X(FrameData_O[15]));
 sg13g2_buf_1 _16_ (.A(FrameData[16]),
    .X(FrameData_O[16]));
 sg13g2_buf_1 _17_ (.A(FrameData[17]),
    .X(FrameData_O[17]));
 sg13g2_buf_1 _18_ (.A(FrameData[18]),
    .X(FrameData_O[18]));
 sg13g2_buf_1 _19_ (.A(FrameData[19]),
    .X(FrameData_O[19]));
 sg13g2_buf_1 _20_ (.A(FrameData[20]),
    .X(FrameData_O[20]));
 sg13g2_buf_1 _21_ (.A(FrameData[21]),
    .X(FrameData_O[21]));
 sg13g2_buf_1 _22_ (.A(FrameData[22]),
    .X(FrameData_O[22]));
 sg13g2_buf_1 _23_ (.A(FrameData[23]),
    .X(FrameData_O[23]));
 sg13g2_buf_1 _24_ (.A(FrameData[24]),
    .X(FrameData_O[24]));
 sg13g2_buf_1 _25_ (.A(FrameData[25]),
    .X(FrameData_O[25]));
 sg13g2_buf_1 _26_ (.A(FrameData[26]),
    .X(FrameData_O[26]));
 sg13g2_buf_1 _27_ (.A(FrameData[27]),
    .X(FrameData_O[27]));
 sg13g2_buf_1 _28_ (.A(FrameData[28]),
    .X(FrameData_O[28]));
 sg13g2_buf_1 _29_ (.A(FrameData[29]),
    .X(FrameData_O[29]));
 sg13g2_buf_1 _30_ (.A(FrameData[30]),
    .X(FrameData_O[30]));
 sg13g2_buf_1 _31_ (.A(FrameData[31]),
    .X(FrameData_O[31]));
 sg13g2_buf_1 _32_ (.A(FrameStrobe[0]),
    .X(FrameStrobe_O[0]));
 sg13g2_buf_1 _33_ (.A(FrameStrobe[1]),
    .X(FrameStrobe_O[1]));
 sg13g2_buf_1 _34_ (.A(FrameStrobe[2]),
    .X(FrameStrobe_O[2]));
 sg13g2_buf_1 _35_ (.A(FrameStrobe[3]),
    .X(FrameStrobe_O[3]));
 sg13g2_buf_1 _36_ (.A(FrameStrobe[4]),
    .X(FrameStrobe_O[4]));
 sg13g2_buf_1 _37_ (.A(FrameStrobe[5]),
    .X(FrameStrobe_O[5]));
 sg13g2_buf_1 _38_ (.A(FrameStrobe[6]),
    .X(FrameStrobe_O[6]));
 sg13g2_buf_1 _39_ (.A(FrameStrobe[7]),
    .X(FrameStrobe_O[7]));
 sg13g2_buf_1 _40_ (.A(FrameStrobe[8]),
    .X(FrameStrobe_O[8]));
 sg13g2_buf_1 _41_ (.A(FrameStrobe[9]),
    .X(FrameStrobe_O[9]));
 sg13g2_buf_1 _42_ (.A(FrameStrobe[10]),
    .X(FrameStrobe_O[10]));
 sg13g2_buf_1 _43_ (.A(FrameStrobe[11]),
    .X(FrameStrobe_O[11]));
 sg13g2_buf_1 _44_ (.A(FrameStrobe[12]),
    .X(FrameStrobe_O[12]));
 sg13g2_buf_1 _45_ (.A(FrameStrobe[13]),
    .X(FrameStrobe_O[13]));
 sg13g2_buf_1 _46_ (.A(FrameStrobe[14]),
    .X(FrameStrobe_O[14]));
 sg13g2_buf_1 _47_ (.A(FrameStrobe[15]),
    .X(FrameStrobe_O[15]));
 sg13g2_buf_1 _48_ (.A(FrameStrobe[16]),
    .X(FrameStrobe_O[16]));
 sg13g2_buf_1 _49_ (.A(FrameStrobe[17]),
    .X(FrameStrobe_O[17]));
 sg13g2_buf_1 _50_ (.A(FrameStrobe[18]),
    .X(FrameStrobe_O[18]));
 sg13g2_buf_1 _51_ (.A(FrameStrobe[19]),
    .X(FrameStrobe_O[19]));
 sg13g2_buf_1 _52_ (.A(S1END[3]),
    .X(N1BEG[0]));
 sg13g2_buf_1 _53_ (.A(S1END[2]),
    .X(N1BEG[1]));
 sg13g2_buf_1 _54_ (.A(S1END[1]),
    .X(N1BEG[2]));
 sg13g2_buf_1 _55_ (.A(S1END[0]),
    .X(N1BEG[3]));
 sg13g2_buf_1 _56_ (.A(S2MID[7]),
    .X(N2BEG[0]));
 sg13g2_buf_1 _57_ (.A(S2MID[6]),
    .X(N2BEG[1]));
 sg13g2_buf_1 _58_ (.A(S2MID[5]),
    .X(N2BEG[2]));
 sg13g2_buf_1 _59_ (.A(S2MID[4]),
    .X(N2BEG[3]));
 sg13g2_buf_1 _60_ (.A(S2MID[3]),
    .X(N2BEG[4]));
 sg13g2_buf_1 _61_ (.A(S2MID[2]),
    .X(N2BEG[5]));
 sg13g2_buf_1 _62_ (.A(S2MID[1]),
    .X(N2BEG[6]));
 sg13g2_buf_1 _63_ (.A(S2MID[0]),
    .X(N2BEG[7]));
 sg13g2_buf_1 _64_ (.A(S2END[7]),
    .X(N2BEGb[0]));
 sg13g2_buf_1 _65_ (.A(S2END[6]),
    .X(N2BEGb[1]));
 sg13g2_buf_1 _66_ (.A(S2END[5]),
    .X(N2BEGb[2]));
 sg13g2_buf_1 _67_ (.A(S2END[4]),
    .X(N2BEGb[3]));
 sg13g2_buf_1 _68_ (.A(S2END[3]),
    .X(N2BEGb[4]));
 sg13g2_buf_1 _69_ (.A(S2END[2]),
    .X(N2BEGb[5]));
 sg13g2_buf_1 _70_ (.A(S2END[1]),
    .X(N2BEGb[6]));
 sg13g2_buf_1 _71_ (.A(S2END[0]),
    .X(N2BEGb[7]));
 sg13g2_buf_1 _72_ (.A(S4END[15]),
    .X(N4BEG[0]));
 sg13g2_buf_1 _73_ (.A(S4END[14]),
    .X(N4BEG[1]));
 sg13g2_buf_1 _74_ (.A(S4END[13]),
    .X(N4BEG[2]));
 sg13g2_buf_1 _75_ (.A(S4END[12]),
    .X(N4BEG[3]));
 sg13g2_buf_1 _76_ (.A(S4END[11]),
    .X(N4BEG[4]));
 sg13g2_buf_1 _77_ (.A(S4END[10]),
    .X(N4BEG[5]));
 sg13g2_buf_1 _78_ (.A(S4END[9]),
    .X(N4BEG[6]));
 sg13g2_buf_1 _79_ (.A(S4END[8]),
    .X(N4BEG[7]));
 sg13g2_buf_1 _80_ (.A(S4END[7]),
    .X(N4BEG[8]));
 sg13g2_buf_1 _81_ (.A(S4END[6]),
    .X(N4BEG[9]));
 sg13g2_buf_1 _82_ (.A(S4END[5]),
    .X(N4BEG[10]));
 sg13g2_buf_1 _83_ (.A(S4END[4]),
    .X(N4BEG[11]));
 sg13g2_buf_1 _84_ (.A(S4END[3]),
    .X(N4BEG[12]));
 sg13g2_buf_1 _85_ (.A(S4END[2]),
    .X(N4BEG[13]));
 sg13g2_buf_1 _86_ (.A(S4END[1]),
    .X(N4BEG[14]));
 sg13g2_buf_1 _87_ (.A(S4END[0]),
    .X(N4BEG[15]));
 sg13g2_buf_1 _88_ (.A(UserCLK),
    .X(UserCLKo));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_4 FILLER_0_196 ();
 sg13g2_fill_2 FILLER_1_0 ();
 sg13g2_fill_1 FILLER_1_2 ();
 sg13g2_decap_4 FILLER_1_15 ();
 sg13g2_fill_2 FILLER_1_19 ();
 sg13g2_fill_2 FILLER_1_25 ();
 sg13g2_fill_1 FILLER_1_27 ();
 sg13g2_decap_4 FILLER_1_40 ();
 sg13g2_fill_2 FILLER_1_44 ();
 sg13g2_decap_8 FILLER_1_58 ();
 sg13g2_decap_8 FILLER_1_65 ();
 sg13g2_fill_2 FILLER_1_72 ();
 sg13g2_decap_8 FILLER_1_78 ();
 sg13g2_decap_4 FILLER_1_85 ();
 sg13g2_decap_4 FILLER_1_93 ();
 sg13g2_decap_8 FILLER_1_101 ();
 sg13g2_fill_2 FILLER_1_108 ();
 sg13g2_fill_1 FILLER_1_110 ();
 sg13g2_decap_8 FILLER_1_115 ();
 sg13g2_fill_1 FILLER_1_122 ();
 sg13g2_decap_8 FILLER_1_127 ();
 sg13g2_fill_2 FILLER_1_134 ();
 sg13g2_fill_1 FILLER_1_136 ();
 sg13g2_decap_4 FILLER_1_141 ();
 sg13g2_fill_2 FILLER_1_149 ();
 sg13g2_fill_1 FILLER_1_155 ();
 sg13g2_decap_8 FILLER_1_160 ();
 sg13g2_fill_2 FILLER_1_167 ();
 sg13g2_decap_8 FILLER_1_177 ();
 sg13g2_fill_2 FILLER_1_184 ();
 sg13g2_fill_2 FILLER_1_198 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_4 FILLER_2_133 ();
 sg13g2_fill_1 FILLER_2_137 ();
 sg13g2_decap_8 FILLER_2_142 ();
 sg13g2_decap_8 FILLER_2_149 ();
 sg13g2_decap_8 FILLER_2_156 ();
 sg13g2_decap_8 FILLER_2_163 ();
 sg13g2_decap_8 FILLER_2_170 ();
 sg13g2_decap_8 FILLER_2_177 ();
 sg13g2_decap_8 FILLER_2_184 ();
 sg13g2_decap_8 FILLER_2_191 ();
 sg13g2_fill_2 FILLER_2_198 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_fill_2 FILLER_3_7 ();
 sg13g2_fill_1 FILLER_3_9 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_4 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_19 ();
 sg13g2_decap_8 FILLER_4_26 ();
 sg13g2_decap_8 FILLER_4_33 ();
 sg13g2_decap_8 FILLER_4_40 ();
 sg13g2_decap_8 FILLER_4_47 ();
 sg13g2_decap_8 FILLER_4_54 ();
 sg13g2_decap_8 FILLER_4_61 ();
 sg13g2_decap_8 FILLER_4_68 ();
 sg13g2_decap_8 FILLER_4_75 ();
 sg13g2_decap_8 FILLER_4_82 ();
 sg13g2_decap_8 FILLER_4_93 ();
 sg13g2_decap_8 FILLER_4_100 ();
 sg13g2_decap_8 FILLER_4_107 ();
 sg13g2_decap_8 FILLER_4_114 ();
 sg13g2_fill_1 FILLER_4_121 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_4 FILLER_4_182 ();
 sg13g2_decap_4 FILLER_4_194 ();
 sg13g2_fill_2 FILLER_4_198 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_4 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_15 ();
 sg13g2_decap_8 FILLER_5_22 ();
 sg13g2_decap_8 FILLER_5_29 ();
 sg13g2_decap_8 FILLER_5_36 ();
 sg13g2_decap_8 FILLER_5_43 ();
 sg13g2_decap_8 FILLER_5_50 ();
 sg13g2_decap_8 FILLER_5_57 ();
 sg13g2_decap_8 FILLER_5_64 ();
 sg13g2_decap_8 FILLER_5_71 ();
 sg13g2_decap_8 FILLER_5_78 ();
 sg13g2_fill_1 FILLER_5_85 ();
 sg13g2_decap_8 FILLER_5_90 ();
 sg13g2_decap_8 FILLER_5_97 ();
 sg13g2_decap_8 FILLER_5_104 ();
 sg13g2_decap_8 FILLER_5_111 ();
 sg13g2_decap_8 FILLER_5_118 ();
 sg13g2_decap_8 FILLER_5_125 ();
 sg13g2_decap_8 FILLER_5_132 ();
 sg13g2_decap_8 FILLER_5_139 ();
 sg13g2_decap_8 FILLER_5_146 ();
 sg13g2_decap_8 FILLER_5_153 ();
 sg13g2_decap_8 FILLER_5_160 ();
 sg13g2_decap_8 FILLER_5_167 ();
 sg13g2_decap_8 FILLER_5_174 ();
 sg13g2_decap_8 FILLER_5_181 ();
 sg13g2_decap_8 FILLER_5_188 ();
 sg13g2_decap_4 FILLER_5_195 ();
 sg13g2_fill_1 FILLER_5_199 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_fill_2 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_118 ();
 sg13g2_decap_8 FILLER_6_125 ();
 sg13g2_decap_8 FILLER_6_132 ();
 sg13g2_decap_8 FILLER_6_139 ();
 sg13g2_decap_8 FILLER_6_146 ();
 sg13g2_decap_8 FILLER_6_153 ();
 sg13g2_fill_2 FILLER_6_160 ();
 sg13g2_decap_8 FILLER_6_166 ();
 sg13g2_decap_8 FILLER_6_173 ();
 sg13g2_decap_4 FILLER_6_184 ();
 sg13g2_fill_1 FILLER_6_188 ();
 sg13g2_decap_8 FILLER_6_193 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_fill_1 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_12 ();
 sg13g2_decap_8 FILLER_7_19 ();
 sg13g2_decap_8 FILLER_7_26 ();
 sg13g2_decap_8 FILLER_7_33 ();
 sg13g2_decap_8 FILLER_7_40 ();
 sg13g2_decap_8 FILLER_7_47 ();
 sg13g2_decap_8 FILLER_7_54 ();
 sg13g2_decap_8 FILLER_7_61 ();
 sg13g2_decap_8 FILLER_7_68 ();
 sg13g2_decap_8 FILLER_7_75 ();
 sg13g2_decap_8 FILLER_7_82 ();
 sg13g2_decap_8 FILLER_7_89 ();
 sg13g2_decap_8 FILLER_7_96 ();
 sg13g2_decap_8 FILLER_7_103 ();
 sg13g2_decap_8 FILLER_7_110 ();
 sg13g2_decap_8 FILLER_7_117 ();
 sg13g2_decap_8 FILLER_7_124 ();
 sg13g2_decap_8 FILLER_7_131 ();
 sg13g2_decap_8 FILLER_7_138 ();
 sg13g2_decap_8 FILLER_7_145 ();
 sg13g2_decap_4 FILLER_7_152 ();
 sg13g2_fill_1 FILLER_7_156 ();
 sg13g2_decap_8 FILLER_7_161 ();
 sg13g2_decap_4 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_176 ();
 sg13g2_fill_2 FILLER_7_183 ();
 sg13g2_decap_8 FILLER_7_193 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_11 ();
 sg13g2_decap_8 FILLER_8_18 ();
 sg13g2_decap_8 FILLER_8_25 ();
 sg13g2_decap_8 FILLER_8_32 ();
 sg13g2_decap_8 FILLER_8_39 ();
 sg13g2_decap_8 FILLER_8_46 ();
 sg13g2_decap_8 FILLER_8_53 ();
 sg13g2_decap_8 FILLER_8_60 ();
 sg13g2_decap_8 FILLER_8_67 ();
 sg13g2_decap_8 FILLER_8_74 ();
 sg13g2_decap_8 FILLER_8_81 ();
 sg13g2_decap_8 FILLER_8_88 ();
 sg13g2_decap_8 FILLER_8_95 ();
 sg13g2_decap_8 FILLER_8_102 ();
 sg13g2_decap_8 FILLER_8_109 ();
 sg13g2_decap_8 FILLER_8_116 ();
 sg13g2_decap_8 FILLER_8_123 ();
 sg13g2_decap_8 FILLER_8_130 ();
 sg13g2_decap_8 FILLER_8_137 ();
 sg13g2_decap_8 FILLER_8_144 ();
 sg13g2_decap_8 FILLER_8_151 ();
 sg13g2_decap_8 FILLER_8_158 ();
 sg13g2_decap_8 FILLER_8_165 ();
 sg13g2_decap_8 FILLER_8_172 ();
 sg13g2_decap_8 FILLER_8_179 ();
 sg13g2_decap_8 FILLER_8_186 ();
 sg13g2_decap_8 FILLER_8_193 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_11 ();
 sg13g2_fill_1 FILLER_9_13 ();
 sg13g2_decap_4 FILLER_9_18 ();
 sg13g2_decap_4 FILLER_9_26 ();
 sg13g2_decap_8 FILLER_9_34 ();
 sg13g2_decap_8 FILLER_9_41 ();
 sg13g2_decap_8 FILLER_9_48 ();
 sg13g2_decap_4 FILLER_9_55 ();
 sg13g2_fill_2 FILLER_9_59 ();
 sg13g2_fill_2 FILLER_9_65 ();
 sg13g2_decap_8 FILLER_9_79 ();
 sg13g2_fill_1 FILLER_9_86 ();
 sg13g2_decap_8 FILLER_9_95 ();
 sg13g2_decap_4 FILLER_9_102 ();
 sg13g2_decap_8 FILLER_9_110 ();
 sg13g2_fill_2 FILLER_9_117 ();
 sg13g2_fill_1 FILLER_9_119 ();
 sg13g2_fill_1 FILLER_9_124 ();
 sg13g2_fill_1 FILLER_9_129 ();
 sg13g2_decap_8 FILLER_9_134 ();
 sg13g2_decap_8 FILLER_9_141 ();
 sg13g2_decap_8 FILLER_9_148 ();
 sg13g2_fill_1 FILLER_9_155 ();
 sg13g2_decap_4 FILLER_9_160 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_4 FILLER_9_182 ();
 sg13g2_fill_1 FILLER_9_186 ();
 sg13g2_decap_8 FILLER_9_191 ();
 sg13g2_fill_2 FILLER_9_198 ();
 sg13g2_decap_4 FILLER_10_0 ();
 sg13g2_fill_2 FILLER_10_4 ();
 sg13g2_decap_8 FILLER_10_18 ();
 sg13g2_decap_8 FILLER_10_25 ();
 sg13g2_fill_1 FILLER_10_32 ();
 sg13g2_fill_1 FILLER_10_45 ();
 sg13g2_fill_1 FILLER_10_50 ();
 sg13g2_decap_4 FILLER_10_55 ();
 sg13g2_fill_2 FILLER_10_59 ();
 sg13g2_fill_2 FILLER_10_69 ();
 sg13g2_decap_8 FILLER_10_75 ();
 sg13g2_decap_8 FILLER_10_82 ();
 sg13g2_fill_2 FILLER_10_89 ();
 sg13g2_fill_1 FILLER_10_91 ();
 sg13g2_fill_2 FILLER_10_96 ();
 sg13g2_decap_8 FILLER_10_114 ();
 sg13g2_decap_8 FILLER_10_121 ();
 sg13g2_decap_8 FILLER_10_128 ();
 sg13g2_fill_1 FILLER_10_135 ();
 sg13g2_fill_2 FILLER_10_144 ();
 sg13g2_decap_4 FILLER_10_150 ();
 sg13g2_fill_1 FILLER_10_154 ();
 sg13g2_fill_2 FILLER_10_163 ();
 sg13g2_fill_2 FILLER_10_169 ();
 sg13g2_fill_1 FILLER_10_171 ();
 sg13g2_decap_8 FILLER_10_176 ();
 sg13g2_decap_4 FILLER_10_195 ();
 sg13g2_fill_1 FILLER_10_199 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_4 FILLER_11_182 ();
 sg13g2_fill_1 FILLER_11_186 ();
 sg13g2_decap_8 FILLER_11_191 ();
 sg13g2_fill_2 FILLER_11_198 ();
endmodule
