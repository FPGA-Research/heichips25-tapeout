module eFPGA
    #(
        parameter MaxFramesPerCol=20,
        parameter FrameBitsPerRow=32
    )
    (
        input  Tile_X1Y0_A_O_top, //EXTERNAL
        output  Tile_X1Y0_A_I_top, //EXTERNAL
        output  Tile_X1Y0_A_T_top, //EXTERNAL
        input  Tile_X1Y0_B_O_top, //EXTERNAL
        output  Tile_X1Y0_B_I_top, //EXTERNAL
        output  Tile_X1Y0_B_T_top, //EXTERNAL
        input  Tile_X1Y0_C_O_top, //EXTERNAL
        output  Tile_X1Y0_C_I_top, //EXTERNAL
        output  Tile_X1Y0_C_T_top, //EXTERNAL
        input  Tile_X1Y0_D_O_top, //EXTERNAL
        output  Tile_X1Y0_D_I_top, //EXTERNAL
        output  Tile_X1Y0_D_T_top, //EXTERNAL
        input  Tile_X2Y0_A_O_top, //EXTERNAL
        output  Tile_X2Y0_A_I_top, //EXTERNAL
        output  Tile_X2Y0_A_T_top, //EXTERNAL
        input  Tile_X2Y0_B_O_top, //EXTERNAL
        output  Tile_X2Y0_B_I_top, //EXTERNAL
        output  Tile_X2Y0_B_T_top, //EXTERNAL
        input  Tile_X2Y0_C_O_top, //EXTERNAL
        output  Tile_X2Y0_C_I_top, //EXTERNAL
        output  Tile_X2Y0_C_T_top, //EXTERNAL
        input  Tile_X2Y0_D_O_top, //EXTERNAL
        output  Tile_X2Y0_D_I_top, //EXTERNAL
        output  Tile_X2Y0_D_T_top, //EXTERNAL
        input  Tile_X3Y0_A_O_top, //EXTERNAL
        output  Tile_X3Y0_A_I_top, //EXTERNAL
        output  Tile_X3Y0_A_T_top, //EXTERNAL
        input  Tile_X3Y0_B_O_top, //EXTERNAL
        output  Tile_X3Y0_B_I_top, //EXTERNAL
        output  Tile_X3Y0_B_T_top, //EXTERNAL
        input  Tile_X3Y0_C_O_top, //EXTERNAL
        output  Tile_X3Y0_C_I_top, //EXTERNAL
        output  Tile_X3Y0_C_T_top, //EXTERNAL
        input  Tile_X3Y0_D_O_top, //EXTERNAL
        output  Tile_X3Y0_D_I_top, //EXTERNAL
        output  Tile_X3Y0_D_T_top, //EXTERNAL
        input  Tile_X4Y0_A_O_top, //EXTERNAL
        output  Tile_X4Y0_A_I_top, //EXTERNAL
        output  Tile_X4Y0_A_T_top, //EXTERNAL
        input  Tile_X4Y0_B_O_top, //EXTERNAL
        output  Tile_X4Y0_B_I_top, //EXTERNAL
        output  Tile_X4Y0_B_T_top, //EXTERNAL
        input  Tile_X4Y0_C_O_top, //EXTERNAL
        output  Tile_X4Y0_C_I_top, //EXTERNAL
        output  Tile_X4Y0_C_T_top, //EXTERNAL
        input  Tile_X4Y0_D_O_top, //EXTERNAL
        output  Tile_X4Y0_D_I_top, //EXTERNAL
        output  Tile_X4Y0_D_T_top, //EXTERNAL
        input  Tile_X0Y2_UO_OUT_TT_PROJECT0, //EXTERNAL
        input  Tile_X0Y2_UO_OUT_TT_PROJECT1, //EXTERNAL
        input  Tile_X0Y2_UO_OUT_TT_PROJECT2, //EXTERNAL
        input  Tile_X0Y2_UO_OUT_TT_PROJECT3, //EXTERNAL
        input  Tile_X0Y2_UO_OUT_TT_PROJECT4, //EXTERNAL
        input  Tile_X0Y2_UO_OUT_TT_PROJECT5, //EXTERNAL
        input  Tile_X0Y2_UO_OUT_TT_PROJECT6, //EXTERNAL
        input  Tile_X0Y2_UO_OUT_TT_PROJECT7, //EXTERNAL
        input  Tile_X0Y2_UIO_OUT_TT_PROJECT0, //EXTERNAL
        input  Tile_X0Y2_UIO_OUT_TT_PROJECT1, //EXTERNAL
        input  Tile_X0Y2_UIO_OUT_TT_PROJECT2, //EXTERNAL
        input  Tile_X0Y2_UIO_OUT_TT_PROJECT3, //EXTERNAL
        input  Tile_X0Y2_UIO_OUT_TT_PROJECT4, //EXTERNAL
        input  Tile_X0Y2_UIO_OUT_TT_PROJECT5, //EXTERNAL
        input  Tile_X0Y2_UIO_OUT_TT_PROJECT6, //EXTERNAL
        input  Tile_X0Y2_UIO_OUT_TT_PROJECT7, //EXTERNAL
        input  Tile_X0Y2_UIO_OE_TT_PROJECT0, //EXTERNAL
        input  Tile_X0Y2_UIO_OE_TT_PROJECT1, //EXTERNAL
        input  Tile_X0Y2_UIO_OE_TT_PROJECT2, //EXTERNAL
        input  Tile_X0Y2_UIO_OE_TT_PROJECT3, //EXTERNAL
        input  Tile_X0Y2_UIO_OE_TT_PROJECT4, //EXTERNAL
        input  Tile_X0Y2_UIO_OE_TT_PROJECT5, //EXTERNAL
        input  Tile_X0Y2_UIO_OE_TT_PROJECT6, //EXTERNAL
        input  Tile_X0Y2_UIO_OE_TT_PROJECT7, //EXTERNAL
        output  Tile_X0Y2_UI_IN_TT_PROJECT0, //EXTERNAL
        output  Tile_X0Y2_UI_IN_TT_PROJECT1, //EXTERNAL
        output  Tile_X0Y2_UI_IN_TT_PROJECT2, //EXTERNAL
        output  Tile_X0Y2_UI_IN_TT_PROJECT3, //EXTERNAL
        output  Tile_X0Y2_UI_IN_TT_PROJECT4, //EXTERNAL
        output  Tile_X0Y2_UI_IN_TT_PROJECT5, //EXTERNAL
        output  Tile_X0Y2_UI_IN_TT_PROJECT6, //EXTERNAL
        output  Tile_X0Y2_UI_IN_TT_PROJECT7, //EXTERNAL
        output  Tile_X0Y2_UIO_IN_TT_PROJECT0, //EXTERNAL
        output  Tile_X0Y2_UIO_IN_TT_PROJECT1, //EXTERNAL
        output  Tile_X0Y2_UIO_IN_TT_PROJECT2, //EXTERNAL
        output  Tile_X0Y2_UIO_IN_TT_PROJECT3, //EXTERNAL
        output  Tile_X0Y2_UIO_IN_TT_PROJECT4, //EXTERNAL
        output  Tile_X0Y2_UIO_IN_TT_PROJECT5, //EXTERNAL
        output  Tile_X0Y2_UIO_IN_TT_PROJECT6, //EXTERNAL
        output  Tile_X0Y2_UIO_IN_TT_PROJECT7, //EXTERNAL
        output  Tile_X0Y2_ENA_TT_PROJECT, //EXTERNAL
        output  Tile_X0Y2_CLK_TT_PROJECT, //EXTERNAL
        output  Tile_X0Y2_RST_N_TT_PROJECT, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM0, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM1, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM2, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM3, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM4, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM5, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM6, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM7, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM8, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM9, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM10, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM11, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM12, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM13, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM14, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM15, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM16, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM17, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM18, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM19, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM20, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM21, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM22, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM23, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM24, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM25, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM26, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM27, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM28, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM29, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM30, //EXTERNAL
        input  Tile_X5Y2_DOUT_SRAM31, //EXTERNAL
        input  Tile_X5Y2_CONFIGURED_top, //EXTERNAL
        output  Tile_X5Y2_ADDR_SRAM0, //EXTERNAL
        output  Tile_X5Y2_ADDR_SRAM1, //EXTERNAL
        output  Tile_X5Y2_ADDR_SRAM2, //EXTERNAL
        output  Tile_X5Y2_ADDR_SRAM3, //EXTERNAL
        output  Tile_X5Y2_ADDR_SRAM4, //EXTERNAL
        output  Tile_X5Y2_ADDR_SRAM5, //EXTERNAL
        output  Tile_X5Y2_ADDR_SRAM6, //EXTERNAL
        output  Tile_X5Y2_ADDR_SRAM7, //EXTERNAL
        output  Tile_X5Y2_ADDR_SRAM8, //EXTERNAL
        output  Tile_X5Y2_ADDR_SRAM9, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM0, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM1, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM2, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM3, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM4, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM5, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM6, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM7, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM8, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM9, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM10, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM11, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM12, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM13, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM14, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM15, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM16, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM17, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM18, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM19, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM20, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM21, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM22, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM23, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM24, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM25, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM26, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM27, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM28, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM29, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM30, //EXTERNAL
        output  Tile_X5Y2_DIN_SRAM31, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM0, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM1, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM2, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM3, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM4, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM5, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM6, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM7, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM8, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM9, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM10, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM11, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM12, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM13, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM14, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM15, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM16, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM17, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM18, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM19, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM20, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM21, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM22, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM23, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM24, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM25, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM26, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM27, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM28, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM29, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM30, //EXTERNAL
        output  Tile_X5Y2_BM_SRAM31, //EXTERNAL
        output  Tile_X5Y2_WEN_SRAM, //EXTERNAL
        output  Tile_X5Y2_MEN_SRAM, //EXTERNAL
        output  Tile_X5Y2_REN_SRAM, //EXTERNAL
        output  Tile_X5Y2_CLK_SRAM, //EXTERNAL
        output  Tile_X5Y2_TIE_HIGH_SRAM, //EXTERNAL
        output  Tile_X5Y2_TIE_LOW_SRAM, //EXTERNAL
        input  Tile_X0Y3_UO_OUT_TT_PROJECT0, //EXTERNAL
        input  Tile_X0Y3_UO_OUT_TT_PROJECT1, //EXTERNAL
        input  Tile_X0Y3_UO_OUT_TT_PROJECT2, //EXTERNAL
        input  Tile_X0Y3_UO_OUT_TT_PROJECT3, //EXTERNAL
        input  Tile_X0Y3_UO_OUT_TT_PROJECT4, //EXTERNAL
        input  Tile_X0Y3_UO_OUT_TT_PROJECT5, //EXTERNAL
        input  Tile_X0Y3_UO_OUT_TT_PROJECT6, //EXTERNAL
        input  Tile_X0Y3_UO_OUT_TT_PROJECT7, //EXTERNAL
        input  Tile_X0Y3_UIO_OUT_TT_PROJECT0, //EXTERNAL
        input  Tile_X0Y3_UIO_OUT_TT_PROJECT1, //EXTERNAL
        input  Tile_X0Y3_UIO_OUT_TT_PROJECT2, //EXTERNAL
        input  Tile_X0Y3_UIO_OUT_TT_PROJECT3, //EXTERNAL
        input  Tile_X0Y3_UIO_OUT_TT_PROJECT4, //EXTERNAL
        input  Tile_X0Y3_UIO_OUT_TT_PROJECT5, //EXTERNAL
        input  Tile_X0Y3_UIO_OUT_TT_PROJECT6, //EXTERNAL
        input  Tile_X0Y3_UIO_OUT_TT_PROJECT7, //EXTERNAL
        input  Tile_X0Y3_UIO_OE_TT_PROJECT0, //EXTERNAL
        input  Tile_X0Y3_UIO_OE_TT_PROJECT1, //EXTERNAL
        input  Tile_X0Y3_UIO_OE_TT_PROJECT2, //EXTERNAL
        input  Tile_X0Y3_UIO_OE_TT_PROJECT3, //EXTERNAL
        input  Tile_X0Y3_UIO_OE_TT_PROJECT4, //EXTERNAL
        input  Tile_X0Y3_UIO_OE_TT_PROJECT5, //EXTERNAL
        input  Tile_X0Y3_UIO_OE_TT_PROJECT6, //EXTERNAL
        input  Tile_X0Y3_UIO_OE_TT_PROJECT7, //EXTERNAL
        output  Tile_X0Y3_UI_IN_TT_PROJECT0, //EXTERNAL
        output  Tile_X0Y3_UI_IN_TT_PROJECT1, //EXTERNAL
        output  Tile_X0Y3_UI_IN_TT_PROJECT2, //EXTERNAL
        output  Tile_X0Y3_UI_IN_TT_PROJECT3, //EXTERNAL
        output  Tile_X0Y3_UI_IN_TT_PROJECT4, //EXTERNAL
        output  Tile_X0Y3_UI_IN_TT_PROJECT5, //EXTERNAL
        output  Tile_X0Y3_UI_IN_TT_PROJECT6, //EXTERNAL
        output  Tile_X0Y3_UI_IN_TT_PROJECT7, //EXTERNAL
        output  Tile_X0Y3_UIO_IN_TT_PROJECT0, //EXTERNAL
        output  Tile_X0Y3_UIO_IN_TT_PROJECT1, //EXTERNAL
        output  Tile_X0Y3_UIO_IN_TT_PROJECT2, //EXTERNAL
        output  Tile_X0Y3_UIO_IN_TT_PROJECT3, //EXTERNAL
        output  Tile_X0Y3_UIO_IN_TT_PROJECT4, //EXTERNAL
        output  Tile_X0Y3_UIO_IN_TT_PROJECT5, //EXTERNAL
        output  Tile_X0Y3_UIO_IN_TT_PROJECT6, //EXTERNAL
        output  Tile_X0Y3_UIO_IN_TT_PROJECT7, //EXTERNAL
        output  Tile_X0Y3_ENA_TT_PROJECT, //EXTERNAL
        output  Tile_X0Y3_CLK_TT_PROJECT, //EXTERNAL
        output  Tile_X0Y3_RST_N_TT_PROJECT, //EXTERNAL
        input  Tile_X0Y4_UO_OUT_TT_PROJECT0, //EXTERNAL
        input  Tile_X0Y4_UO_OUT_TT_PROJECT1, //EXTERNAL
        input  Tile_X0Y4_UO_OUT_TT_PROJECT2, //EXTERNAL
        input  Tile_X0Y4_UO_OUT_TT_PROJECT3, //EXTERNAL
        input  Tile_X0Y4_UO_OUT_TT_PROJECT4, //EXTERNAL
        input  Tile_X0Y4_UO_OUT_TT_PROJECT5, //EXTERNAL
        input  Tile_X0Y4_UO_OUT_TT_PROJECT6, //EXTERNAL
        input  Tile_X0Y4_UO_OUT_TT_PROJECT7, //EXTERNAL
        input  Tile_X0Y4_UIO_OUT_TT_PROJECT0, //EXTERNAL
        input  Tile_X0Y4_UIO_OUT_TT_PROJECT1, //EXTERNAL
        input  Tile_X0Y4_UIO_OUT_TT_PROJECT2, //EXTERNAL
        input  Tile_X0Y4_UIO_OUT_TT_PROJECT3, //EXTERNAL
        input  Tile_X0Y4_UIO_OUT_TT_PROJECT4, //EXTERNAL
        input  Tile_X0Y4_UIO_OUT_TT_PROJECT5, //EXTERNAL
        input  Tile_X0Y4_UIO_OUT_TT_PROJECT6, //EXTERNAL
        input  Tile_X0Y4_UIO_OUT_TT_PROJECT7, //EXTERNAL
        input  Tile_X0Y4_UIO_OE_TT_PROJECT0, //EXTERNAL
        input  Tile_X0Y4_UIO_OE_TT_PROJECT1, //EXTERNAL
        input  Tile_X0Y4_UIO_OE_TT_PROJECT2, //EXTERNAL
        input  Tile_X0Y4_UIO_OE_TT_PROJECT3, //EXTERNAL
        input  Tile_X0Y4_UIO_OE_TT_PROJECT4, //EXTERNAL
        input  Tile_X0Y4_UIO_OE_TT_PROJECT5, //EXTERNAL
        input  Tile_X0Y4_UIO_OE_TT_PROJECT6, //EXTERNAL
        input  Tile_X0Y4_UIO_OE_TT_PROJECT7, //EXTERNAL
        output  Tile_X0Y4_UI_IN_TT_PROJECT0, //EXTERNAL
        output  Tile_X0Y4_UI_IN_TT_PROJECT1, //EXTERNAL
        output  Tile_X0Y4_UI_IN_TT_PROJECT2, //EXTERNAL
        output  Tile_X0Y4_UI_IN_TT_PROJECT3, //EXTERNAL
        output  Tile_X0Y4_UI_IN_TT_PROJECT4, //EXTERNAL
        output  Tile_X0Y4_UI_IN_TT_PROJECT5, //EXTERNAL
        output  Tile_X0Y4_UI_IN_TT_PROJECT6, //EXTERNAL
        output  Tile_X0Y4_UI_IN_TT_PROJECT7, //EXTERNAL
        output  Tile_X0Y4_UIO_IN_TT_PROJECT0, //EXTERNAL
        output  Tile_X0Y4_UIO_IN_TT_PROJECT1, //EXTERNAL
        output  Tile_X0Y4_UIO_IN_TT_PROJECT2, //EXTERNAL
        output  Tile_X0Y4_UIO_IN_TT_PROJECT3, //EXTERNAL
        output  Tile_X0Y4_UIO_IN_TT_PROJECT4, //EXTERNAL
        output  Tile_X0Y4_UIO_IN_TT_PROJECT5, //EXTERNAL
        output  Tile_X0Y4_UIO_IN_TT_PROJECT6, //EXTERNAL
        output  Tile_X0Y4_UIO_IN_TT_PROJECT7, //EXTERNAL
        output  Tile_X0Y4_ENA_TT_PROJECT, //EXTERNAL
        output  Tile_X0Y4_CLK_TT_PROJECT, //EXTERNAL
        output  Tile_X0Y4_RST_N_TT_PROJECT, //EXTERNAL
        input  Tile_X5Y4_UO_OUT_TT_PROJECT0, //EXTERNAL
        input  Tile_X5Y4_UO_OUT_TT_PROJECT1, //EXTERNAL
        input  Tile_X5Y4_UO_OUT_TT_PROJECT2, //EXTERNAL
        input  Tile_X5Y4_UO_OUT_TT_PROJECT3, //EXTERNAL
        input  Tile_X5Y4_UO_OUT_TT_PROJECT4, //EXTERNAL
        input  Tile_X5Y4_UO_OUT_TT_PROJECT5, //EXTERNAL
        input  Tile_X5Y4_UO_OUT_TT_PROJECT6, //EXTERNAL
        input  Tile_X5Y4_UO_OUT_TT_PROJECT7, //EXTERNAL
        input  Tile_X5Y4_UIO_OUT_TT_PROJECT0, //EXTERNAL
        input  Tile_X5Y4_UIO_OUT_TT_PROJECT1, //EXTERNAL
        input  Tile_X5Y4_UIO_OUT_TT_PROJECT2, //EXTERNAL
        input  Tile_X5Y4_UIO_OUT_TT_PROJECT3, //EXTERNAL
        input  Tile_X5Y4_UIO_OUT_TT_PROJECT4, //EXTERNAL
        input  Tile_X5Y4_UIO_OUT_TT_PROJECT5, //EXTERNAL
        input  Tile_X5Y4_UIO_OUT_TT_PROJECT6, //EXTERNAL
        input  Tile_X5Y4_UIO_OUT_TT_PROJECT7, //EXTERNAL
        input  Tile_X5Y4_UIO_OE_TT_PROJECT0, //EXTERNAL
        input  Tile_X5Y4_UIO_OE_TT_PROJECT1, //EXTERNAL
        input  Tile_X5Y4_UIO_OE_TT_PROJECT2, //EXTERNAL
        input  Tile_X5Y4_UIO_OE_TT_PROJECT3, //EXTERNAL
        input  Tile_X5Y4_UIO_OE_TT_PROJECT4, //EXTERNAL
        input  Tile_X5Y4_UIO_OE_TT_PROJECT5, //EXTERNAL
        input  Tile_X5Y4_UIO_OE_TT_PROJECT6, //EXTERNAL
        input  Tile_X5Y4_UIO_OE_TT_PROJECT7, //EXTERNAL
        output  Tile_X5Y4_UI_IN_TT_PROJECT0, //EXTERNAL
        output  Tile_X5Y4_UI_IN_TT_PROJECT1, //EXTERNAL
        output  Tile_X5Y4_UI_IN_TT_PROJECT2, //EXTERNAL
        output  Tile_X5Y4_UI_IN_TT_PROJECT3, //EXTERNAL
        output  Tile_X5Y4_UI_IN_TT_PROJECT4, //EXTERNAL
        output  Tile_X5Y4_UI_IN_TT_PROJECT5, //EXTERNAL
        output  Tile_X5Y4_UI_IN_TT_PROJECT6, //EXTERNAL
        output  Tile_X5Y4_UI_IN_TT_PROJECT7, //EXTERNAL
        output  Tile_X5Y4_UIO_IN_TT_PROJECT0, //EXTERNAL
        output  Tile_X5Y4_UIO_IN_TT_PROJECT1, //EXTERNAL
        output  Tile_X5Y4_UIO_IN_TT_PROJECT2, //EXTERNAL
        output  Tile_X5Y4_UIO_IN_TT_PROJECT3, //EXTERNAL
        output  Tile_X5Y4_UIO_IN_TT_PROJECT4, //EXTERNAL
        output  Tile_X5Y4_UIO_IN_TT_PROJECT5, //EXTERNAL
        output  Tile_X5Y4_UIO_IN_TT_PROJECT6, //EXTERNAL
        output  Tile_X5Y4_UIO_IN_TT_PROJECT7, //EXTERNAL
        output  Tile_X5Y4_ENA_TT_PROJECT, //EXTERNAL
        output  Tile_X5Y4_CLK_TT_PROJECT, //EXTERNAL
        output  Tile_X5Y4_RST_N_TT_PROJECT, //EXTERNAL
        input  Tile_X0Y5_UO_OUT_TT_PROJECT0, //EXTERNAL
        input  Tile_X0Y5_UO_OUT_TT_PROJECT1, //EXTERNAL
        input  Tile_X0Y5_UO_OUT_TT_PROJECT2, //EXTERNAL
        input  Tile_X0Y5_UO_OUT_TT_PROJECT3, //EXTERNAL
        input  Tile_X0Y5_UO_OUT_TT_PROJECT4, //EXTERNAL
        input  Tile_X0Y5_UO_OUT_TT_PROJECT5, //EXTERNAL
        input  Tile_X0Y5_UO_OUT_TT_PROJECT6, //EXTERNAL
        input  Tile_X0Y5_UO_OUT_TT_PROJECT7, //EXTERNAL
        input  Tile_X0Y5_UIO_OUT_TT_PROJECT0, //EXTERNAL
        input  Tile_X0Y5_UIO_OUT_TT_PROJECT1, //EXTERNAL
        input  Tile_X0Y5_UIO_OUT_TT_PROJECT2, //EXTERNAL
        input  Tile_X0Y5_UIO_OUT_TT_PROJECT3, //EXTERNAL
        input  Tile_X0Y5_UIO_OUT_TT_PROJECT4, //EXTERNAL
        input  Tile_X0Y5_UIO_OUT_TT_PROJECT5, //EXTERNAL
        input  Tile_X0Y5_UIO_OUT_TT_PROJECT6, //EXTERNAL
        input  Tile_X0Y5_UIO_OUT_TT_PROJECT7, //EXTERNAL
        input  Tile_X0Y5_UIO_OE_TT_PROJECT0, //EXTERNAL
        input  Tile_X0Y5_UIO_OE_TT_PROJECT1, //EXTERNAL
        input  Tile_X0Y5_UIO_OE_TT_PROJECT2, //EXTERNAL
        input  Tile_X0Y5_UIO_OE_TT_PROJECT3, //EXTERNAL
        input  Tile_X0Y5_UIO_OE_TT_PROJECT4, //EXTERNAL
        input  Tile_X0Y5_UIO_OE_TT_PROJECT5, //EXTERNAL
        input  Tile_X0Y5_UIO_OE_TT_PROJECT6, //EXTERNAL
        input  Tile_X0Y5_UIO_OE_TT_PROJECT7, //EXTERNAL
        output  Tile_X0Y5_UI_IN_TT_PROJECT0, //EXTERNAL
        output  Tile_X0Y5_UI_IN_TT_PROJECT1, //EXTERNAL
        output  Tile_X0Y5_UI_IN_TT_PROJECT2, //EXTERNAL
        output  Tile_X0Y5_UI_IN_TT_PROJECT3, //EXTERNAL
        output  Tile_X0Y5_UI_IN_TT_PROJECT4, //EXTERNAL
        output  Tile_X0Y5_UI_IN_TT_PROJECT5, //EXTERNAL
        output  Tile_X0Y5_UI_IN_TT_PROJECT6, //EXTERNAL
        output  Tile_X0Y5_UI_IN_TT_PROJECT7, //EXTERNAL
        output  Tile_X0Y5_UIO_IN_TT_PROJECT0, //EXTERNAL
        output  Tile_X0Y5_UIO_IN_TT_PROJECT1, //EXTERNAL
        output  Tile_X0Y5_UIO_IN_TT_PROJECT2, //EXTERNAL
        output  Tile_X0Y5_UIO_IN_TT_PROJECT3, //EXTERNAL
        output  Tile_X0Y5_UIO_IN_TT_PROJECT4, //EXTERNAL
        output  Tile_X0Y5_UIO_IN_TT_PROJECT5, //EXTERNAL
        output  Tile_X0Y5_UIO_IN_TT_PROJECT6, //EXTERNAL
        output  Tile_X0Y5_UIO_IN_TT_PROJECT7, //EXTERNAL
        output  Tile_X0Y5_ENA_TT_PROJECT, //EXTERNAL
        output  Tile_X0Y5_CLK_TT_PROJECT, //EXTERNAL
        output  Tile_X0Y5_RST_N_TT_PROJECT, //EXTERNAL
        input  Tile_X5Y5_UO_OUT_TT_PROJECT0, //EXTERNAL
        input  Tile_X5Y5_UO_OUT_TT_PROJECT1, //EXTERNAL
        input  Tile_X5Y5_UO_OUT_TT_PROJECT2, //EXTERNAL
        input  Tile_X5Y5_UO_OUT_TT_PROJECT3, //EXTERNAL
        input  Tile_X5Y5_UO_OUT_TT_PROJECT4, //EXTERNAL
        input  Tile_X5Y5_UO_OUT_TT_PROJECT5, //EXTERNAL
        input  Tile_X5Y5_UO_OUT_TT_PROJECT6, //EXTERNAL
        input  Tile_X5Y5_UO_OUT_TT_PROJECT7, //EXTERNAL
        input  Tile_X5Y5_UIO_OUT_TT_PROJECT0, //EXTERNAL
        input  Tile_X5Y5_UIO_OUT_TT_PROJECT1, //EXTERNAL
        input  Tile_X5Y5_UIO_OUT_TT_PROJECT2, //EXTERNAL
        input  Tile_X5Y5_UIO_OUT_TT_PROJECT3, //EXTERNAL
        input  Tile_X5Y5_UIO_OUT_TT_PROJECT4, //EXTERNAL
        input  Tile_X5Y5_UIO_OUT_TT_PROJECT5, //EXTERNAL
        input  Tile_X5Y5_UIO_OUT_TT_PROJECT6, //EXTERNAL
        input  Tile_X5Y5_UIO_OUT_TT_PROJECT7, //EXTERNAL
        input  Tile_X5Y5_UIO_OE_TT_PROJECT0, //EXTERNAL
        input  Tile_X5Y5_UIO_OE_TT_PROJECT1, //EXTERNAL
        input  Tile_X5Y5_UIO_OE_TT_PROJECT2, //EXTERNAL
        input  Tile_X5Y5_UIO_OE_TT_PROJECT3, //EXTERNAL
        input  Tile_X5Y5_UIO_OE_TT_PROJECT4, //EXTERNAL
        input  Tile_X5Y5_UIO_OE_TT_PROJECT5, //EXTERNAL
        input  Tile_X5Y5_UIO_OE_TT_PROJECT6, //EXTERNAL
        input  Tile_X5Y5_UIO_OE_TT_PROJECT7, //EXTERNAL
        output  Tile_X5Y5_UI_IN_TT_PROJECT0, //EXTERNAL
        output  Tile_X5Y5_UI_IN_TT_PROJECT1, //EXTERNAL
        output  Tile_X5Y5_UI_IN_TT_PROJECT2, //EXTERNAL
        output  Tile_X5Y5_UI_IN_TT_PROJECT3, //EXTERNAL
        output  Tile_X5Y5_UI_IN_TT_PROJECT4, //EXTERNAL
        output  Tile_X5Y5_UI_IN_TT_PROJECT5, //EXTERNAL
        output  Tile_X5Y5_UI_IN_TT_PROJECT6, //EXTERNAL
        output  Tile_X5Y5_UI_IN_TT_PROJECT7, //EXTERNAL
        output  Tile_X5Y5_UIO_IN_TT_PROJECT0, //EXTERNAL
        output  Tile_X5Y5_UIO_IN_TT_PROJECT1, //EXTERNAL
        output  Tile_X5Y5_UIO_IN_TT_PROJECT2, //EXTERNAL
        output  Tile_X5Y5_UIO_IN_TT_PROJECT3, //EXTERNAL
        output  Tile_X5Y5_UIO_IN_TT_PROJECT4, //EXTERNAL
        output  Tile_X5Y5_UIO_IN_TT_PROJECT5, //EXTERNAL
        output  Tile_X5Y5_UIO_IN_TT_PROJECT6, //EXTERNAL
        output  Tile_X5Y5_UIO_IN_TT_PROJECT7, //EXTERNAL
        output  Tile_X5Y5_ENA_TT_PROJECT, //EXTERNAL
        output  Tile_X5Y5_CLK_TT_PROJECT, //EXTERNAL
        output  Tile_X5Y5_RST_N_TT_PROJECT, //EXTERNAL
        input  Tile_X0Y6_UO_OUT_TT_PROJECT0, //EXTERNAL
        input  Tile_X0Y6_UO_OUT_TT_PROJECT1, //EXTERNAL
        input  Tile_X0Y6_UO_OUT_TT_PROJECT2, //EXTERNAL
        input  Tile_X0Y6_UO_OUT_TT_PROJECT3, //EXTERNAL
        input  Tile_X0Y6_UO_OUT_TT_PROJECT4, //EXTERNAL
        input  Tile_X0Y6_UO_OUT_TT_PROJECT5, //EXTERNAL
        input  Tile_X0Y6_UO_OUT_TT_PROJECT6, //EXTERNAL
        input  Tile_X0Y6_UO_OUT_TT_PROJECT7, //EXTERNAL
        input  Tile_X0Y6_UIO_OUT_TT_PROJECT0, //EXTERNAL
        input  Tile_X0Y6_UIO_OUT_TT_PROJECT1, //EXTERNAL
        input  Tile_X0Y6_UIO_OUT_TT_PROJECT2, //EXTERNAL
        input  Tile_X0Y6_UIO_OUT_TT_PROJECT3, //EXTERNAL
        input  Tile_X0Y6_UIO_OUT_TT_PROJECT4, //EXTERNAL
        input  Tile_X0Y6_UIO_OUT_TT_PROJECT5, //EXTERNAL
        input  Tile_X0Y6_UIO_OUT_TT_PROJECT6, //EXTERNAL
        input  Tile_X0Y6_UIO_OUT_TT_PROJECT7, //EXTERNAL
        input  Tile_X0Y6_UIO_OE_TT_PROJECT0, //EXTERNAL
        input  Tile_X0Y6_UIO_OE_TT_PROJECT1, //EXTERNAL
        input  Tile_X0Y6_UIO_OE_TT_PROJECT2, //EXTERNAL
        input  Tile_X0Y6_UIO_OE_TT_PROJECT3, //EXTERNAL
        input  Tile_X0Y6_UIO_OE_TT_PROJECT4, //EXTERNAL
        input  Tile_X0Y6_UIO_OE_TT_PROJECT5, //EXTERNAL
        input  Tile_X0Y6_UIO_OE_TT_PROJECT6, //EXTERNAL
        input  Tile_X0Y6_UIO_OE_TT_PROJECT7, //EXTERNAL
        output  Tile_X0Y6_UI_IN_TT_PROJECT0, //EXTERNAL
        output  Tile_X0Y6_UI_IN_TT_PROJECT1, //EXTERNAL
        output  Tile_X0Y6_UI_IN_TT_PROJECT2, //EXTERNAL
        output  Tile_X0Y6_UI_IN_TT_PROJECT3, //EXTERNAL
        output  Tile_X0Y6_UI_IN_TT_PROJECT4, //EXTERNAL
        output  Tile_X0Y6_UI_IN_TT_PROJECT5, //EXTERNAL
        output  Tile_X0Y6_UI_IN_TT_PROJECT6, //EXTERNAL
        output  Tile_X0Y6_UI_IN_TT_PROJECT7, //EXTERNAL
        output  Tile_X0Y6_UIO_IN_TT_PROJECT0, //EXTERNAL
        output  Tile_X0Y6_UIO_IN_TT_PROJECT1, //EXTERNAL
        output  Tile_X0Y6_UIO_IN_TT_PROJECT2, //EXTERNAL
        output  Tile_X0Y6_UIO_IN_TT_PROJECT3, //EXTERNAL
        output  Tile_X0Y6_UIO_IN_TT_PROJECT4, //EXTERNAL
        output  Tile_X0Y6_UIO_IN_TT_PROJECT5, //EXTERNAL
        output  Tile_X0Y6_UIO_IN_TT_PROJECT6, //EXTERNAL
        output  Tile_X0Y6_UIO_IN_TT_PROJECT7, //EXTERNAL
        output  Tile_X0Y6_ENA_TT_PROJECT, //EXTERNAL
        output  Tile_X0Y6_CLK_TT_PROJECT, //EXTERNAL
        output  Tile_X0Y6_RST_N_TT_PROJECT, //EXTERNAL
        input  Tile_X5Y6_UO_OUT_TT_PROJECT0, //EXTERNAL
        input  Tile_X5Y6_UO_OUT_TT_PROJECT1, //EXTERNAL
        input  Tile_X5Y6_UO_OUT_TT_PROJECT2, //EXTERNAL
        input  Tile_X5Y6_UO_OUT_TT_PROJECT3, //EXTERNAL
        input  Tile_X5Y6_UO_OUT_TT_PROJECT4, //EXTERNAL
        input  Tile_X5Y6_UO_OUT_TT_PROJECT5, //EXTERNAL
        input  Tile_X5Y6_UO_OUT_TT_PROJECT6, //EXTERNAL
        input  Tile_X5Y6_UO_OUT_TT_PROJECT7, //EXTERNAL
        input  Tile_X5Y6_UIO_OUT_TT_PROJECT0, //EXTERNAL
        input  Tile_X5Y6_UIO_OUT_TT_PROJECT1, //EXTERNAL
        input  Tile_X5Y6_UIO_OUT_TT_PROJECT2, //EXTERNAL
        input  Tile_X5Y6_UIO_OUT_TT_PROJECT3, //EXTERNAL
        input  Tile_X5Y6_UIO_OUT_TT_PROJECT4, //EXTERNAL
        input  Tile_X5Y6_UIO_OUT_TT_PROJECT5, //EXTERNAL
        input  Tile_X5Y6_UIO_OUT_TT_PROJECT6, //EXTERNAL
        input  Tile_X5Y6_UIO_OUT_TT_PROJECT7, //EXTERNAL
        input  Tile_X5Y6_UIO_OE_TT_PROJECT0, //EXTERNAL
        input  Tile_X5Y6_UIO_OE_TT_PROJECT1, //EXTERNAL
        input  Tile_X5Y6_UIO_OE_TT_PROJECT2, //EXTERNAL
        input  Tile_X5Y6_UIO_OE_TT_PROJECT3, //EXTERNAL
        input  Tile_X5Y6_UIO_OE_TT_PROJECT4, //EXTERNAL
        input  Tile_X5Y6_UIO_OE_TT_PROJECT5, //EXTERNAL
        input  Tile_X5Y6_UIO_OE_TT_PROJECT6, //EXTERNAL
        input  Tile_X5Y6_UIO_OE_TT_PROJECT7, //EXTERNAL
        output  Tile_X5Y6_UI_IN_TT_PROJECT0, //EXTERNAL
        output  Tile_X5Y6_UI_IN_TT_PROJECT1, //EXTERNAL
        output  Tile_X5Y6_UI_IN_TT_PROJECT2, //EXTERNAL
        output  Tile_X5Y6_UI_IN_TT_PROJECT3, //EXTERNAL
        output  Tile_X5Y6_UI_IN_TT_PROJECT4, //EXTERNAL
        output  Tile_X5Y6_UI_IN_TT_PROJECT5, //EXTERNAL
        output  Tile_X5Y6_UI_IN_TT_PROJECT6, //EXTERNAL
        output  Tile_X5Y6_UI_IN_TT_PROJECT7, //EXTERNAL
        output  Tile_X5Y6_UIO_IN_TT_PROJECT0, //EXTERNAL
        output  Tile_X5Y6_UIO_IN_TT_PROJECT1, //EXTERNAL
        output  Tile_X5Y6_UIO_IN_TT_PROJECT2, //EXTERNAL
        output  Tile_X5Y6_UIO_IN_TT_PROJECT3, //EXTERNAL
        output  Tile_X5Y6_UIO_IN_TT_PROJECT4, //EXTERNAL
        output  Tile_X5Y6_UIO_IN_TT_PROJECT5, //EXTERNAL
        output  Tile_X5Y6_UIO_IN_TT_PROJECT6, //EXTERNAL
        output  Tile_X5Y6_UIO_IN_TT_PROJECT7, //EXTERNAL
        output  Tile_X5Y6_ENA_TT_PROJECT, //EXTERNAL
        output  Tile_X5Y6_CLK_TT_PROJECT, //EXTERNAL
        output  Tile_X5Y6_RST_N_TT_PROJECT, //EXTERNAL
        input  Tile_X0Y7_UO_OUT_TT_PROJECT0, //EXTERNAL
        input  Tile_X0Y7_UO_OUT_TT_PROJECT1, //EXTERNAL
        input  Tile_X0Y7_UO_OUT_TT_PROJECT2, //EXTERNAL
        input  Tile_X0Y7_UO_OUT_TT_PROJECT3, //EXTERNAL
        input  Tile_X0Y7_UO_OUT_TT_PROJECT4, //EXTERNAL
        input  Tile_X0Y7_UO_OUT_TT_PROJECT5, //EXTERNAL
        input  Tile_X0Y7_UO_OUT_TT_PROJECT6, //EXTERNAL
        input  Tile_X0Y7_UO_OUT_TT_PROJECT7, //EXTERNAL
        input  Tile_X0Y7_UIO_OUT_TT_PROJECT0, //EXTERNAL
        input  Tile_X0Y7_UIO_OUT_TT_PROJECT1, //EXTERNAL
        input  Tile_X0Y7_UIO_OUT_TT_PROJECT2, //EXTERNAL
        input  Tile_X0Y7_UIO_OUT_TT_PROJECT3, //EXTERNAL
        input  Tile_X0Y7_UIO_OUT_TT_PROJECT4, //EXTERNAL
        input  Tile_X0Y7_UIO_OUT_TT_PROJECT5, //EXTERNAL
        input  Tile_X0Y7_UIO_OUT_TT_PROJECT6, //EXTERNAL
        input  Tile_X0Y7_UIO_OUT_TT_PROJECT7, //EXTERNAL
        input  Tile_X0Y7_UIO_OE_TT_PROJECT0, //EXTERNAL
        input  Tile_X0Y7_UIO_OE_TT_PROJECT1, //EXTERNAL
        input  Tile_X0Y7_UIO_OE_TT_PROJECT2, //EXTERNAL
        input  Tile_X0Y7_UIO_OE_TT_PROJECT3, //EXTERNAL
        input  Tile_X0Y7_UIO_OE_TT_PROJECT4, //EXTERNAL
        input  Tile_X0Y7_UIO_OE_TT_PROJECT5, //EXTERNAL
        input  Tile_X0Y7_UIO_OE_TT_PROJECT6, //EXTERNAL
        input  Tile_X0Y7_UIO_OE_TT_PROJECT7, //EXTERNAL
        output  Tile_X0Y7_UI_IN_TT_PROJECT0, //EXTERNAL
        output  Tile_X0Y7_UI_IN_TT_PROJECT1, //EXTERNAL
        output  Tile_X0Y7_UI_IN_TT_PROJECT2, //EXTERNAL
        output  Tile_X0Y7_UI_IN_TT_PROJECT3, //EXTERNAL
        output  Tile_X0Y7_UI_IN_TT_PROJECT4, //EXTERNAL
        output  Tile_X0Y7_UI_IN_TT_PROJECT5, //EXTERNAL
        output  Tile_X0Y7_UI_IN_TT_PROJECT6, //EXTERNAL
        output  Tile_X0Y7_UI_IN_TT_PROJECT7, //EXTERNAL
        output  Tile_X0Y7_UIO_IN_TT_PROJECT0, //EXTERNAL
        output  Tile_X0Y7_UIO_IN_TT_PROJECT1, //EXTERNAL
        output  Tile_X0Y7_UIO_IN_TT_PROJECT2, //EXTERNAL
        output  Tile_X0Y7_UIO_IN_TT_PROJECT3, //EXTERNAL
        output  Tile_X0Y7_UIO_IN_TT_PROJECT4, //EXTERNAL
        output  Tile_X0Y7_UIO_IN_TT_PROJECT5, //EXTERNAL
        output  Tile_X0Y7_UIO_IN_TT_PROJECT6, //EXTERNAL
        output  Tile_X0Y7_UIO_IN_TT_PROJECT7, //EXTERNAL
        output  Tile_X0Y7_ENA_TT_PROJECT, //EXTERNAL
        output  Tile_X0Y7_CLK_TT_PROJECT, //EXTERNAL
        output  Tile_X0Y7_RST_N_TT_PROJECT, //EXTERNAL
        input  Tile_X5Y7_UO_OUT_TT_PROJECT0, //EXTERNAL
        input  Tile_X5Y7_UO_OUT_TT_PROJECT1, //EXTERNAL
        input  Tile_X5Y7_UO_OUT_TT_PROJECT2, //EXTERNAL
        input  Tile_X5Y7_UO_OUT_TT_PROJECT3, //EXTERNAL
        input  Tile_X5Y7_UO_OUT_TT_PROJECT4, //EXTERNAL
        input  Tile_X5Y7_UO_OUT_TT_PROJECT5, //EXTERNAL
        input  Tile_X5Y7_UO_OUT_TT_PROJECT6, //EXTERNAL
        input  Tile_X5Y7_UO_OUT_TT_PROJECT7, //EXTERNAL
        input  Tile_X5Y7_UIO_OUT_TT_PROJECT0, //EXTERNAL
        input  Tile_X5Y7_UIO_OUT_TT_PROJECT1, //EXTERNAL
        input  Tile_X5Y7_UIO_OUT_TT_PROJECT2, //EXTERNAL
        input  Tile_X5Y7_UIO_OUT_TT_PROJECT3, //EXTERNAL
        input  Tile_X5Y7_UIO_OUT_TT_PROJECT4, //EXTERNAL
        input  Tile_X5Y7_UIO_OUT_TT_PROJECT5, //EXTERNAL
        input  Tile_X5Y7_UIO_OUT_TT_PROJECT6, //EXTERNAL
        input  Tile_X5Y7_UIO_OUT_TT_PROJECT7, //EXTERNAL
        input  Tile_X5Y7_UIO_OE_TT_PROJECT0, //EXTERNAL
        input  Tile_X5Y7_UIO_OE_TT_PROJECT1, //EXTERNAL
        input  Tile_X5Y7_UIO_OE_TT_PROJECT2, //EXTERNAL
        input  Tile_X5Y7_UIO_OE_TT_PROJECT3, //EXTERNAL
        input  Tile_X5Y7_UIO_OE_TT_PROJECT4, //EXTERNAL
        input  Tile_X5Y7_UIO_OE_TT_PROJECT5, //EXTERNAL
        input  Tile_X5Y7_UIO_OE_TT_PROJECT6, //EXTERNAL
        input  Tile_X5Y7_UIO_OE_TT_PROJECT7, //EXTERNAL
        output  Tile_X5Y7_UI_IN_TT_PROJECT0, //EXTERNAL
        output  Tile_X5Y7_UI_IN_TT_PROJECT1, //EXTERNAL
        output  Tile_X5Y7_UI_IN_TT_PROJECT2, //EXTERNAL
        output  Tile_X5Y7_UI_IN_TT_PROJECT3, //EXTERNAL
        output  Tile_X5Y7_UI_IN_TT_PROJECT4, //EXTERNAL
        output  Tile_X5Y7_UI_IN_TT_PROJECT5, //EXTERNAL
        output  Tile_X5Y7_UI_IN_TT_PROJECT6, //EXTERNAL
        output  Tile_X5Y7_UI_IN_TT_PROJECT7, //EXTERNAL
        output  Tile_X5Y7_UIO_IN_TT_PROJECT0, //EXTERNAL
        output  Tile_X5Y7_UIO_IN_TT_PROJECT1, //EXTERNAL
        output  Tile_X5Y7_UIO_IN_TT_PROJECT2, //EXTERNAL
        output  Tile_X5Y7_UIO_IN_TT_PROJECT3, //EXTERNAL
        output  Tile_X5Y7_UIO_IN_TT_PROJECT4, //EXTERNAL
        output  Tile_X5Y7_UIO_IN_TT_PROJECT5, //EXTERNAL
        output  Tile_X5Y7_UIO_IN_TT_PROJECT6, //EXTERNAL
        output  Tile_X5Y7_UIO_IN_TT_PROJECT7, //EXTERNAL
        output  Tile_X5Y7_ENA_TT_PROJECT, //EXTERNAL
        output  Tile_X5Y7_CLK_TT_PROJECT, //EXTERNAL
        output  Tile_X5Y7_RST_N_TT_PROJECT, //EXTERNAL
        input  Tile_X0Y8_UO_OUT_TT_PROJECT0, //EXTERNAL
        input  Tile_X0Y8_UO_OUT_TT_PROJECT1, //EXTERNAL
        input  Tile_X0Y8_UO_OUT_TT_PROJECT2, //EXTERNAL
        input  Tile_X0Y8_UO_OUT_TT_PROJECT3, //EXTERNAL
        input  Tile_X0Y8_UO_OUT_TT_PROJECT4, //EXTERNAL
        input  Tile_X0Y8_UO_OUT_TT_PROJECT5, //EXTERNAL
        input  Tile_X0Y8_UO_OUT_TT_PROJECT6, //EXTERNAL
        input  Tile_X0Y8_UO_OUT_TT_PROJECT7, //EXTERNAL
        input  Tile_X0Y8_UIO_OUT_TT_PROJECT0, //EXTERNAL
        input  Tile_X0Y8_UIO_OUT_TT_PROJECT1, //EXTERNAL
        input  Tile_X0Y8_UIO_OUT_TT_PROJECT2, //EXTERNAL
        input  Tile_X0Y8_UIO_OUT_TT_PROJECT3, //EXTERNAL
        input  Tile_X0Y8_UIO_OUT_TT_PROJECT4, //EXTERNAL
        input  Tile_X0Y8_UIO_OUT_TT_PROJECT5, //EXTERNAL
        input  Tile_X0Y8_UIO_OUT_TT_PROJECT6, //EXTERNAL
        input  Tile_X0Y8_UIO_OUT_TT_PROJECT7, //EXTERNAL
        input  Tile_X0Y8_UIO_OE_TT_PROJECT0, //EXTERNAL
        input  Tile_X0Y8_UIO_OE_TT_PROJECT1, //EXTERNAL
        input  Tile_X0Y8_UIO_OE_TT_PROJECT2, //EXTERNAL
        input  Tile_X0Y8_UIO_OE_TT_PROJECT3, //EXTERNAL
        input  Tile_X0Y8_UIO_OE_TT_PROJECT4, //EXTERNAL
        input  Tile_X0Y8_UIO_OE_TT_PROJECT5, //EXTERNAL
        input  Tile_X0Y8_UIO_OE_TT_PROJECT6, //EXTERNAL
        input  Tile_X0Y8_UIO_OE_TT_PROJECT7, //EXTERNAL
        output  Tile_X0Y8_UI_IN_TT_PROJECT0, //EXTERNAL
        output  Tile_X0Y8_UI_IN_TT_PROJECT1, //EXTERNAL
        output  Tile_X0Y8_UI_IN_TT_PROJECT2, //EXTERNAL
        output  Tile_X0Y8_UI_IN_TT_PROJECT3, //EXTERNAL
        output  Tile_X0Y8_UI_IN_TT_PROJECT4, //EXTERNAL
        output  Tile_X0Y8_UI_IN_TT_PROJECT5, //EXTERNAL
        output  Tile_X0Y8_UI_IN_TT_PROJECT6, //EXTERNAL
        output  Tile_X0Y8_UI_IN_TT_PROJECT7, //EXTERNAL
        output  Tile_X0Y8_UIO_IN_TT_PROJECT0, //EXTERNAL
        output  Tile_X0Y8_UIO_IN_TT_PROJECT1, //EXTERNAL
        output  Tile_X0Y8_UIO_IN_TT_PROJECT2, //EXTERNAL
        output  Tile_X0Y8_UIO_IN_TT_PROJECT3, //EXTERNAL
        output  Tile_X0Y8_UIO_IN_TT_PROJECT4, //EXTERNAL
        output  Tile_X0Y8_UIO_IN_TT_PROJECT5, //EXTERNAL
        output  Tile_X0Y8_UIO_IN_TT_PROJECT6, //EXTERNAL
        output  Tile_X0Y8_UIO_IN_TT_PROJECT7, //EXTERNAL
        output  Tile_X0Y8_ENA_TT_PROJECT, //EXTERNAL
        output  Tile_X0Y8_CLK_TT_PROJECT, //EXTERNAL
        output  Tile_X0Y8_RST_N_TT_PROJECT, //EXTERNAL
        input  Tile_X5Y8_UO_OUT_TT_PROJECT0, //EXTERNAL
        input  Tile_X5Y8_UO_OUT_TT_PROJECT1, //EXTERNAL
        input  Tile_X5Y8_UO_OUT_TT_PROJECT2, //EXTERNAL
        input  Tile_X5Y8_UO_OUT_TT_PROJECT3, //EXTERNAL
        input  Tile_X5Y8_UO_OUT_TT_PROJECT4, //EXTERNAL
        input  Tile_X5Y8_UO_OUT_TT_PROJECT5, //EXTERNAL
        input  Tile_X5Y8_UO_OUT_TT_PROJECT6, //EXTERNAL
        input  Tile_X5Y8_UO_OUT_TT_PROJECT7, //EXTERNAL
        input  Tile_X5Y8_UIO_OUT_TT_PROJECT0, //EXTERNAL
        input  Tile_X5Y8_UIO_OUT_TT_PROJECT1, //EXTERNAL
        input  Tile_X5Y8_UIO_OUT_TT_PROJECT2, //EXTERNAL
        input  Tile_X5Y8_UIO_OUT_TT_PROJECT3, //EXTERNAL
        input  Tile_X5Y8_UIO_OUT_TT_PROJECT4, //EXTERNAL
        input  Tile_X5Y8_UIO_OUT_TT_PROJECT5, //EXTERNAL
        input  Tile_X5Y8_UIO_OUT_TT_PROJECT6, //EXTERNAL
        input  Tile_X5Y8_UIO_OUT_TT_PROJECT7, //EXTERNAL
        input  Tile_X5Y8_UIO_OE_TT_PROJECT0, //EXTERNAL
        input  Tile_X5Y8_UIO_OE_TT_PROJECT1, //EXTERNAL
        input  Tile_X5Y8_UIO_OE_TT_PROJECT2, //EXTERNAL
        input  Tile_X5Y8_UIO_OE_TT_PROJECT3, //EXTERNAL
        input  Tile_X5Y8_UIO_OE_TT_PROJECT4, //EXTERNAL
        input  Tile_X5Y8_UIO_OE_TT_PROJECT5, //EXTERNAL
        input  Tile_X5Y8_UIO_OE_TT_PROJECT6, //EXTERNAL
        input  Tile_X5Y8_UIO_OE_TT_PROJECT7, //EXTERNAL
        output  Tile_X5Y8_UI_IN_TT_PROJECT0, //EXTERNAL
        output  Tile_X5Y8_UI_IN_TT_PROJECT1, //EXTERNAL
        output  Tile_X5Y8_UI_IN_TT_PROJECT2, //EXTERNAL
        output  Tile_X5Y8_UI_IN_TT_PROJECT3, //EXTERNAL
        output  Tile_X5Y8_UI_IN_TT_PROJECT4, //EXTERNAL
        output  Tile_X5Y8_UI_IN_TT_PROJECT5, //EXTERNAL
        output  Tile_X5Y8_UI_IN_TT_PROJECT6, //EXTERNAL
        output  Tile_X5Y8_UI_IN_TT_PROJECT7, //EXTERNAL
        output  Tile_X5Y8_UIO_IN_TT_PROJECT0, //EXTERNAL
        output  Tile_X5Y8_UIO_IN_TT_PROJECT1, //EXTERNAL
        output  Tile_X5Y8_UIO_IN_TT_PROJECT2, //EXTERNAL
        output  Tile_X5Y8_UIO_IN_TT_PROJECT3, //EXTERNAL
        output  Tile_X5Y8_UIO_IN_TT_PROJECT4, //EXTERNAL
        output  Tile_X5Y8_UIO_IN_TT_PROJECT5, //EXTERNAL
        output  Tile_X5Y8_UIO_IN_TT_PROJECT6, //EXTERNAL
        output  Tile_X5Y8_UIO_IN_TT_PROJECT7, //EXTERNAL
        output  Tile_X5Y8_ENA_TT_PROJECT, //EXTERNAL
        output  Tile_X5Y8_CLK_TT_PROJECT, //EXTERNAL
        output  Tile_X5Y8_RST_N_TT_PROJECT, //EXTERNAL
        input  Tile_X1Y9_A_O_top, //EXTERNAL
        output  Tile_X1Y9_A_I_top, //EXTERNAL
        output  Tile_X1Y9_A_T_top, //EXTERNAL
        input  Tile_X1Y9_B_O_top, //EXTERNAL
        output  Tile_X1Y9_B_I_top, //EXTERNAL
        output  Tile_X1Y9_B_T_top, //EXTERNAL
        input  Tile_X1Y9_C_O_top, //EXTERNAL
        output  Tile_X1Y9_C_I_top, //EXTERNAL
        output  Tile_X1Y9_C_T_top, //EXTERNAL
        input  Tile_X1Y9_D_O_top, //EXTERNAL
        output  Tile_X1Y9_D_I_top, //EXTERNAL
        output  Tile_X1Y9_D_T_top, //EXTERNAL
        input  Tile_X2Y9_A_O_top, //EXTERNAL
        output  Tile_X2Y9_A_I_top, //EXTERNAL
        output  Tile_X2Y9_A_T_top, //EXTERNAL
        input  Tile_X2Y9_B_O_top, //EXTERNAL
        output  Tile_X2Y9_B_I_top, //EXTERNAL
        output  Tile_X2Y9_B_T_top, //EXTERNAL
        input  Tile_X2Y9_C_O_top, //EXTERNAL
        output  Tile_X2Y9_C_I_top, //EXTERNAL
        output  Tile_X2Y9_C_T_top, //EXTERNAL
        input  Tile_X2Y9_D_O_top, //EXTERNAL
        output  Tile_X2Y9_D_I_top, //EXTERNAL
        output  Tile_X2Y9_D_T_top, //EXTERNAL
        input  Tile_X3Y9_A_O_top, //EXTERNAL
        output  Tile_X3Y9_A_I_top, //EXTERNAL
        output  Tile_X3Y9_A_T_top, //EXTERNAL
        input  Tile_X3Y9_B_O_top, //EXTERNAL
        output  Tile_X3Y9_B_I_top, //EXTERNAL
        output  Tile_X3Y9_B_T_top, //EXTERNAL
        input  Tile_X3Y9_C_O_top, //EXTERNAL
        output  Tile_X3Y9_C_I_top, //EXTERNAL
        output  Tile_X3Y9_C_T_top, //EXTERNAL
        input  Tile_X3Y9_D_O_top, //EXTERNAL
        output  Tile_X3Y9_D_I_top, //EXTERNAL
        output  Tile_X3Y9_D_T_top, //EXTERNAL
        input  Tile_X4Y9_A_O_top, //EXTERNAL
        output  Tile_X4Y9_A_I_top, //EXTERNAL
        output  Tile_X4Y9_A_T_top, //EXTERNAL
        input  Tile_X4Y9_B_O_top, //EXTERNAL
        output  Tile_X4Y9_B_I_top, //EXTERNAL
        output  Tile_X4Y9_B_T_top, //EXTERNAL
        input  Tile_X4Y9_C_O_top, //EXTERNAL
        output  Tile_X4Y9_C_I_top, //EXTERNAL
        output  Tile_X4Y9_C_T_top, //EXTERNAL
        input  Tile_X4Y9_D_O_top, //EXTERNAL
        output  Tile_X4Y9_D_I_top, //EXTERNAL
        output  Tile_X4Y9_D_T_top, //EXTERNAL
        input  [(FrameBitsPerRow*10)-1:0] FrameData, //CONFIG_PORT
        input  [(MaxFramesPerCol*6)-1:0] FrameStrobe, //CONFIG_PORT
        input  UserCLK
);

 //signal declarations

wire Tile_X0Y0_UserCLKo;
wire Tile_X1Y0_UserCLKo;
wire Tile_X2Y0_UserCLKo;
wire Tile_X3Y0_UserCLKo;
wire Tile_X4Y0_UserCLKo;
wire Tile_X5Y0_UserCLKo;
wire Tile_X0Y1_UserCLKo;
wire Tile_X1Y1_UserCLKo;
wire Tile_X2Y1_UserCLKo;
wire Tile_X3Y1_UserCLKo;
wire Tile_X4Y1_UserCLKo;
wire Tile_X5Y1_UserCLKo;
wire Tile_X0Y2_UserCLKo;
wire Tile_X1Y2_UserCLKo;
wire Tile_X2Y2_UserCLKo;
wire Tile_X3Y2_UserCLKo;
wire Tile_X4Y2_UserCLKo;
wire Tile_X5Y2_UserCLKo;
wire Tile_X0Y3_UserCLKo;
wire Tile_X1Y3_UserCLKo;
wire Tile_X2Y3_UserCLKo;
wire Tile_X3Y3_UserCLKo;
wire Tile_X4Y3_UserCLKo;
wire Tile_X5Y3_UserCLKo;
wire Tile_X0Y4_UserCLKo;
wire Tile_X1Y4_UserCLKo;
wire Tile_X2Y4_UserCLKo;
wire Tile_X3Y4_UserCLKo;
wire Tile_X4Y4_UserCLKo;
wire Tile_X5Y4_UserCLKo;
wire Tile_X0Y5_UserCLKo;
wire Tile_X1Y5_UserCLKo;
wire Tile_X2Y5_UserCLKo;
wire Tile_X3Y5_UserCLKo;
wire Tile_X4Y5_UserCLKo;
wire Tile_X5Y5_UserCLKo;
wire Tile_X0Y6_UserCLKo;
wire Tile_X1Y6_UserCLKo;
wire Tile_X2Y6_UserCLKo;
wire Tile_X3Y6_UserCLKo;
wire Tile_X4Y6_UserCLKo;
wire Tile_X5Y6_UserCLKo;
wire Tile_X0Y7_UserCLKo;
wire Tile_X1Y7_UserCLKo;
wire Tile_X2Y7_UserCLKo;
wire Tile_X3Y7_UserCLKo;
wire Tile_X4Y7_UserCLKo;
wire Tile_X5Y7_UserCLKo;
wire Tile_X0Y8_UserCLKo;
wire Tile_X1Y8_UserCLKo;
wire Tile_X2Y8_UserCLKo;
wire Tile_X3Y8_UserCLKo;
wire Tile_X4Y8_UserCLKo;
wire Tile_X5Y8_UserCLKo;
wire Tile_X0Y9_UserCLKo;
wire Tile_X1Y9_UserCLKo;
wire Tile_X2Y9_UserCLKo;
wire Tile_X3Y9_UserCLKo;
wire Tile_X4Y9_UserCLKo;
wire Tile_X5Y9_UserCLKo;
 //configuration signal declarations

wire[FrameBitsPerRow -1:0] Row_Y0_FrameData;
wire[FrameBitsPerRow -1:0] Row_Y1_FrameData;
wire[FrameBitsPerRow -1:0] Row_Y2_FrameData;
wire[FrameBitsPerRow -1:0] Row_Y3_FrameData;
wire[FrameBitsPerRow -1:0] Row_Y4_FrameData;
wire[FrameBitsPerRow -1:0] Row_Y5_FrameData;
wire[FrameBitsPerRow -1:0] Row_Y6_FrameData;
wire[FrameBitsPerRow -1:0] Row_Y7_FrameData;
wire[FrameBitsPerRow -1:0] Row_Y8_FrameData;
wire[FrameBitsPerRow -1:0] Row_Y9_FrameData;
wire[MaxFramesPerCol - 1:0] Column_X0_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Column_X1_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Column_X2_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Column_X3_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Column_X4_FrameStrobe;
wire[MaxFramesPerCol - 1:0] Column_X5_FrameStrobe;
wire[FrameBitsPerRow - 1:0] Tile_X0Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y0_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y1_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y2_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y3_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y4_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y5_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y6_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y7_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y8_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y8_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y8_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y8_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y8_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y8_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X0Y9_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X1Y9_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X2Y9_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X3Y9_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X4Y9_FrameData_O;
wire[FrameBitsPerRow - 1:0] Tile_X5Y9_FrameData_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y0_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y1_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y2_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y3_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y4_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y5_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y6_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y7_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y8_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y9_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y9_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y9_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y9_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y9_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y9_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X0Y10_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X1Y10_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X2Y10_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X3Y10_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X4Y10_FrameStrobe_O;
wire[MaxFramesPerCol - 1:0] Tile_X5Y10_FrameStrobe_O;
 //tile-to-tile signal declarations
wire[3:0] Tile_X0Y0_S1BEG;
wire[7:0] Tile_X0Y0_S2BEG;
wire[7:0] Tile_X0Y0_S2BEGb;
wire[15:0] Tile_X0Y0_S4BEG;
wire[3:0] Tile_X1Y0_S1BEG;
wire[7:0] Tile_X1Y0_S2BEG;
wire[7:0] Tile_X1Y0_S2BEGb;
wire[15:0] Tile_X1Y0_S4BEG;
wire[15:0] Tile_X1Y0_SS4BEG;
wire[3:0] Tile_X2Y0_S1BEG;
wire[7:0] Tile_X2Y0_S2BEG;
wire[7:0] Tile_X2Y0_S2BEGb;
wire[15:0] Tile_X2Y0_S4BEG;
wire[15:0] Tile_X2Y0_SS4BEG;
wire[3:0] Tile_X3Y0_S1BEG;
wire[7:0] Tile_X3Y0_S2BEG;
wire[7:0] Tile_X3Y0_S2BEGb;
wire[15:0] Tile_X3Y0_S4BEG;
wire[15:0] Tile_X3Y0_SS4BEG;
wire[3:0] Tile_X4Y0_S1BEG;
wire[7:0] Tile_X4Y0_S2BEG;
wire[7:0] Tile_X4Y0_S2BEGb;
wire[15:0] Tile_X4Y0_S4BEG;
wire[15:0] Tile_X4Y0_SS4BEG;
wire[3:0] Tile_X5Y0_S1BEG;
wire[7:0] Tile_X5Y0_S2BEG;
wire[7:0] Tile_X5Y0_S2BEGb;
wire[15:0] Tile_X5Y0_S4BEG;
wire[3:0] Tile_X0Y1_N1BEG;
wire[7:0] Tile_X0Y1_N2BEG;
wire[7:0] Tile_X0Y1_N2BEGb;
wire[15:0] Tile_X0Y1_N4BEG;
wire[3:0] Tile_X0Y1_S1BEG;
wire[7:0] Tile_X0Y1_S2BEG;
wire[7:0] Tile_X0Y1_S2BEGb;
wire[15:0] Tile_X0Y1_S4BEG;
wire[3:0] Tile_X0Y1_E1BEG;
wire[7:0] Tile_X0Y1_E2BEG;
wire[7:0] Tile_X0Y1_E2BEGb;
wire[15:0] Tile_X0Y1_EE4BEG;
wire[11:0] Tile_X0Y1_E6BEG;
wire[7:0] Tile_X0Y1_top2bot_UIO_IN;
wire[3:0] Tile_X1Y1_N1BEG;
wire[7:0] Tile_X1Y1_N2BEG;
wire[7:0] Tile_X1Y1_N2BEGb;
wire[15:0] Tile_X1Y1_N4BEG;
wire[15:0] Tile_X1Y1_NN4BEG;
wire[3:0] Tile_X1Y1_E1BEG;
wire[7:0] Tile_X1Y1_E2BEG;
wire[7:0] Tile_X1Y1_E2BEGb;
wire[15:0] Tile_X1Y1_EE4BEG;
wire[11:0] Tile_X1Y1_E6BEG;
wire[3:0] Tile_X1Y1_S1BEG;
wire[7:0] Tile_X1Y1_S2BEG;
wire[7:0] Tile_X1Y1_S2BEGb;
wire[15:0] Tile_X1Y1_S4BEG;
wire[15:0] Tile_X1Y1_SS4BEG;
wire[3:0] Tile_X1Y1_W1BEG;
wire[7:0] Tile_X1Y1_W2BEG;
wire[7:0] Tile_X1Y1_W2BEGb;
wire[15:0] Tile_X1Y1_WW4BEG;
wire[11:0] Tile_X1Y1_W6BEG;
wire[0:0] Tile_X1Y1_Co;
wire[3:0] Tile_X2Y1_N1BEG;
wire[7:0] Tile_X2Y1_N2BEG;
wire[7:0] Tile_X2Y1_N2BEGb;
wire[15:0] Tile_X2Y1_N4BEG;
wire[15:0] Tile_X2Y1_NN4BEG;
wire[3:0] Tile_X2Y1_E1BEG;
wire[7:0] Tile_X2Y1_E2BEG;
wire[7:0] Tile_X2Y1_E2BEGb;
wire[15:0] Tile_X2Y1_EE4BEG;
wire[11:0] Tile_X2Y1_E6BEG;
wire[3:0] Tile_X2Y1_S1BEG;
wire[7:0] Tile_X2Y1_S2BEG;
wire[7:0] Tile_X2Y1_S2BEGb;
wire[15:0] Tile_X2Y1_S4BEG;
wire[15:0] Tile_X2Y1_SS4BEG;
wire[3:0] Tile_X2Y1_W1BEG;
wire[7:0] Tile_X2Y1_W2BEG;
wire[7:0] Tile_X2Y1_W2BEGb;
wire[15:0] Tile_X2Y1_WW4BEG;
wire[11:0] Tile_X2Y1_W6BEG;
wire[0:0] Tile_X2Y1_Co;
wire[3:0] Tile_X3Y1_N1BEG;
wire[7:0] Tile_X3Y1_N2BEG;
wire[7:0] Tile_X3Y1_N2BEGb;
wire[15:0] Tile_X3Y1_N4BEG;
wire[15:0] Tile_X3Y1_NN4BEG;
wire[3:0] Tile_X3Y1_E1BEG;
wire[7:0] Tile_X3Y1_E2BEG;
wire[7:0] Tile_X3Y1_E2BEGb;
wire[15:0] Tile_X3Y1_EE4BEG;
wire[11:0] Tile_X3Y1_E6BEG;
wire[3:0] Tile_X3Y1_S1BEG;
wire[7:0] Tile_X3Y1_S2BEG;
wire[7:0] Tile_X3Y1_S2BEGb;
wire[15:0] Tile_X3Y1_S4BEG;
wire[15:0] Tile_X3Y1_SS4BEG;
wire[3:0] Tile_X3Y1_W1BEG;
wire[7:0] Tile_X3Y1_W2BEG;
wire[7:0] Tile_X3Y1_W2BEGb;
wire[15:0] Tile_X3Y1_WW4BEG;
wire[11:0] Tile_X3Y1_W6BEG;
wire[0:0] Tile_X3Y1_Co;
wire[3:0] Tile_X4Y1_N1BEG;
wire[7:0] Tile_X4Y1_N2BEG;
wire[7:0] Tile_X4Y1_N2BEGb;
wire[15:0] Tile_X4Y1_N4BEG;
wire[15:0] Tile_X4Y1_NN4BEG;
wire[3:0] Tile_X4Y1_E1BEG;
wire[7:0] Tile_X4Y1_E2BEG;
wire[7:0] Tile_X4Y1_E2BEGb;
wire[15:0] Tile_X4Y1_EE4BEG;
wire[11:0] Tile_X4Y1_E6BEG;
wire[3:0] Tile_X4Y1_S1BEG;
wire[7:0] Tile_X4Y1_S2BEG;
wire[7:0] Tile_X4Y1_S2BEGb;
wire[15:0] Tile_X4Y1_S4BEG;
wire[15:0] Tile_X4Y1_SS4BEG;
wire[3:0] Tile_X4Y1_W1BEG;
wire[7:0] Tile_X4Y1_W2BEG;
wire[7:0] Tile_X4Y1_W2BEGb;
wire[15:0] Tile_X4Y1_WW4BEG;
wire[11:0] Tile_X4Y1_W6BEG;
wire[0:0] Tile_X4Y1_Co;
wire[3:0] Tile_X5Y1_N1BEG;
wire[7:0] Tile_X5Y1_N2BEG;
wire[7:0] Tile_X5Y1_N2BEGb;
wire[15:0] Tile_X5Y1_N4BEG;
wire[3:0] Tile_X5Y1_S1BEG;
wire[7:0] Tile_X5Y1_S2BEG;
wire[7:0] Tile_X5Y1_S2BEGb;
wire[15:0] Tile_X5Y1_S4BEG;
wire[3:0] Tile_X5Y1_W1BEG;
wire[7:0] Tile_X5Y1_W2BEG;
wire[7:0] Tile_X5Y1_W2BEGb;
wire[15:0] Tile_X5Y1_WW4BEG;
wire[11:0] Tile_X5Y1_W6BEG;
wire[15:0] Tile_X5Y1_top2bot_DIN;
wire[15:0] Tile_X5Y1_top2bot_BM;
wire[4:0] Tile_X5Y1_top2bot_ADDR;
wire[3:0] Tile_X0Y2_N1BEG;
wire[7:0] Tile_X0Y2_N2BEG;
wire[7:0] Tile_X0Y2_N2BEGb;
wire[15:0] Tile_X0Y2_N4BEG;
wire[3:0] Tile_X0Y2_S1BEG;
wire[7:0] Tile_X0Y2_S2BEG;
wire[7:0] Tile_X0Y2_S2BEGb;
wire[15:0] Tile_X0Y2_S4BEG;
wire[3:0] Tile_X0Y2_E1BEG;
wire[7:0] Tile_X0Y2_E2BEG;
wire[7:0] Tile_X0Y2_E2BEGb;
wire[15:0] Tile_X0Y2_EE4BEG;
wire[11:0] Tile_X0Y2_E6BEG;
wire[7:0] Tile_X0Y2_bot2top_UIO_OUT;
wire[7:0] Tile_X0Y2_bot2top_UIO_OE;
wire[3:0] Tile_X1Y2_N1BEG;
wire[7:0] Tile_X1Y2_N2BEG;
wire[7:0] Tile_X1Y2_N2BEGb;
wire[15:0] Tile_X1Y2_N4BEG;
wire[15:0] Tile_X1Y2_NN4BEG;
wire[3:0] Tile_X1Y2_E1BEG;
wire[7:0] Tile_X1Y2_E2BEG;
wire[7:0] Tile_X1Y2_E2BEGb;
wire[15:0] Tile_X1Y2_EE4BEG;
wire[11:0] Tile_X1Y2_E6BEG;
wire[3:0] Tile_X1Y2_S1BEG;
wire[7:0] Tile_X1Y2_S2BEG;
wire[7:0] Tile_X1Y2_S2BEGb;
wire[15:0] Tile_X1Y2_S4BEG;
wire[15:0] Tile_X1Y2_SS4BEG;
wire[3:0] Tile_X1Y2_W1BEG;
wire[7:0] Tile_X1Y2_W2BEG;
wire[7:0] Tile_X1Y2_W2BEGb;
wire[15:0] Tile_X1Y2_WW4BEG;
wire[11:0] Tile_X1Y2_W6BEG;
wire[0:0] Tile_X1Y2_Co;
wire[3:0] Tile_X2Y2_N1BEG;
wire[7:0] Tile_X2Y2_N2BEG;
wire[7:0] Tile_X2Y2_N2BEGb;
wire[15:0] Tile_X2Y2_N4BEG;
wire[15:0] Tile_X2Y2_NN4BEG;
wire[3:0] Tile_X2Y2_E1BEG;
wire[7:0] Tile_X2Y2_E2BEG;
wire[7:0] Tile_X2Y2_E2BEGb;
wire[15:0] Tile_X2Y2_EE4BEG;
wire[11:0] Tile_X2Y2_E6BEG;
wire[3:0] Tile_X2Y2_S1BEG;
wire[7:0] Tile_X2Y2_S2BEG;
wire[7:0] Tile_X2Y2_S2BEGb;
wire[15:0] Tile_X2Y2_S4BEG;
wire[15:0] Tile_X2Y2_SS4BEG;
wire[3:0] Tile_X2Y2_W1BEG;
wire[7:0] Tile_X2Y2_W2BEG;
wire[7:0] Tile_X2Y2_W2BEGb;
wire[15:0] Tile_X2Y2_WW4BEG;
wire[11:0] Tile_X2Y2_W6BEG;
wire[0:0] Tile_X2Y2_Co;
wire[3:0] Tile_X3Y2_N1BEG;
wire[7:0] Tile_X3Y2_N2BEG;
wire[7:0] Tile_X3Y2_N2BEGb;
wire[15:0] Tile_X3Y2_N4BEG;
wire[15:0] Tile_X3Y2_NN4BEG;
wire[3:0] Tile_X3Y2_E1BEG;
wire[7:0] Tile_X3Y2_E2BEG;
wire[7:0] Tile_X3Y2_E2BEGb;
wire[15:0] Tile_X3Y2_EE4BEG;
wire[11:0] Tile_X3Y2_E6BEG;
wire[3:0] Tile_X3Y2_S1BEG;
wire[7:0] Tile_X3Y2_S2BEG;
wire[7:0] Tile_X3Y2_S2BEGb;
wire[15:0] Tile_X3Y2_S4BEG;
wire[15:0] Tile_X3Y2_SS4BEG;
wire[3:0] Tile_X3Y2_W1BEG;
wire[7:0] Tile_X3Y2_W2BEG;
wire[7:0] Tile_X3Y2_W2BEGb;
wire[15:0] Tile_X3Y2_WW4BEG;
wire[11:0] Tile_X3Y2_W6BEG;
wire[0:0] Tile_X3Y2_Co;
wire[3:0] Tile_X4Y2_N1BEG;
wire[7:0] Tile_X4Y2_N2BEG;
wire[7:0] Tile_X4Y2_N2BEGb;
wire[15:0] Tile_X4Y2_N4BEG;
wire[15:0] Tile_X4Y2_NN4BEG;
wire[3:0] Tile_X4Y2_E1BEG;
wire[7:0] Tile_X4Y2_E2BEG;
wire[7:0] Tile_X4Y2_E2BEGb;
wire[15:0] Tile_X4Y2_EE4BEG;
wire[11:0] Tile_X4Y2_E6BEG;
wire[3:0] Tile_X4Y2_S1BEG;
wire[7:0] Tile_X4Y2_S2BEG;
wire[7:0] Tile_X4Y2_S2BEGb;
wire[15:0] Tile_X4Y2_S4BEG;
wire[15:0] Tile_X4Y2_SS4BEG;
wire[3:0] Tile_X4Y2_W1BEG;
wire[7:0] Tile_X4Y2_W2BEG;
wire[7:0] Tile_X4Y2_W2BEGb;
wire[15:0] Tile_X4Y2_WW4BEG;
wire[11:0] Tile_X4Y2_W6BEG;
wire[0:0] Tile_X4Y2_Co;
wire[3:0] Tile_X5Y2_N1BEG;
wire[7:0] Tile_X5Y2_N2BEG;
wire[7:0] Tile_X5Y2_N2BEGb;
wire[15:0] Tile_X5Y2_N4BEG;
wire[3:0] Tile_X5Y2_S1BEG;
wire[7:0] Tile_X5Y2_S2BEG;
wire[7:0] Tile_X5Y2_S2BEGb;
wire[15:0] Tile_X5Y2_S4BEG;
wire[3:0] Tile_X5Y2_W1BEG;
wire[7:0] Tile_X5Y2_W2BEG;
wire[7:0] Tile_X5Y2_W2BEGb;
wire[15:0] Tile_X5Y2_WW4BEG;
wire[11:0] Tile_X5Y2_W6BEG;
wire[15:0] Tile_X5Y2_bot2top_DOUT;
wire[3:0] Tile_X0Y3_N1BEG;
wire[7:0] Tile_X0Y3_N2BEG;
wire[7:0] Tile_X0Y3_N2BEGb;
wire[15:0] Tile_X0Y3_N4BEG;
wire[3:0] Tile_X0Y3_S1BEG;
wire[7:0] Tile_X0Y3_S2BEG;
wire[7:0] Tile_X0Y3_S2BEGb;
wire[15:0] Tile_X0Y3_S4BEG;
wire[3:0] Tile_X0Y3_E1BEG;
wire[7:0] Tile_X0Y3_E2BEG;
wire[7:0] Tile_X0Y3_E2BEGb;
wire[15:0] Tile_X0Y3_EE4BEG;
wire[11:0] Tile_X0Y3_E6BEG;
wire[3:0] Tile_X1Y3_N1BEG;
wire[7:0] Tile_X1Y3_N2BEG;
wire[7:0] Tile_X1Y3_N2BEGb;
wire[15:0] Tile_X1Y3_N4BEG;
wire[15:0] Tile_X1Y3_NN4BEG;
wire[3:0] Tile_X1Y3_E1BEG;
wire[7:0] Tile_X1Y3_E2BEG;
wire[7:0] Tile_X1Y3_E2BEGb;
wire[15:0] Tile_X1Y3_EE4BEG;
wire[11:0] Tile_X1Y3_E6BEG;
wire[3:0] Tile_X1Y3_S1BEG;
wire[7:0] Tile_X1Y3_S2BEG;
wire[7:0] Tile_X1Y3_S2BEGb;
wire[15:0] Tile_X1Y3_S4BEG;
wire[15:0] Tile_X1Y3_SS4BEG;
wire[3:0] Tile_X1Y3_W1BEG;
wire[7:0] Tile_X1Y3_W2BEG;
wire[7:0] Tile_X1Y3_W2BEGb;
wire[15:0] Tile_X1Y3_WW4BEG;
wire[11:0] Tile_X1Y3_W6BEG;
wire[0:0] Tile_X1Y3_Co;
wire[3:0] Tile_X2Y3_N1BEG;
wire[7:0] Tile_X2Y3_N2BEG;
wire[7:0] Tile_X2Y3_N2BEGb;
wire[15:0] Tile_X2Y3_N4BEG;
wire[15:0] Tile_X2Y3_NN4BEG;
wire[3:0] Tile_X2Y3_E1BEG;
wire[7:0] Tile_X2Y3_E2BEG;
wire[7:0] Tile_X2Y3_E2BEGb;
wire[15:0] Tile_X2Y3_EE4BEG;
wire[11:0] Tile_X2Y3_E6BEG;
wire[3:0] Tile_X2Y3_S1BEG;
wire[7:0] Tile_X2Y3_S2BEG;
wire[7:0] Tile_X2Y3_S2BEGb;
wire[15:0] Tile_X2Y3_S4BEG;
wire[15:0] Tile_X2Y3_SS4BEG;
wire[3:0] Tile_X2Y3_W1BEG;
wire[7:0] Tile_X2Y3_W2BEG;
wire[7:0] Tile_X2Y3_W2BEGb;
wire[15:0] Tile_X2Y3_WW4BEG;
wire[11:0] Tile_X2Y3_W6BEG;
wire[0:0] Tile_X2Y3_Co;
wire[3:0] Tile_X3Y3_N1BEG;
wire[7:0] Tile_X3Y3_N2BEG;
wire[7:0] Tile_X3Y3_N2BEGb;
wire[15:0] Tile_X3Y3_N4BEG;
wire[15:0] Tile_X3Y3_NN4BEG;
wire[3:0] Tile_X3Y3_E1BEG;
wire[7:0] Tile_X3Y3_E2BEG;
wire[7:0] Tile_X3Y3_E2BEGb;
wire[15:0] Tile_X3Y3_EE4BEG;
wire[11:0] Tile_X3Y3_E6BEG;
wire[3:0] Tile_X3Y3_S1BEG;
wire[7:0] Tile_X3Y3_S2BEG;
wire[7:0] Tile_X3Y3_S2BEGb;
wire[15:0] Tile_X3Y3_S4BEG;
wire[15:0] Tile_X3Y3_SS4BEG;
wire[3:0] Tile_X3Y3_W1BEG;
wire[7:0] Tile_X3Y3_W2BEG;
wire[7:0] Tile_X3Y3_W2BEGb;
wire[15:0] Tile_X3Y3_WW4BEG;
wire[11:0] Tile_X3Y3_W6BEG;
wire[0:0] Tile_X3Y3_Co;
wire[3:0] Tile_X4Y3_N1BEG;
wire[7:0] Tile_X4Y3_N2BEG;
wire[7:0] Tile_X4Y3_N2BEGb;
wire[15:0] Tile_X4Y3_N4BEG;
wire[15:0] Tile_X4Y3_NN4BEG;
wire[3:0] Tile_X4Y3_E1BEG;
wire[7:0] Tile_X4Y3_E2BEG;
wire[7:0] Tile_X4Y3_E2BEGb;
wire[15:0] Tile_X4Y3_EE4BEG;
wire[11:0] Tile_X4Y3_E6BEG;
wire[3:0] Tile_X4Y3_S1BEG;
wire[7:0] Tile_X4Y3_S2BEG;
wire[7:0] Tile_X4Y3_S2BEGb;
wire[15:0] Tile_X4Y3_S4BEG;
wire[15:0] Tile_X4Y3_SS4BEG;
wire[3:0] Tile_X4Y3_W1BEG;
wire[7:0] Tile_X4Y3_W2BEG;
wire[7:0] Tile_X4Y3_W2BEGb;
wire[15:0] Tile_X4Y3_WW4BEG;
wire[11:0] Tile_X4Y3_W6BEG;
wire[0:0] Tile_X4Y3_Co;
wire[3:0] Tile_X5Y3_N1BEG;
wire[7:0] Tile_X5Y3_N2BEG;
wire[7:0] Tile_X5Y3_N2BEGb;
wire[15:0] Tile_X5Y3_N4BEG;
wire[3:0] Tile_X5Y3_S1BEG;
wire[7:0] Tile_X5Y3_S2BEG;
wire[7:0] Tile_X5Y3_S2BEGb;
wire[15:0] Tile_X5Y3_S4BEG;
wire[3:0] Tile_X5Y3_W1BEG;
wire[7:0] Tile_X5Y3_W2BEG;
wire[7:0] Tile_X5Y3_W2BEGb;
wire[15:0] Tile_X5Y3_WW4BEG;
wire[11:0] Tile_X5Y3_W6BEG;
wire[7:0] Tile_X5Y3_top2bot_UIO_IN;
wire[3:0] Tile_X0Y4_N1BEG;
wire[7:0] Tile_X0Y4_N2BEG;
wire[7:0] Tile_X0Y4_N2BEGb;
wire[15:0] Tile_X0Y4_N4BEG;
wire[3:0] Tile_X0Y4_S1BEG;
wire[7:0] Tile_X0Y4_S2BEG;
wire[7:0] Tile_X0Y4_S2BEGb;
wire[15:0] Tile_X0Y4_S4BEG;
wire[3:0] Tile_X0Y4_E1BEG;
wire[7:0] Tile_X0Y4_E2BEG;
wire[7:0] Tile_X0Y4_E2BEGb;
wire[15:0] Tile_X0Y4_EE4BEG;
wire[11:0] Tile_X0Y4_E6BEG;
wire[3:0] Tile_X1Y4_N1BEG;
wire[7:0] Tile_X1Y4_N2BEG;
wire[7:0] Tile_X1Y4_N2BEGb;
wire[15:0] Tile_X1Y4_N4BEG;
wire[15:0] Tile_X1Y4_NN4BEG;
wire[3:0] Tile_X1Y4_E1BEG;
wire[7:0] Tile_X1Y4_E2BEG;
wire[7:0] Tile_X1Y4_E2BEGb;
wire[15:0] Tile_X1Y4_EE4BEG;
wire[11:0] Tile_X1Y4_E6BEG;
wire[3:0] Tile_X1Y4_S1BEG;
wire[7:0] Tile_X1Y4_S2BEG;
wire[7:0] Tile_X1Y4_S2BEGb;
wire[15:0] Tile_X1Y4_S4BEG;
wire[15:0] Tile_X1Y4_SS4BEG;
wire[3:0] Tile_X1Y4_W1BEG;
wire[7:0] Tile_X1Y4_W2BEG;
wire[7:0] Tile_X1Y4_W2BEGb;
wire[15:0] Tile_X1Y4_WW4BEG;
wire[11:0] Tile_X1Y4_W6BEG;
wire[0:0] Tile_X1Y4_Co;
wire[3:0] Tile_X2Y4_N1BEG;
wire[7:0] Tile_X2Y4_N2BEG;
wire[7:0] Tile_X2Y4_N2BEGb;
wire[15:0] Tile_X2Y4_N4BEG;
wire[15:0] Tile_X2Y4_NN4BEG;
wire[3:0] Tile_X2Y4_E1BEG;
wire[7:0] Tile_X2Y4_E2BEG;
wire[7:0] Tile_X2Y4_E2BEGb;
wire[15:0] Tile_X2Y4_EE4BEG;
wire[11:0] Tile_X2Y4_E6BEG;
wire[3:0] Tile_X2Y4_S1BEG;
wire[7:0] Tile_X2Y4_S2BEG;
wire[7:0] Tile_X2Y4_S2BEGb;
wire[15:0] Tile_X2Y4_S4BEG;
wire[15:0] Tile_X2Y4_SS4BEG;
wire[3:0] Tile_X2Y4_W1BEG;
wire[7:0] Tile_X2Y4_W2BEG;
wire[7:0] Tile_X2Y4_W2BEGb;
wire[15:0] Tile_X2Y4_WW4BEG;
wire[11:0] Tile_X2Y4_W6BEG;
wire[0:0] Tile_X2Y4_Co;
wire[3:0] Tile_X3Y4_N1BEG;
wire[7:0] Tile_X3Y4_N2BEG;
wire[7:0] Tile_X3Y4_N2BEGb;
wire[15:0] Tile_X3Y4_N4BEG;
wire[15:0] Tile_X3Y4_NN4BEG;
wire[3:0] Tile_X3Y4_E1BEG;
wire[7:0] Tile_X3Y4_E2BEG;
wire[7:0] Tile_X3Y4_E2BEGb;
wire[15:0] Tile_X3Y4_EE4BEG;
wire[11:0] Tile_X3Y4_E6BEG;
wire[3:0] Tile_X3Y4_S1BEG;
wire[7:0] Tile_X3Y4_S2BEG;
wire[7:0] Tile_X3Y4_S2BEGb;
wire[15:0] Tile_X3Y4_S4BEG;
wire[15:0] Tile_X3Y4_SS4BEG;
wire[3:0] Tile_X3Y4_W1BEG;
wire[7:0] Tile_X3Y4_W2BEG;
wire[7:0] Tile_X3Y4_W2BEGb;
wire[15:0] Tile_X3Y4_WW4BEG;
wire[11:0] Tile_X3Y4_W6BEG;
wire[0:0] Tile_X3Y4_Co;
wire[3:0] Tile_X4Y4_N1BEG;
wire[7:0] Tile_X4Y4_N2BEG;
wire[7:0] Tile_X4Y4_N2BEGb;
wire[15:0] Tile_X4Y4_N4BEG;
wire[15:0] Tile_X4Y4_NN4BEG;
wire[3:0] Tile_X4Y4_E1BEG;
wire[7:0] Tile_X4Y4_E2BEG;
wire[7:0] Tile_X4Y4_E2BEGb;
wire[15:0] Tile_X4Y4_EE4BEG;
wire[11:0] Tile_X4Y4_E6BEG;
wire[3:0] Tile_X4Y4_S1BEG;
wire[7:0] Tile_X4Y4_S2BEG;
wire[7:0] Tile_X4Y4_S2BEGb;
wire[15:0] Tile_X4Y4_S4BEG;
wire[15:0] Tile_X4Y4_SS4BEG;
wire[3:0] Tile_X4Y4_W1BEG;
wire[7:0] Tile_X4Y4_W2BEG;
wire[7:0] Tile_X4Y4_W2BEGb;
wire[15:0] Tile_X4Y4_WW4BEG;
wire[11:0] Tile_X4Y4_W6BEG;
wire[0:0] Tile_X4Y4_Co;
wire[3:0] Tile_X5Y4_N1BEG;
wire[7:0] Tile_X5Y4_N2BEG;
wire[7:0] Tile_X5Y4_N2BEGb;
wire[15:0] Tile_X5Y4_N4BEG;
wire[3:0] Tile_X5Y4_S1BEG;
wire[7:0] Tile_X5Y4_S2BEG;
wire[7:0] Tile_X5Y4_S2BEGb;
wire[15:0] Tile_X5Y4_S4BEG;
wire[3:0] Tile_X5Y4_W1BEG;
wire[7:0] Tile_X5Y4_W2BEG;
wire[7:0] Tile_X5Y4_W2BEGb;
wire[15:0] Tile_X5Y4_WW4BEG;
wire[11:0] Tile_X5Y4_W6BEG;
wire[7:0] Tile_X5Y4_bot2top_UIO_OUT;
wire[7:0] Tile_X5Y4_bot2top_UIO_OE;
wire[3:0] Tile_X0Y5_N1BEG;
wire[7:0] Tile_X0Y5_N2BEG;
wire[7:0] Tile_X0Y5_N2BEGb;
wire[15:0] Tile_X0Y5_N4BEG;
wire[3:0] Tile_X0Y5_S1BEG;
wire[7:0] Tile_X0Y5_S2BEG;
wire[7:0] Tile_X0Y5_S2BEGb;
wire[15:0] Tile_X0Y5_S4BEG;
wire[3:0] Tile_X0Y5_E1BEG;
wire[7:0] Tile_X0Y5_E2BEG;
wire[7:0] Tile_X0Y5_E2BEGb;
wire[15:0] Tile_X0Y5_EE4BEG;
wire[11:0] Tile_X0Y5_E6BEG;
wire[3:0] Tile_X1Y5_N1BEG;
wire[7:0] Tile_X1Y5_N2BEG;
wire[7:0] Tile_X1Y5_N2BEGb;
wire[15:0] Tile_X1Y5_N4BEG;
wire[15:0] Tile_X1Y5_NN4BEG;
wire[3:0] Tile_X1Y5_E1BEG;
wire[7:0] Tile_X1Y5_E2BEG;
wire[7:0] Tile_X1Y5_E2BEGb;
wire[15:0] Tile_X1Y5_EE4BEG;
wire[11:0] Tile_X1Y5_E6BEG;
wire[3:0] Tile_X1Y5_S1BEG;
wire[7:0] Tile_X1Y5_S2BEG;
wire[7:0] Tile_X1Y5_S2BEGb;
wire[15:0] Tile_X1Y5_S4BEG;
wire[15:0] Tile_X1Y5_SS4BEG;
wire[3:0] Tile_X1Y5_W1BEG;
wire[7:0] Tile_X1Y5_W2BEG;
wire[7:0] Tile_X1Y5_W2BEGb;
wire[15:0] Tile_X1Y5_WW4BEG;
wire[11:0] Tile_X1Y5_W6BEG;
wire[0:0] Tile_X1Y5_Co;
wire[3:0] Tile_X2Y5_N1BEG;
wire[7:0] Tile_X2Y5_N2BEG;
wire[7:0] Tile_X2Y5_N2BEGb;
wire[15:0] Tile_X2Y5_N4BEG;
wire[15:0] Tile_X2Y5_NN4BEG;
wire[3:0] Tile_X2Y5_E1BEG;
wire[7:0] Tile_X2Y5_E2BEG;
wire[7:0] Tile_X2Y5_E2BEGb;
wire[15:0] Tile_X2Y5_EE4BEG;
wire[11:0] Tile_X2Y5_E6BEG;
wire[3:0] Tile_X2Y5_S1BEG;
wire[7:0] Tile_X2Y5_S2BEG;
wire[7:0] Tile_X2Y5_S2BEGb;
wire[15:0] Tile_X2Y5_S4BEG;
wire[15:0] Tile_X2Y5_SS4BEG;
wire[3:0] Tile_X2Y5_W1BEG;
wire[7:0] Tile_X2Y5_W2BEG;
wire[7:0] Tile_X2Y5_W2BEGb;
wire[15:0] Tile_X2Y5_WW4BEG;
wire[11:0] Tile_X2Y5_W6BEG;
wire[0:0] Tile_X2Y5_Co;
wire[3:0] Tile_X3Y5_N1BEG;
wire[7:0] Tile_X3Y5_N2BEG;
wire[7:0] Tile_X3Y5_N2BEGb;
wire[15:0] Tile_X3Y5_N4BEG;
wire[15:0] Tile_X3Y5_NN4BEG;
wire[3:0] Tile_X3Y5_E1BEG;
wire[7:0] Tile_X3Y5_E2BEG;
wire[7:0] Tile_X3Y5_E2BEGb;
wire[15:0] Tile_X3Y5_EE4BEG;
wire[11:0] Tile_X3Y5_E6BEG;
wire[3:0] Tile_X3Y5_S1BEG;
wire[7:0] Tile_X3Y5_S2BEG;
wire[7:0] Tile_X3Y5_S2BEGb;
wire[15:0] Tile_X3Y5_S4BEG;
wire[15:0] Tile_X3Y5_SS4BEG;
wire[3:0] Tile_X3Y5_W1BEG;
wire[7:0] Tile_X3Y5_W2BEG;
wire[7:0] Tile_X3Y5_W2BEGb;
wire[15:0] Tile_X3Y5_WW4BEG;
wire[11:0] Tile_X3Y5_W6BEG;
wire[0:0] Tile_X3Y5_Co;
wire[3:0] Tile_X4Y5_N1BEG;
wire[7:0] Tile_X4Y5_N2BEG;
wire[7:0] Tile_X4Y5_N2BEGb;
wire[15:0] Tile_X4Y5_N4BEG;
wire[15:0] Tile_X4Y5_NN4BEG;
wire[3:0] Tile_X4Y5_E1BEG;
wire[7:0] Tile_X4Y5_E2BEG;
wire[7:0] Tile_X4Y5_E2BEGb;
wire[15:0] Tile_X4Y5_EE4BEG;
wire[11:0] Tile_X4Y5_E6BEG;
wire[3:0] Tile_X4Y5_S1BEG;
wire[7:0] Tile_X4Y5_S2BEG;
wire[7:0] Tile_X4Y5_S2BEGb;
wire[15:0] Tile_X4Y5_S4BEG;
wire[15:0] Tile_X4Y5_SS4BEG;
wire[3:0] Tile_X4Y5_W1BEG;
wire[7:0] Tile_X4Y5_W2BEG;
wire[7:0] Tile_X4Y5_W2BEGb;
wire[15:0] Tile_X4Y5_WW4BEG;
wire[11:0] Tile_X4Y5_W6BEG;
wire[0:0] Tile_X4Y5_Co;
wire[3:0] Tile_X5Y5_N1BEG;
wire[7:0] Tile_X5Y5_N2BEG;
wire[7:0] Tile_X5Y5_N2BEGb;
wire[15:0] Tile_X5Y5_N4BEG;
wire[3:0] Tile_X5Y5_S1BEG;
wire[7:0] Tile_X5Y5_S2BEG;
wire[7:0] Tile_X5Y5_S2BEGb;
wire[15:0] Tile_X5Y5_S4BEG;
wire[3:0] Tile_X5Y5_W1BEG;
wire[7:0] Tile_X5Y5_W2BEG;
wire[7:0] Tile_X5Y5_W2BEGb;
wire[15:0] Tile_X5Y5_WW4BEG;
wire[11:0] Tile_X5Y5_W6BEG;
wire[3:0] Tile_X0Y6_N1BEG;
wire[7:0] Tile_X0Y6_N2BEG;
wire[7:0] Tile_X0Y6_N2BEGb;
wire[15:0] Tile_X0Y6_N4BEG;
wire[3:0] Tile_X0Y6_S1BEG;
wire[7:0] Tile_X0Y6_S2BEG;
wire[7:0] Tile_X0Y6_S2BEGb;
wire[15:0] Tile_X0Y6_S4BEG;
wire[3:0] Tile_X0Y6_E1BEG;
wire[7:0] Tile_X0Y6_E2BEG;
wire[7:0] Tile_X0Y6_E2BEGb;
wire[15:0] Tile_X0Y6_EE4BEG;
wire[11:0] Tile_X0Y6_E6BEG;
wire[3:0] Tile_X1Y6_N1BEG;
wire[7:0] Tile_X1Y6_N2BEG;
wire[7:0] Tile_X1Y6_N2BEGb;
wire[15:0] Tile_X1Y6_N4BEG;
wire[15:0] Tile_X1Y6_NN4BEG;
wire[3:0] Tile_X1Y6_E1BEG;
wire[7:0] Tile_X1Y6_E2BEG;
wire[7:0] Tile_X1Y6_E2BEGb;
wire[15:0] Tile_X1Y6_EE4BEG;
wire[11:0] Tile_X1Y6_E6BEG;
wire[3:0] Tile_X1Y6_S1BEG;
wire[7:0] Tile_X1Y6_S2BEG;
wire[7:0] Tile_X1Y6_S2BEGb;
wire[15:0] Tile_X1Y6_S4BEG;
wire[15:0] Tile_X1Y6_SS4BEG;
wire[3:0] Tile_X1Y6_W1BEG;
wire[7:0] Tile_X1Y6_W2BEG;
wire[7:0] Tile_X1Y6_W2BEGb;
wire[15:0] Tile_X1Y6_WW4BEG;
wire[11:0] Tile_X1Y6_W6BEG;
wire[0:0] Tile_X1Y6_Co;
wire[3:0] Tile_X2Y6_N1BEG;
wire[7:0] Tile_X2Y6_N2BEG;
wire[7:0] Tile_X2Y6_N2BEGb;
wire[15:0] Tile_X2Y6_N4BEG;
wire[15:0] Tile_X2Y6_NN4BEG;
wire[3:0] Tile_X2Y6_E1BEG;
wire[7:0] Tile_X2Y6_E2BEG;
wire[7:0] Tile_X2Y6_E2BEGb;
wire[15:0] Tile_X2Y6_EE4BEG;
wire[11:0] Tile_X2Y6_E6BEG;
wire[3:0] Tile_X2Y6_S1BEG;
wire[7:0] Tile_X2Y6_S2BEG;
wire[7:0] Tile_X2Y6_S2BEGb;
wire[15:0] Tile_X2Y6_S4BEG;
wire[15:0] Tile_X2Y6_SS4BEG;
wire[3:0] Tile_X2Y6_W1BEG;
wire[7:0] Tile_X2Y6_W2BEG;
wire[7:0] Tile_X2Y6_W2BEGb;
wire[15:0] Tile_X2Y6_WW4BEG;
wire[11:0] Tile_X2Y6_W6BEG;
wire[0:0] Tile_X2Y6_Co;
wire[3:0] Tile_X3Y6_N1BEG;
wire[7:0] Tile_X3Y6_N2BEG;
wire[7:0] Tile_X3Y6_N2BEGb;
wire[15:0] Tile_X3Y6_N4BEG;
wire[15:0] Tile_X3Y6_NN4BEG;
wire[3:0] Tile_X3Y6_E1BEG;
wire[7:0] Tile_X3Y6_E2BEG;
wire[7:0] Tile_X3Y6_E2BEGb;
wire[15:0] Tile_X3Y6_EE4BEG;
wire[11:0] Tile_X3Y6_E6BEG;
wire[3:0] Tile_X3Y6_S1BEG;
wire[7:0] Tile_X3Y6_S2BEG;
wire[7:0] Tile_X3Y6_S2BEGb;
wire[15:0] Tile_X3Y6_S4BEG;
wire[15:0] Tile_X3Y6_SS4BEG;
wire[3:0] Tile_X3Y6_W1BEG;
wire[7:0] Tile_X3Y6_W2BEG;
wire[7:0] Tile_X3Y6_W2BEGb;
wire[15:0] Tile_X3Y6_WW4BEG;
wire[11:0] Tile_X3Y6_W6BEG;
wire[0:0] Tile_X3Y6_Co;
wire[3:0] Tile_X4Y6_N1BEG;
wire[7:0] Tile_X4Y6_N2BEG;
wire[7:0] Tile_X4Y6_N2BEGb;
wire[15:0] Tile_X4Y6_N4BEG;
wire[15:0] Tile_X4Y6_NN4BEG;
wire[3:0] Tile_X4Y6_E1BEG;
wire[7:0] Tile_X4Y6_E2BEG;
wire[7:0] Tile_X4Y6_E2BEGb;
wire[15:0] Tile_X4Y6_EE4BEG;
wire[11:0] Tile_X4Y6_E6BEG;
wire[3:0] Tile_X4Y6_S1BEG;
wire[7:0] Tile_X4Y6_S2BEG;
wire[7:0] Tile_X4Y6_S2BEGb;
wire[15:0] Tile_X4Y6_S4BEG;
wire[15:0] Tile_X4Y6_SS4BEG;
wire[3:0] Tile_X4Y6_W1BEG;
wire[7:0] Tile_X4Y6_W2BEG;
wire[7:0] Tile_X4Y6_W2BEGb;
wire[15:0] Tile_X4Y6_WW4BEG;
wire[11:0] Tile_X4Y6_W6BEG;
wire[0:0] Tile_X4Y6_Co;
wire[3:0] Tile_X5Y6_N1BEG;
wire[7:0] Tile_X5Y6_N2BEG;
wire[7:0] Tile_X5Y6_N2BEGb;
wire[15:0] Tile_X5Y6_N4BEG;
wire[3:0] Tile_X5Y6_S1BEG;
wire[7:0] Tile_X5Y6_S2BEG;
wire[7:0] Tile_X5Y6_S2BEGb;
wire[15:0] Tile_X5Y6_S4BEG;
wire[3:0] Tile_X5Y6_W1BEG;
wire[7:0] Tile_X5Y6_W2BEG;
wire[7:0] Tile_X5Y6_W2BEGb;
wire[15:0] Tile_X5Y6_WW4BEG;
wire[11:0] Tile_X5Y6_W6BEG;
wire[3:0] Tile_X0Y7_N1BEG;
wire[7:0] Tile_X0Y7_N2BEG;
wire[7:0] Tile_X0Y7_N2BEGb;
wire[15:0] Tile_X0Y7_N4BEG;
wire[3:0] Tile_X0Y7_S1BEG;
wire[7:0] Tile_X0Y7_S2BEG;
wire[7:0] Tile_X0Y7_S2BEGb;
wire[15:0] Tile_X0Y7_S4BEG;
wire[3:0] Tile_X0Y7_E1BEG;
wire[7:0] Tile_X0Y7_E2BEG;
wire[7:0] Tile_X0Y7_E2BEGb;
wire[15:0] Tile_X0Y7_EE4BEG;
wire[11:0] Tile_X0Y7_E6BEG;
wire[3:0] Tile_X1Y7_N1BEG;
wire[7:0] Tile_X1Y7_N2BEG;
wire[7:0] Tile_X1Y7_N2BEGb;
wire[15:0] Tile_X1Y7_N4BEG;
wire[15:0] Tile_X1Y7_NN4BEG;
wire[3:0] Tile_X1Y7_E1BEG;
wire[7:0] Tile_X1Y7_E2BEG;
wire[7:0] Tile_X1Y7_E2BEGb;
wire[15:0] Tile_X1Y7_EE4BEG;
wire[11:0] Tile_X1Y7_E6BEG;
wire[3:0] Tile_X1Y7_S1BEG;
wire[7:0] Tile_X1Y7_S2BEG;
wire[7:0] Tile_X1Y7_S2BEGb;
wire[15:0] Tile_X1Y7_S4BEG;
wire[15:0] Tile_X1Y7_SS4BEG;
wire[3:0] Tile_X1Y7_W1BEG;
wire[7:0] Tile_X1Y7_W2BEG;
wire[7:0] Tile_X1Y7_W2BEGb;
wire[15:0] Tile_X1Y7_WW4BEG;
wire[11:0] Tile_X1Y7_W6BEG;
wire[0:0] Tile_X1Y7_Co;
wire[3:0] Tile_X2Y7_N1BEG;
wire[7:0] Tile_X2Y7_N2BEG;
wire[7:0] Tile_X2Y7_N2BEGb;
wire[15:0] Tile_X2Y7_N4BEG;
wire[15:0] Tile_X2Y7_NN4BEG;
wire[3:0] Tile_X2Y7_E1BEG;
wire[7:0] Tile_X2Y7_E2BEG;
wire[7:0] Tile_X2Y7_E2BEGb;
wire[15:0] Tile_X2Y7_EE4BEG;
wire[11:0] Tile_X2Y7_E6BEG;
wire[3:0] Tile_X2Y7_S1BEG;
wire[7:0] Tile_X2Y7_S2BEG;
wire[7:0] Tile_X2Y7_S2BEGb;
wire[15:0] Tile_X2Y7_S4BEG;
wire[15:0] Tile_X2Y7_SS4BEG;
wire[3:0] Tile_X2Y7_W1BEG;
wire[7:0] Tile_X2Y7_W2BEG;
wire[7:0] Tile_X2Y7_W2BEGb;
wire[15:0] Tile_X2Y7_WW4BEG;
wire[11:0] Tile_X2Y7_W6BEG;
wire[0:0] Tile_X2Y7_Co;
wire[3:0] Tile_X3Y7_N1BEG;
wire[7:0] Tile_X3Y7_N2BEG;
wire[7:0] Tile_X3Y7_N2BEGb;
wire[15:0] Tile_X3Y7_N4BEG;
wire[15:0] Tile_X3Y7_NN4BEG;
wire[3:0] Tile_X3Y7_E1BEG;
wire[7:0] Tile_X3Y7_E2BEG;
wire[7:0] Tile_X3Y7_E2BEGb;
wire[15:0] Tile_X3Y7_EE4BEG;
wire[11:0] Tile_X3Y7_E6BEG;
wire[3:0] Tile_X3Y7_S1BEG;
wire[7:0] Tile_X3Y7_S2BEG;
wire[7:0] Tile_X3Y7_S2BEGb;
wire[15:0] Tile_X3Y7_S4BEG;
wire[15:0] Tile_X3Y7_SS4BEG;
wire[3:0] Tile_X3Y7_W1BEG;
wire[7:0] Tile_X3Y7_W2BEG;
wire[7:0] Tile_X3Y7_W2BEGb;
wire[15:0] Tile_X3Y7_WW4BEG;
wire[11:0] Tile_X3Y7_W6BEG;
wire[0:0] Tile_X3Y7_Co;
wire[3:0] Tile_X4Y7_N1BEG;
wire[7:0] Tile_X4Y7_N2BEG;
wire[7:0] Tile_X4Y7_N2BEGb;
wire[15:0] Tile_X4Y7_N4BEG;
wire[15:0] Tile_X4Y7_NN4BEG;
wire[3:0] Tile_X4Y7_E1BEG;
wire[7:0] Tile_X4Y7_E2BEG;
wire[7:0] Tile_X4Y7_E2BEGb;
wire[15:0] Tile_X4Y7_EE4BEG;
wire[11:0] Tile_X4Y7_E6BEG;
wire[3:0] Tile_X4Y7_S1BEG;
wire[7:0] Tile_X4Y7_S2BEG;
wire[7:0] Tile_X4Y7_S2BEGb;
wire[15:0] Tile_X4Y7_S4BEG;
wire[15:0] Tile_X4Y7_SS4BEG;
wire[3:0] Tile_X4Y7_W1BEG;
wire[7:0] Tile_X4Y7_W2BEG;
wire[7:0] Tile_X4Y7_W2BEGb;
wire[15:0] Tile_X4Y7_WW4BEG;
wire[11:0] Tile_X4Y7_W6BEG;
wire[0:0] Tile_X4Y7_Co;
wire[3:0] Tile_X5Y7_N1BEG;
wire[7:0] Tile_X5Y7_N2BEG;
wire[7:0] Tile_X5Y7_N2BEGb;
wire[15:0] Tile_X5Y7_N4BEG;
wire[3:0] Tile_X5Y7_S1BEG;
wire[7:0] Tile_X5Y7_S2BEG;
wire[7:0] Tile_X5Y7_S2BEGb;
wire[15:0] Tile_X5Y7_S4BEG;
wire[3:0] Tile_X5Y7_W1BEG;
wire[7:0] Tile_X5Y7_W2BEG;
wire[7:0] Tile_X5Y7_W2BEGb;
wire[15:0] Tile_X5Y7_WW4BEG;
wire[11:0] Tile_X5Y7_W6BEG;
wire[3:0] Tile_X0Y8_N1BEG;
wire[7:0] Tile_X0Y8_N2BEG;
wire[7:0] Tile_X0Y8_N2BEGb;
wire[15:0] Tile_X0Y8_N4BEG;
wire[3:0] Tile_X0Y8_S1BEG;
wire[7:0] Tile_X0Y8_S2BEG;
wire[7:0] Tile_X0Y8_S2BEGb;
wire[15:0] Tile_X0Y8_S4BEG;
wire[3:0] Tile_X0Y8_E1BEG;
wire[7:0] Tile_X0Y8_E2BEG;
wire[7:0] Tile_X0Y8_E2BEGb;
wire[15:0] Tile_X0Y8_EE4BEG;
wire[11:0] Tile_X0Y8_E6BEG;
wire[3:0] Tile_X1Y8_N1BEG;
wire[7:0] Tile_X1Y8_N2BEG;
wire[7:0] Tile_X1Y8_N2BEGb;
wire[15:0] Tile_X1Y8_N4BEG;
wire[15:0] Tile_X1Y8_NN4BEG;
wire[3:0] Tile_X1Y8_E1BEG;
wire[7:0] Tile_X1Y8_E2BEG;
wire[7:0] Tile_X1Y8_E2BEGb;
wire[15:0] Tile_X1Y8_EE4BEG;
wire[11:0] Tile_X1Y8_E6BEG;
wire[3:0] Tile_X1Y8_S1BEG;
wire[7:0] Tile_X1Y8_S2BEG;
wire[7:0] Tile_X1Y8_S2BEGb;
wire[15:0] Tile_X1Y8_S4BEG;
wire[15:0] Tile_X1Y8_SS4BEG;
wire[3:0] Tile_X1Y8_W1BEG;
wire[7:0] Tile_X1Y8_W2BEG;
wire[7:0] Tile_X1Y8_W2BEGb;
wire[15:0] Tile_X1Y8_WW4BEG;
wire[11:0] Tile_X1Y8_W6BEG;
wire[0:0] Tile_X1Y8_Co;
wire[3:0] Tile_X2Y8_N1BEG;
wire[7:0] Tile_X2Y8_N2BEG;
wire[7:0] Tile_X2Y8_N2BEGb;
wire[15:0] Tile_X2Y8_N4BEG;
wire[15:0] Tile_X2Y8_NN4BEG;
wire[3:0] Tile_X2Y8_E1BEG;
wire[7:0] Tile_X2Y8_E2BEG;
wire[7:0] Tile_X2Y8_E2BEGb;
wire[15:0] Tile_X2Y8_EE4BEG;
wire[11:0] Tile_X2Y8_E6BEG;
wire[3:0] Tile_X2Y8_S1BEG;
wire[7:0] Tile_X2Y8_S2BEG;
wire[7:0] Tile_X2Y8_S2BEGb;
wire[15:0] Tile_X2Y8_S4BEG;
wire[15:0] Tile_X2Y8_SS4BEG;
wire[3:0] Tile_X2Y8_W1BEG;
wire[7:0] Tile_X2Y8_W2BEG;
wire[7:0] Tile_X2Y8_W2BEGb;
wire[15:0] Tile_X2Y8_WW4BEG;
wire[11:0] Tile_X2Y8_W6BEG;
wire[0:0] Tile_X2Y8_Co;
wire[3:0] Tile_X3Y8_N1BEG;
wire[7:0] Tile_X3Y8_N2BEG;
wire[7:0] Tile_X3Y8_N2BEGb;
wire[15:0] Tile_X3Y8_N4BEG;
wire[15:0] Tile_X3Y8_NN4BEG;
wire[3:0] Tile_X3Y8_E1BEG;
wire[7:0] Tile_X3Y8_E2BEG;
wire[7:0] Tile_X3Y8_E2BEGb;
wire[15:0] Tile_X3Y8_EE4BEG;
wire[11:0] Tile_X3Y8_E6BEG;
wire[3:0] Tile_X3Y8_S1BEG;
wire[7:0] Tile_X3Y8_S2BEG;
wire[7:0] Tile_X3Y8_S2BEGb;
wire[15:0] Tile_X3Y8_S4BEG;
wire[15:0] Tile_X3Y8_SS4BEG;
wire[3:0] Tile_X3Y8_W1BEG;
wire[7:0] Tile_X3Y8_W2BEG;
wire[7:0] Tile_X3Y8_W2BEGb;
wire[15:0] Tile_X3Y8_WW4BEG;
wire[11:0] Tile_X3Y8_W6BEG;
wire[0:0] Tile_X3Y8_Co;
wire[3:0] Tile_X4Y8_N1BEG;
wire[7:0] Tile_X4Y8_N2BEG;
wire[7:0] Tile_X4Y8_N2BEGb;
wire[15:0] Tile_X4Y8_N4BEG;
wire[15:0] Tile_X4Y8_NN4BEG;
wire[3:0] Tile_X4Y8_E1BEG;
wire[7:0] Tile_X4Y8_E2BEG;
wire[7:0] Tile_X4Y8_E2BEGb;
wire[15:0] Tile_X4Y8_EE4BEG;
wire[11:0] Tile_X4Y8_E6BEG;
wire[3:0] Tile_X4Y8_S1BEG;
wire[7:0] Tile_X4Y8_S2BEG;
wire[7:0] Tile_X4Y8_S2BEGb;
wire[15:0] Tile_X4Y8_S4BEG;
wire[15:0] Tile_X4Y8_SS4BEG;
wire[3:0] Tile_X4Y8_W1BEG;
wire[7:0] Tile_X4Y8_W2BEG;
wire[7:0] Tile_X4Y8_W2BEGb;
wire[15:0] Tile_X4Y8_WW4BEG;
wire[11:0] Tile_X4Y8_W6BEG;
wire[0:0] Tile_X4Y8_Co;
wire[3:0] Tile_X5Y8_N1BEG;
wire[7:0] Tile_X5Y8_N2BEG;
wire[7:0] Tile_X5Y8_N2BEGb;
wire[15:0] Tile_X5Y8_N4BEG;
wire[3:0] Tile_X5Y8_S1BEG;
wire[7:0] Tile_X5Y8_S2BEG;
wire[7:0] Tile_X5Y8_S2BEGb;
wire[15:0] Tile_X5Y8_S4BEG;
wire[3:0] Tile_X5Y8_W1BEG;
wire[7:0] Tile_X5Y8_W2BEG;
wire[7:0] Tile_X5Y8_W2BEGb;
wire[15:0] Tile_X5Y8_WW4BEG;
wire[11:0] Tile_X5Y8_W6BEG;
wire[3:0] Tile_X0Y9_N1BEG;
wire[7:0] Tile_X0Y9_N2BEG;
wire[7:0] Tile_X0Y9_N2BEGb;
wire[15:0] Tile_X0Y9_N4BEG;
wire[3:0] Tile_X1Y9_N1BEG;
wire[7:0] Tile_X1Y9_N2BEG;
wire[7:0] Tile_X1Y9_N2BEGb;
wire[15:0] Tile_X1Y9_N4BEG;
wire[15:0] Tile_X1Y9_NN4BEG;
wire[0:0] Tile_X1Y9_Co;
wire[3:0] Tile_X2Y9_N1BEG;
wire[7:0] Tile_X2Y9_N2BEG;
wire[7:0] Tile_X2Y9_N2BEGb;
wire[15:0] Tile_X2Y9_N4BEG;
wire[15:0] Tile_X2Y9_NN4BEG;
wire[0:0] Tile_X2Y9_Co;
wire[3:0] Tile_X3Y9_N1BEG;
wire[7:0] Tile_X3Y9_N2BEG;
wire[7:0] Tile_X3Y9_N2BEGb;
wire[15:0] Tile_X3Y9_N4BEG;
wire[15:0] Tile_X3Y9_NN4BEG;
wire[0:0] Tile_X3Y9_Co;
wire[3:0] Tile_X4Y9_N1BEG;
wire[7:0] Tile_X4Y9_N2BEG;
wire[7:0] Tile_X4Y9_N2BEGb;
wire[15:0] Tile_X4Y9_N4BEG;
wire[15:0] Tile_X4Y9_NN4BEG;
wire[0:0] Tile_X4Y9_Co;
wire[3:0] Tile_X5Y9_N1BEG;
wire[7:0] Tile_X5Y9_N2BEG;
wire[7:0] Tile_X5Y9_N2BEGb;
wire[15:0] Tile_X5Y9_N4BEG;

assign Row_Y0_FrameData = FrameData[FrameBitsPerRow*(0+1)-1:FrameBitsPerRow*0];
assign Row_Y1_FrameData = FrameData[FrameBitsPerRow*(1+1)-1:FrameBitsPerRow*1];
assign Row_Y2_FrameData = FrameData[FrameBitsPerRow*(2+1)-1:FrameBitsPerRow*2];
assign Row_Y3_FrameData = FrameData[FrameBitsPerRow*(3+1)-1:FrameBitsPerRow*3];
assign Row_Y4_FrameData = FrameData[FrameBitsPerRow*(4+1)-1:FrameBitsPerRow*4];
assign Row_Y5_FrameData = FrameData[FrameBitsPerRow*(5+1)-1:FrameBitsPerRow*5];
assign Row_Y6_FrameData = FrameData[FrameBitsPerRow*(6+1)-1:FrameBitsPerRow*6];
assign Row_Y7_FrameData = FrameData[FrameBitsPerRow*(7+1)-1:FrameBitsPerRow*7];
assign Row_Y8_FrameData = FrameData[FrameBitsPerRow*(8+1)-1:FrameBitsPerRow*8];
assign Row_Y9_FrameData = FrameData[FrameBitsPerRow*(9+1)-1:FrameBitsPerRow*9];
assign Column_X0_FrameStrobe = FrameStrobe[MaxFramesPerCol*(0+1)-1:MaxFramesPerCol*0];
assign Column_X1_FrameStrobe = FrameStrobe[MaxFramesPerCol*(1+1)-1:MaxFramesPerCol*1];
assign Column_X2_FrameStrobe = FrameStrobe[MaxFramesPerCol*(2+1)-1:MaxFramesPerCol*2];
assign Column_X3_FrameStrobe = FrameStrobe[MaxFramesPerCol*(3+1)-1:MaxFramesPerCol*3];
assign Column_X4_FrameStrobe = FrameStrobe[MaxFramesPerCol*(4+1)-1:MaxFramesPerCol*4];
assign Column_X5_FrameStrobe = FrameStrobe[MaxFramesPerCol*(5+1)-1:MaxFramesPerCol*5];

 //tile IO port will get directly connected to top-level tile module
NW_term Tile_X0Y0_NW_term (
    .N1END(Tile_X0Y1_N1BEG),
    .N2MID(Tile_X0Y1_N2BEG),
    .N2END(Tile_X0Y1_N2BEGb),
    .N4END(Tile_X0Y1_N4BEG),
    .S1BEG(Tile_X0Y0_S1BEG),
    .S2BEG(Tile_X0Y0_S2BEG),
    .S2BEGb(Tile_X0Y0_S2BEGb),
    .S4BEG(Tile_X0Y0_S4BEG),
    .UserCLK(Tile_X0Y1_UserCLKo),
    .UserCLKo(Tile_X0Y0_UserCLKo),
    .FrameData(Row_Y0_FrameData),
    .FrameData_O(Tile_X0Y0_FrameData_O),
    .FrameStrobe(Tile_X0Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
N_IO4 Tile_X1Y0_N_IO4 (
    .N1END(Tile_X1Y1_N1BEG),
    .N2MID(Tile_X1Y1_N2BEG),
    .N2END(Tile_X1Y1_N2BEGb),
    .N4END(Tile_X1Y1_N4BEG),
    .NN4END(Tile_X1Y1_NN4BEG),
    .Ci(Tile_X1Y1_Co),
    .S1BEG(Tile_X1Y0_S1BEG),
    .S2BEG(Tile_X1Y0_S2BEG),
    .S2BEGb(Tile_X1Y0_S2BEGb),
    .S4BEG(Tile_X1Y0_S4BEG),
    .SS4BEG(Tile_X1Y0_SS4BEG),
    .A_O_top(Tile_X1Y0_A_O_top),
    .A_I_top(Tile_X1Y0_A_I_top),
    .A_T_top(Tile_X1Y0_A_T_top),
    .B_O_top(Tile_X1Y0_B_O_top),
    .B_I_top(Tile_X1Y0_B_I_top),
    .B_T_top(Tile_X1Y0_B_T_top),
    .C_O_top(Tile_X1Y0_C_O_top),
    .C_I_top(Tile_X1Y0_C_I_top),
    .C_T_top(Tile_X1Y0_C_T_top),
    .D_O_top(Tile_X1Y0_D_O_top),
    .D_I_top(Tile_X1Y0_D_I_top),
    .D_T_top(Tile_X1Y0_D_T_top),
    .UserCLK(Tile_X1Y1_UserCLKo),
    .UserCLKo(Tile_X1Y0_UserCLKo),
    .FrameData(Tile_X0Y0_FrameData_O),
    .FrameData_O(Tile_X1Y0_FrameData_O),
    .FrameStrobe(Tile_X1Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
N_IO4 Tile_X2Y0_N_IO4 (
    .N1END(Tile_X2Y1_N1BEG),
    .N2MID(Tile_X2Y1_N2BEG),
    .N2END(Tile_X2Y1_N2BEGb),
    .N4END(Tile_X2Y1_N4BEG),
    .NN4END(Tile_X2Y1_NN4BEG),
    .Ci(Tile_X2Y1_Co),
    .S1BEG(Tile_X2Y0_S1BEG),
    .S2BEG(Tile_X2Y0_S2BEG),
    .S2BEGb(Tile_X2Y0_S2BEGb),
    .S4BEG(Tile_X2Y0_S4BEG),
    .SS4BEG(Tile_X2Y0_SS4BEG),
    .A_O_top(Tile_X2Y0_A_O_top),
    .A_I_top(Tile_X2Y0_A_I_top),
    .A_T_top(Tile_X2Y0_A_T_top),
    .B_O_top(Tile_X2Y0_B_O_top),
    .B_I_top(Tile_X2Y0_B_I_top),
    .B_T_top(Tile_X2Y0_B_T_top),
    .C_O_top(Tile_X2Y0_C_O_top),
    .C_I_top(Tile_X2Y0_C_I_top),
    .C_T_top(Tile_X2Y0_C_T_top),
    .D_O_top(Tile_X2Y0_D_O_top),
    .D_I_top(Tile_X2Y0_D_I_top),
    .D_T_top(Tile_X2Y0_D_T_top),
    .UserCLK(Tile_X2Y1_UserCLKo),
    .UserCLKo(Tile_X2Y0_UserCLKo),
    .FrameData(Tile_X1Y0_FrameData_O),
    .FrameData_O(Tile_X2Y0_FrameData_O),
    .FrameStrobe(Tile_X2Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
N_IO4 Tile_X3Y0_N_IO4 (
    .N1END(Tile_X3Y1_N1BEG),
    .N2MID(Tile_X3Y1_N2BEG),
    .N2END(Tile_X3Y1_N2BEGb),
    .N4END(Tile_X3Y1_N4BEG),
    .NN4END(Tile_X3Y1_NN4BEG),
    .Ci(Tile_X3Y1_Co),
    .S1BEG(Tile_X3Y0_S1BEG),
    .S2BEG(Tile_X3Y0_S2BEG),
    .S2BEGb(Tile_X3Y0_S2BEGb),
    .S4BEG(Tile_X3Y0_S4BEG),
    .SS4BEG(Tile_X3Y0_SS4BEG),
    .A_O_top(Tile_X3Y0_A_O_top),
    .A_I_top(Tile_X3Y0_A_I_top),
    .A_T_top(Tile_X3Y0_A_T_top),
    .B_O_top(Tile_X3Y0_B_O_top),
    .B_I_top(Tile_X3Y0_B_I_top),
    .B_T_top(Tile_X3Y0_B_T_top),
    .C_O_top(Tile_X3Y0_C_O_top),
    .C_I_top(Tile_X3Y0_C_I_top),
    .C_T_top(Tile_X3Y0_C_T_top),
    .D_O_top(Tile_X3Y0_D_O_top),
    .D_I_top(Tile_X3Y0_D_I_top),
    .D_T_top(Tile_X3Y0_D_T_top),
    .UserCLK(Tile_X3Y1_UserCLKo),
    .UserCLKo(Tile_X3Y0_UserCLKo),
    .FrameData(Tile_X2Y0_FrameData_O),
    .FrameData_O(Tile_X3Y0_FrameData_O),
    .FrameStrobe(Tile_X3Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
N_IO4 Tile_X4Y0_N_IO4 (
    .N1END(Tile_X4Y1_N1BEG),
    .N2MID(Tile_X4Y1_N2BEG),
    .N2END(Tile_X4Y1_N2BEGb),
    .N4END(Tile_X4Y1_N4BEG),
    .NN4END(Tile_X4Y1_NN4BEG),
    .Ci(Tile_X4Y1_Co),
    .S1BEG(Tile_X4Y0_S1BEG),
    .S2BEG(Tile_X4Y0_S2BEG),
    .S2BEGb(Tile_X4Y0_S2BEGb),
    .S4BEG(Tile_X4Y0_S4BEG),
    .SS4BEG(Tile_X4Y0_SS4BEG),
    .A_O_top(Tile_X4Y0_A_O_top),
    .A_I_top(Tile_X4Y0_A_I_top),
    .A_T_top(Tile_X4Y0_A_T_top),
    .B_O_top(Tile_X4Y0_B_O_top),
    .B_I_top(Tile_X4Y0_B_I_top),
    .B_T_top(Tile_X4Y0_B_T_top),
    .C_O_top(Tile_X4Y0_C_O_top),
    .C_I_top(Tile_X4Y0_C_I_top),
    .C_T_top(Tile_X4Y0_C_T_top),
    .D_O_top(Tile_X4Y0_D_O_top),
    .D_I_top(Tile_X4Y0_D_I_top),
    .D_T_top(Tile_X4Y0_D_T_top),
    .UserCLK(Tile_X4Y1_UserCLKo),
    .UserCLKo(Tile_X4Y0_UserCLKo),
    .FrameData(Tile_X3Y0_FrameData_O),
    .FrameData_O(Tile_X4Y0_FrameData_O),
    .FrameStrobe(Tile_X4Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
NE_term Tile_X5Y0_NE_term (
    .N1END(Tile_X5Y1_N1BEG),
    .N2MID(Tile_X5Y1_N2BEG),
    .N2END(Tile_X5Y1_N2BEGb),
    .N4END(Tile_X5Y1_N4BEG),
    .S1BEG(Tile_X5Y0_S1BEG),
    .S2BEG(Tile_X5Y0_S2BEG),
    .S2BEGb(Tile_X5Y0_S2BEGb),
    .S4BEG(Tile_X5Y0_S4BEG),
    .UserCLK(Tile_X5Y1_UserCLKo),
    .UserCLKo(Tile_X5Y0_UserCLKo),
    .FrameData(Tile_X4Y0_FrameData_O),
    .FrameData_O(Tile_X5Y0_FrameData_O),
    .FrameStrobe(Tile_X5Y1_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y0_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_TT_IF2
`ifdef EMULATION
    #(
    .Tile_X0Y0_Emulate_Bitstream(`Tile_X0Y1_Emulate_Bitstream),
    .Tile_X0Y1_Emulate_Bitstream(`Tile_X0Y2_Emulate_Bitstream)
    )
`endif
    Tile_X0Y1_W_TT_IF2
    (
    .Tile_X0Y0_S1END(Tile_X0Y0_S1BEG),
    .Tile_X0Y0_S2MID(Tile_X0Y0_S2BEG),
    .Tile_X0Y0_S2END(Tile_X0Y0_S2BEGb),
    .Tile_X0Y0_S4END(Tile_X0Y0_S4BEG),
    .Tile_X0Y0_W1END(Tile_X1Y1_W1BEG),
    .Tile_X0Y0_W2MID(Tile_X1Y1_W2BEG),
    .Tile_X0Y0_W2END(Tile_X1Y1_W2BEGb),
    .Tile_X0Y0_WW4END(Tile_X1Y1_WW4BEG),
    .Tile_X0Y0_W6END(Tile_X1Y1_W6BEG),
    .Tile_X0Y1_N1END(Tile_X0Y3_N1BEG),
    .Tile_X0Y1_N2MID(Tile_X0Y3_N2BEG),
    .Tile_X0Y1_N2END(Tile_X0Y3_N2BEGb),
    .Tile_X0Y1_N4END(Tile_X0Y3_N4BEG),
    .Tile_X0Y1_W1END(Tile_X1Y2_W1BEG),
    .Tile_X0Y1_W2MID(Tile_X1Y2_W2BEG),
    .Tile_X0Y1_W2END(Tile_X1Y2_W2BEGb),
    .Tile_X0Y1_WW4END(Tile_X1Y2_WW4BEG),
    .Tile_X0Y1_W6END(Tile_X1Y2_W6BEG),
    .Tile_X0Y0_N1BEG(Tile_X0Y1_N1BEG),
    .Tile_X0Y0_N2BEG(Tile_X0Y1_N2BEG),
    .Tile_X0Y0_N2BEGb(Tile_X0Y1_N2BEGb),
    .Tile_X0Y0_N4BEG(Tile_X0Y1_N4BEG),
    .Tile_X0Y0_E1BEG(Tile_X0Y1_E1BEG),
    .Tile_X0Y0_E2BEG(Tile_X0Y1_E2BEG),
    .Tile_X0Y0_E2BEGb(Tile_X0Y1_E2BEGb),
    .Tile_X0Y0_EE4BEG(Tile_X0Y1_EE4BEG),
    .Tile_X0Y0_E6BEG(Tile_X0Y1_E6BEG),
    .Tile_X0Y1_E1BEG(Tile_X0Y2_E1BEG),
    .Tile_X0Y1_E2BEG(Tile_X0Y2_E2BEG),
    .Tile_X0Y1_E2BEGb(Tile_X0Y2_E2BEGb),
    .Tile_X0Y1_EE4BEG(Tile_X0Y2_EE4BEG),
    .Tile_X0Y1_E6BEG(Tile_X0Y2_E6BEG),
    .Tile_X0Y1_S1BEG(Tile_X0Y2_S1BEG),
    .Tile_X0Y1_S2BEG(Tile_X0Y2_S2BEG),
    .Tile_X0Y1_S2BEGb(Tile_X0Y2_S2BEGb),
    .Tile_X0Y1_S4BEG(Tile_X0Y2_S4BEG),
    .UO_OUT_TT_PROJECT0(Tile_X0Y2_UO_OUT_TT_PROJECT0),
    .UO_OUT_TT_PROJECT1(Tile_X0Y2_UO_OUT_TT_PROJECT1),
    .UO_OUT_TT_PROJECT2(Tile_X0Y2_UO_OUT_TT_PROJECT2),
    .UO_OUT_TT_PROJECT3(Tile_X0Y2_UO_OUT_TT_PROJECT3),
    .UO_OUT_TT_PROJECT4(Tile_X0Y2_UO_OUT_TT_PROJECT4),
    .UO_OUT_TT_PROJECT5(Tile_X0Y2_UO_OUT_TT_PROJECT5),
    .UO_OUT_TT_PROJECT6(Tile_X0Y2_UO_OUT_TT_PROJECT6),
    .UO_OUT_TT_PROJECT7(Tile_X0Y2_UO_OUT_TT_PROJECT7),
    .UIO_OUT_TT_PROJECT0(Tile_X0Y2_UIO_OUT_TT_PROJECT0),
    .UIO_OUT_TT_PROJECT1(Tile_X0Y2_UIO_OUT_TT_PROJECT1),
    .UIO_OUT_TT_PROJECT2(Tile_X0Y2_UIO_OUT_TT_PROJECT2),
    .UIO_OUT_TT_PROJECT3(Tile_X0Y2_UIO_OUT_TT_PROJECT3),
    .UIO_OUT_TT_PROJECT4(Tile_X0Y2_UIO_OUT_TT_PROJECT4),
    .UIO_OUT_TT_PROJECT5(Tile_X0Y2_UIO_OUT_TT_PROJECT5),
    .UIO_OUT_TT_PROJECT6(Tile_X0Y2_UIO_OUT_TT_PROJECT6),
    .UIO_OUT_TT_PROJECT7(Tile_X0Y2_UIO_OUT_TT_PROJECT7),
    .UIO_OE_TT_PROJECT0(Tile_X0Y2_UIO_OE_TT_PROJECT0),
    .UIO_OE_TT_PROJECT1(Tile_X0Y2_UIO_OE_TT_PROJECT1),
    .UIO_OE_TT_PROJECT2(Tile_X0Y2_UIO_OE_TT_PROJECT2),
    .UIO_OE_TT_PROJECT3(Tile_X0Y2_UIO_OE_TT_PROJECT3),
    .UIO_OE_TT_PROJECT4(Tile_X0Y2_UIO_OE_TT_PROJECT4),
    .UIO_OE_TT_PROJECT5(Tile_X0Y2_UIO_OE_TT_PROJECT5),
    .UIO_OE_TT_PROJECT6(Tile_X0Y2_UIO_OE_TT_PROJECT6),
    .UIO_OE_TT_PROJECT7(Tile_X0Y2_UIO_OE_TT_PROJECT7),
    .UI_IN_TT_PROJECT0(Tile_X0Y2_UI_IN_TT_PROJECT0),
    .UI_IN_TT_PROJECT1(Tile_X0Y2_UI_IN_TT_PROJECT1),
    .UI_IN_TT_PROJECT2(Tile_X0Y2_UI_IN_TT_PROJECT2),
    .UI_IN_TT_PROJECT3(Tile_X0Y2_UI_IN_TT_PROJECT3),
    .UI_IN_TT_PROJECT4(Tile_X0Y2_UI_IN_TT_PROJECT4),
    .UI_IN_TT_PROJECT5(Tile_X0Y2_UI_IN_TT_PROJECT5),
    .UI_IN_TT_PROJECT6(Tile_X0Y2_UI_IN_TT_PROJECT6),
    .UI_IN_TT_PROJECT7(Tile_X0Y2_UI_IN_TT_PROJECT7),
    .UIO_IN_TT_PROJECT0(Tile_X0Y2_UIO_IN_TT_PROJECT0),
    .UIO_IN_TT_PROJECT1(Tile_X0Y2_UIO_IN_TT_PROJECT1),
    .UIO_IN_TT_PROJECT2(Tile_X0Y2_UIO_IN_TT_PROJECT2),
    .UIO_IN_TT_PROJECT3(Tile_X0Y2_UIO_IN_TT_PROJECT3),
    .UIO_IN_TT_PROJECT4(Tile_X0Y2_UIO_IN_TT_PROJECT4),
    .UIO_IN_TT_PROJECT5(Tile_X0Y2_UIO_IN_TT_PROJECT5),
    .UIO_IN_TT_PROJECT6(Tile_X0Y2_UIO_IN_TT_PROJECT6),
    .UIO_IN_TT_PROJECT7(Tile_X0Y2_UIO_IN_TT_PROJECT7),
    .ENA_TT_PROJECT(Tile_X0Y2_ENA_TT_PROJECT),
    .CLK_TT_PROJECT(Tile_X0Y2_CLK_TT_PROJECT),
    .RST_N_TT_PROJECT(Tile_X0Y2_RST_N_TT_PROJECT),
    .Tile_X0Y0_UserCLKo(Tile_X0Y1_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X0Y3_UserCLKo),
    .Tile_X0Y0_FrameData(Row_Y1_FrameData),
    .Tile_X0Y0_FrameData_O(Tile_X0Y1_FrameData_O),
    .Tile_X0Y0_FrameStrobe_O(Tile_X0Y1_FrameStrobe_O),
    .Tile_X0Y1_FrameData(Row_Y2_FrameData),
    .Tile_X0Y1_FrameData_O(Tile_X0Y2_FrameData_O),
    .Tile_X0Y1_FrameStrobe(Tile_X0Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y1_Emulate_Bitstream)
    )
`endif
    Tile_X1Y1_LUT4AB
    (
    .N1END(Tile_X1Y2_N1BEG),
    .N2MID(Tile_X1Y2_N2BEG),
    .N2END(Tile_X1Y2_N2BEGb),
    .N4END(Tile_X1Y2_N4BEG),
    .NN4END(Tile_X1Y2_NN4BEG),
    .Ci(Tile_X1Y2_Co),
    .E1END(Tile_X0Y1_E1BEG),
    .E2MID(Tile_X0Y1_E2BEG),
    .E2END(Tile_X0Y1_E2BEGb),
    .EE4END(Tile_X0Y1_EE4BEG),
    .E6END(Tile_X0Y1_E6BEG),
    .S1END(Tile_X1Y0_S1BEG),
    .S2MID(Tile_X1Y0_S2BEG),
    .S2END(Tile_X1Y0_S2BEGb),
    .S4END(Tile_X1Y0_S4BEG),
    .SS4END(Tile_X1Y0_SS4BEG),
    .W1END(Tile_X2Y1_W1BEG),
    .W2MID(Tile_X2Y1_W2BEG),
    .W2END(Tile_X2Y1_W2BEGb),
    .WW4END(Tile_X2Y1_WW4BEG),
    .W6END(Tile_X2Y1_W6BEG),
    .N1BEG(Tile_X1Y1_N1BEG),
    .N2BEG(Tile_X1Y1_N2BEG),
    .N2BEGb(Tile_X1Y1_N2BEGb),
    .N4BEG(Tile_X1Y1_N4BEG),
    .NN4BEG(Tile_X1Y1_NN4BEG),
    .E1BEG(Tile_X1Y1_E1BEG),
    .E2BEG(Tile_X1Y1_E2BEG),
    .E2BEGb(Tile_X1Y1_E2BEGb),
    .EE4BEG(Tile_X1Y1_EE4BEG),
    .E6BEG(Tile_X1Y1_E6BEG),
    .S1BEG(Tile_X1Y1_S1BEG),
    .S2BEG(Tile_X1Y1_S2BEG),
    .S2BEGb(Tile_X1Y1_S2BEGb),
    .S4BEG(Tile_X1Y1_S4BEG),
    .SS4BEG(Tile_X1Y1_SS4BEG),
    .W1BEG(Tile_X1Y1_W1BEG),
    .W2BEG(Tile_X1Y1_W2BEG),
    .W2BEGb(Tile_X1Y1_W2BEGb),
    .WW4BEG(Tile_X1Y1_WW4BEG),
    .W6BEG(Tile_X1Y1_W6BEG),
    .Co(Tile_X1Y1_Co),
    .UserCLK(Tile_X1Y2_UserCLKo),
    .UserCLKo(Tile_X1Y1_UserCLKo),
    .FrameData(Tile_X0Y1_FrameData_O),
    .FrameData_O(Tile_X1Y1_FrameData_O),
    .FrameStrobe(Tile_X1Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y1_Emulate_Bitstream)
    )
`endif
    Tile_X2Y1_LUT4AB
    (
    .N1END(Tile_X2Y2_N1BEG),
    .N2MID(Tile_X2Y2_N2BEG),
    .N2END(Tile_X2Y2_N2BEGb),
    .N4END(Tile_X2Y2_N4BEG),
    .NN4END(Tile_X2Y2_NN4BEG),
    .Ci(Tile_X2Y2_Co),
    .E1END(Tile_X1Y1_E1BEG),
    .E2MID(Tile_X1Y1_E2BEG),
    .E2END(Tile_X1Y1_E2BEGb),
    .EE4END(Tile_X1Y1_EE4BEG),
    .E6END(Tile_X1Y1_E6BEG),
    .S1END(Tile_X2Y0_S1BEG),
    .S2MID(Tile_X2Y0_S2BEG),
    .S2END(Tile_X2Y0_S2BEGb),
    .S4END(Tile_X2Y0_S4BEG),
    .SS4END(Tile_X2Y0_SS4BEG),
    .W1END(Tile_X3Y1_W1BEG),
    .W2MID(Tile_X3Y1_W2BEG),
    .W2END(Tile_X3Y1_W2BEGb),
    .WW4END(Tile_X3Y1_WW4BEG),
    .W6END(Tile_X3Y1_W6BEG),
    .N1BEG(Tile_X2Y1_N1BEG),
    .N2BEG(Tile_X2Y1_N2BEG),
    .N2BEGb(Tile_X2Y1_N2BEGb),
    .N4BEG(Tile_X2Y1_N4BEG),
    .NN4BEG(Tile_X2Y1_NN4BEG),
    .E1BEG(Tile_X2Y1_E1BEG),
    .E2BEG(Tile_X2Y1_E2BEG),
    .E2BEGb(Tile_X2Y1_E2BEGb),
    .EE4BEG(Tile_X2Y1_EE4BEG),
    .E6BEG(Tile_X2Y1_E6BEG),
    .S1BEG(Tile_X2Y1_S1BEG),
    .S2BEG(Tile_X2Y1_S2BEG),
    .S2BEGb(Tile_X2Y1_S2BEGb),
    .S4BEG(Tile_X2Y1_S4BEG),
    .SS4BEG(Tile_X2Y1_SS4BEG),
    .W1BEG(Tile_X2Y1_W1BEG),
    .W2BEG(Tile_X2Y1_W2BEG),
    .W2BEGb(Tile_X2Y1_W2BEGb),
    .WW4BEG(Tile_X2Y1_WW4BEG),
    .W6BEG(Tile_X2Y1_W6BEG),
    .Co(Tile_X2Y1_Co),
    .UserCLK(Tile_X2Y2_UserCLKo),
    .UserCLKo(Tile_X2Y1_UserCLKo),
    .FrameData(Tile_X1Y1_FrameData_O),
    .FrameData_O(Tile_X2Y1_FrameData_O),
    .FrameStrobe(Tile_X2Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y1_Emulate_Bitstream)
    )
`endif
    Tile_X3Y1_LUT4AB
    (
    .N1END(Tile_X3Y2_N1BEG),
    .N2MID(Tile_X3Y2_N2BEG),
    .N2END(Tile_X3Y2_N2BEGb),
    .N4END(Tile_X3Y2_N4BEG),
    .NN4END(Tile_X3Y2_NN4BEG),
    .Ci(Tile_X3Y2_Co),
    .E1END(Tile_X2Y1_E1BEG),
    .E2MID(Tile_X2Y1_E2BEG),
    .E2END(Tile_X2Y1_E2BEGb),
    .EE4END(Tile_X2Y1_EE4BEG),
    .E6END(Tile_X2Y1_E6BEG),
    .S1END(Tile_X3Y0_S1BEG),
    .S2MID(Tile_X3Y0_S2BEG),
    .S2END(Tile_X3Y0_S2BEGb),
    .S4END(Tile_X3Y0_S4BEG),
    .SS4END(Tile_X3Y0_SS4BEG),
    .W1END(Tile_X4Y1_W1BEG),
    .W2MID(Tile_X4Y1_W2BEG),
    .W2END(Tile_X4Y1_W2BEGb),
    .WW4END(Tile_X4Y1_WW4BEG),
    .W6END(Tile_X4Y1_W6BEG),
    .N1BEG(Tile_X3Y1_N1BEG),
    .N2BEG(Tile_X3Y1_N2BEG),
    .N2BEGb(Tile_X3Y1_N2BEGb),
    .N4BEG(Tile_X3Y1_N4BEG),
    .NN4BEG(Tile_X3Y1_NN4BEG),
    .E1BEG(Tile_X3Y1_E1BEG),
    .E2BEG(Tile_X3Y1_E2BEG),
    .E2BEGb(Tile_X3Y1_E2BEGb),
    .EE4BEG(Tile_X3Y1_EE4BEG),
    .E6BEG(Tile_X3Y1_E6BEG),
    .S1BEG(Tile_X3Y1_S1BEG),
    .S2BEG(Tile_X3Y1_S2BEG),
    .S2BEGb(Tile_X3Y1_S2BEGb),
    .S4BEG(Tile_X3Y1_S4BEG),
    .SS4BEG(Tile_X3Y1_SS4BEG),
    .W1BEG(Tile_X3Y1_W1BEG),
    .W2BEG(Tile_X3Y1_W2BEG),
    .W2BEGb(Tile_X3Y1_W2BEGb),
    .WW4BEG(Tile_X3Y1_WW4BEG),
    .W6BEG(Tile_X3Y1_W6BEG),
    .Co(Tile_X3Y1_Co),
    .UserCLK(Tile_X3Y2_UserCLKo),
    .UserCLKo(Tile_X3Y1_UserCLKo),
    .FrameData(Tile_X2Y1_FrameData_O),
    .FrameData_O(Tile_X3Y1_FrameData_O),
    .FrameStrobe(Tile_X3Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y1_Emulate_Bitstream)
    )
`endif
    Tile_X4Y1_LUT4AB
    (
    .N1END(Tile_X4Y2_N1BEG),
    .N2MID(Tile_X4Y2_N2BEG),
    .N2END(Tile_X4Y2_N2BEGb),
    .N4END(Tile_X4Y2_N4BEG),
    .NN4END(Tile_X4Y2_NN4BEG),
    .Ci(Tile_X4Y2_Co),
    .E1END(Tile_X3Y1_E1BEG),
    .E2MID(Tile_X3Y1_E2BEG),
    .E2END(Tile_X3Y1_E2BEGb),
    .EE4END(Tile_X3Y1_EE4BEG),
    .E6END(Tile_X3Y1_E6BEG),
    .S1END(Tile_X4Y0_S1BEG),
    .S2MID(Tile_X4Y0_S2BEG),
    .S2END(Tile_X4Y0_S2BEGb),
    .S4END(Tile_X4Y0_S4BEG),
    .SS4END(Tile_X4Y0_SS4BEG),
    .W1END(Tile_X5Y1_W1BEG),
    .W2MID(Tile_X5Y1_W2BEG),
    .W2END(Tile_X5Y1_W2BEGb),
    .WW4END(Tile_X5Y1_WW4BEG),
    .W6END(Tile_X5Y1_W6BEG),
    .N1BEG(Tile_X4Y1_N1BEG),
    .N2BEG(Tile_X4Y1_N2BEG),
    .N2BEGb(Tile_X4Y1_N2BEGb),
    .N4BEG(Tile_X4Y1_N4BEG),
    .NN4BEG(Tile_X4Y1_NN4BEG),
    .E1BEG(Tile_X4Y1_E1BEG),
    .E2BEG(Tile_X4Y1_E2BEG),
    .E2BEGb(Tile_X4Y1_E2BEGb),
    .EE4BEG(Tile_X4Y1_EE4BEG),
    .E6BEG(Tile_X4Y1_E6BEG),
    .S1BEG(Tile_X4Y1_S1BEG),
    .S2BEG(Tile_X4Y1_S2BEG),
    .S2BEGb(Tile_X4Y1_S2BEGb),
    .S4BEG(Tile_X4Y1_S4BEG),
    .SS4BEG(Tile_X4Y1_SS4BEG),
    .W1BEG(Tile_X4Y1_W1BEG),
    .W2BEG(Tile_X4Y1_W2BEG),
    .W2BEGb(Tile_X4Y1_W2BEGb),
    .WW4BEG(Tile_X4Y1_WW4BEG),
    .W6BEG(Tile_X4Y1_W6BEG),
    .Co(Tile_X4Y1_Co),
    .UserCLK(Tile_X4Y2_UserCLKo),
    .UserCLKo(Tile_X4Y1_UserCLKo),
    .FrameData(Tile_X3Y1_FrameData_O),
    .FrameData_O(Tile_X4Y1_FrameData_O),
    .FrameStrobe(Tile_X4Y2_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y1_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
IHP_SRAM
`ifdef EMULATION
    #(
    .Tile_X0Y0_Emulate_Bitstream(`Tile_X5Y1_Emulate_Bitstream),
    .Tile_X0Y1_Emulate_Bitstream(`Tile_X5Y2_Emulate_Bitstream)
    )
`endif
    Tile_X5Y1_IHP_SRAM
    (
    .Tile_X0Y0_E1END(Tile_X4Y1_E1BEG),
    .Tile_X0Y0_E2MID(Tile_X4Y1_E2BEG),
    .Tile_X0Y0_E2END(Tile_X4Y1_E2BEGb),
    .Tile_X0Y0_EE4END(Tile_X4Y1_EE4BEG),
    .Tile_X0Y0_E6END(Tile_X4Y1_E6BEG),
    .Tile_X0Y0_S1END(Tile_X5Y0_S1BEG),
    .Tile_X0Y0_S2MID(Tile_X5Y0_S2BEG),
    .Tile_X0Y0_S2END(Tile_X5Y0_S2BEGb),
    .Tile_X0Y0_S4END(Tile_X5Y0_S4BEG),
    .Tile_X0Y1_N1END(Tile_X5Y3_N1BEG),
    .Tile_X0Y1_N2MID(Tile_X5Y3_N2BEG),
    .Tile_X0Y1_N2END(Tile_X5Y3_N2BEGb),
    .Tile_X0Y1_N4END(Tile_X5Y3_N4BEG),
    .Tile_X0Y1_E1END(Tile_X4Y2_E1BEG),
    .Tile_X0Y1_E2MID(Tile_X4Y2_E2BEG),
    .Tile_X0Y1_E2END(Tile_X4Y2_E2BEGb),
    .Tile_X0Y1_EE4END(Tile_X4Y2_EE4BEG),
    .Tile_X0Y1_E6END(Tile_X4Y2_E6BEG),
    .Tile_X0Y0_N1BEG(Tile_X5Y1_N1BEG),
    .Tile_X0Y0_N2BEG(Tile_X5Y1_N2BEG),
    .Tile_X0Y0_N2BEGb(Tile_X5Y1_N2BEGb),
    .Tile_X0Y0_N4BEG(Tile_X5Y1_N4BEG),
    .Tile_X0Y0_W1BEG(Tile_X5Y1_W1BEG),
    .Tile_X0Y0_W2BEG(Tile_X5Y1_W2BEG),
    .Tile_X0Y0_W2BEGb(Tile_X5Y1_W2BEGb),
    .Tile_X0Y0_WW4BEG(Tile_X5Y1_WW4BEG),
    .Tile_X0Y0_W6BEG(Tile_X5Y1_W6BEG),
    .Tile_X0Y1_S1BEG(Tile_X5Y2_S1BEG),
    .Tile_X0Y1_S2BEG(Tile_X5Y2_S2BEG),
    .Tile_X0Y1_S2BEGb(Tile_X5Y2_S2BEGb),
    .Tile_X0Y1_S4BEG(Tile_X5Y2_S4BEG),
    .Tile_X0Y1_W1BEG(Tile_X5Y2_W1BEG),
    .Tile_X0Y1_W2BEG(Tile_X5Y2_W2BEG),
    .Tile_X0Y1_W2BEGb(Tile_X5Y2_W2BEGb),
    .Tile_X0Y1_WW4BEG(Tile_X5Y2_WW4BEG),
    .Tile_X0Y1_W6BEG(Tile_X5Y2_W6BEG),
    .DOUT_SRAM0(Tile_X5Y2_DOUT_SRAM0),
    .DOUT_SRAM1(Tile_X5Y2_DOUT_SRAM1),
    .DOUT_SRAM2(Tile_X5Y2_DOUT_SRAM2),
    .DOUT_SRAM3(Tile_X5Y2_DOUT_SRAM3),
    .DOUT_SRAM4(Tile_X5Y2_DOUT_SRAM4),
    .DOUT_SRAM5(Tile_X5Y2_DOUT_SRAM5),
    .DOUT_SRAM6(Tile_X5Y2_DOUT_SRAM6),
    .DOUT_SRAM7(Tile_X5Y2_DOUT_SRAM7),
    .DOUT_SRAM8(Tile_X5Y2_DOUT_SRAM8),
    .DOUT_SRAM9(Tile_X5Y2_DOUT_SRAM9),
    .DOUT_SRAM10(Tile_X5Y2_DOUT_SRAM10),
    .DOUT_SRAM11(Tile_X5Y2_DOUT_SRAM11),
    .DOUT_SRAM12(Tile_X5Y2_DOUT_SRAM12),
    .DOUT_SRAM13(Tile_X5Y2_DOUT_SRAM13),
    .DOUT_SRAM14(Tile_X5Y2_DOUT_SRAM14),
    .DOUT_SRAM15(Tile_X5Y2_DOUT_SRAM15),
    .DOUT_SRAM16(Tile_X5Y2_DOUT_SRAM16),
    .DOUT_SRAM17(Tile_X5Y2_DOUT_SRAM17),
    .DOUT_SRAM18(Tile_X5Y2_DOUT_SRAM18),
    .DOUT_SRAM19(Tile_X5Y2_DOUT_SRAM19),
    .DOUT_SRAM20(Tile_X5Y2_DOUT_SRAM20),
    .DOUT_SRAM21(Tile_X5Y2_DOUT_SRAM21),
    .DOUT_SRAM22(Tile_X5Y2_DOUT_SRAM22),
    .DOUT_SRAM23(Tile_X5Y2_DOUT_SRAM23),
    .DOUT_SRAM24(Tile_X5Y2_DOUT_SRAM24),
    .DOUT_SRAM25(Tile_X5Y2_DOUT_SRAM25),
    .DOUT_SRAM26(Tile_X5Y2_DOUT_SRAM26),
    .DOUT_SRAM27(Tile_X5Y2_DOUT_SRAM27),
    .DOUT_SRAM28(Tile_X5Y2_DOUT_SRAM28),
    .DOUT_SRAM29(Tile_X5Y2_DOUT_SRAM29),
    .DOUT_SRAM30(Tile_X5Y2_DOUT_SRAM30),
    .DOUT_SRAM31(Tile_X5Y2_DOUT_SRAM31),
    .CONFIGURED_top(Tile_X5Y2_CONFIGURED_top),
    .ADDR_SRAM0(Tile_X5Y2_ADDR_SRAM0),
    .ADDR_SRAM1(Tile_X5Y2_ADDR_SRAM1),
    .ADDR_SRAM2(Tile_X5Y2_ADDR_SRAM2),
    .ADDR_SRAM3(Tile_X5Y2_ADDR_SRAM3),
    .ADDR_SRAM4(Tile_X5Y2_ADDR_SRAM4),
    .ADDR_SRAM5(Tile_X5Y2_ADDR_SRAM5),
    .ADDR_SRAM6(Tile_X5Y2_ADDR_SRAM6),
    .ADDR_SRAM7(Tile_X5Y2_ADDR_SRAM7),
    .ADDR_SRAM8(Tile_X5Y2_ADDR_SRAM8),
    .ADDR_SRAM9(Tile_X5Y2_ADDR_SRAM9),
    .DIN_SRAM0(Tile_X5Y2_DIN_SRAM0),
    .DIN_SRAM1(Tile_X5Y2_DIN_SRAM1),
    .DIN_SRAM2(Tile_X5Y2_DIN_SRAM2),
    .DIN_SRAM3(Tile_X5Y2_DIN_SRAM3),
    .DIN_SRAM4(Tile_X5Y2_DIN_SRAM4),
    .DIN_SRAM5(Tile_X5Y2_DIN_SRAM5),
    .DIN_SRAM6(Tile_X5Y2_DIN_SRAM6),
    .DIN_SRAM7(Tile_X5Y2_DIN_SRAM7),
    .DIN_SRAM8(Tile_X5Y2_DIN_SRAM8),
    .DIN_SRAM9(Tile_X5Y2_DIN_SRAM9),
    .DIN_SRAM10(Tile_X5Y2_DIN_SRAM10),
    .DIN_SRAM11(Tile_X5Y2_DIN_SRAM11),
    .DIN_SRAM12(Tile_X5Y2_DIN_SRAM12),
    .DIN_SRAM13(Tile_X5Y2_DIN_SRAM13),
    .DIN_SRAM14(Tile_X5Y2_DIN_SRAM14),
    .DIN_SRAM15(Tile_X5Y2_DIN_SRAM15),
    .DIN_SRAM16(Tile_X5Y2_DIN_SRAM16),
    .DIN_SRAM17(Tile_X5Y2_DIN_SRAM17),
    .DIN_SRAM18(Tile_X5Y2_DIN_SRAM18),
    .DIN_SRAM19(Tile_X5Y2_DIN_SRAM19),
    .DIN_SRAM20(Tile_X5Y2_DIN_SRAM20),
    .DIN_SRAM21(Tile_X5Y2_DIN_SRAM21),
    .DIN_SRAM22(Tile_X5Y2_DIN_SRAM22),
    .DIN_SRAM23(Tile_X5Y2_DIN_SRAM23),
    .DIN_SRAM24(Tile_X5Y2_DIN_SRAM24),
    .DIN_SRAM25(Tile_X5Y2_DIN_SRAM25),
    .DIN_SRAM26(Tile_X5Y2_DIN_SRAM26),
    .DIN_SRAM27(Tile_X5Y2_DIN_SRAM27),
    .DIN_SRAM28(Tile_X5Y2_DIN_SRAM28),
    .DIN_SRAM29(Tile_X5Y2_DIN_SRAM29),
    .DIN_SRAM30(Tile_X5Y2_DIN_SRAM30),
    .DIN_SRAM31(Tile_X5Y2_DIN_SRAM31),
    .BM_SRAM0(Tile_X5Y2_BM_SRAM0),
    .BM_SRAM1(Tile_X5Y2_BM_SRAM1),
    .BM_SRAM2(Tile_X5Y2_BM_SRAM2),
    .BM_SRAM3(Tile_X5Y2_BM_SRAM3),
    .BM_SRAM4(Tile_X5Y2_BM_SRAM4),
    .BM_SRAM5(Tile_X5Y2_BM_SRAM5),
    .BM_SRAM6(Tile_X5Y2_BM_SRAM6),
    .BM_SRAM7(Tile_X5Y2_BM_SRAM7),
    .BM_SRAM8(Tile_X5Y2_BM_SRAM8),
    .BM_SRAM9(Tile_X5Y2_BM_SRAM9),
    .BM_SRAM10(Tile_X5Y2_BM_SRAM10),
    .BM_SRAM11(Tile_X5Y2_BM_SRAM11),
    .BM_SRAM12(Tile_X5Y2_BM_SRAM12),
    .BM_SRAM13(Tile_X5Y2_BM_SRAM13),
    .BM_SRAM14(Tile_X5Y2_BM_SRAM14),
    .BM_SRAM15(Tile_X5Y2_BM_SRAM15),
    .BM_SRAM16(Tile_X5Y2_BM_SRAM16),
    .BM_SRAM17(Tile_X5Y2_BM_SRAM17),
    .BM_SRAM18(Tile_X5Y2_BM_SRAM18),
    .BM_SRAM19(Tile_X5Y2_BM_SRAM19),
    .BM_SRAM20(Tile_X5Y2_BM_SRAM20),
    .BM_SRAM21(Tile_X5Y2_BM_SRAM21),
    .BM_SRAM22(Tile_X5Y2_BM_SRAM22),
    .BM_SRAM23(Tile_X5Y2_BM_SRAM23),
    .BM_SRAM24(Tile_X5Y2_BM_SRAM24),
    .BM_SRAM25(Tile_X5Y2_BM_SRAM25),
    .BM_SRAM26(Tile_X5Y2_BM_SRAM26),
    .BM_SRAM27(Tile_X5Y2_BM_SRAM27),
    .BM_SRAM28(Tile_X5Y2_BM_SRAM28),
    .BM_SRAM29(Tile_X5Y2_BM_SRAM29),
    .BM_SRAM30(Tile_X5Y2_BM_SRAM30),
    .BM_SRAM31(Tile_X5Y2_BM_SRAM31),
    .WEN_SRAM(Tile_X5Y2_WEN_SRAM),
    .MEN_SRAM(Tile_X5Y2_MEN_SRAM),
    .REN_SRAM(Tile_X5Y2_REN_SRAM),
    .CLK_SRAM(Tile_X5Y2_CLK_SRAM),
    .TIE_HIGH_SRAM(Tile_X5Y2_TIE_HIGH_SRAM),
    .TIE_LOW_SRAM(Tile_X5Y2_TIE_LOW_SRAM),
    .Tile_X0Y0_UserCLKo(Tile_X5Y1_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X5Y3_UserCLKo),
    .Tile_X0Y0_FrameData(Tile_X4Y1_FrameData_O),
    .Tile_X0Y0_FrameData_O(Tile_X5Y1_FrameData_O),
    .Tile_X0Y0_FrameStrobe_O(Tile_X5Y1_FrameStrobe_O),
    .Tile_X0Y1_FrameData(Tile_X4Y2_FrameData_O),
    .Tile_X0Y1_FrameData_O(Tile_X5Y2_FrameData_O),
    .Tile_X0Y1_FrameStrobe(Tile_X5Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y2_Emulate_Bitstream)
    )
`endif
    Tile_X1Y2_LUT4AB
    (
    .N1END(Tile_X1Y3_N1BEG),
    .N2MID(Tile_X1Y3_N2BEG),
    .N2END(Tile_X1Y3_N2BEGb),
    .N4END(Tile_X1Y3_N4BEG),
    .NN4END(Tile_X1Y3_NN4BEG),
    .Ci(Tile_X1Y3_Co),
    .E1END(Tile_X0Y2_E1BEG),
    .E2MID(Tile_X0Y2_E2BEG),
    .E2END(Tile_X0Y2_E2BEGb),
    .EE4END(Tile_X0Y2_EE4BEG),
    .E6END(Tile_X0Y2_E6BEG),
    .S1END(Tile_X1Y1_S1BEG),
    .S2MID(Tile_X1Y1_S2BEG),
    .S2END(Tile_X1Y1_S2BEGb),
    .S4END(Tile_X1Y1_S4BEG),
    .SS4END(Tile_X1Y1_SS4BEG),
    .W1END(Tile_X2Y2_W1BEG),
    .W2MID(Tile_X2Y2_W2BEG),
    .W2END(Tile_X2Y2_W2BEGb),
    .WW4END(Tile_X2Y2_WW4BEG),
    .W6END(Tile_X2Y2_W6BEG),
    .N1BEG(Tile_X1Y2_N1BEG),
    .N2BEG(Tile_X1Y2_N2BEG),
    .N2BEGb(Tile_X1Y2_N2BEGb),
    .N4BEG(Tile_X1Y2_N4BEG),
    .NN4BEG(Tile_X1Y2_NN4BEG),
    .E1BEG(Tile_X1Y2_E1BEG),
    .E2BEG(Tile_X1Y2_E2BEG),
    .E2BEGb(Tile_X1Y2_E2BEGb),
    .EE4BEG(Tile_X1Y2_EE4BEG),
    .E6BEG(Tile_X1Y2_E6BEG),
    .S1BEG(Tile_X1Y2_S1BEG),
    .S2BEG(Tile_X1Y2_S2BEG),
    .S2BEGb(Tile_X1Y2_S2BEGb),
    .S4BEG(Tile_X1Y2_S4BEG),
    .SS4BEG(Tile_X1Y2_SS4BEG),
    .W1BEG(Tile_X1Y2_W1BEG),
    .W2BEG(Tile_X1Y2_W2BEG),
    .W2BEGb(Tile_X1Y2_W2BEGb),
    .WW4BEG(Tile_X1Y2_WW4BEG),
    .W6BEG(Tile_X1Y2_W6BEG),
    .Co(Tile_X1Y2_Co),
    .UserCLK(Tile_X1Y3_UserCLKo),
    .UserCLKo(Tile_X1Y2_UserCLKo),
    .FrameData(Tile_X0Y2_FrameData_O),
    .FrameData_O(Tile_X1Y2_FrameData_O),
    .FrameStrobe(Tile_X1Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y2_Emulate_Bitstream)
    )
`endif
    Tile_X2Y2_LUT4AB
    (
    .N1END(Tile_X2Y3_N1BEG),
    .N2MID(Tile_X2Y3_N2BEG),
    .N2END(Tile_X2Y3_N2BEGb),
    .N4END(Tile_X2Y3_N4BEG),
    .NN4END(Tile_X2Y3_NN4BEG),
    .Ci(Tile_X2Y3_Co),
    .E1END(Tile_X1Y2_E1BEG),
    .E2MID(Tile_X1Y2_E2BEG),
    .E2END(Tile_X1Y2_E2BEGb),
    .EE4END(Tile_X1Y2_EE4BEG),
    .E6END(Tile_X1Y2_E6BEG),
    .S1END(Tile_X2Y1_S1BEG),
    .S2MID(Tile_X2Y1_S2BEG),
    .S2END(Tile_X2Y1_S2BEGb),
    .S4END(Tile_X2Y1_S4BEG),
    .SS4END(Tile_X2Y1_SS4BEG),
    .W1END(Tile_X3Y2_W1BEG),
    .W2MID(Tile_X3Y2_W2BEG),
    .W2END(Tile_X3Y2_W2BEGb),
    .WW4END(Tile_X3Y2_WW4BEG),
    .W6END(Tile_X3Y2_W6BEG),
    .N1BEG(Tile_X2Y2_N1BEG),
    .N2BEG(Tile_X2Y2_N2BEG),
    .N2BEGb(Tile_X2Y2_N2BEGb),
    .N4BEG(Tile_X2Y2_N4BEG),
    .NN4BEG(Tile_X2Y2_NN4BEG),
    .E1BEG(Tile_X2Y2_E1BEG),
    .E2BEG(Tile_X2Y2_E2BEG),
    .E2BEGb(Tile_X2Y2_E2BEGb),
    .EE4BEG(Tile_X2Y2_EE4BEG),
    .E6BEG(Tile_X2Y2_E6BEG),
    .S1BEG(Tile_X2Y2_S1BEG),
    .S2BEG(Tile_X2Y2_S2BEG),
    .S2BEGb(Tile_X2Y2_S2BEGb),
    .S4BEG(Tile_X2Y2_S4BEG),
    .SS4BEG(Tile_X2Y2_SS4BEG),
    .W1BEG(Tile_X2Y2_W1BEG),
    .W2BEG(Tile_X2Y2_W2BEG),
    .W2BEGb(Tile_X2Y2_W2BEGb),
    .WW4BEG(Tile_X2Y2_WW4BEG),
    .W6BEG(Tile_X2Y2_W6BEG),
    .Co(Tile_X2Y2_Co),
    .UserCLK(Tile_X2Y3_UserCLKo),
    .UserCLKo(Tile_X2Y2_UserCLKo),
    .FrameData(Tile_X1Y2_FrameData_O),
    .FrameData_O(Tile_X2Y2_FrameData_O),
    .FrameStrobe(Tile_X2Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y2_Emulate_Bitstream)
    )
`endif
    Tile_X3Y2_LUT4AB
    (
    .N1END(Tile_X3Y3_N1BEG),
    .N2MID(Tile_X3Y3_N2BEG),
    .N2END(Tile_X3Y3_N2BEGb),
    .N4END(Tile_X3Y3_N4BEG),
    .NN4END(Tile_X3Y3_NN4BEG),
    .Ci(Tile_X3Y3_Co),
    .E1END(Tile_X2Y2_E1BEG),
    .E2MID(Tile_X2Y2_E2BEG),
    .E2END(Tile_X2Y2_E2BEGb),
    .EE4END(Tile_X2Y2_EE4BEG),
    .E6END(Tile_X2Y2_E6BEG),
    .S1END(Tile_X3Y1_S1BEG),
    .S2MID(Tile_X3Y1_S2BEG),
    .S2END(Tile_X3Y1_S2BEGb),
    .S4END(Tile_X3Y1_S4BEG),
    .SS4END(Tile_X3Y1_SS4BEG),
    .W1END(Tile_X4Y2_W1BEG),
    .W2MID(Tile_X4Y2_W2BEG),
    .W2END(Tile_X4Y2_W2BEGb),
    .WW4END(Tile_X4Y2_WW4BEG),
    .W6END(Tile_X4Y2_W6BEG),
    .N1BEG(Tile_X3Y2_N1BEG),
    .N2BEG(Tile_X3Y2_N2BEG),
    .N2BEGb(Tile_X3Y2_N2BEGb),
    .N4BEG(Tile_X3Y2_N4BEG),
    .NN4BEG(Tile_X3Y2_NN4BEG),
    .E1BEG(Tile_X3Y2_E1BEG),
    .E2BEG(Tile_X3Y2_E2BEG),
    .E2BEGb(Tile_X3Y2_E2BEGb),
    .EE4BEG(Tile_X3Y2_EE4BEG),
    .E6BEG(Tile_X3Y2_E6BEG),
    .S1BEG(Tile_X3Y2_S1BEG),
    .S2BEG(Tile_X3Y2_S2BEG),
    .S2BEGb(Tile_X3Y2_S2BEGb),
    .S4BEG(Tile_X3Y2_S4BEG),
    .SS4BEG(Tile_X3Y2_SS4BEG),
    .W1BEG(Tile_X3Y2_W1BEG),
    .W2BEG(Tile_X3Y2_W2BEG),
    .W2BEGb(Tile_X3Y2_W2BEGb),
    .WW4BEG(Tile_X3Y2_WW4BEG),
    .W6BEG(Tile_X3Y2_W6BEG),
    .Co(Tile_X3Y2_Co),
    .UserCLK(Tile_X3Y3_UserCLKo),
    .UserCLKo(Tile_X3Y2_UserCLKo),
    .FrameData(Tile_X2Y2_FrameData_O),
    .FrameData_O(Tile_X3Y2_FrameData_O),
    .FrameStrobe(Tile_X3Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y2_Emulate_Bitstream)
    )
`endif
    Tile_X4Y2_LUT4AB
    (
    .N1END(Tile_X4Y3_N1BEG),
    .N2MID(Tile_X4Y3_N2BEG),
    .N2END(Tile_X4Y3_N2BEGb),
    .N4END(Tile_X4Y3_N4BEG),
    .NN4END(Tile_X4Y3_NN4BEG),
    .Ci(Tile_X4Y3_Co),
    .E1END(Tile_X3Y2_E1BEG),
    .E2MID(Tile_X3Y2_E2BEG),
    .E2END(Tile_X3Y2_E2BEGb),
    .EE4END(Tile_X3Y2_EE4BEG),
    .E6END(Tile_X3Y2_E6BEG),
    .S1END(Tile_X4Y1_S1BEG),
    .S2MID(Tile_X4Y1_S2BEG),
    .S2END(Tile_X4Y1_S2BEGb),
    .S4END(Tile_X4Y1_S4BEG),
    .SS4END(Tile_X4Y1_SS4BEG),
    .W1END(Tile_X5Y2_W1BEG),
    .W2MID(Tile_X5Y2_W2BEG),
    .W2END(Tile_X5Y2_W2BEGb),
    .WW4END(Tile_X5Y2_WW4BEG),
    .W6END(Tile_X5Y2_W6BEG),
    .N1BEG(Tile_X4Y2_N1BEG),
    .N2BEG(Tile_X4Y2_N2BEG),
    .N2BEGb(Tile_X4Y2_N2BEGb),
    .N4BEG(Tile_X4Y2_N4BEG),
    .NN4BEG(Tile_X4Y2_NN4BEG),
    .E1BEG(Tile_X4Y2_E1BEG),
    .E2BEG(Tile_X4Y2_E2BEG),
    .E2BEGb(Tile_X4Y2_E2BEGb),
    .EE4BEG(Tile_X4Y2_EE4BEG),
    .E6BEG(Tile_X4Y2_E6BEG),
    .S1BEG(Tile_X4Y2_S1BEG),
    .S2BEG(Tile_X4Y2_S2BEG),
    .S2BEGb(Tile_X4Y2_S2BEGb),
    .S4BEG(Tile_X4Y2_S4BEG),
    .SS4BEG(Tile_X4Y2_SS4BEG),
    .W1BEG(Tile_X4Y2_W1BEG),
    .W2BEG(Tile_X4Y2_W2BEG),
    .W2BEGb(Tile_X4Y2_W2BEGb),
    .WW4BEG(Tile_X4Y2_WW4BEG),
    .W6BEG(Tile_X4Y2_W6BEG),
    .Co(Tile_X4Y2_Co),
    .UserCLK(Tile_X4Y3_UserCLKo),
    .UserCLKo(Tile_X4Y2_UserCLKo),
    .FrameData(Tile_X3Y2_FrameData_O),
    .FrameData_O(Tile_X4Y2_FrameData_O),
    .FrameStrobe(Tile_X4Y3_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y2_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_TT_IF
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y3_Emulate_Bitstream)
    )
`endif
    Tile_X0Y3_W_TT_IF
    (
    .N1END(Tile_X0Y4_N1BEG),
    .N2MID(Tile_X0Y4_N2BEG),
    .N2END(Tile_X0Y4_N2BEGb),
    .N4END(Tile_X0Y4_N4BEG),
    .S1END(Tile_X0Y2_S1BEG),
    .S2MID(Tile_X0Y2_S2BEG),
    .S2END(Tile_X0Y2_S2BEGb),
    .S4END(Tile_X0Y2_S4BEG),
    .W1END(Tile_X1Y3_W1BEG),
    .W2MID(Tile_X1Y3_W2BEG),
    .W2END(Tile_X1Y3_W2BEGb),
    .WW4END(Tile_X1Y3_WW4BEG),
    .W6END(Tile_X1Y3_W6BEG),
    .N1BEG(Tile_X0Y3_N1BEG),
    .N2BEG(Tile_X0Y3_N2BEG),
    .N2BEGb(Tile_X0Y3_N2BEGb),
    .N4BEG(Tile_X0Y3_N4BEG),
    .S1BEG(Tile_X0Y3_S1BEG),
    .S2BEG(Tile_X0Y3_S2BEG),
    .S2BEGb(Tile_X0Y3_S2BEGb),
    .S4BEG(Tile_X0Y3_S4BEG),
    .E1BEG(Tile_X0Y3_E1BEG),
    .E2BEG(Tile_X0Y3_E2BEG),
    .E2BEGb(Tile_X0Y3_E2BEGb),
    .EE4BEG(Tile_X0Y3_EE4BEG),
    .E6BEG(Tile_X0Y3_E6BEG),
    .UO_OUT_TT_PROJECT0(Tile_X0Y3_UO_OUT_TT_PROJECT0),
    .UO_OUT_TT_PROJECT1(Tile_X0Y3_UO_OUT_TT_PROJECT1),
    .UO_OUT_TT_PROJECT2(Tile_X0Y3_UO_OUT_TT_PROJECT2),
    .UO_OUT_TT_PROJECT3(Tile_X0Y3_UO_OUT_TT_PROJECT3),
    .UO_OUT_TT_PROJECT4(Tile_X0Y3_UO_OUT_TT_PROJECT4),
    .UO_OUT_TT_PROJECT5(Tile_X0Y3_UO_OUT_TT_PROJECT5),
    .UO_OUT_TT_PROJECT6(Tile_X0Y3_UO_OUT_TT_PROJECT6),
    .UO_OUT_TT_PROJECT7(Tile_X0Y3_UO_OUT_TT_PROJECT7),
    .UIO_OUT_TT_PROJECT0(Tile_X0Y3_UIO_OUT_TT_PROJECT0),
    .UIO_OUT_TT_PROJECT1(Tile_X0Y3_UIO_OUT_TT_PROJECT1),
    .UIO_OUT_TT_PROJECT2(Tile_X0Y3_UIO_OUT_TT_PROJECT2),
    .UIO_OUT_TT_PROJECT3(Tile_X0Y3_UIO_OUT_TT_PROJECT3),
    .UIO_OUT_TT_PROJECT4(Tile_X0Y3_UIO_OUT_TT_PROJECT4),
    .UIO_OUT_TT_PROJECT5(Tile_X0Y3_UIO_OUT_TT_PROJECT5),
    .UIO_OUT_TT_PROJECT6(Tile_X0Y3_UIO_OUT_TT_PROJECT6),
    .UIO_OUT_TT_PROJECT7(Tile_X0Y3_UIO_OUT_TT_PROJECT7),
    .UIO_OE_TT_PROJECT0(Tile_X0Y3_UIO_OE_TT_PROJECT0),
    .UIO_OE_TT_PROJECT1(Tile_X0Y3_UIO_OE_TT_PROJECT1),
    .UIO_OE_TT_PROJECT2(Tile_X0Y3_UIO_OE_TT_PROJECT2),
    .UIO_OE_TT_PROJECT3(Tile_X0Y3_UIO_OE_TT_PROJECT3),
    .UIO_OE_TT_PROJECT4(Tile_X0Y3_UIO_OE_TT_PROJECT4),
    .UIO_OE_TT_PROJECT5(Tile_X0Y3_UIO_OE_TT_PROJECT5),
    .UIO_OE_TT_PROJECT6(Tile_X0Y3_UIO_OE_TT_PROJECT6),
    .UIO_OE_TT_PROJECT7(Tile_X0Y3_UIO_OE_TT_PROJECT7),
    .UI_IN_TT_PROJECT0(Tile_X0Y3_UI_IN_TT_PROJECT0),
    .UI_IN_TT_PROJECT1(Tile_X0Y3_UI_IN_TT_PROJECT1),
    .UI_IN_TT_PROJECT2(Tile_X0Y3_UI_IN_TT_PROJECT2),
    .UI_IN_TT_PROJECT3(Tile_X0Y3_UI_IN_TT_PROJECT3),
    .UI_IN_TT_PROJECT4(Tile_X0Y3_UI_IN_TT_PROJECT4),
    .UI_IN_TT_PROJECT5(Tile_X0Y3_UI_IN_TT_PROJECT5),
    .UI_IN_TT_PROJECT6(Tile_X0Y3_UI_IN_TT_PROJECT6),
    .UI_IN_TT_PROJECT7(Tile_X0Y3_UI_IN_TT_PROJECT7),
    .UIO_IN_TT_PROJECT0(Tile_X0Y3_UIO_IN_TT_PROJECT0),
    .UIO_IN_TT_PROJECT1(Tile_X0Y3_UIO_IN_TT_PROJECT1),
    .UIO_IN_TT_PROJECT2(Tile_X0Y3_UIO_IN_TT_PROJECT2),
    .UIO_IN_TT_PROJECT3(Tile_X0Y3_UIO_IN_TT_PROJECT3),
    .UIO_IN_TT_PROJECT4(Tile_X0Y3_UIO_IN_TT_PROJECT4),
    .UIO_IN_TT_PROJECT5(Tile_X0Y3_UIO_IN_TT_PROJECT5),
    .UIO_IN_TT_PROJECT6(Tile_X0Y3_UIO_IN_TT_PROJECT6),
    .UIO_IN_TT_PROJECT7(Tile_X0Y3_UIO_IN_TT_PROJECT7),
    .ENA_TT_PROJECT(Tile_X0Y3_ENA_TT_PROJECT),
    .CLK_TT_PROJECT(Tile_X0Y3_CLK_TT_PROJECT),
    .RST_N_TT_PROJECT(Tile_X0Y3_RST_N_TT_PROJECT),
    .UserCLK(Tile_X0Y4_UserCLKo),
    .UserCLKo(Tile_X0Y3_UserCLKo),
    .FrameData(Row_Y3_FrameData),
    .FrameData_O(Tile_X0Y3_FrameData_O),
    .FrameStrobe(Tile_X0Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y3_Emulate_Bitstream)
    )
`endif
    Tile_X1Y3_LUT4AB
    (
    .N1END(Tile_X1Y4_N1BEG),
    .N2MID(Tile_X1Y4_N2BEG),
    .N2END(Tile_X1Y4_N2BEGb),
    .N4END(Tile_X1Y4_N4BEG),
    .NN4END(Tile_X1Y4_NN4BEG),
    .Ci(Tile_X1Y4_Co),
    .E1END(Tile_X0Y3_E1BEG),
    .E2MID(Tile_X0Y3_E2BEG),
    .E2END(Tile_X0Y3_E2BEGb),
    .EE4END(Tile_X0Y3_EE4BEG),
    .E6END(Tile_X0Y3_E6BEG),
    .S1END(Tile_X1Y2_S1BEG),
    .S2MID(Tile_X1Y2_S2BEG),
    .S2END(Tile_X1Y2_S2BEGb),
    .S4END(Tile_X1Y2_S4BEG),
    .SS4END(Tile_X1Y2_SS4BEG),
    .W1END(Tile_X2Y3_W1BEG),
    .W2MID(Tile_X2Y3_W2BEG),
    .W2END(Tile_X2Y3_W2BEGb),
    .WW4END(Tile_X2Y3_WW4BEG),
    .W6END(Tile_X2Y3_W6BEG),
    .N1BEG(Tile_X1Y3_N1BEG),
    .N2BEG(Tile_X1Y3_N2BEG),
    .N2BEGb(Tile_X1Y3_N2BEGb),
    .N4BEG(Tile_X1Y3_N4BEG),
    .NN4BEG(Tile_X1Y3_NN4BEG),
    .E1BEG(Tile_X1Y3_E1BEG),
    .E2BEG(Tile_X1Y3_E2BEG),
    .E2BEGb(Tile_X1Y3_E2BEGb),
    .EE4BEG(Tile_X1Y3_EE4BEG),
    .E6BEG(Tile_X1Y3_E6BEG),
    .S1BEG(Tile_X1Y3_S1BEG),
    .S2BEG(Tile_X1Y3_S2BEG),
    .S2BEGb(Tile_X1Y3_S2BEGb),
    .S4BEG(Tile_X1Y3_S4BEG),
    .SS4BEG(Tile_X1Y3_SS4BEG),
    .W1BEG(Tile_X1Y3_W1BEG),
    .W2BEG(Tile_X1Y3_W2BEG),
    .W2BEGb(Tile_X1Y3_W2BEGb),
    .WW4BEG(Tile_X1Y3_WW4BEG),
    .W6BEG(Tile_X1Y3_W6BEG),
    .Co(Tile_X1Y3_Co),
    .UserCLK(Tile_X1Y4_UserCLKo),
    .UserCLKo(Tile_X1Y3_UserCLKo),
    .FrameData(Tile_X0Y3_FrameData_O),
    .FrameData_O(Tile_X1Y3_FrameData_O),
    .FrameStrobe(Tile_X1Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y3_Emulate_Bitstream)
    )
`endif
    Tile_X2Y3_LUT4AB
    (
    .N1END(Tile_X2Y4_N1BEG),
    .N2MID(Tile_X2Y4_N2BEG),
    .N2END(Tile_X2Y4_N2BEGb),
    .N4END(Tile_X2Y4_N4BEG),
    .NN4END(Tile_X2Y4_NN4BEG),
    .Ci(Tile_X2Y4_Co),
    .E1END(Tile_X1Y3_E1BEG),
    .E2MID(Tile_X1Y3_E2BEG),
    .E2END(Tile_X1Y3_E2BEGb),
    .EE4END(Tile_X1Y3_EE4BEG),
    .E6END(Tile_X1Y3_E6BEG),
    .S1END(Tile_X2Y2_S1BEG),
    .S2MID(Tile_X2Y2_S2BEG),
    .S2END(Tile_X2Y2_S2BEGb),
    .S4END(Tile_X2Y2_S4BEG),
    .SS4END(Tile_X2Y2_SS4BEG),
    .W1END(Tile_X3Y3_W1BEG),
    .W2MID(Tile_X3Y3_W2BEG),
    .W2END(Tile_X3Y3_W2BEGb),
    .WW4END(Tile_X3Y3_WW4BEG),
    .W6END(Tile_X3Y3_W6BEG),
    .N1BEG(Tile_X2Y3_N1BEG),
    .N2BEG(Tile_X2Y3_N2BEG),
    .N2BEGb(Tile_X2Y3_N2BEGb),
    .N4BEG(Tile_X2Y3_N4BEG),
    .NN4BEG(Tile_X2Y3_NN4BEG),
    .E1BEG(Tile_X2Y3_E1BEG),
    .E2BEG(Tile_X2Y3_E2BEG),
    .E2BEGb(Tile_X2Y3_E2BEGb),
    .EE4BEG(Tile_X2Y3_EE4BEG),
    .E6BEG(Tile_X2Y3_E6BEG),
    .S1BEG(Tile_X2Y3_S1BEG),
    .S2BEG(Tile_X2Y3_S2BEG),
    .S2BEGb(Tile_X2Y3_S2BEGb),
    .S4BEG(Tile_X2Y3_S4BEG),
    .SS4BEG(Tile_X2Y3_SS4BEG),
    .W1BEG(Tile_X2Y3_W1BEG),
    .W2BEG(Tile_X2Y3_W2BEG),
    .W2BEGb(Tile_X2Y3_W2BEGb),
    .WW4BEG(Tile_X2Y3_WW4BEG),
    .W6BEG(Tile_X2Y3_W6BEG),
    .Co(Tile_X2Y3_Co),
    .UserCLK(Tile_X2Y4_UserCLKo),
    .UserCLKo(Tile_X2Y3_UserCLKo),
    .FrameData(Tile_X1Y3_FrameData_O),
    .FrameData_O(Tile_X2Y3_FrameData_O),
    .FrameStrobe(Tile_X2Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y3_Emulate_Bitstream)
    )
`endif
    Tile_X3Y3_LUT4AB
    (
    .N1END(Tile_X3Y4_N1BEG),
    .N2MID(Tile_X3Y4_N2BEG),
    .N2END(Tile_X3Y4_N2BEGb),
    .N4END(Tile_X3Y4_N4BEG),
    .NN4END(Tile_X3Y4_NN4BEG),
    .Ci(Tile_X3Y4_Co),
    .E1END(Tile_X2Y3_E1BEG),
    .E2MID(Tile_X2Y3_E2BEG),
    .E2END(Tile_X2Y3_E2BEGb),
    .EE4END(Tile_X2Y3_EE4BEG),
    .E6END(Tile_X2Y3_E6BEG),
    .S1END(Tile_X3Y2_S1BEG),
    .S2MID(Tile_X3Y2_S2BEG),
    .S2END(Tile_X3Y2_S2BEGb),
    .S4END(Tile_X3Y2_S4BEG),
    .SS4END(Tile_X3Y2_SS4BEG),
    .W1END(Tile_X4Y3_W1BEG),
    .W2MID(Tile_X4Y3_W2BEG),
    .W2END(Tile_X4Y3_W2BEGb),
    .WW4END(Tile_X4Y3_WW4BEG),
    .W6END(Tile_X4Y3_W6BEG),
    .N1BEG(Tile_X3Y3_N1BEG),
    .N2BEG(Tile_X3Y3_N2BEG),
    .N2BEGb(Tile_X3Y3_N2BEGb),
    .N4BEG(Tile_X3Y3_N4BEG),
    .NN4BEG(Tile_X3Y3_NN4BEG),
    .E1BEG(Tile_X3Y3_E1BEG),
    .E2BEG(Tile_X3Y3_E2BEG),
    .E2BEGb(Tile_X3Y3_E2BEGb),
    .EE4BEG(Tile_X3Y3_EE4BEG),
    .E6BEG(Tile_X3Y3_E6BEG),
    .S1BEG(Tile_X3Y3_S1BEG),
    .S2BEG(Tile_X3Y3_S2BEG),
    .S2BEGb(Tile_X3Y3_S2BEGb),
    .S4BEG(Tile_X3Y3_S4BEG),
    .SS4BEG(Tile_X3Y3_SS4BEG),
    .W1BEG(Tile_X3Y3_W1BEG),
    .W2BEG(Tile_X3Y3_W2BEG),
    .W2BEGb(Tile_X3Y3_W2BEGb),
    .WW4BEG(Tile_X3Y3_WW4BEG),
    .W6BEG(Tile_X3Y3_W6BEG),
    .Co(Tile_X3Y3_Co),
    .UserCLK(Tile_X3Y4_UserCLKo),
    .UserCLKo(Tile_X3Y3_UserCLKo),
    .FrameData(Tile_X2Y3_FrameData_O),
    .FrameData_O(Tile_X3Y3_FrameData_O),
    .FrameStrobe(Tile_X3Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y3_Emulate_Bitstream)
    )
`endif
    Tile_X4Y3_LUT4AB
    (
    .N1END(Tile_X4Y4_N1BEG),
    .N2MID(Tile_X4Y4_N2BEG),
    .N2END(Tile_X4Y4_N2BEGb),
    .N4END(Tile_X4Y4_N4BEG),
    .NN4END(Tile_X4Y4_NN4BEG),
    .Ci(Tile_X4Y4_Co),
    .E1END(Tile_X3Y3_E1BEG),
    .E2MID(Tile_X3Y3_E2BEG),
    .E2END(Tile_X3Y3_E2BEGb),
    .EE4END(Tile_X3Y3_EE4BEG),
    .E6END(Tile_X3Y3_E6BEG),
    .S1END(Tile_X4Y2_S1BEG),
    .S2MID(Tile_X4Y2_S2BEG),
    .S2END(Tile_X4Y2_S2BEGb),
    .S4END(Tile_X4Y2_S4BEG),
    .SS4END(Tile_X4Y2_SS4BEG),
    .W1END(Tile_X5Y3_W1BEG),
    .W2MID(Tile_X5Y3_W2BEG),
    .W2END(Tile_X5Y3_W2BEGb),
    .WW4END(Tile_X5Y3_WW4BEG),
    .W6END(Tile_X5Y3_W6BEG),
    .N1BEG(Tile_X4Y3_N1BEG),
    .N2BEG(Tile_X4Y3_N2BEG),
    .N2BEGb(Tile_X4Y3_N2BEGb),
    .N4BEG(Tile_X4Y3_N4BEG),
    .NN4BEG(Tile_X4Y3_NN4BEG),
    .E1BEG(Tile_X4Y3_E1BEG),
    .E2BEG(Tile_X4Y3_E2BEG),
    .E2BEGb(Tile_X4Y3_E2BEGb),
    .EE4BEG(Tile_X4Y3_EE4BEG),
    .E6BEG(Tile_X4Y3_E6BEG),
    .S1BEG(Tile_X4Y3_S1BEG),
    .S2BEG(Tile_X4Y3_S2BEG),
    .S2BEGb(Tile_X4Y3_S2BEGb),
    .S4BEG(Tile_X4Y3_S4BEG),
    .SS4BEG(Tile_X4Y3_SS4BEG),
    .W1BEG(Tile_X4Y3_W1BEG),
    .W2BEG(Tile_X4Y3_W2BEG),
    .W2BEGb(Tile_X4Y3_W2BEGb),
    .WW4BEG(Tile_X4Y3_WW4BEG),
    .W6BEG(Tile_X4Y3_W6BEG),
    .Co(Tile_X4Y3_Co),
    .UserCLK(Tile_X4Y4_UserCLKo),
    .UserCLKo(Tile_X4Y3_UserCLKo),
    .FrameData(Tile_X3Y3_FrameData_O),
    .FrameData_O(Tile_X4Y3_FrameData_O),
    .FrameStrobe(Tile_X4Y4_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y3_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
E_TT_IF2
`ifdef EMULATION
    #(
    .Tile_X0Y0_Emulate_Bitstream(`Tile_X5Y3_Emulate_Bitstream),
    .Tile_X0Y1_Emulate_Bitstream(`Tile_X5Y4_Emulate_Bitstream)
    )
`endif
    Tile_X5Y3_E_TT_IF2
    (
    .Tile_X0Y0_E1END(Tile_X4Y3_E1BEG),
    .Tile_X0Y0_E2MID(Tile_X4Y3_E2BEG),
    .Tile_X0Y0_E2END(Tile_X4Y3_E2BEGb),
    .Tile_X0Y0_EE4END(Tile_X4Y3_EE4BEG),
    .Tile_X0Y0_E6END(Tile_X4Y3_E6BEG),
    .Tile_X0Y0_S1END(Tile_X5Y2_S1BEG),
    .Tile_X0Y0_S2MID(Tile_X5Y2_S2BEG),
    .Tile_X0Y0_S2END(Tile_X5Y2_S2BEGb),
    .Tile_X0Y0_S4END(Tile_X5Y2_S4BEG),
    .Tile_X0Y1_N1END(Tile_X5Y5_N1BEG),
    .Tile_X0Y1_N2MID(Tile_X5Y5_N2BEG),
    .Tile_X0Y1_N2END(Tile_X5Y5_N2BEGb),
    .Tile_X0Y1_N4END(Tile_X5Y5_N4BEG),
    .Tile_X0Y1_E1END(Tile_X4Y4_E1BEG),
    .Tile_X0Y1_E2MID(Tile_X4Y4_E2BEG),
    .Tile_X0Y1_E2END(Tile_X4Y4_E2BEGb),
    .Tile_X0Y1_EE4END(Tile_X4Y4_EE4BEG),
    .Tile_X0Y1_E6END(Tile_X4Y4_E6BEG),
    .Tile_X0Y0_N1BEG(Tile_X5Y3_N1BEG),
    .Tile_X0Y0_N2BEG(Tile_X5Y3_N2BEG),
    .Tile_X0Y0_N2BEGb(Tile_X5Y3_N2BEGb),
    .Tile_X0Y0_N4BEG(Tile_X5Y3_N4BEG),
    .Tile_X0Y0_W1BEG(Tile_X5Y3_W1BEG),
    .Tile_X0Y0_W2BEG(Tile_X5Y3_W2BEG),
    .Tile_X0Y0_W2BEGb(Tile_X5Y3_W2BEGb),
    .Tile_X0Y0_WW4BEG(Tile_X5Y3_WW4BEG),
    .Tile_X0Y0_W6BEG(Tile_X5Y3_W6BEG),
    .Tile_X0Y1_S1BEG(Tile_X5Y4_S1BEG),
    .Tile_X0Y1_S2BEG(Tile_X5Y4_S2BEG),
    .Tile_X0Y1_S2BEGb(Tile_X5Y4_S2BEGb),
    .Tile_X0Y1_S4BEG(Tile_X5Y4_S4BEG),
    .Tile_X0Y1_W1BEG(Tile_X5Y4_W1BEG),
    .Tile_X0Y1_W2BEG(Tile_X5Y4_W2BEG),
    .Tile_X0Y1_W2BEGb(Tile_X5Y4_W2BEGb),
    .Tile_X0Y1_WW4BEG(Tile_X5Y4_WW4BEG),
    .Tile_X0Y1_W6BEG(Tile_X5Y4_W6BEG),
    .UO_OUT_TT_PROJECT0(Tile_X5Y4_UO_OUT_TT_PROJECT0),
    .UO_OUT_TT_PROJECT1(Tile_X5Y4_UO_OUT_TT_PROJECT1),
    .UO_OUT_TT_PROJECT2(Tile_X5Y4_UO_OUT_TT_PROJECT2),
    .UO_OUT_TT_PROJECT3(Tile_X5Y4_UO_OUT_TT_PROJECT3),
    .UO_OUT_TT_PROJECT4(Tile_X5Y4_UO_OUT_TT_PROJECT4),
    .UO_OUT_TT_PROJECT5(Tile_X5Y4_UO_OUT_TT_PROJECT5),
    .UO_OUT_TT_PROJECT6(Tile_X5Y4_UO_OUT_TT_PROJECT6),
    .UO_OUT_TT_PROJECT7(Tile_X5Y4_UO_OUT_TT_PROJECT7),
    .UIO_OUT_TT_PROJECT0(Tile_X5Y4_UIO_OUT_TT_PROJECT0),
    .UIO_OUT_TT_PROJECT1(Tile_X5Y4_UIO_OUT_TT_PROJECT1),
    .UIO_OUT_TT_PROJECT2(Tile_X5Y4_UIO_OUT_TT_PROJECT2),
    .UIO_OUT_TT_PROJECT3(Tile_X5Y4_UIO_OUT_TT_PROJECT3),
    .UIO_OUT_TT_PROJECT4(Tile_X5Y4_UIO_OUT_TT_PROJECT4),
    .UIO_OUT_TT_PROJECT5(Tile_X5Y4_UIO_OUT_TT_PROJECT5),
    .UIO_OUT_TT_PROJECT6(Tile_X5Y4_UIO_OUT_TT_PROJECT6),
    .UIO_OUT_TT_PROJECT7(Tile_X5Y4_UIO_OUT_TT_PROJECT7),
    .UIO_OE_TT_PROJECT0(Tile_X5Y4_UIO_OE_TT_PROJECT0),
    .UIO_OE_TT_PROJECT1(Tile_X5Y4_UIO_OE_TT_PROJECT1),
    .UIO_OE_TT_PROJECT2(Tile_X5Y4_UIO_OE_TT_PROJECT2),
    .UIO_OE_TT_PROJECT3(Tile_X5Y4_UIO_OE_TT_PROJECT3),
    .UIO_OE_TT_PROJECT4(Tile_X5Y4_UIO_OE_TT_PROJECT4),
    .UIO_OE_TT_PROJECT5(Tile_X5Y4_UIO_OE_TT_PROJECT5),
    .UIO_OE_TT_PROJECT6(Tile_X5Y4_UIO_OE_TT_PROJECT6),
    .UIO_OE_TT_PROJECT7(Tile_X5Y4_UIO_OE_TT_PROJECT7),
    .UI_IN_TT_PROJECT0(Tile_X5Y4_UI_IN_TT_PROJECT0),
    .UI_IN_TT_PROJECT1(Tile_X5Y4_UI_IN_TT_PROJECT1),
    .UI_IN_TT_PROJECT2(Tile_X5Y4_UI_IN_TT_PROJECT2),
    .UI_IN_TT_PROJECT3(Tile_X5Y4_UI_IN_TT_PROJECT3),
    .UI_IN_TT_PROJECT4(Tile_X5Y4_UI_IN_TT_PROJECT4),
    .UI_IN_TT_PROJECT5(Tile_X5Y4_UI_IN_TT_PROJECT5),
    .UI_IN_TT_PROJECT6(Tile_X5Y4_UI_IN_TT_PROJECT6),
    .UI_IN_TT_PROJECT7(Tile_X5Y4_UI_IN_TT_PROJECT7),
    .UIO_IN_TT_PROJECT0(Tile_X5Y4_UIO_IN_TT_PROJECT0),
    .UIO_IN_TT_PROJECT1(Tile_X5Y4_UIO_IN_TT_PROJECT1),
    .UIO_IN_TT_PROJECT2(Tile_X5Y4_UIO_IN_TT_PROJECT2),
    .UIO_IN_TT_PROJECT3(Tile_X5Y4_UIO_IN_TT_PROJECT3),
    .UIO_IN_TT_PROJECT4(Tile_X5Y4_UIO_IN_TT_PROJECT4),
    .UIO_IN_TT_PROJECT5(Tile_X5Y4_UIO_IN_TT_PROJECT5),
    .UIO_IN_TT_PROJECT6(Tile_X5Y4_UIO_IN_TT_PROJECT6),
    .UIO_IN_TT_PROJECT7(Tile_X5Y4_UIO_IN_TT_PROJECT7),
    .ENA_TT_PROJECT(Tile_X5Y4_ENA_TT_PROJECT),
    .CLK_TT_PROJECT(Tile_X5Y4_CLK_TT_PROJECT),
    .RST_N_TT_PROJECT(Tile_X5Y4_RST_N_TT_PROJECT),
    .Tile_X0Y0_UserCLKo(Tile_X5Y3_UserCLKo),
    .Tile_X0Y1_UserCLK(Tile_X5Y5_UserCLKo),
    .Tile_X0Y0_FrameData(Tile_X4Y3_FrameData_O),
    .Tile_X0Y0_FrameData_O(Tile_X5Y3_FrameData_O),
    .Tile_X0Y0_FrameStrobe_O(Tile_X5Y3_FrameStrobe_O),
    .Tile_X0Y1_FrameData(Tile_X4Y4_FrameData_O),
    .Tile_X0Y1_FrameData_O(Tile_X5Y4_FrameData_O),
    .Tile_X0Y1_FrameStrobe(Tile_X5Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_TT_IF
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y4_Emulate_Bitstream)
    )
`endif
    Tile_X0Y4_W_TT_IF
    (
    .N1END(Tile_X0Y5_N1BEG),
    .N2MID(Tile_X0Y5_N2BEG),
    .N2END(Tile_X0Y5_N2BEGb),
    .N4END(Tile_X0Y5_N4BEG),
    .S1END(Tile_X0Y3_S1BEG),
    .S2MID(Tile_X0Y3_S2BEG),
    .S2END(Tile_X0Y3_S2BEGb),
    .S4END(Tile_X0Y3_S4BEG),
    .W1END(Tile_X1Y4_W1BEG),
    .W2MID(Tile_X1Y4_W2BEG),
    .W2END(Tile_X1Y4_W2BEGb),
    .WW4END(Tile_X1Y4_WW4BEG),
    .W6END(Tile_X1Y4_W6BEG),
    .N1BEG(Tile_X0Y4_N1BEG),
    .N2BEG(Tile_X0Y4_N2BEG),
    .N2BEGb(Tile_X0Y4_N2BEGb),
    .N4BEG(Tile_X0Y4_N4BEG),
    .S1BEG(Tile_X0Y4_S1BEG),
    .S2BEG(Tile_X0Y4_S2BEG),
    .S2BEGb(Tile_X0Y4_S2BEGb),
    .S4BEG(Tile_X0Y4_S4BEG),
    .E1BEG(Tile_X0Y4_E1BEG),
    .E2BEG(Tile_X0Y4_E2BEG),
    .E2BEGb(Tile_X0Y4_E2BEGb),
    .EE4BEG(Tile_X0Y4_EE4BEG),
    .E6BEG(Tile_X0Y4_E6BEG),
    .UO_OUT_TT_PROJECT0(Tile_X0Y4_UO_OUT_TT_PROJECT0),
    .UO_OUT_TT_PROJECT1(Tile_X0Y4_UO_OUT_TT_PROJECT1),
    .UO_OUT_TT_PROJECT2(Tile_X0Y4_UO_OUT_TT_PROJECT2),
    .UO_OUT_TT_PROJECT3(Tile_X0Y4_UO_OUT_TT_PROJECT3),
    .UO_OUT_TT_PROJECT4(Tile_X0Y4_UO_OUT_TT_PROJECT4),
    .UO_OUT_TT_PROJECT5(Tile_X0Y4_UO_OUT_TT_PROJECT5),
    .UO_OUT_TT_PROJECT6(Tile_X0Y4_UO_OUT_TT_PROJECT6),
    .UO_OUT_TT_PROJECT7(Tile_X0Y4_UO_OUT_TT_PROJECT7),
    .UIO_OUT_TT_PROJECT0(Tile_X0Y4_UIO_OUT_TT_PROJECT0),
    .UIO_OUT_TT_PROJECT1(Tile_X0Y4_UIO_OUT_TT_PROJECT1),
    .UIO_OUT_TT_PROJECT2(Tile_X0Y4_UIO_OUT_TT_PROJECT2),
    .UIO_OUT_TT_PROJECT3(Tile_X0Y4_UIO_OUT_TT_PROJECT3),
    .UIO_OUT_TT_PROJECT4(Tile_X0Y4_UIO_OUT_TT_PROJECT4),
    .UIO_OUT_TT_PROJECT5(Tile_X0Y4_UIO_OUT_TT_PROJECT5),
    .UIO_OUT_TT_PROJECT6(Tile_X0Y4_UIO_OUT_TT_PROJECT6),
    .UIO_OUT_TT_PROJECT7(Tile_X0Y4_UIO_OUT_TT_PROJECT7),
    .UIO_OE_TT_PROJECT0(Tile_X0Y4_UIO_OE_TT_PROJECT0),
    .UIO_OE_TT_PROJECT1(Tile_X0Y4_UIO_OE_TT_PROJECT1),
    .UIO_OE_TT_PROJECT2(Tile_X0Y4_UIO_OE_TT_PROJECT2),
    .UIO_OE_TT_PROJECT3(Tile_X0Y4_UIO_OE_TT_PROJECT3),
    .UIO_OE_TT_PROJECT4(Tile_X0Y4_UIO_OE_TT_PROJECT4),
    .UIO_OE_TT_PROJECT5(Tile_X0Y4_UIO_OE_TT_PROJECT5),
    .UIO_OE_TT_PROJECT6(Tile_X0Y4_UIO_OE_TT_PROJECT6),
    .UIO_OE_TT_PROJECT7(Tile_X0Y4_UIO_OE_TT_PROJECT7),
    .UI_IN_TT_PROJECT0(Tile_X0Y4_UI_IN_TT_PROJECT0),
    .UI_IN_TT_PROJECT1(Tile_X0Y4_UI_IN_TT_PROJECT1),
    .UI_IN_TT_PROJECT2(Tile_X0Y4_UI_IN_TT_PROJECT2),
    .UI_IN_TT_PROJECT3(Tile_X0Y4_UI_IN_TT_PROJECT3),
    .UI_IN_TT_PROJECT4(Tile_X0Y4_UI_IN_TT_PROJECT4),
    .UI_IN_TT_PROJECT5(Tile_X0Y4_UI_IN_TT_PROJECT5),
    .UI_IN_TT_PROJECT6(Tile_X0Y4_UI_IN_TT_PROJECT6),
    .UI_IN_TT_PROJECT7(Tile_X0Y4_UI_IN_TT_PROJECT7),
    .UIO_IN_TT_PROJECT0(Tile_X0Y4_UIO_IN_TT_PROJECT0),
    .UIO_IN_TT_PROJECT1(Tile_X0Y4_UIO_IN_TT_PROJECT1),
    .UIO_IN_TT_PROJECT2(Tile_X0Y4_UIO_IN_TT_PROJECT2),
    .UIO_IN_TT_PROJECT3(Tile_X0Y4_UIO_IN_TT_PROJECT3),
    .UIO_IN_TT_PROJECT4(Tile_X0Y4_UIO_IN_TT_PROJECT4),
    .UIO_IN_TT_PROJECT5(Tile_X0Y4_UIO_IN_TT_PROJECT5),
    .UIO_IN_TT_PROJECT6(Tile_X0Y4_UIO_IN_TT_PROJECT6),
    .UIO_IN_TT_PROJECT7(Tile_X0Y4_UIO_IN_TT_PROJECT7),
    .ENA_TT_PROJECT(Tile_X0Y4_ENA_TT_PROJECT),
    .CLK_TT_PROJECT(Tile_X0Y4_CLK_TT_PROJECT),
    .RST_N_TT_PROJECT(Tile_X0Y4_RST_N_TT_PROJECT),
    .UserCLK(Tile_X0Y5_UserCLKo),
    .UserCLKo(Tile_X0Y4_UserCLKo),
    .FrameData(Row_Y4_FrameData),
    .FrameData_O(Tile_X0Y4_FrameData_O),
    .FrameStrobe(Tile_X0Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y4_Emulate_Bitstream)
    )
`endif
    Tile_X1Y4_LUT4AB
    (
    .N1END(Tile_X1Y5_N1BEG),
    .N2MID(Tile_X1Y5_N2BEG),
    .N2END(Tile_X1Y5_N2BEGb),
    .N4END(Tile_X1Y5_N4BEG),
    .NN4END(Tile_X1Y5_NN4BEG),
    .Ci(Tile_X1Y5_Co),
    .E1END(Tile_X0Y4_E1BEG),
    .E2MID(Tile_X0Y4_E2BEG),
    .E2END(Tile_X0Y4_E2BEGb),
    .EE4END(Tile_X0Y4_EE4BEG),
    .E6END(Tile_X0Y4_E6BEG),
    .S1END(Tile_X1Y3_S1BEG),
    .S2MID(Tile_X1Y3_S2BEG),
    .S2END(Tile_X1Y3_S2BEGb),
    .S4END(Tile_X1Y3_S4BEG),
    .SS4END(Tile_X1Y3_SS4BEG),
    .W1END(Tile_X2Y4_W1BEG),
    .W2MID(Tile_X2Y4_W2BEG),
    .W2END(Tile_X2Y4_W2BEGb),
    .WW4END(Tile_X2Y4_WW4BEG),
    .W6END(Tile_X2Y4_W6BEG),
    .N1BEG(Tile_X1Y4_N1BEG),
    .N2BEG(Tile_X1Y4_N2BEG),
    .N2BEGb(Tile_X1Y4_N2BEGb),
    .N4BEG(Tile_X1Y4_N4BEG),
    .NN4BEG(Tile_X1Y4_NN4BEG),
    .E1BEG(Tile_X1Y4_E1BEG),
    .E2BEG(Tile_X1Y4_E2BEG),
    .E2BEGb(Tile_X1Y4_E2BEGb),
    .EE4BEG(Tile_X1Y4_EE4BEG),
    .E6BEG(Tile_X1Y4_E6BEG),
    .S1BEG(Tile_X1Y4_S1BEG),
    .S2BEG(Tile_X1Y4_S2BEG),
    .S2BEGb(Tile_X1Y4_S2BEGb),
    .S4BEG(Tile_X1Y4_S4BEG),
    .SS4BEG(Tile_X1Y4_SS4BEG),
    .W1BEG(Tile_X1Y4_W1BEG),
    .W2BEG(Tile_X1Y4_W2BEG),
    .W2BEGb(Tile_X1Y4_W2BEGb),
    .WW4BEG(Tile_X1Y4_WW4BEG),
    .W6BEG(Tile_X1Y4_W6BEG),
    .Co(Tile_X1Y4_Co),
    .UserCLK(Tile_X1Y5_UserCLKo),
    .UserCLKo(Tile_X1Y4_UserCLKo),
    .FrameData(Tile_X0Y4_FrameData_O),
    .FrameData_O(Tile_X1Y4_FrameData_O),
    .FrameStrobe(Tile_X1Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y4_Emulate_Bitstream)
    )
`endif
    Tile_X2Y4_LUT4AB
    (
    .N1END(Tile_X2Y5_N1BEG),
    .N2MID(Tile_X2Y5_N2BEG),
    .N2END(Tile_X2Y5_N2BEGb),
    .N4END(Tile_X2Y5_N4BEG),
    .NN4END(Tile_X2Y5_NN4BEG),
    .Ci(Tile_X2Y5_Co),
    .E1END(Tile_X1Y4_E1BEG),
    .E2MID(Tile_X1Y4_E2BEG),
    .E2END(Tile_X1Y4_E2BEGb),
    .EE4END(Tile_X1Y4_EE4BEG),
    .E6END(Tile_X1Y4_E6BEG),
    .S1END(Tile_X2Y3_S1BEG),
    .S2MID(Tile_X2Y3_S2BEG),
    .S2END(Tile_X2Y3_S2BEGb),
    .S4END(Tile_X2Y3_S4BEG),
    .SS4END(Tile_X2Y3_SS4BEG),
    .W1END(Tile_X3Y4_W1BEG),
    .W2MID(Tile_X3Y4_W2BEG),
    .W2END(Tile_X3Y4_W2BEGb),
    .WW4END(Tile_X3Y4_WW4BEG),
    .W6END(Tile_X3Y4_W6BEG),
    .N1BEG(Tile_X2Y4_N1BEG),
    .N2BEG(Tile_X2Y4_N2BEG),
    .N2BEGb(Tile_X2Y4_N2BEGb),
    .N4BEG(Tile_X2Y4_N4BEG),
    .NN4BEG(Tile_X2Y4_NN4BEG),
    .E1BEG(Tile_X2Y4_E1BEG),
    .E2BEG(Tile_X2Y4_E2BEG),
    .E2BEGb(Tile_X2Y4_E2BEGb),
    .EE4BEG(Tile_X2Y4_EE4BEG),
    .E6BEG(Tile_X2Y4_E6BEG),
    .S1BEG(Tile_X2Y4_S1BEG),
    .S2BEG(Tile_X2Y4_S2BEG),
    .S2BEGb(Tile_X2Y4_S2BEGb),
    .S4BEG(Tile_X2Y4_S4BEG),
    .SS4BEG(Tile_X2Y4_SS4BEG),
    .W1BEG(Tile_X2Y4_W1BEG),
    .W2BEG(Tile_X2Y4_W2BEG),
    .W2BEGb(Tile_X2Y4_W2BEGb),
    .WW4BEG(Tile_X2Y4_WW4BEG),
    .W6BEG(Tile_X2Y4_W6BEG),
    .Co(Tile_X2Y4_Co),
    .UserCLK(Tile_X2Y5_UserCLKo),
    .UserCLKo(Tile_X2Y4_UserCLKo),
    .FrameData(Tile_X1Y4_FrameData_O),
    .FrameData_O(Tile_X2Y4_FrameData_O),
    .FrameStrobe(Tile_X2Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y4_Emulate_Bitstream)
    )
`endif
    Tile_X3Y4_LUT4AB
    (
    .N1END(Tile_X3Y5_N1BEG),
    .N2MID(Tile_X3Y5_N2BEG),
    .N2END(Tile_X3Y5_N2BEGb),
    .N4END(Tile_X3Y5_N4BEG),
    .NN4END(Tile_X3Y5_NN4BEG),
    .Ci(Tile_X3Y5_Co),
    .E1END(Tile_X2Y4_E1BEG),
    .E2MID(Tile_X2Y4_E2BEG),
    .E2END(Tile_X2Y4_E2BEGb),
    .EE4END(Tile_X2Y4_EE4BEG),
    .E6END(Tile_X2Y4_E6BEG),
    .S1END(Tile_X3Y3_S1BEG),
    .S2MID(Tile_X3Y3_S2BEG),
    .S2END(Tile_X3Y3_S2BEGb),
    .S4END(Tile_X3Y3_S4BEG),
    .SS4END(Tile_X3Y3_SS4BEG),
    .W1END(Tile_X4Y4_W1BEG),
    .W2MID(Tile_X4Y4_W2BEG),
    .W2END(Tile_X4Y4_W2BEGb),
    .WW4END(Tile_X4Y4_WW4BEG),
    .W6END(Tile_X4Y4_W6BEG),
    .N1BEG(Tile_X3Y4_N1BEG),
    .N2BEG(Tile_X3Y4_N2BEG),
    .N2BEGb(Tile_X3Y4_N2BEGb),
    .N4BEG(Tile_X3Y4_N4BEG),
    .NN4BEG(Tile_X3Y4_NN4BEG),
    .E1BEG(Tile_X3Y4_E1BEG),
    .E2BEG(Tile_X3Y4_E2BEG),
    .E2BEGb(Tile_X3Y4_E2BEGb),
    .EE4BEG(Tile_X3Y4_EE4BEG),
    .E6BEG(Tile_X3Y4_E6BEG),
    .S1BEG(Tile_X3Y4_S1BEG),
    .S2BEG(Tile_X3Y4_S2BEG),
    .S2BEGb(Tile_X3Y4_S2BEGb),
    .S4BEG(Tile_X3Y4_S4BEG),
    .SS4BEG(Tile_X3Y4_SS4BEG),
    .W1BEG(Tile_X3Y4_W1BEG),
    .W2BEG(Tile_X3Y4_W2BEG),
    .W2BEGb(Tile_X3Y4_W2BEGb),
    .WW4BEG(Tile_X3Y4_WW4BEG),
    .W6BEG(Tile_X3Y4_W6BEG),
    .Co(Tile_X3Y4_Co),
    .UserCLK(Tile_X3Y5_UserCLKo),
    .UserCLKo(Tile_X3Y4_UserCLKo),
    .FrameData(Tile_X2Y4_FrameData_O),
    .FrameData_O(Tile_X3Y4_FrameData_O),
    .FrameStrobe(Tile_X3Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y4_Emulate_Bitstream)
    )
`endif
    Tile_X4Y4_LUT4AB
    (
    .N1END(Tile_X4Y5_N1BEG),
    .N2MID(Tile_X4Y5_N2BEG),
    .N2END(Tile_X4Y5_N2BEGb),
    .N4END(Tile_X4Y5_N4BEG),
    .NN4END(Tile_X4Y5_NN4BEG),
    .Ci(Tile_X4Y5_Co),
    .E1END(Tile_X3Y4_E1BEG),
    .E2MID(Tile_X3Y4_E2BEG),
    .E2END(Tile_X3Y4_E2BEGb),
    .EE4END(Tile_X3Y4_EE4BEG),
    .E6END(Tile_X3Y4_E6BEG),
    .S1END(Tile_X4Y3_S1BEG),
    .S2MID(Tile_X4Y3_S2BEG),
    .S2END(Tile_X4Y3_S2BEGb),
    .S4END(Tile_X4Y3_S4BEG),
    .SS4END(Tile_X4Y3_SS4BEG),
    .W1END(Tile_X5Y4_W1BEG),
    .W2MID(Tile_X5Y4_W2BEG),
    .W2END(Tile_X5Y4_W2BEGb),
    .WW4END(Tile_X5Y4_WW4BEG),
    .W6END(Tile_X5Y4_W6BEG),
    .N1BEG(Tile_X4Y4_N1BEG),
    .N2BEG(Tile_X4Y4_N2BEG),
    .N2BEGb(Tile_X4Y4_N2BEGb),
    .N4BEG(Tile_X4Y4_N4BEG),
    .NN4BEG(Tile_X4Y4_NN4BEG),
    .E1BEG(Tile_X4Y4_E1BEG),
    .E2BEG(Tile_X4Y4_E2BEG),
    .E2BEGb(Tile_X4Y4_E2BEGb),
    .EE4BEG(Tile_X4Y4_EE4BEG),
    .E6BEG(Tile_X4Y4_E6BEG),
    .S1BEG(Tile_X4Y4_S1BEG),
    .S2BEG(Tile_X4Y4_S2BEG),
    .S2BEGb(Tile_X4Y4_S2BEGb),
    .S4BEG(Tile_X4Y4_S4BEG),
    .SS4BEG(Tile_X4Y4_SS4BEG),
    .W1BEG(Tile_X4Y4_W1BEG),
    .W2BEG(Tile_X4Y4_W2BEG),
    .W2BEGb(Tile_X4Y4_W2BEGb),
    .WW4BEG(Tile_X4Y4_WW4BEG),
    .W6BEG(Tile_X4Y4_W6BEG),
    .Co(Tile_X4Y4_Co),
    .UserCLK(Tile_X4Y5_UserCLKo),
    .UserCLKo(Tile_X4Y4_UserCLKo),
    .FrameData(Tile_X3Y4_FrameData_O),
    .FrameData_O(Tile_X4Y4_FrameData_O),
    .FrameStrobe(Tile_X4Y5_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y4_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_TT_IF
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y5_Emulate_Bitstream)
    )
`endif
    Tile_X0Y5_W_TT_IF
    (
    .N1END(Tile_X0Y6_N1BEG),
    .N2MID(Tile_X0Y6_N2BEG),
    .N2END(Tile_X0Y6_N2BEGb),
    .N4END(Tile_X0Y6_N4BEG),
    .S1END(Tile_X0Y4_S1BEG),
    .S2MID(Tile_X0Y4_S2BEG),
    .S2END(Tile_X0Y4_S2BEGb),
    .S4END(Tile_X0Y4_S4BEG),
    .W1END(Tile_X1Y5_W1BEG),
    .W2MID(Tile_X1Y5_W2BEG),
    .W2END(Tile_X1Y5_W2BEGb),
    .WW4END(Tile_X1Y5_WW4BEG),
    .W6END(Tile_X1Y5_W6BEG),
    .N1BEG(Tile_X0Y5_N1BEG),
    .N2BEG(Tile_X0Y5_N2BEG),
    .N2BEGb(Tile_X0Y5_N2BEGb),
    .N4BEG(Tile_X0Y5_N4BEG),
    .S1BEG(Tile_X0Y5_S1BEG),
    .S2BEG(Tile_X0Y5_S2BEG),
    .S2BEGb(Tile_X0Y5_S2BEGb),
    .S4BEG(Tile_X0Y5_S4BEG),
    .E1BEG(Tile_X0Y5_E1BEG),
    .E2BEG(Tile_X0Y5_E2BEG),
    .E2BEGb(Tile_X0Y5_E2BEGb),
    .EE4BEG(Tile_X0Y5_EE4BEG),
    .E6BEG(Tile_X0Y5_E6BEG),
    .UO_OUT_TT_PROJECT0(Tile_X0Y5_UO_OUT_TT_PROJECT0),
    .UO_OUT_TT_PROJECT1(Tile_X0Y5_UO_OUT_TT_PROJECT1),
    .UO_OUT_TT_PROJECT2(Tile_X0Y5_UO_OUT_TT_PROJECT2),
    .UO_OUT_TT_PROJECT3(Tile_X0Y5_UO_OUT_TT_PROJECT3),
    .UO_OUT_TT_PROJECT4(Tile_X0Y5_UO_OUT_TT_PROJECT4),
    .UO_OUT_TT_PROJECT5(Tile_X0Y5_UO_OUT_TT_PROJECT5),
    .UO_OUT_TT_PROJECT6(Tile_X0Y5_UO_OUT_TT_PROJECT6),
    .UO_OUT_TT_PROJECT7(Tile_X0Y5_UO_OUT_TT_PROJECT7),
    .UIO_OUT_TT_PROJECT0(Tile_X0Y5_UIO_OUT_TT_PROJECT0),
    .UIO_OUT_TT_PROJECT1(Tile_X0Y5_UIO_OUT_TT_PROJECT1),
    .UIO_OUT_TT_PROJECT2(Tile_X0Y5_UIO_OUT_TT_PROJECT2),
    .UIO_OUT_TT_PROJECT3(Tile_X0Y5_UIO_OUT_TT_PROJECT3),
    .UIO_OUT_TT_PROJECT4(Tile_X0Y5_UIO_OUT_TT_PROJECT4),
    .UIO_OUT_TT_PROJECT5(Tile_X0Y5_UIO_OUT_TT_PROJECT5),
    .UIO_OUT_TT_PROJECT6(Tile_X0Y5_UIO_OUT_TT_PROJECT6),
    .UIO_OUT_TT_PROJECT7(Tile_X0Y5_UIO_OUT_TT_PROJECT7),
    .UIO_OE_TT_PROJECT0(Tile_X0Y5_UIO_OE_TT_PROJECT0),
    .UIO_OE_TT_PROJECT1(Tile_X0Y5_UIO_OE_TT_PROJECT1),
    .UIO_OE_TT_PROJECT2(Tile_X0Y5_UIO_OE_TT_PROJECT2),
    .UIO_OE_TT_PROJECT3(Tile_X0Y5_UIO_OE_TT_PROJECT3),
    .UIO_OE_TT_PROJECT4(Tile_X0Y5_UIO_OE_TT_PROJECT4),
    .UIO_OE_TT_PROJECT5(Tile_X0Y5_UIO_OE_TT_PROJECT5),
    .UIO_OE_TT_PROJECT6(Tile_X0Y5_UIO_OE_TT_PROJECT6),
    .UIO_OE_TT_PROJECT7(Tile_X0Y5_UIO_OE_TT_PROJECT7),
    .UI_IN_TT_PROJECT0(Tile_X0Y5_UI_IN_TT_PROJECT0),
    .UI_IN_TT_PROJECT1(Tile_X0Y5_UI_IN_TT_PROJECT1),
    .UI_IN_TT_PROJECT2(Tile_X0Y5_UI_IN_TT_PROJECT2),
    .UI_IN_TT_PROJECT3(Tile_X0Y5_UI_IN_TT_PROJECT3),
    .UI_IN_TT_PROJECT4(Tile_X0Y5_UI_IN_TT_PROJECT4),
    .UI_IN_TT_PROJECT5(Tile_X0Y5_UI_IN_TT_PROJECT5),
    .UI_IN_TT_PROJECT6(Tile_X0Y5_UI_IN_TT_PROJECT6),
    .UI_IN_TT_PROJECT7(Tile_X0Y5_UI_IN_TT_PROJECT7),
    .UIO_IN_TT_PROJECT0(Tile_X0Y5_UIO_IN_TT_PROJECT0),
    .UIO_IN_TT_PROJECT1(Tile_X0Y5_UIO_IN_TT_PROJECT1),
    .UIO_IN_TT_PROJECT2(Tile_X0Y5_UIO_IN_TT_PROJECT2),
    .UIO_IN_TT_PROJECT3(Tile_X0Y5_UIO_IN_TT_PROJECT3),
    .UIO_IN_TT_PROJECT4(Tile_X0Y5_UIO_IN_TT_PROJECT4),
    .UIO_IN_TT_PROJECT5(Tile_X0Y5_UIO_IN_TT_PROJECT5),
    .UIO_IN_TT_PROJECT6(Tile_X0Y5_UIO_IN_TT_PROJECT6),
    .UIO_IN_TT_PROJECT7(Tile_X0Y5_UIO_IN_TT_PROJECT7),
    .ENA_TT_PROJECT(Tile_X0Y5_ENA_TT_PROJECT),
    .CLK_TT_PROJECT(Tile_X0Y5_CLK_TT_PROJECT),
    .RST_N_TT_PROJECT(Tile_X0Y5_RST_N_TT_PROJECT),
    .UserCLK(Tile_X0Y6_UserCLKo),
    .UserCLKo(Tile_X0Y5_UserCLKo),
    .FrameData(Row_Y5_FrameData),
    .FrameData_O(Tile_X0Y5_FrameData_O),
    .FrameStrobe(Tile_X0Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y5_Emulate_Bitstream)
    )
`endif
    Tile_X1Y5_LUT4AB
    (
    .N1END(Tile_X1Y6_N1BEG),
    .N2MID(Tile_X1Y6_N2BEG),
    .N2END(Tile_X1Y6_N2BEGb),
    .N4END(Tile_X1Y6_N4BEG),
    .NN4END(Tile_X1Y6_NN4BEG),
    .Ci(Tile_X1Y6_Co),
    .E1END(Tile_X0Y5_E1BEG),
    .E2MID(Tile_X0Y5_E2BEG),
    .E2END(Tile_X0Y5_E2BEGb),
    .EE4END(Tile_X0Y5_EE4BEG),
    .E6END(Tile_X0Y5_E6BEG),
    .S1END(Tile_X1Y4_S1BEG),
    .S2MID(Tile_X1Y4_S2BEG),
    .S2END(Tile_X1Y4_S2BEGb),
    .S4END(Tile_X1Y4_S4BEG),
    .SS4END(Tile_X1Y4_SS4BEG),
    .W1END(Tile_X2Y5_W1BEG),
    .W2MID(Tile_X2Y5_W2BEG),
    .W2END(Tile_X2Y5_W2BEGb),
    .WW4END(Tile_X2Y5_WW4BEG),
    .W6END(Tile_X2Y5_W6BEG),
    .N1BEG(Tile_X1Y5_N1BEG),
    .N2BEG(Tile_X1Y5_N2BEG),
    .N2BEGb(Tile_X1Y5_N2BEGb),
    .N4BEG(Tile_X1Y5_N4BEG),
    .NN4BEG(Tile_X1Y5_NN4BEG),
    .E1BEG(Tile_X1Y5_E1BEG),
    .E2BEG(Tile_X1Y5_E2BEG),
    .E2BEGb(Tile_X1Y5_E2BEGb),
    .EE4BEG(Tile_X1Y5_EE4BEG),
    .E6BEG(Tile_X1Y5_E6BEG),
    .S1BEG(Tile_X1Y5_S1BEG),
    .S2BEG(Tile_X1Y5_S2BEG),
    .S2BEGb(Tile_X1Y5_S2BEGb),
    .S4BEG(Tile_X1Y5_S4BEG),
    .SS4BEG(Tile_X1Y5_SS4BEG),
    .W1BEG(Tile_X1Y5_W1BEG),
    .W2BEG(Tile_X1Y5_W2BEG),
    .W2BEGb(Tile_X1Y5_W2BEGb),
    .WW4BEG(Tile_X1Y5_WW4BEG),
    .W6BEG(Tile_X1Y5_W6BEG),
    .Co(Tile_X1Y5_Co),
    .UserCLK(Tile_X1Y6_UserCLKo),
    .UserCLKo(Tile_X1Y5_UserCLKo),
    .FrameData(Tile_X0Y5_FrameData_O),
    .FrameData_O(Tile_X1Y5_FrameData_O),
    .FrameStrobe(Tile_X1Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y5_Emulate_Bitstream)
    )
`endif
    Tile_X2Y5_LUT4AB
    (
    .N1END(Tile_X2Y6_N1BEG),
    .N2MID(Tile_X2Y6_N2BEG),
    .N2END(Tile_X2Y6_N2BEGb),
    .N4END(Tile_X2Y6_N4BEG),
    .NN4END(Tile_X2Y6_NN4BEG),
    .Ci(Tile_X2Y6_Co),
    .E1END(Tile_X1Y5_E1BEG),
    .E2MID(Tile_X1Y5_E2BEG),
    .E2END(Tile_X1Y5_E2BEGb),
    .EE4END(Tile_X1Y5_EE4BEG),
    .E6END(Tile_X1Y5_E6BEG),
    .S1END(Tile_X2Y4_S1BEG),
    .S2MID(Tile_X2Y4_S2BEG),
    .S2END(Tile_X2Y4_S2BEGb),
    .S4END(Tile_X2Y4_S4BEG),
    .SS4END(Tile_X2Y4_SS4BEG),
    .W1END(Tile_X3Y5_W1BEG),
    .W2MID(Tile_X3Y5_W2BEG),
    .W2END(Tile_X3Y5_W2BEGb),
    .WW4END(Tile_X3Y5_WW4BEG),
    .W6END(Tile_X3Y5_W6BEG),
    .N1BEG(Tile_X2Y5_N1BEG),
    .N2BEG(Tile_X2Y5_N2BEG),
    .N2BEGb(Tile_X2Y5_N2BEGb),
    .N4BEG(Tile_X2Y5_N4BEG),
    .NN4BEG(Tile_X2Y5_NN4BEG),
    .E1BEG(Tile_X2Y5_E1BEG),
    .E2BEG(Tile_X2Y5_E2BEG),
    .E2BEGb(Tile_X2Y5_E2BEGb),
    .EE4BEG(Tile_X2Y5_EE4BEG),
    .E6BEG(Tile_X2Y5_E6BEG),
    .S1BEG(Tile_X2Y5_S1BEG),
    .S2BEG(Tile_X2Y5_S2BEG),
    .S2BEGb(Tile_X2Y5_S2BEGb),
    .S4BEG(Tile_X2Y5_S4BEG),
    .SS4BEG(Tile_X2Y5_SS4BEG),
    .W1BEG(Tile_X2Y5_W1BEG),
    .W2BEG(Tile_X2Y5_W2BEG),
    .W2BEGb(Tile_X2Y5_W2BEGb),
    .WW4BEG(Tile_X2Y5_WW4BEG),
    .W6BEG(Tile_X2Y5_W6BEG),
    .Co(Tile_X2Y5_Co),
    .UserCLK(Tile_X2Y6_UserCLKo),
    .UserCLKo(Tile_X2Y5_UserCLKo),
    .FrameData(Tile_X1Y5_FrameData_O),
    .FrameData_O(Tile_X2Y5_FrameData_O),
    .FrameStrobe(Tile_X2Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y5_Emulate_Bitstream)
    )
`endif
    Tile_X3Y5_LUT4AB
    (
    .N1END(Tile_X3Y6_N1BEG),
    .N2MID(Tile_X3Y6_N2BEG),
    .N2END(Tile_X3Y6_N2BEGb),
    .N4END(Tile_X3Y6_N4BEG),
    .NN4END(Tile_X3Y6_NN4BEG),
    .Ci(Tile_X3Y6_Co),
    .E1END(Tile_X2Y5_E1BEG),
    .E2MID(Tile_X2Y5_E2BEG),
    .E2END(Tile_X2Y5_E2BEGb),
    .EE4END(Tile_X2Y5_EE4BEG),
    .E6END(Tile_X2Y5_E6BEG),
    .S1END(Tile_X3Y4_S1BEG),
    .S2MID(Tile_X3Y4_S2BEG),
    .S2END(Tile_X3Y4_S2BEGb),
    .S4END(Tile_X3Y4_S4BEG),
    .SS4END(Tile_X3Y4_SS4BEG),
    .W1END(Tile_X4Y5_W1BEG),
    .W2MID(Tile_X4Y5_W2BEG),
    .W2END(Tile_X4Y5_W2BEGb),
    .WW4END(Tile_X4Y5_WW4BEG),
    .W6END(Tile_X4Y5_W6BEG),
    .N1BEG(Tile_X3Y5_N1BEG),
    .N2BEG(Tile_X3Y5_N2BEG),
    .N2BEGb(Tile_X3Y5_N2BEGb),
    .N4BEG(Tile_X3Y5_N4BEG),
    .NN4BEG(Tile_X3Y5_NN4BEG),
    .E1BEG(Tile_X3Y5_E1BEG),
    .E2BEG(Tile_X3Y5_E2BEG),
    .E2BEGb(Tile_X3Y5_E2BEGb),
    .EE4BEG(Tile_X3Y5_EE4BEG),
    .E6BEG(Tile_X3Y5_E6BEG),
    .S1BEG(Tile_X3Y5_S1BEG),
    .S2BEG(Tile_X3Y5_S2BEG),
    .S2BEGb(Tile_X3Y5_S2BEGb),
    .S4BEG(Tile_X3Y5_S4BEG),
    .SS4BEG(Tile_X3Y5_SS4BEG),
    .W1BEG(Tile_X3Y5_W1BEG),
    .W2BEG(Tile_X3Y5_W2BEG),
    .W2BEGb(Tile_X3Y5_W2BEGb),
    .WW4BEG(Tile_X3Y5_WW4BEG),
    .W6BEG(Tile_X3Y5_W6BEG),
    .Co(Tile_X3Y5_Co),
    .UserCLK(Tile_X3Y6_UserCLKo),
    .UserCLKo(Tile_X3Y5_UserCLKo),
    .FrameData(Tile_X2Y5_FrameData_O),
    .FrameData_O(Tile_X3Y5_FrameData_O),
    .FrameStrobe(Tile_X3Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y5_Emulate_Bitstream)
    )
`endif
    Tile_X4Y5_LUT4AB
    (
    .N1END(Tile_X4Y6_N1BEG),
    .N2MID(Tile_X4Y6_N2BEG),
    .N2END(Tile_X4Y6_N2BEGb),
    .N4END(Tile_X4Y6_N4BEG),
    .NN4END(Tile_X4Y6_NN4BEG),
    .Ci(Tile_X4Y6_Co),
    .E1END(Tile_X3Y5_E1BEG),
    .E2MID(Tile_X3Y5_E2BEG),
    .E2END(Tile_X3Y5_E2BEGb),
    .EE4END(Tile_X3Y5_EE4BEG),
    .E6END(Tile_X3Y5_E6BEG),
    .S1END(Tile_X4Y4_S1BEG),
    .S2MID(Tile_X4Y4_S2BEG),
    .S2END(Tile_X4Y4_S2BEGb),
    .S4END(Tile_X4Y4_S4BEG),
    .SS4END(Tile_X4Y4_SS4BEG),
    .W1END(Tile_X5Y5_W1BEG),
    .W2MID(Tile_X5Y5_W2BEG),
    .W2END(Tile_X5Y5_W2BEGb),
    .WW4END(Tile_X5Y5_WW4BEG),
    .W6END(Tile_X5Y5_W6BEG),
    .N1BEG(Tile_X4Y5_N1BEG),
    .N2BEG(Tile_X4Y5_N2BEG),
    .N2BEGb(Tile_X4Y5_N2BEGb),
    .N4BEG(Tile_X4Y5_N4BEG),
    .NN4BEG(Tile_X4Y5_NN4BEG),
    .E1BEG(Tile_X4Y5_E1BEG),
    .E2BEG(Tile_X4Y5_E2BEG),
    .E2BEGb(Tile_X4Y5_E2BEGb),
    .EE4BEG(Tile_X4Y5_EE4BEG),
    .E6BEG(Tile_X4Y5_E6BEG),
    .S1BEG(Tile_X4Y5_S1BEG),
    .S2BEG(Tile_X4Y5_S2BEG),
    .S2BEGb(Tile_X4Y5_S2BEGb),
    .S4BEG(Tile_X4Y5_S4BEG),
    .SS4BEG(Tile_X4Y5_SS4BEG),
    .W1BEG(Tile_X4Y5_W1BEG),
    .W2BEG(Tile_X4Y5_W2BEG),
    .W2BEGb(Tile_X4Y5_W2BEGb),
    .WW4BEG(Tile_X4Y5_WW4BEG),
    .W6BEG(Tile_X4Y5_W6BEG),
    .Co(Tile_X4Y5_Co),
    .UserCLK(Tile_X4Y6_UserCLKo),
    .UserCLKo(Tile_X4Y5_UserCLKo),
    .FrameData(Tile_X3Y5_FrameData_O),
    .FrameData_O(Tile_X4Y5_FrameData_O),
    .FrameStrobe(Tile_X4Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
E_TT_IF
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y5_Emulate_Bitstream)
    )
`endif
    Tile_X5Y5_E_TT_IF
    (
    .N1END(Tile_X5Y6_N1BEG),
    .N2MID(Tile_X5Y6_N2BEG),
    .N2END(Tile_X5Y6_N2BEGb),
    .N4END(Tile_X5Y6_N4BEG),
    .E1END(Tile_X4Y5_E1BEG),
    .E2MID(Tile_X4Y5_E2BEG),
    .E2END(Tile_X4Y5_E2BEGb),
    .EE4END(Tile_X4Y5_EE4BEG),
    .E6END(Tile_X4Y5_E6BEG),
    .S1END(Tile_X5Y4_S1BEG),
    .S2MID(Tile_X5Y4_S2BEG),
    .S2END(Tile_X5Y4_S2BEGb),
    .S4END(Tile_X5Y4_S4BEG),
    .N1BEG(Tile_X5Y5_N1BEG),
    .N2BEG(Tile_X5Y5_N2BEG),
    .N2BEGb(Tile_X5Y5_N2BEGb),
    .N4BEG(Tile_X5Y5_N4BEG),
    .S1BEG(Tile_X5Y5_S1BEG),
    .S2BEG(Tile_X5Y5_S2BEG),
    .S2BEGb(Tile_X5Y5_S2BEGb),
    .S4BEG(Tile_X5Y5_S4BEG),
    .W1BEG(Tile_X5Y5_W1BEG),
    .W2BEG(Tile_X5Y5_W2BEG),
    .W2BEGb(Tile_X5Y5_W2BEGb),
    .WW4BEG(Tile_X5Y5_WW4BEG),
    .W6BEG(Tile_X5Y5_W6BEG),
    .UO_OUT_TT_PROJECT0(Tile_X5Y5_UO_OUT_TT_PROJECT0),
    .UO_OUT_TT_PROJECT1(Tile_X5Y5_UO_OUT_TT_PROJECT1),
    .UO_OUT_TT_PROJECT2(Tile_X5Y5_UO_OUT_TT_PROJECT2),
    .UO_OUT_TT_PROJECT3(Tile_X5Y5_UO_OUT_TT_PROJECT3),
    .UO_OUT_TT_PROJECT4(Tile_X5Y5_UO_OUT_TT_PROJECT4),
    .UO_OUT_TT_PROJECT5(Tile_X5Y5_UO_OUT_TT_PROJECT5),
    .UO_OUT_TT_PROJECT6(Tile_X5Y5_UO_OUT_TT_PROJECT6),
    .UO_OUT_TT_PROJECT7(Tile_X5Y5_UO_OUT_TT_PROJECT7),
    .UIO_OUT_TT_PROJECT0(Tile_X5Y5_UIO_OUT_TT_PROJECT0),
    .UIO_OUT_TT_PROJECT1(Tile_X5Y5_UIO_OUT_TT_PROJECT1),
    .UIO_OUT_TT_PROJECT2(Tile_X5Y5_UIO_OUT_TT_PROJECT2),
    .UIO_OUT_TT_PROJECT3(Tile_X5Y5_UIO_OUT_TT_PROJECT3),
    .UIO_OUT_TT_PROJECT4(Tile_X5Y5_UIO_OUT_TT_PROJECT4),
    .UIO_OUT_TT_PROJECT5(Tile_X5Y5_UIO_OUT_TT_PROJECT5),
    .UIO_OUT_TT_PROJECT6(Tile_X5Y5_UIO_OUT_TT_PROJECT6),
    .UIO_OUT_TT_PROJECT7(Tile_X5Y5_UIO_OUT_TT_PROJECT7),
    .UIO_OE_TT_PROJECT0(Tile_X5Y5_UIO_OE_TT_PROJECT0),
    .UIO_OE_TT_PROJECT1(Tile_X5Y5_UIO_OE_TT_PROJECT1),
    .UIO_OE_TT_PROJECT2(Tile_X5Y5_UIO_OE_TT_PROJECT2),
    .UIO_OE_TT_PROJECT3(Tile_X5Y5_UIO_OE_TT_PROJECT3),
    .UIO_OE_TT_PROJECT4(Tile_X5Y5_UIO_OE_TT_PROJECT4),
    .UIO_OE_TT_PROJECT5(Tile_X5Y5_UIO_OE_TT_PROJECT5),
    .UIO_OE_TT_PROJECT6(Tile_X5Y5_UIO_OE_TT_PROJECT6),
    .UIO_OE_TT_PROJECT7(Tile_X5Y5_UIO_OE_TT_PROJECT7),
    .UI_IN_TT_PROJECT0(Tile_X5Y5_UI_IN_TT_PROJECT0),
    .UI_IN_TT_PROJECT1(Tile_X5Y5_UI_IN_TT_PROJECT1),
    .UI_IN_TT_PROJECT2(Tile_X5Y5_UI_IN_TT_PROJECT2),
    .UI_IN_TT_PROJECT3(Tile_X5Y5_UI_IN_TT_PROJECT3),
    .UI_IN_TT_PROJECT4(Tile_X5Y5_UI_IN_TT_PROJECT4),
    .UI_IN_TT_PROJECT5(Tile_X5Y5_UI_IN_TT_PROJECT5),
    .UI_IN_TT_PROJECT6(Tile_X5Y5_UI_IN_TT_PROJECT6),
    .UI_IN_TT_PROJECT7(Tile_X5Y5_UI_IN_TT_PROJECT7),
    .UIO_IN_TT_PROJECT0(Tile_X5Y5_UIO_IN_TT_PROJECT0),
    .UIO_IN_TT_PROJECT1(Tile_X5Y5_UIO_IN_TT_PROJECT1),
    .UIO_IN_TT_PROJECT2(Tile_X5Y5_UIO_IN_TT_PROJECT2),
    .UIO_IN_TT_PROJECT3(Tile_X5Y5_UIO_IN_TT_PROJECT3),
    .UIO_IN_TT_PROJECT4(Tile_X5Y5_UIO_IN_TT_PROJECT4),
    .UIO_IN_TT_PROJECT5(Tile_X5Y5_UIO_IN_TT_PROJECT5),
    .UIO_IN_TT_PROJECT6(Tile_X5Y5_UIO_IN_TT_PROJECT6),
    .UIO_IN_TT_PROJECT7(Tile_X5Y5_UIO_IN_TT_PROJECT7),
    .ENA_TT_PROJECT(Tile_X5Y5_ENA_TT_PROJECT),
    .CLK_TT_PROJECT(Tile_X5Y5_CLK_TT_PROJECT),
    .RST_N_TT_PROJECT(Tile_X5Y5_RST_N_TT_PROJECT),
    .UserCLK(Tile_X5Y6_UserCLKo),
    .UserCLKo(Tile_X5Y5_UserCLKo),
    .FrameData(Tile_X4Y5_FrameData_O),
    .FrameData_O(Tile_X5Y5_FrameData_O),
    .FrameStrobe(Tile_X5Y6_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y5_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_TT_IF
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y6_Emulate_Bitstream)
    )
`endif
    Tile_X0Y6_W_TT_IF
    (
    .N1END(Tile_X0Y7_N1BEG),
    .N2MID(Tile_X0Y7_N2BEG),
    .N2END(Tile_X0Y7_N2BEGb),
    .N4END(Tile_X0Y7_N4BEG),
    .S1END(Tile_X0Y5_S1BEG),
    .S2MID(Tile_X0Y5_S2BEG),
    .S2END(Tile_X0Y5_S2BEGb),
    .S4END(Tile_X0Y5_S4BEG),
    .W1END(Tile_X1Y6_W1BEG),
    .W2MID(Tile_X1Y6_W2BEG),
    .W2END(Tile_X1Y6_W2BEGb),
    .WW4END(Tile_X1Y6_WW4BEG),
    .W6END(Tile_X1Y6_W6BEG),
    .N1BEG(Tile_X0Y6_N1BEG),
    .N2BEG(Tile_X0Y6_N2BEG),
    .N2BEGb(Tile_X0Y6_N2BEGb),
    .N4BEG(Tile_X0Y6_N4BEG),
    .S1BEG(Tile_X0Y6_S1BEG),
    .S2BEG(Tile_X0Y6_S2BEG),
    .S2BEGb(Tile_X0Y6_S2BEGb),
    .S4BEG(Tile_X0Y6_S4BEG),
    .E1BEG(Tile_X0Y6_E1BEG),
    .E2BEG(Tile_X0Y6_E2BEG),
    .E2BEGb(Tile_X0Y6_E2BEGb),
    .EE4BEG(Tile_X0Y6_EE4BEG),
    .E6BEG(Tile_X0Y6_E6BEG),
    .UO_OUT_TT_PROJECT0(Tile_X0Y6_UO_OUT_TT_PROJECT0),
    .UO_OUT_TT_PROJECT1(Tile_X0Y6_UO_OUT_TT_PROJECT1),
    .UO_OUT_TT_PROJECT2(Tile_X0Y6_UO_OUT_TT_PROJECT2),
    .UO_OUT_TT_PROJECT3(Tile_X0Y6_UO_OUT_TT_PROJECT3),
    .UO_OUT_TT_PROJECT4(Tile_X0Y6_UO_OUT_TT_PROJECT4),
    .UO_OUT_TT_PROJECT5(Tile_X0Y6_UO_OUT_TT_PROJECT5),
    .UO_OUT_TT_PROJECT6(Tile_X0Y6_UO_OUT_TT_PROJECT6),
    .UO_OUT_TT_PROJECT7(Tile_X0Y6_UO_OUT_TT_PROJECT7),
    .UIO_OUT_TT_PROJECT0(Tile_X0Y6_UIO_OUT_TT_PROJECT0),
    .UIO_OUT_TT_PROJECT1(Tile_X0Y6_UIO_OUT_TT_PROJECT1),
    .UIO_OUT_TT_PROJECT2(Tile_X0Y6_UIO_OUT_TT_PROJECT2),
    .UIO_OUT_TT_PROJECT3(Tile_X0Y6_UIO_OUT_TT_PROJECT3),
    .UIO_OUT_TT_PROJECT4(Tile_X0Y6_UIO_OUT_TT_PROJECT4),
    .UIO_OUT_TT_PROJECT5(Tile_X0Y6_UIO_OUT_TT_PROJECT5),
    .UIO_OUT_TT_PROJECT6(Tile_X0Y6_UIO_OUT_TT_PROJECT6),
    .UIO_OUT_TT_PROJECT7(Tile_X0Y6_UIO_OUT_TT_PROJECT7),
    .UIO_OE_TT_PROJECT0(Tile_X0Y6_UIO_OE_TT_PROJECT0),
    .UIO_OE_TT_PROJECT1(Tile_X0Y6_UIO_OE_TT_PROJECT1),
    .UIO_OE_TT_PROJECT2(Tile_X0Y6_UIO_OE_TT_PROJECT2),
    .UIO_OE_TT_PROJECT3(Tile_X0Y6_UIO_OE_TT_PROJECT3),
    .UIO_OE_TT_PROJECT4(Tile_X0Y6_UIO_OE_TT_PROJECT4),
    .UIO_OE_TT_PROJECT5(Tile_X0Y6_UIO_OE_TT_PROJECT5),
    .UIO_OE_TT_PROJECT6(Tile_X0Y6_UIO_OE_TT_PROJECT6),
    .UIO_OE_TT_PROJECT7(Tile_X0Y6_UIO_OE_TT_PROJECT7),
    .UI_IN_TT_PROJECT0(Tile_X0Y6_UI_IN_TT_PROJECT0),
    .UI_IN_TT_PROJECT1(Tile_X0Y6_UI_IN_TT_PROJECT1),
    .UI_IN_TT_PROJECT2(Tile_X0Y6_UI_IN_TT_PROJECT2),
    .UI_IN_TT_PROJECT3(Tile_X0Y6_UI_IN_TT_PROJECT3),
    .UI_IN_TT_PROJECT4(Tile_X0Y6_UI_IN_TT_PROJECT4),
    .UI_IN_TT_PROJECT5(Tile_X0Y6_UI_IN_TT_PROJECT5),
    .UI_IN_TT_PROJECT6(Tile_X0Y6_UI_IN_TT_PROJECT6),
    .UI_IN_TT_PROJECT7(Tile_X0Y6_UI_IN_TT_PROJECT7),
    .UIO_IN_TT_PROJECT0(Tile_X0Y6_UIO_IN_TT_PROJECT0),
    .UIO_IN_TT_PROJECT1(Tile_X0Y6_UIO_IN_TT_PROJECT1),
    .UIO_IN_TT_PROJECT2(Tile_X0Y6_UIO_IN_TT_PROJECT2),
    .UIO_IN_TT_PROJECT3(Tile_X0Y6_UIO_IN_TT_PROJECT3),
    .UIO_IN_TT_PROJECT4(Tile_X0Y6_UIO_IN_TT_PROJECT4),
    .UIO_IN_TT_PROJECT5(Tile_X0Y6_UIO_IN_TT_PROJECT5),
    .UIO_IN_TT_PROJECT6(Tile_X0Y6_UIO_IN_TT_PROJECT6),
    .UIO_IN_TT_PROJECT7(Tile_X0Y6_UIO_IN_TT_PROJECT7),
    .ENA_TT_PROJECT(Tile_X0Y6_ENA_TT_PROJECT),
    .CLK_TT_PROJECT(Tile_X0Y6_CLK_TT_PROJECT),
    .RST_N_TT_PROJECT(Tile_X0Y6_RST_N_TT_PROJECT),
    .UserCLK(Tile_X0Y7_UserCLKo),
    .UserCLKo(Tile_X0Y6_UserCLKo),
    .FrameData(Row_Y6_FrameData),
    .FrameData_O(Tile_X0Y6_FrameData_O),
    .FrameStrobe(Tile_X0Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y6_Emulate_Bitstream)
    )
`endif
    Tile_X1Y6_LUT4AB
    (
    .N1END(Tile_X1Y7_N1BEG),
    .N2MID(Tile_X1Y7_N2BEG),
    .N2END(Tile_X1Y7_N2BEGb),
    .N4END(Tile_X1Y7_N4BEG),
    .NN4END(Tile_X1Y7_NN4BEG),
    .Ci(Tile_X1Y7_Co),
    .E1END(Tile_X0Y6_E1BEG),
    .E2MID(Tile_X0Y6_E2BEG),
    .E2END(Tile_X0Y6_E2BEGb),
    .EE4END(Tile_X0Y6_EE4BEG),
    .E6END(Tile_X0Y6_E6BEG),
    .S1END(Tile_X1Y5_S1BEG),
    .S2MID(Tile_X1Y5_S2BEG),
    .S2END(Tile_X1Y5_S2BEGb),
    .S4END(Tile_X1Y5_S4BEG),
    .SS4END(Tile_X1Y5_SS4BEG),
    .W1END(Tile_X2Y6_W1BEG),
    .W2MID(Tile_X2Y6_W2BEG),
    .W2END(Tile_X2Y6_W2BEGb),
    .WW4END(Tile_X2Y6_WW4BEG),
    .W6END(Tile_X2Y6_W6BEG),
    .N1BEG(Tile_X1Y6_N1BEG),
    .N2BEG(Tile_X1Y6_N2BEG),
    .N2BEGb(Tile_X1Y6_N2BEGb),
    .N4BEG(Tile_X1Y6_N4BEG),
    .NN4BEG(Tile_X1Y6_NN4BEG),
    .E1BEG(Tile_X1Y6_E1BEG),
    .E2BEG(Tile_X1Y6_E2BEG),
    .E2BEGb(Tile_X1Y6_E2BEGb),
    .EE4BEG(Tile_X1Y6_EE4BEG),
    .E6BEG(Tile_X1Y6_E6BEG),
    .S1BEG(Tile_X1Y6_S1BEG),
    .S2BEG(Tile_X1Y6_S2BEG),
    .S2BEGb(Tile_X1Y6_S2BEGb),
    .S4BEG(Tile_X1Y6_S4BEG),
    .SS4BEG(Tile_X1Y6_SS4BEG),
    .W1BEG(Tile_X1Y6_W1BEG),
    .W2BEG(Tile_X1Y6_W2BEG),
    .W2BEGb(Tile_X1Y6_W2BEGb),
    .WW4BEG(Tile_X1Y6_WW4BEG),
    .W6BEG(Tile_X1Y6_W6BEG),
    .Co(Tile_X1Y6_Co),
    .UserCLK(Tile_X1Y7_UserCLKo),
    .UserCLKo(Tile_X1Y6_UserCLKo),
    .FrameData(Tile_X0Y6_FrameData_O),
    .FrameData_O(Tile_X1Y6_FrameData_O),
    .FrameStrobe(Tile_X1Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y6_Emulate_Bitstream)
    )
`endif
    Tile_X2Y6_LUT4AB
    (
    .N1END(Tile_X2Y7_N1BEG),
    .N2MID(Tile_X2Y7_N2BEG),
    .N2END(Tile_X2Y7_N2BEGb),
    .N4END(Tile_X2Y7_N4BEG),
    .NN4END(Tile_X2Y7_NN4BEG),
    .Ci(Tile_X2Y7_Co),
    .E1END(Tile_X1Y6_E1BEG),
    .E2MID(Tile_X1Y6_E2BEG),
    .E2END(Tile_X1Y6_E2BEGb),
    .EE4END(Tile_X1Y6_EE4BEG),
    .E6END(Tile_X1Y6_E6BEG),
    .S1END(Tile_X2Y5_S1BEG),
    .S2MID(Tile_X2Y5_S2BEG),
    .S2END(Tile_X2Y5_S2BEGb),
    .S4END(Tile_X2Y5_S4BEG),
    .SS4END(Tile_X2Y5_SS4BEG),
    .W1END(Tile_X3Y6_W1BEG),
    .W2MID(Tile_X3Y6_W2BEG),
    .W2END(Tile_X3Y6_W2BEGb),
    .WW4END(Tile_X3Y6_WW4BEG),
    .W6END(Tile_X3Y6_W6BEG),
    .N1BEG(Tile_X2Y6_N1BEG),
    .N2BEG(Tile_X2Y6_N2BEG),
    .N2BEGb(Tile_X2Y6_N2BEGb),
    .N4BEG(Tile_X2Y6_N4BEG),
    .NN4BEG(Tile_X2Y6_NN4BEG),
    .E1BEG(Tile_X2Y6_E1BEG),
    .E2BEG(Tile_X2Y6_E2BEG),
    .E2BEGb(Tile_X2Y6_E2BEGb),
    .EE4BEG(Tile_X2Y6_EE4BEG),
    .E6BEG(Tile_X2Y6_E6BEG),
    .S1BEG(Tile_X2Y6_S1BEG),
    .S2BEG(Tile_X2Y6_S2BEG),
    .S2BEGb(Tile_X2Y6_S2BEGb),
    .S4BEG(Tile_X2Y6_S4BEG),
    .SS4BEG(Tile_X2Y6_SS4BEG),
    .W1BEG(Tile_X2Y6_W1BEG),
    .W2BEG(Tile_X2Y6_W2BEG),
    .W2BEGb(Tile_X2Y6_W2BEGb),
    .WW4BEG(Tile_X2Y6_WW4BEG),
    .W6BEG(Tile_X2Y6_W6BEG),
    .Co(Tile_X2Y6_Co),
    .UserCLK(Tile_X2Y7_UserCLKo),
    .UserCLKo(Tile_X2Y6_UserCLKo),
    .FrameData(Tile_X1Y6_FrameData_O),
    .FrameData_O(Tile_X2Y6_FrameData_O),
    .FrameStrobe(Tile_X2Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y6_Emulate_Bitstream)
    )
`endif
    Tile_X3Y6_LUT4AB
    (
    .N1END(Tile_X3Y7_N1BEG),
    .N2MID(Tile_X3Y7_N2BEG),
    .N2END(Tile_X3Y7_N2BEGb),
    .N4END(Tile_X3Y7_N4BEG),
    .NN4END(Tile_X3Y7_NN4BEG),
    .Ci(Tile_X3Y7_Co),
    .E1END(Tile_X2Y6_E1BEG),
    .E2MID(Tile_X2Y6_E2BEG),
    .E2END(Tile_X2Y6_E2BEGb),
    .EE4END(Tile_X2Y6_EE4BEG),
    .E6END(Tile_X2Y6_E6BEG),
    .S1END(Tile_X3Y5_S1BEG),
    .S2MID(Tile_X3Y5_S2BEG),
    .S2END(Tile_X3Y5_S2BEGb),
    .S4END(Tile_X3Y5_S4BEG),
    .SS4END(Tile_X3Y5_SS4BEG),
    .W1END(Tile_X4Y6_W1BEG),
    .W2MID(Tile_X4Y6_W2BEG),
    .W2END(Tile_X4Y6_W2BEGb),
    .WW4END(Tile_X4Y6_WW4BEG),
    .W6END(Tile_X4Y6_W6BEG),
    .N1BEG(Tile_X3Y6_N1BEG),
    .N2BEG(Tile_X3Y6_N2BEG),
    .N2BEGb(Tile_X3Y6_N2BEGb),
    .N4BEG(Tile_X3Y6_N4BEG),
    .NN4BEG(Tile_X3Y6_NN4BEG),
    .E1BEG(Tile_X3Y6_E1BEG),
    .E2BEG(Tile_X3Y6_E2BEG),
    .E2BEGb(Tile_X3Y6_E2BEGb),
    .EE4BEG(Tile_X3Y6_EE4BEG),
    .E6BEG(Tile_X3Y6_E6BEG),
    .S1BEG(Tile_X3Y6_S1BEG),
    .S2BEG(Tile_X3Y6_S2BEG),
    .S2BEGb(Tile_X3Y6_S2BEGb),
    .S4BEG(Tile_X3Y6_S4BEG),
    .SS4BEG(Tile_X3Y6_SS4BEG),
    .W1BEG(Tile_X3Y6_W1BEG),
    .W2BEG(Tile_X3Y6_W2BEG),
    .W2BEGb(Tile_X3Y6_W2BEGb),
    .WW4BEG(Tile_X3Y6_WW4BEG),
    .W6BEG(Tile_X3Y6_W6BEG),
    .Co(Tile_X3Y6_Co),
    .UserCLK(Tile_X3Y7_UserCLKo),
    .UserCLKo(Tile_X3Y6_UserCLKo),
    .FrameData(Tile_X2Y6_FrameData_O),
    .FrameData_O(Tile_X3Y6_FrameData_O),
    .FrameStrobe(Tile_X3Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y6_Emulate_Bitstream)
    )
`endif
    Tile_X4Y6_LUT4AB
    (
    .N1END(Tile_X4Y7_N1BEG),
    .N2MID(Tile_X4Y7_N2BEG),
    .N2END(Tile_X4Y7_N2BEGb),
    .N4END(Tile_X4Y7_N4BEG),
    .NN4END(Tile_X4Y7_NN4BEG),
    .Ci(Tile_X4Y7_Co),
    .E1END(Tile_X3Y6_E1BEG),
    .E2MID(Tile_X3Y6_E2BEG),
    .E2END(Tile_X3Y6_E2BEGb),
    .EE4END(Tile_X3Y6_EE4BEG),
    .E6END(Tile_X3Y6_E6BEG),
    .S1END(Tile_X4Y5_S1BEG),
    .S2MID(Tile_X4Y5_S2BEG),
    .S2END(Tile_X4Y5_S2BEGb),
    .S4END(Tile_X4Y5_S4BEG),
    .SS4END(Tile_X4Y5_SS4BEG),
    .W1END(Tile_X5Y6_W1BEG),
    .W2MID(Tile_X5Y6_W2BEG),
    .W2END(Tile_X5Y6_W2BEGb),
    .WW4END(Tile_X5Y6_WW4BEG),
    .W6END(Tile_X5Y6_W6BEG),
    .N1BEG(Tile_X4Y6_N1BEG),
    .N2BEG(Tile_X4Y6_N2BEG),
    .N2BEGb(Tile_X4Y6_N2BEGb),
    .N4BEG(Tile_X4Y6_N4BEG),
    .NN4BEG(Tile_X4Y6_NN4BEG),
    .E1BEG(Tile_X4Y6_E1BEG),
    .E2BEG(Tile_X4Y6_E2BEG),
    .E2BEGb(Tile_X4Y6_E2BEGb),
    .EE4BEG(Tile_X4Y6_EE4BEG),
    .E6BEG(Tile_X4Y6_E6BEG),
    .S1BEG(Tile_X4Y6_S1BEG),
    .S2BEG(Tile_X4Y6_S2BEG),
    .S2BEGb(Tile_X4Y6_S2BEGb),
    .S4BEG(Tile_X4Y6_S4BEG),
    .SS4BEG(Tile_X4Y6_SS4BEG),
    .W1BEG(Tile_X4Y6_W1BEG),
    .W2BEG(Tile_X4Y6_W2BEG),
    .W2BEGb(Tile_X4Y6_W2BEGb),
    .WW4BEG(Tile_X4Y6_WW4BEG),
    .W6BEG(Tile_X4Y6_W6BEG),
    .Co(Tile_X4Y6_Co),
    .UserCLK(Tile_X4Y7_UserCLKo),
    .UserCLKo(Tile_X4Y6_UserCLKo),
    .FrameData(Tile_X3Y6_FrameData_O),
    .FrameData_O(Tile_X4Y6_FrameData_O),
    .FrameStrobe(Tile_X4Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
E_TT_IF
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y6_Emulate_Bitstream)
    )
`endif
    Tile_X5Y6_E_TT_IF
    (
    .N1END(Tile_X5Y7_N1BEG),
    .N2MID(Tile_X5Y7_N2BEG),
    .N2END(Tile_X5Y7_N2BEGb),
    .N4END(Tile_X5Y7_N4BEG),
    .E1END(Tile_X4Y6_E1BEG),
    .E2MID(Tile_X4Y6_E2BEG),
    .E2END(Tile_X4Y6_E2BEGb),
    .EE4END(Tile_X4Y6_EE4BEG),
    .E6END(Tile_X4Y6_E6BEG),
    .S1END(Tile_X5Y5_S1BEG),
    .S2MID(Tile_X5Y5_S2BEG),
    .S2END(Tile_X5Y5_S2BEGb),
    .S4END(Tile_X5Y5_S4BEG),
    .N1BEG(Tile_X5Y6_N1BEG),
    .N2BEG(Tile_X5Y6_N2BEG),
    .N2BEGb(Tile_X5Y6_N2BEGb),
    .N4BEG(Tile_X5Y6_N4BEG),
    .S1BEG(Tile_X5Y6_S1BEG),
    .S2BEG(Tile_X5Y6_S2BEG),
    .S2BEGb(Tile_X5Y6_S2BEGb),
    .S4BEG(Tile_X5Y6_S4BEG),
    .W1BEG(Tile_X5Y6_W1BEG),
    .W2BEG(Tile_X5Y6_W2BEG),
    .W2BEGb(Tile_X5Y6_W2BEGb),
    .WW4BEG(Tile_X5Y6_WW4BEG),
    .W6BEG(Tile_X5Y6_W6BEG),
    .UO_OUT_TT_PROJECT0(Tile_X5Y6_UO_OUT_TT_PROJECT0),
    .UO_OUT_TT_PROJECT1(Tile_X5Y6_UO_OUT_TT_PROJECT1),
    .UO_OUT_TT_PROJECT2(Tile_X5Y6_UO_OUT_TT_PROJECT2),
    .UO_OUT_TT_PROJECT3(Tile_X5Y6_UO_OUT_TT_PROJECT3),
    .UO_OUT_TT_PROJECT4(Tile_X5Y6_UO_OUT_TT_PROJECT4),
    .UO_OUT_TT_PROJECT5(Tile_X5Y6_UO_OUT_TT_PROJECT5),
    .UO_OUT_TT_PROJECT6(Tile_X5Y6_UO_OUT_TT_PROJECT6),
    .UO_OUT_TT_PROJECT7(Tile_X5Y6_UO_OUT_TT_PROJECT7),
    .UIO_OUT_TT_PROJECT0(Tile_X5Y6_UIO_OUT_TT_PROJECT0),
    .UIO_OUT_TT_PROJECT1(Tile_X5Y6_UIO_OUT_TT_PROJECT1),
    .UIO_OUT_TT_PROJECT2(Tile_X5Y6_UIO_OUT_TT_PROJECT2),
    .UIO_OUT_TT_PROJECT3(Tile_X5Y6_UIO_OUT_TT_PROJECT3),
    .UIO_OUT_TT_PROJECT4(Tile_X5Y6_UIO_OUT_TT_PROJECT4),
    .UIO_OUT_TT_PROJECT5(Tile_X5Y6_UIO_OUT_TT_PROJECT5),
    .UIO_OUT_TT_PROJECT6(Tile_X5Y6_UIO_OUT_TT_PROJECT6),
    .UIO_OUT_TT_PROJECT7(Tile_X5Y6_UIO_OUT_TT_PROJECT7),
    .UIO_OE_TT_PROJECT0(Tile_X5Y6_UIO_OE_TT_PROJECT0),
    .UIO_OE_TT_PROJECT1(Tile_X5Y6_UIO_OE_TT_PROJECT1),
    .UIO_OE_TT_PROJECT2(Tile_X5Y6_UIO_OE_TT_PROJECT2),
    .UIO_OE_TT_PROJECT3(Tile_X5Y6_UIO_OE_TT_PROJECT3),
    .UIO_OE_TT_PROJECT4(Tile_X5Y6_UIO_OE_TT_PROJECT4),
    .UIO_OE_TT_PROJECT5(Tile_X5Y6_UIO_OE_TT_PROJECT5),
    .UIO_OE_TT_PROJECT6(Tile_X5Y6_UIO_OE_TT_PROJECT6),
    .UIO_OE_TT_PROJECT7(Tile_X5Y6_UIO_OE_TT_PROJECT7),
    .UI_IN_TT_PROJECT0(Tile_X5Y6_UI_IN_TT_PROJECT0),
    .UI_IN_TT_PROJECT1(Tile_X5Y6_UI_IN_TT_PROJECT1),
    .UI_IN_TT_PROJECT2(Tile_X5Y6_UI_IN_TT_PROJECT2),
    .UI_IN_TT_PROJECT3(Tile_X5Y6_UI_IN_TT_PROJECT3),
    .UI_IN_TT_PROJECT4(Tile_X5Y6_UI_IN_TT_PROJECT4),
    .UI_IN_TT_PROJECT5(Tile_X5Y6_UI_IN_TT_PROJECT5),
    .UI_IN_TT_PROJECT6(Tile_X5Y6_UI_IN_TT_PROJECT6),
    .UI_IN_TT_PROJECT7(Tile_X5Y6_UI_IN_TT_PROJECT7),
    .UIO_IN_TT_PROJECT0(Tile_X5Y6_UIO_IN_TT_PROJECT0),
    .UIO_IN_TT_PROJECT1(Tile_X5Y6_UIO_IN_TT_PROJECT1),
    .UIO_IN_TT_PROJECT2(Tile_X5Y6_UIO_IN_TT_PROJECT2),
    .UIO_IN_TT_PROJECT3(Tile_X5Y6_UIO_IN_TT_PROJECT3),
    .UIO_IN_TT_PROJECT4(Tile_X5Y6_UIO_IN_TT_PROJECT4),
    .UIO_IN_TT_PROJECT5(Tile_X5Y6_UIO_IN_TT_PROJECT5),
    .UIO_IN_TT_PROJECT6(Tile_X5Y6_UIO_IN_TT_PROJECT6),
    .UIO_IN_TT_PROJECT7(Tile_X5Y6_UIO_IN_TT_PROJECT7),
    .ENA_TT_PROJECT(Tile_X5Y6_ENA_TT_PROJECT),
    .CLK_TT_PROJECT(Tile_X5Y6_CLK_TT_PROJECT),
    .RST_N_TT_PROJECT(Tile_X5Y6_RST_N_TT_PROJECT),
    .UserCLK(Tile_X5Y7_UserCLKo),
    .UserCLKo(Tile_X5Y6_UserCLKo),
    .FrameData(Tile_X4Y6_FrameData_O),
    .FrameData_O(Tile_X5Y6_FrameData_O),
    .FrameStrobe(Tile_X5Y7_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y6_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_TT_IF
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y7_Emulate_Bitstream)
    )
`endif
    Tile_X0Y7_W_TT_IF
    (
    .N1END(Tile_X0Y8_N1BEG),
    .N2MID(Tile_X0Y8_N2BEG),
    .N2END(Tile_X0Y8_N2BEGb),
    .N4END(Tile_X0Y8_N4BEG),
    .S1END(Tile_X0Y6_S1BEG),
    .S2MID(Tile_X0Y6_S2BEG),
    .S2END(Tile_X0Y6_S2BEGb),
    .S4END(Tile_X0Y6_S4BEG),
    .W1END(Tile_X1Y7_W1BEG),
    .W2MID(Tile_X1Y7_W2BEG),
    .W2END(Tile_X1Y7_W2BEGb),
    .WW4END(Tile_X1Y7_WW4BEG),
    .W6END(Tile_X1Y7_W6BEG),
    .N1BEG(Tile_X0Y7_N1BEG),
    .N2BEG(Tile_X0Y7_N2BEG),
    .N2BEGb(Tile_X0Y7_N2BEGb),
    .N4BEG(Tile_X0Y7_N4BEG),
    .S1BEG(Tile_X0Y7_S1BEG),
    .S2BEG(Tile_X0Y7_S2BEG),
    .S2BEGb(Tile_X0Y7_S2BEGb),
    .S4BEG(Tile_X0Y7_S4BEG),
    .E1BEG(Tile_X0Y7_E1BEG),
    .E2BEG(Tile_X0Y7_E2BEG),
    .E2BEGb(Tile_X0Y7_E2BEGb),
    .EE4BEG(Tile_X0Y7_EE4BEG),
    .E6BEG(Tile_X0Y7_E6BEG),
    .UO_OUT_TT_PROJECT0(Tile_X0Y7_UO_OUT_TT_PROJECT0),
    .UO_OUT_TT_PROJECT1(Tile_X0Y7_UO_OUT_TT_PROJECT1),
    .UO_OUT_TT_PROJECT2(Tile_X0Y7_UO_OUT_TT_PROJECT2),
    .UO_OUT_TT_PROJECT3(Tile_X0Y7_UO_OUT_TT_PROJECT3),
    .UO_OUT_TT_PROJECT4(Tile_X0Y7_UO_OUT_TT_PROJECT4),
    .UO_OUT_TT_PROJECT5(Tile_X0Y7_UO_OUT_TT_PROJECT5),
    .UO_OUT_TT_PROJECT6(Tile_X0Y7_UO_OUT_TT_PROJECT6),
    .UO_OUT_TT_PROJECT7(Tile_X0Y7_UO_OUT_TT_PROJECT7),
    .UIO_OUT_TT_PROJECT0(Tile_X0Y7_UIO_OUT_TT_PROJECT0),
    .UIO_OUT_TT_PROJECT1(Tile_X0Y7_UIO_OUT_TT_PROJECT1),
    .UIO_OUT_TT_PROJECT2(Tile_X0Y7_UIO_OUT_TT_PROJECT2),
    .UIO_OUT_TT_PROJECT3(Tile_X0Y7_UIO_OUT_TT_PROJECT3),
    .UIO_OUT_TT_PROJECT4(Tile_X0Y7_UIO_OUT_TT_PROJECT4),
    .UIO_OUT_TT_PROJECT5(Tile_X0Y7_UIO_OUT_TT_PROJECT5),
    .UIO_OUT_TT_PROJECT6(Tile_X0Y7_UIO_OUT_TT_PROJECT6),
    .UIO_OUT_TT_PROJECT7(Tile_X0Y7_UIO_OUT_TT_PROJECT7),
    .UIO_OE_TT_PROJECT0(Tile_X0Y7_UIO_OE_TT_PROJECT0),
    .UIO_OE_TT_PROJECT1(Tile_X0Y7_UIO_OE_TT_PROJECT1),
    .UIO_OE_TT_PROJECT2(Tile_X0Y7_UIO_OE_TT_PROJECT2),
    .UIO_OE_TT_PROJECT3(Tile_X0Y7_UIO_OE_TT_PROJECT3),
    .UIO_OE_TT_PROJECT4(Tile_X0Y7_UIO_OE_TT_PROJECT4),
    .UIO_OE_TT_PROJECT5(Tile_X0Y7_UIO_OE_TT_PROJECT5),
    .UIO_OE_TT_PROJECT6(Tile_X0Y7_UIO_OE_TT_PROJECT6),
    .UIO_OE_TT_PROJECT7(Tile_X0Y7_UIO_OE_TT_PROJECT7),
    .UI_IN_TT_PROJECT0(Tile_X0Y7_UI_IN_TT_PROJECT0),
    .UI_IN_TT_PROJECT1(Tile_X0Y7_UI_IN_TT_PROJECT1),
    .UI_IN_TT_PROJECT2(Tile_X0Y7_UI_IN_TT_PROJECT2),
    .UI_IN_TT_PROJECT3(Tile_X0Y7_UI_IN_TT_PROJECT3),
    .UI_IN_TT_PROJECT4(Tile_X0Y7_UI_IN_TT_PROJECT4),
    .UI_IN_TT_PROJECT5(Tile_X0Y7_UI_IN_TT_PROJECT5),
    .UI_IN_TT_PROJECT6(Tile_X0Y7_UI_IN_TT_PROJECT6),
    .UI_IN_TT_PROJECT7(Tile_X0Y7_UI_IN_TT_PROJECT7),
    .UIO_IN_TT_PROJECT0(Tile_X0Y7_UIO_IN_TT_PROJECT0),
    .UIO_IN_TT_PROJECT1(Tile_X0Y7_UIO_IN_TT_PROJECT1),
    .UIO_IN_TT_PROJECT2(Tile_X0Y7_UIO_IN_TT_PROJECT2),
    .UIO_IN_TT_PROJECT3(Tile_X0Y7_UIO_IN_TT_PROJECT3),
    .UIO_IN_TT_PROJECT4(Tile_X0Y7_UIO_IN_TT_PROJECT4),
    .UIO_IN_TT_PROJECT5(Tile_X0Y7_UIO_IN_TT_PROJECT5),
    .UIO_IN_TT_PROJECT6(Tile_X0Y7_UIO_IN_TT_PROJECT6),
    .UIO_IN_TT_PROJECT7(Tile_X0Y7_UIO_IN_TT_PROJECT7),
    .ENA_TT_PROJECT(Tile_X0Y7_ENA_TT_PROJECT),
    .CLK_TT_PROJECT(Tile_X0Y7_CLK_TT_PROJECT),
    .RST_N_TT_PROJECT(Tile_X0Y7_RST_N_TT_PROJECT),
    .UserCLK(Tile_X0Y8_UserCLKo),
    .UserCLKo(Tile_X0Y7_UserCLKo),
    .FrameData(Row_Y7_FrameData),
    .FrameData_O(Tile_X0Y7_FrameData_O),
    .FrameStrobe(Tile_X0Y8_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y7_Emulate_Bitstream)
    )
`endif
    Tile_X1Y7_LUT4AB
    (
    .N1END(Tile_X1Y8_N1BEG),
    .N2MID(Tile_X1Y8_N2BEG),
    .N2END(Tile_X1Y8_N2BEGb),
    .N4END(Tile_X1Y8_N4BEG),
    .NN4END(Tile_X1Y8_NN4BEG),
    .Ci(Tile_X1Y8_Co),
    .E1END(Tile_X0Y7_E1BEG),
    .E2MID(Tile_X0Y7_E2BEG),
    .E2END(Tile_X0Y7_E2BEGb),
    .EE4END(Tile_X0Y7_EE4BEG),
    .E6END(Tile_X0Y7_E6BEG),
    .S1END(Tile_X1Y6_S1BEG),
    .S2MID(Tile_X1Y6_S2BEG),
    .S2END(Tile_X1Y6_S2BEGb),
    .S4END(Tile_X1Y6_S4BEG),
    .SS4END(Tile_X1Y6_SS4BEG),
    .W1END(Tile_X2Y7_W1BEG),
    .W2MID(Tile_X2Y7_W2BEG),
    .W2END(Tile_X2Y7_W2BEGb),
    .WW4END(Tile_X2Y7_WW4BEG),
    .W6END(Tile_X2Y7_W6BEG),
    .N1BEG(Tile_X1Y7_N1BEG),
    .N2BEG(Tile_X1Y7_N2BEG),
    .N2BEGb(Tile_X1Y7_N2BEGb),
    .N4BEG(Tile_X1Y7_N4BEG),
    .NN4BEG(Tile_X1Y7_NN4BEG),
    .E1BEG(Tile_X1Y7_E1BEG),
    .E2BEG(Tile_X1Y7_E2BEG),
    .E2BEGb(Tile_X1Y7_E2BEGb),
    .EE4BEG(Tile_X1Y7_EE4BEG),
    .E6BEG(Tile_X1Y7_E6BEG),
    .S1BEG(Tile_X1Y7_S1BEG),
    .S2BEG(Tile_X1Y7_S2BEG),
    .S2BEGb(Tile_X1Y7_S2BEGb),
    .S4BEG(Tile_X1Y7_S4BEG),
    .SS4BEG(Tile_X1Y7_SS4BEG),
    .W1BEG(Tile_X1Y7_W1BEG),
    .W2BEG(Tile_X1Y7_W2BEG),
    .W2BEGb(Tile_X1Y7_W2BEGb),
    .WW4BEG(Tile_X1Y7_WW4BEG),
    .W6BEG(Tile_X1Y7_W6BEG),
    .Co(Tile_X1Y7_Co),
    .UserCLK(Tile_X1Y8_UserCLKo),
    .UserCLKo(Tile_X1Y7_UserCLKo),
    .FrameData(Tile_X0Y7_FrameData_O),
    .FrameData_O(Tile_X1Y7_FrameData_O),
    .FrameStrobe(Tile_X1Y8_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y7_Emulate_Bitstream)
    )
`endif
    Tile_X2Y7_LUT4AB
    (
    .N1END(Tile_X2Y8_N1BEG),
    .N2MID(Tile_X2Y8_N2BEG),
    .N2END(Tile_X2Y8_N2BEGb),
    .N4END(Tile_X2Y8_N4BEG),
    .NN4END(Tile_X2Y8_NN4BEG),
    .Ci(Tile_X2Y8_Co),
    .E1END(Tile_X1Y7_E1BEG),
    .E2MID(Tile_X1Y7_E2BEG),
    .E2END(Tile_X1Y7_E2BEGb),
    .EE4END(Tile_X1Y7_EE4BEG),
    .E6END(Tile_X1Y7_E6BEG),
    .S1END(Tile_X2Y6_S1BEG),
    .S2MID(Tile_X2Y6_S2BEG),
    .S2END(Tile_X2Y6_S2BEGb),
    .S4END(Tile_X2Y6_S4BEG),
    .SS4END(Tile_X2Y6_SS4BEG),
    .W1END(Tile_X3Y7_W1BEG),
    .W2MID(Tile_X3Y7_W2BEG),
    .W2END(Tile_X3Y7_W2BEGb),
    .WW4END(Tile_X3Y7_WW4BEG),
    .W6END(Tile_X3Y7_W6BEG),
    .N1BEG(Tile_X2Y7_N1BEG),
    .N2BEG(Tile_X2Y7_N2BEG),
    .N2BEGb(Tile_X2Y7_N2BEGb),
    .N4BEG(Tile_X2Y7_N4BEG),
    .NN4BEG(Tile_X2Y7_NN4BEG),
    .E1BEG(Tile_X2Y7_E1BEG),
    .E2BEG(Tile_X2Y7_E2BEG),
    .E2BEGb(Tile_X2Y7_E2BEGb),
    .EE4BEG(Tile_X2Y7_EE4BEG),
    .E6BEG(Tile_X2Y7_E6BEG),
    .S1BEG(Tile_X2Y7_S1BEG),
    .S2BEG(Tile_X2Y7_S2BEG),
    .S2BEGb(Tile_X2Y7_S2BEGb),
    .S4BEG(Tile_X2Y7_S4BEG),
    .SS4BEG(Tile_X2Y7_SS4BEG),
    .W1BEG(Tile_X2Y7_W1BEG),
    .W2BEG(Tile_X2Y7_W2BEG),
    .W2BEGb(Tile_X2Y7_W2BEGb),
    .WW4BEG(Tile_X2Y7_WW4BEG),
    .W6BEG(Tile_X2Y7_W6BEG),
    .Co(Tile_X2Y7_Co),
    .UserCLK(Tile_X2Y8_UserCLKo),
    .UserCLKo(Tile_X2Y7_UserCLKo),
    .FrameData(Tile_X1Y7_FrameData_O),
    .FrameData_O(Tile_X2Y7_FrameData_O),
    .FrameStrobe(Tile_X2Y8_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y7_Emulate_Bitstream)
    )
`endif
    Tile_X3Y7_LUT4AB
    (
    .N1END(Tile_X3Y8_N1BEG),
    .N2MID(Tile_X3Y8_N2BEG),
    .N2END(Tile_X3Y8_N2BEGb),
    .N4END(Tile_X3Y8_N4BEG),
    .NN4END(Tile_X3Y8_NN4BEG),
    .Ci(Tile_X3Y8_Co),
    .E1END(Tile_X2Y7_E1BEG),
    .E2MID(Tile_X2Y7_E2BEG),
    .E2END(Tile_X2Y7_E2BEGb),
    .EE4END(Tile_X2Y7_EE4BEG),
    .E6END(Tile_X2Y7_E6BEG),
    .S1END(Tile_X3Y6_S1BEG),
    .S2MID(Tile_X3Y6_S2BEG),
    .S2END(Tile_X3Y6_S2BEGb),
    .S4END(Tile_X3Y6_S4BEG),
    .SS4END(Tile_X3Y6_SS4BEG),
    .W1END(Tile_X4Y7_W1BEG),
    .W2MID(Tile_X4Y7_W2BEG),
    .W2END(Tile_X4Y7_W2BEGb),
    .WW4END(Tile_X4Y7_WW4BEG),
    .W6END(Tile_X4Y7_W6BEG),
    .N1BEG(Tile_X3Y7_N1BEG),
    .N2BEG(Tile_X3Y7_N2BEG),
    .N2BEGb(Tile_X3Y7_N2BEGb),
    .N4BEG(Tile_X3Y7_N4BEG),
    .NN4BEG(Tile_X3Y7_NN4BEG),
    .E1BEG(Tile_X3Y7_E1BEG),
    .E2BEG(Tile_X3Y7_E2BEG),
    .E2BEGb(Tile_X3Y7_E2BEGb),
    .EE4BEG(Tile_X3Y7_EE4BEG),
    .E6BEG(Tile_X3Y7_E6BEG),
    .S1BEG(Tile_X3Y7_S1BEG),
    .S2BEG(Tile_X3Y7_S2BEG),
    .S2BEGb(Tile_X3Y7_S2BEGb),
    .S4BEG(Tile_X3Y7_S4BEG),
    .SS4BEG(Tile_X3Y7_SS4BEG),
    .W1BEG(Tile_X3Y7_W1BEG),
    .W2BEG(Tile_X3Y7_W2BEG),
    .W2BEGb(Tile_X3Y7_W2BEGb),
    .WW4BEG(Tile_X3Y7_WW4BEG),
    .W6BEG(Tile_X3Y7_W6BEG),
    .Co(Tile_X3Y7_Co),
    .UserCLK(Tile_X3Y8_UserCLKo),
    .UserCLKo(Tile_X3Y7_UserCLKo),
    .FrameData(Tile_X2Y7_FrameData_O),
    .FrameData_O(Tile_X3Y7_FrameData_O),
    .FrameStrobe(Tile_X3Y8_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y7_Emulate_Bitstream)
    )
`endif
    Tile_X4Y7_LUT4AB
    (
    .N1END(Tile_X4Y8_N1BEG),
    .N2MID(Tile_X4Y8_N2BEG),
    .N2END(Tile_X4Y8_N2BEGb),
    .N4END(Tile_X4Y8_N4BEG),
    .NN4END(Tile_X4Y8_NN4BEG),
    .Ci(Tile_X4Y8_Co),
    .E1END(Tile_X3Y7_E1BEG),
    .E2MID(Tile_X3Y7_E2BEG),
    .E2END(Tile_X3Y7_E2BEGb),
    .EE4END(Tile_X3Y7_EE4BEG),
    .E6END(Tile_X3Y7_E6BEG),
    .S1END(Tile_X4Y6_S1BEG),
    .S2MID(Tile_X4Y6_S2BEG),
    .S2END(Tile_X4Y6_S2BEGb),
    .S4END(Tile_X4Y6_S4BEG),
    .SS4END(Tile_X4Y6_SS4BEG),
    .W1END(Tile_X5Y7_W1BEG),
    .W2MID(Tile_X5Y7_W2BEG),
    .W2END(Tile_X5Y7_W2BEGb),
    .WW4END(Tile_X5Y7_WW4BEG),
    .W6END(Tile_X5Y7_W6BEG),
    .N1BEG(Tile_X4Y7_N1BEG),
    .N2BEG(Tile_X4Y7_N2BEG),
    .N2BEGb(Tile_X4Y7_N2BEGb),
    .N4BEG(Tile_X4Y7_N4BEG),
    .NN4BEG(Tile_X4Y7_NN4BEG),
    .E1BEG(Tile_X4Y7_E1BEG),
    .E2BEG(Tile_X4Y7_E2BEG),
    .E2BEGb(Tile_X4Y7_E2BEGb),
    .EE4BEG(Tile_X4Y7_EE4BEG),
    .E6BEG(Tile_X4Y7_E6BEG),
    .S1BEG(Tile_X4Y7_S1BEG),
    .S2BEG(Tile_X4Y7_S2BEG),
    .S2BEGb(Tile_X4Y7_S2BEGb),
    .S4BEG(Tile_X4Y7_S4BEG),
    .SS4BEG(Tile_X4Y7_SS4BEG),
    .W1BEG(Tile_X4Y7_W1BEG),
    .W2BEG(Tile_X4Y7_W2BEG),
    .W2BEGb(Tile_X4Y7_W2BEGb),
    .WW4BEG(Tile_X4Y7_WW4BEG),
    .W6BEG(Tile_X4Y7_W6BEG),
    .Co(Tile_X4Y7_Co),
    .UserCLK(Tile_X4Y8_UserCLKo),
    .UserCLKo(Tile_X4Y7_UserCLKo),
    .FrameData(Tile_X3Y7_FrameData_O),
    .FrameData_O(Tile_X4Y7_FrameData_O),
    .FrameStrobe(Tile_X4Y8_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
E_TT_IF
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y7_Emulate_Bitstream)
    )
`endif
    Tile_X5Y7_E_TT_IF
    (
    .N1END(Tile_X5Y8_N1BEG),
    .N2MID(Tile_X5Y8_N2BEG),
    .N2END(Tile_X5Y8_N2BEGb),
    .N4END(Tile_X5Y8_N4BEG),
    .E1END(Tile_X4Y7_E1BEG),
    .E2MID(Tile_X4Y7_E2BEG),
    .E2END(Tile_X4Y7_E2BEGb),
    .EE4END(Tile_X4Y7_EE4BEG),
    .E6END(Tile_X4Y7_E6BEG),
    .S1END(Tile_X5Y6_S1BEG),
    .S2MID(Tile_X5Y6_S2BEG),
    .S2END(Tile_X5Y6_S2BEGb),
    .S4END(Tile_X5Y6_S4BEG),
    .N1BEG(Tile_X5Y7_N1BEG),
    .N2BEG(Tile_X5Y7_N2BEG),
    .N2BEGb(Tile_X5Y7_N2BEGb),
    .N4BEG(Tile_X5Y7_N4BEG),
    .S1BEG(Tile_X5Y7_S1BEG),
    .S2BEG(Tile_X5Y7_S2BEG),
    .S2BEGb(Tile_X5Y7_S2BEGb),
    .S4BEG(Tile_X5Y7_S4BEG),
    .W1BEG(Tile_X5Y7_W1BEG),
    .W2BEG(Tile_X5Y7_W2BEG),
    .W2BEGb(Tile_X5Y7_W2BEGb),
    .WW4BEG(Tile_X5Y7_WW4BEG),
    .W6BEG(Tile_X5Y7_W6BEG),
    .UO_OUT_TT_PROJECT0(Tile_X5Y7_UO_OUT_TT_PROJECT0),
    .UO_OUT_TT_PROJECT1(Tile_X5Y7_UO_OUT_TT_PROJECT1),
    .UO_OUT_TT_PROJECT2(Tile_X5Y7_UO_OUT_TT_PROJECT2),
    .UO_OUT_TT_PROJECT3(Tile_X5Y7_UO_OUT_TT_PROJECT3),
    .UO_OUT_TT_PROJECT4(Tile_X5Y7_UO_OUT_TT_PROJECT4),
    .UO_OUT_TT_PROJECT5(Tile_X5Y7_UO_OUT_TT_PROJECT5),
    .UO_OUT_TT_PROJECT6(Tile_X5Y7_UO_OUT_TT_PROJECT6),
    .UO_OUT_TT_PROJECT7(Tile_X5Y7_UO_OUT_TT_PROJECT7),
    .UIO_OUT_TT_PROJECT0(Tile_X5Y7_UIO_OUT_TT_PROJECT0),
    .UIO_OUT_TT_PROJECT1(Tile_X5Y7_UIO_OUT_TT_PROJECT1),
    .UIO_OUT_TT_PROJECT2(Tile_X5Y7_UIO_OUT_TT_PROJECT2),
    .UIO_OUT_TT_PROJECT3(Tile_X5Y7_UIO_OUT_TT_PROJECT3),
    .UIO_OUT_TT_PROJECT4(Tile_X5Y7_UIO_OUT_TT_PROJECT4),
    .UIO_OUT_TT_PROJECT5(Tile_X5Y7_UIO_OUT_TT_PROJECT5),
    .UIO_OUT_TT_PROJECT6(Tile_X5Y7_UIO_OUT_TT_PROJECT6),
    .UIO_OUT_TT_PROJECT7(Tile_X5Y7_UIO_OUT_TT_PROJECT7),
    .UIO_OE_TT_PROJECT0(Tile_X5Y7_UIO_OE_TT_PROJECT0),
    .UIO_OE_TT_PROJECT1(Tile_X5Y7_UIO_OE_TT_PROJECT1),
    .UIO_OE_TT_PROJECT2(Tile_X5Y7_UIO_OE_TT_PROJECT2),
    .UIO_OE_TT_PROJECT3(Tile_X5Y7_UIO_OE_TT_PROJECT3),
    .UIO_OE_TT_PROJECT4(Tile_X5Y7_UIO_OE_TT_PROJECT4),
    .UIO_OE_TT_PROJECT5(Tile_X5Y7_UIO_OE_TT_PROJECT5),
    .UIO_OE_TT_PROJECT6(Tile_X5Y7_UIO_OE_TT_PROJECT6),
    .UIO_OE_TT_PROJECT7(Tile_X5Y7_UIO_OE_TT_PROJECT7),
    .UI_IN_TT_PROJECT0(Tile_X5Y7_UI_IN_TT_PROJECT0),
    .UI_IN_TT_PROJECT1(Tile_X5Y7_UI_IN_TT_PROJECT1),
    .UI_IN_TT_PROJECT2(Tile_X5Y7_UI_IN_TT_PROJECT2),
    .UI_IN_TT_PROJECT3(Tile_X5Y7_UI_IN_TT_PROJECT3),
    .UI_IN_TT_PROJECT4(Tile_X5Y7_UI_IN_TT_PROJECT4),
    .UI_IN_TT_PROJECT5(Tile_X5Y7_UI_IN_TT_PROJECT5),
    .UI_IN_TT_PROJECT6(Tile_X5Y7_UI_IN_TT_PROJECT6),
    .UI_IN_TT_PROJECT7(Tile_X5Y7_UI_IN_TT_PROJECT7),
    .UIO_IN_TT_PROJECT0(Tile_X5Y7_UIO_IN_TT_PROJECT0),
    .UIO_IN_TT_PROJECT1(Tile_X5Y7_UIO_IN_TT_PROJECT1),
    .UIO_IN_TT_PROJECT2(Tile_X5Y7_UIO_IN_TT_PROJECT2),
    .UIO_IN_TT_PROJECT3(Tile_X5Y7_UIO_IN_TT_PROJECT3),
    .UIO_IN_TT_PROJECT4(Tile_X5Y7_UIO_IN_TT_PROJECT4),
    .UIO_IN_TT_PROJECT5(Tile_X5Y7_UIO_IN_TT_PROJECT5),
    .UIO_IN_TT_PROJECT6(Tile_X5Y7_UIO_IN_TT_PROJECT6),
    .UIO_IN_TT_PROJECT7(Tile_X5Y7_UIO_IN_TT_PROJECT7),
    .ENA_TT_PROJECT(Tile_X5Y7_ENA_TT_PROJECT),
    .CLK_TT_PROJECT(Tile_X5Y7_CLK_TT_PROJECT),
    .RST_N_TT_PROJECT(Tile_X5Y7_RST_N_TT_PROJECT),
    .UserCLK(Tile_X5Y8_UserCLKo),
    .UserCLKo(Tile_X5Y7_UserCLKo),
    .FrameData(Tile_X4Y7_FrameData_O),
    .FrameData_O(Tile_X5Y7_FrameData_O),
    .FrameStrobe(Tile_X5Y8_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y7_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
W_TT_IF
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X0Y8_Emulate_Bitstream)
    )
`endif
    Tile_X0Y8_W_TT_IF
    (
    .N1END(Tile_X0Y9_N1BEG),
    .N2MID(Tile_X0Y9_N2BEG),
    .N2END(Tile_X0Y9_N2BEGb),
    .N4END(Tile_X0Y9_N4BEG),
    .S1END(Tile_X0Y7_S1BEG),
    .S2MID(Tile_X0Y7_S2BEG),
    .S2END(Tile_X0Y7_S2BEGb),
    .S4END(Tile_X0Y7_S4BEG),
    .W1END(Tile_X1Y8_W1BEG),
    .W2MID(Tile_X1Y8_W2BEG),
    .W2END(Tile_X1Y8_W2BEGb),
    .WW4END(Tile_X1Y8_WW4BEG),
    .W6END(Tile_X1Y8_W6BEG),
    .N1BEG(Tile_X0Y8_N1BEG),
    .N2BEG(Tile_X0Y8_N2BEG),
    .N2BEGb(Tile_X0Y8_N2BEGb),
    .N4BEG(Tile_X0Y8_N4BEG),
    .S1BEG(Tile_X0Y8_S1BEG),
    .S2BEG(Tile_X0Y8_S2BEG),
    .S2BEGb(Tile_X0Y8_S2BEGb),
    .S4BEG(Tile_X0Y8_S4BEG),
    .E1BEG(Tile_X0Y8_E1BEG),
    .E2BEG(Tile_X0Y8_E2BEG),
    .E2BEGb(Tile_X0Y8_E2BEGb),
    .EE4BEG(Tile_X0Y8_EE4BEG),
    .E6BEG(Tile_X0Y8_E6BEG),
    .UO_OUT_TT_PROJECT0(Tile_X0Y8_UO_OUT_TT_PROJECT0),
    .UO_OUT_TT_PROJECT1(Tile_X0Y8_UO_OUT_TT_PROJECT1),
    .UO_OUT_TT_PROJECT2(Tile_X0Y8_UO_OUT_TT_PROJECT2),
    .UO_OUT_TT_PROJECT3(Tile_X0Y8_UO_OUT_TT_PROJECT3),
    .UO_OUT_TT_PROJECT4(Tile_X0Y8_UO_OUT_TT_PROJECT4),
    .UO_OUT_TT_PROJECT5(Tile_X0Y8_UO_OUT_TT_PROJECT5),
    .UO_OUT_TT_PROJECT6(Tile_X0Y8_UO_OUT_TT_PROJECT6),
    .UO_OUT_TT_PROJECT7(Tile_X0Y8_UO_OUT_TT_PROJECT7),
    .UIO_OUT_TT_PROJECT0(Tile_X0Y8_UIO_OUT_TT_PROJECT0),
    .UIO_OUT_TT_PROJECT1(Tile_X0Y8_UIO_OUT_TT_PROJECT1),
    .UIO_OUT_TT_PROJECT2(Tile_X0Y8_UIO_OUT_TT_PROJECT2),
    .UIO_OUT_TT_PROJECT3(Tile_X0Y8_UIO_OUT_TT_PROJECT3),
    .UIO_OUT_TT_PROJECT4(Tile_X0Y8_UIO_OUT_TT_PROJECT4),
    .UIO_OUT_TT_PROJECT5(Tile_X0Y8_UIO_OUT_TT_PROJECT5),
    .UIO_OUT_TT_PROJECT6(Tile_X0Y8_UIO_OUT_TT_PROJECT6),
    .UIO_OUT_TT_PROJECT7(Tile_X0Y8_UIO_OUT_TT_PROJECT7),
    .UIO_OE_TT_PROJECT0(Tile_X0Y8_UIO_OE_TT_PROJECT0),
    .UIO_OE_TT_PROJECT1(Tile_X0Y8_UIO_OE_TT_PROJECT1),
    .UIO_OE_TT_PROJECT2(Tile_X0Y8_UIO_OE_TT_PROJECT2),
    .UIO_OE_TT_PROJECT3(Tile_X0Y8_UIO_OE_TT_PROJECT3),
    .UIO_OE_TT_PROJECT4(Tile_X0Y8_UIO_OE_TT_PROJECT4),
    .UIO_OE_TT_PROJECT5(Tile_X0Y8_UIO_OE_TT_PROJECT5),
    .UIO_OE_TT_PROJECT6(Tile_X0Y8_UIO_OE_TT_PROJECT6),
    .UIO_OE_TT_PROJECT7(Tile_X0Y8_UIO_OE_TT_PROJECT7),
    .UI_IN_TT_PROJECT0(Tile_X0Y8_UI_IN_TT_PROJECT0),
    .UI_IN_TT_PROJECT1(Tile_X0Y8_UI_IN_TT_PROJECT1),
    .UI_IN_TT_PROJECT2(Tile_X0Y8_UI_IN_TT_PROJECT2),
    .UI_IN_TT_PROJECT3(Tile_X0Y8_UI_IN_TT_PROJECT3),
    .UI_IN_TT_PROJECT4(Tile_X0Y8_UI_IN_TT_PROJECT4),
    .UI_IN_TT_PROJECT5(Tile_X0Y8_UI_IN_TT_PROJECT5),
    .UI_IN_TT_PROJECT6(Tile_X0Y8_UI_IN_TT_PROJECT6),
    .UI_IN_TT_PROJECT7(Tile_X0Y8_UI_IN_TT_PROJECT7),
    .UIO_IN_TT_PROJECT0(Tile_X0Y8_UIO_IN_TT_PROJECT0),
    .UIO_IN_TT_PROJECT1(Tile_X0Y8_UIO_IN_TT_PROJECT1),
    .UIO_IN_TT_PROJECT2(Tile_X0Y8_UIO_IN_TT_PROJECT2),
    .UIO_IN_TT_PROJECT3(Tile_X0Y8_UIO_IN_TT_PROJECT3),
    .UIO_IN_TT_PROJECT4(Tile_X0Y8_UIO_IN_TT_PROJECT4),
    .UIO_IN_TT_PROJECT5(Tile_X0Y8_UIO_IN_TT_PROJECT5),
    .UIO_IN_TT_PROJECT6(Tile_X0Y8_UIO_IN_TT_PROJECT6),
    .UIO_IN_TT_PROJECT7(Tile_X0Y8_UIO_IN_TT_PROJECT7),
    .ENA_TT_PROJECT(Tile_X0Y8_ENA_TT_PROJECT),
    .CLK_TT_PROJECT(Tile_X0Y8_CLK_TT_PROJECT),
    .RST_N_TT_PROJECT(Tile_X0Y8_RST_N_TT_PROJECT),
    .UserCLK(Tile_X0Y9_UserCLKo),
    .UserCLKo(Tile_X0Y8_UserCLKo),
    .FrameData(Row_Y8_FrameData),
    .FrameData_O(Tile_X0Y8_FrameData_O),
    .FrameStrobe(Tile_X0Y9_FrameStrobe_O),
    .FrameStrobe_O(Tile_X0Y8_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X1Y8_Emulate_Bitstream)
    )
`endif
    Tile_X1Y8_LUT4AB
    (
    .N1END(Tile_X1Y9_N1BEG),
    .N2MID(Tile_X1Y9_N2BEG),
    .N2END(Tile_X1Y9_N2BEGb),
    .N4END(Tile_X1Y9_N4BEG),
    .NN4END(Tile_X1Y9_NN4BEG),
    .Ci(Tile_X1Y9_Co),
    .E1END(Tile_X0Y8_E1BEG),
    .E2MID(Tile_X0Y8_E2BEG),
    .E2END(Tile_X0Y8_E2BEGb),
    .EE4END(Tile_X0Y8_EE4BEG),
    .E6END(Tile_X0Y8_E6BEG),
    .S1END(Tile_X1Y7_S1BEG),
    .S2MID(Tile_X1Y7_S2BEG),
    .S2END(Tile_X1Y7_S2BEGb),
    .S4END(Tile_X1Y7_S4BEG),
    .SS4END(Tile_X1Y7_SS4BEG),
    .W1END(Tile_X2Y8_W1BEG),
    .W2MID(Tile_X2Y8_W2BEG),
    .W2END(Tile_X2Y8_W2BEGb),
    .WW4END(Tile_X2Y8_WW4BEG),
    .W6END(Tile_X2Y8_W6BEG),
    .N1BEG(Tile_X1Y8_N1BEG),
    .N2BEG(Tile_X1Y8_N2BEG),
    .N2BEGb(Tile_X1Y8_N2BEGb),
    .N4BEG(Tile_X1Y8_N4BEG),
    .NN4BEG(Tile_X1Y8_NN4BEG),
    .E1BEG(Tile_X1Y8_E1BEG),
    .E2BEG(Tile_X1Y8_E2BEG),
    .E2BEGb(Tile_X1Y8_E2BEGb),
    .EE4BEG(Tile_X1Y8_EE4BEG),
    .E6BEG(Tile_X1Y8_E6BEG),
    .S1BEG(Tile_X1Y8_S1BEG),
    .S2BEG(Tile_X1Y8_S2BEG),
    .S2BEGb(Tile_X1Y8_S2BEGb),
    .S4BEG(Tile_X1Y8_S4BEG),
    .SS4BEG(Tile_X1Y8_SS4BEG),
    .W1BEG(Tile_X1Y8_W1BEG),
    .W2BEG(Tile_X1Y8_W2BEG),
    .W2BEGb(Tile_X1Y8_W2BEGb),
    .WW4BEG(Tile_X1Y8_WW4BEG),
    .W6BEG(Tile_X1Y8_W6BEG),
    .Co(Tile_X1Y8_Co),
    .UserCLK(Tile_X1Y9_UserCLKo),
    .UserCLKo(Tile_X1Y8_UserCLKo),
    .FrameData(Tile_X0Y8_FrameData_O),
    .FrameData_O(Tile_X1Y8_FrameData_O),
    .FrameStrobe(Tile_X1Y9_FrameStrobe_O),
    .FrameStrobe_O(Tile_X1Y8_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X2Y8_Emulate_Bitstream)
    )
`endif
    Tile_X2Y8_LUT4AB
    (
    .N1END(Tile_X2Y9_N1BEG),
    .N2MID(Tile_X2Y9_N2BEG),
    .N2END(Tile_X2Y9_N2BEGb),
    .N4END(Tile_X2Y9_N4BEG),
    .NN4END(Tile_X2Y9_NN4BEG),
    .Ci(Tile_X2Y9_Co),
    .E1END(Tile_X1Y8_E1BEG),
    .E2MID(Tile_X1Y8_E2BEG),
    .E2END(Tile_X1Y8_E2BEGb),
    .EE4END(Tile_X1Y8_EE4BEG),
    .E6END(Tile_X1Y8_E6BEG),
    .S1END(Tile_X2Y7_S1BEG),
    .S2MID(Tile_X2Y7_S2BEG),
    .S2END(Tile_X2Y7_S2BEGb),
    .S4END(Tile_X2Y7_S4BEG),
    .SS4END(Tile_X2Y7_SS4BEG),
    .W1END(Tile_X3Y8_W1BEG),
    .W2MID(Tile_X3Y8_W2BEG),
    .W2END(Tile_X3Y8_W2BEGb),
    .WW4END(Tile_X3Y8_WW4BEG),
    .W6END(Tile_X3Y8_W6BEG),
    .N1BEG(Tile_X2Y8_N1BEG),
    .N2BEG(Tile_X2Y8_N2BEG),
    .N2BEGb(Tile_X2Y8_N2BEGb),
    .N4BEG(Tile_X2Y8_N4BEG),
    .NN4BEG(Tile_X2Y8_NN4BEG),
    .E1BEG(Tile_X2Y8_E1BEG),
    .E2BEG(Tile_X2Y8_E2BEG),
    .E2BEGb(Tile_X2Y8_E2BEGb),
    .EE4BEG(Tile_X2Y8_EE4BEG),
    .E6BEG(Tile_X2Y8_E6BEG),
    .S1BEG(Tile_X2Y8_S1BEG),
    .S2BEG(Tile_X2Y8_S2BEG),
    .S2BEGb(Tile_X2Y8_S2BEGb),
    .S4BEG(Tile_X2Y8_S4BEG),
    .SS4BEG(Tile_X2Y8_SS4BEG),
    .W1BEG(Tile_X2Y8_W1BEG),
    .W2BEG(Tile_X2Y8_W2BEG),
    .W2BEGb(Tile_X2Y8_W2BEGb),
    .WW4BEG(Tile_X2Y8_WW4BEG),
    .W6BEG(Tile_X2Y8_W6BEG),
    .Co(Tile_X2Y8_Co),
    .UserCLK(Tile_X2Y9_UserCLKo),
    .UserCLKo(Tile_X2Y8_UserCLKo),
    .FrameData(Tile_X1Y8_FrameData_O),
    .FrameData_O(Tile_X2Y8_FrameData_O),
    .FrameStrobe(Tile_X2Y9_FrameStrobe_O),
    .FrameStrobe_O(Tile_X2Y8_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X3Y8_Emulate_Bitstream)
    )
`endif
    Tile_X3Y8_LUT4AB
    (
    .N1END(Tile_X3Y9_N1BEG),
    .N2MID(Tile_X3Y9_N2BEG),
    .N2END(Tile_X3Y9_N2BEGb),
    .N4END(Tile_X3Y9_N4BEG),
    .NN4END(Tile_X3Y9_NN4BEG),
    .Ci(Tile_X3Y9_Co),
    .E1END(Tile_X2Y8_E1BEG),
    .E2MID(Tile_X2Y8_E2BEG),
    .E2END(Tile_X2Y8_E2BEGb),
    .EE4END(Tile_X2Y8_EE4BEG),
    .E6END(Tile_X2Y8_E6BEG),
    .S1END(Tile_X3Y7_S1BEG),
    .S2MID(Tile_X3Y7_S2BEG),
    .S2END(Tile_X3Y7_S2BEGb),
    .S4END(Tile_X3Y7_S4BEG),
    .SS4END(Tile_X3Y7_SS4BEG),
    .W1END(Tile_X4Y8_W1BEG),
    .W2MID(Tile_X4Y8_W2BEG),
    .W2END(Tile_X4Y8_W2BEGb),
    .WW4END(Tile_X4Y8_WW4BEG),
    .W6END(Tile_X4Y8_W6BEG),
    .N1BEG(Tile_X3Y8_N1BEG),
    .N2BEG(Tile_X3Y8_N2BEG),
    .N2BEGb(Tile_X3Y8_N2BEGb),
    .N4BEG(Tile_X3Y8_N4BEG),
    .NN4BEG(Tile_X3Y8_NN4BEG),
    .E1BEG(Tile_X3Y8_E1BEG),
    .E2BEG(Tile_X3Y8_E2BEG),
    .E2BEGb(Tile_X3Y8_E2BEGb),
    .EE4BEG(Tile_X3Y8_EE4BEG),
    .E6BEG(Tile_X3Y8_E6BEG),
    .S1BEG(Tile_X3Y8_S1BEG),
    .S2BEG(Tile_X3Y8_S2BEG),
    .S2BEGb(Tile_X3Y8_S2BEGb),
    .S4BEG(Tile_X3Y8_S4BEG),
    .SS4BEG(Tile_X3Y8_SS4BEG),
    .W1BEG(Tile_X3Y8_W1BEG),
    .W2BEG(Tile_X3Y8_W2BEG),
    .W2BEGb(Tile_X3Y8_W2BEGb),
    .WW4BEG(Tile_X3Y8_WW4BEG),
    .W6BEG(Tile_X3Y8_W6BEG),
    .Co(Tile_X3Y8_Co),
    .UserCLK(Tile_X3Y9_UserCLKo),
    .UserCLKo(Tile_X3Y8_UserCLKo),
    .FrameData(Tile_X2Y8_FrameData_O),
    .FrameData_O(Tile_X3Y8_FrameData_O),
    .FrameStrobe(Tile_X3Y9_FrameStrobe_O),
    .FrameStrobe_O(Tile_X3Y8_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
LUT4AB
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X4Y8_Emulate_Bitstream)
    )
`endif
    Tile_X4Y8_LUT4AB
    (
    .N1END(Tile_X4Y9_N1BEG),
    .N2MID(Tile_X4Y9_N2BEG),
    .N2END(Tile_X4Y9_N2BEGb),
    .N4END(Tile_X4Y9_N4BEG),
    .NN4END(Tile_X4Y9_NN4BEG),
    .Ci(Tile_X4Y9_Co),
    .E1END(Tile_X3Y8_E1BEG),
    .E2MID(Tile_X3Y8_E2BEG),
    .E2END(Tile_X3Y8_E2BEGb),
    .EE4END(Tile_X3Y8_EE4BEG),
    .E6END(Tile_X3Y8_E6BEG),
    .S1END(Tile_X4Y7_S1BEG),
    .S2MID(Tile_X4Y7_S2BEG),
    .S2END(Tile_X4Y7_S2BEGb),
    .S4END(Tile_X4Y7_S4BEG),
    .SS4END(Tile_X4Y7_SS4BEG),
    .W1END(Tile_X5Y8_W1BEG),
    .W2MID(Tile_X5Y8_W2BEG),
    .W2END(Tile_X5Y8_W2BEGb),
    .WW4END(Tile_X5Y8_WW4BEG),
    .W6END(Tile_X5Y8_W6BEG),
    .N1BEG(Tile_X4Y8_N1BEG),
    .N2BEG(Tile_X4Y8_N2BEG),
    .N2BEGb(Tile_X4Y8_N2BEGb),
    .N4BEG(Tile_X4Y8_N4BEG),
    .NN4BEG(Tile_X4Y8_NN4BEG),
    .E1BEG(Tile_X4Y8_E1BEG),
    .E2BEG(Tile_X4Y8_E2BEG),
    .E2BEGb(Tile_X4Y8_E2BEGb),
    .EE4BEG(Tile_X4Y8_EE4BEG),
    .E6BEG(Tile_X4Y8_E6BEG),
    .S1BEG(Tile_X4Y8_S1BEG),
    .S2BEG(Tile_X4Y8_S2BEG),
    .S2BEGb(Tile_X4Y8_S2BEGb),
    .S4BEG(Tile_X4Y8_S4BEG),
    .SS4BEG(Tile_X4Y8_SS4BEG),
    .W1BEG(Tile_X4Y8_W1BEG),
    .W2BEG(Tile_X4Y8_W2BEG),
    .W2BEGb(Tile_X4Y8_W2BEGb),
    .WW4BEG(Tile_X4Y8_WW4BEG),
    .W6BEG(Tile_X4Y8_W6BEG),
    .Co(Tile_X4Y8_Co),
    .UserCLK(Tile_X4Y9_UserCLKo),
    .UserCLKo(Tile_X4Y8_UserCLKo),
    .FrameData(Tile_X3Y8_FrameData_O),
    .FrameData_O(Tile_X4Y8_FrameData_O),
    .FrameStrobe(Tile_X4Y9_FrameStrobe_O),
    .FrameStrobe_O(Tile_X4Y8_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
E_TT_IF
`ifdef EMULATION
    #(
    .Emulate_Bitstream(`Tile_X5Y8_Emulate_Bitstream)
    )
`endif
    Tile_X5Y8_E_TT_IF
    (
    .N1END(Tile_X5Y9_N1BEG),
    .N2MID(Tile_X5Y9_N2BEG),
    .N2END(Tile_X5Y9_N2BEGb),
    .N4END(Tile_X5Y9_N4BEG),
    .E1END(Tile_X4Y8_E1BEG),
    .E2MID(Tile_X4Y8_E2BEG),
    .E2END(Tile_X4Y8_E2BEGb),
    .EE4END(Tile_X4Y8_EE4BEG),
    .E6END(Tile_X4Y8_E6BEG),
    .S1END(Tile_X5Y7_S1BEG),
    .S2MID(Tile_X5Y7_S2BEG),
    .S2END(Tile_X5Y7_S2BEGb),
    .S4END(Tile_X5Y7_S4BEG),
    .N1BEG(Tile_X5Y8_N1BEG),
    .N2BEG(Tile_X5Y8_N2BEG),
    .N2BEGb(Tile_X5Y8_N2BEGb),
    .N4BEG(Tile_X5Y8_N4BEG),
    .S1BEG(Tile_X5Y8_S1BEG),
    .S2BEG(Tile_X5Y8_S2BEG),
    .S2BEGb(Tile_X5Y8_S2BEGb),
    .S4BEG(Tile_X5Y8_S4BEG),
    .W1BEG(Tile_X5Y8_W1BEG),
    .W2BEG(Tile_X5Y8_W2BEG),
    .W2BEGb(Tile_X5Y8_W2BEGb),
    .WW4BEG(Tile_X5Y8_WW4BEG),
    .W6BEG(Tile_X5Y8_W6BEG),
    .UO_OUT_TT_PROJECT0(Tile_X5Y8_UO_OUT_TT_PROJECT0),
    .UO_OUT_TT_PROJECT1(Tile_X5Y8_UO_OUT_TT_PROJECT1),
    .UO_OUT_TT_PROJECT2(Tile_X5Y8_UO_OUT_TT_PROJECT2),
    .UO_OUT_TT_PROJECT3(Tile_X5Y8_UO_OUT_TT_PROJECT3),
    .UO_OUT_TT_PROJECT4(Tile_X5Y8_UO_OUT_TT_PROJECT4),
    .UO_OUT_TT_PROJECT5(Tile_X5Y8_UO_OUT_TT_PROJECT5),
    .UO_OUT_TT_PROJECT6(Tile_X5Y8_UO_OUT_TT_PROJECT6),
    .UO_OUT_TT_PROJECT7(Tile_X5Y8_UO_OUT_TT_PROJECT7),
    .UIO_OUT_TT_PROJECT0(Tile_X5Y8_UIO_OUT_TT_PROJECT0),
    .UIO_OUT_TT_PROJECT1(Tile_X5Y8_UIO_OUT_TT_PROJECT1),
    .UIO_OUT_TT_PROJECT2(Tile_X5Y8_UIO_OUT_TT_PROJECT2),
    .UIO_OUT_TT_PROJECT3(Tile_X5Y8_UIO_OUT_TT_PROJECT3),
    .UIO_OUT_TT_PROJECT4(Tile_X5Y8_UIO_OUT_TT_PROJECT4),
    .UIO_OUT_TT_PROJECT5(Tile_X5Y8_UIO_OUT_TT_PROJECT5),
    .UIO_OUT_TT_PROJECT6(Tile_X5Y8_UIO_OUT_TT_PROJECT6),
    .UIO_OUT_TT_PROJECT7(Tile_X5Y8_UIO_OUT_TT_PROJECT7),
    .UIO_OE_TT_PROJECT0(Tile_X5Y8_UIO_OE_TT_PROJECT0),
    .UIO_OE_TT_PROJECT1(Tile_X5Y8_UIO_OE_TT_PROJECT1),
    .UIO_OE_TT_PROJECT2(Tile_X5Y8_UIO_OE_TT_PROJECT2),
    .UIO_OE_TT_PROJECT3(Tile_X5Y8_UIO_OE_TT_PROJECT3),
    .UIO_OE_TT_PROJECT4(Tile_X5Y8_UIO_OE_TT_PROJECT4),
    .UIO_OE_TT_PROJECT5(Tile_X5Y8_UIO_OE_TT_PROJECT5),
    .UIO_OE_TT_PROJECT6(Tile_X5Y8_UIO_OE_TT_PROJECT6),
    .UIO_OE_TT_PROJECT7(Tile_X5Y8_UIO_OE_TT_PROJECT7),
    .UI_IN_TT_PROJECT0(Tile_X5Y8_UI_IN_TT_PROJECT0),
    .UI_IN_TT_PROJECT1(Tile_X5Y8_UI_IN_TT_PROJECT1),
    .UI_IN_TT_PROJECT2(Tile_X5Y8_UI_IN_TT_PROJECT2),
    .UI_IN_TT_PROJECT3(Tile_X5Y8_UI_IN_TT_PROJECT3),
    .UI_IN_TT_PROJECT4(Tile_X5Y8_UI_IN_TT_PROJECT4),
    .UI_IN_TT_PROJECT5(Tile_X5Y8_UI_IN_TT_PROJECT5),
    .UI_IN_TT_PROJECT6(Tile_X5Y8_UI_IN_TT_PROJECT6),
    .UI_IN_TT_PROJECT7(Tile_X5Y8_UI_IN_TT_PROJECT7),
    .UIO_IN_TT_PROJECT0(Tile_X5Y8_UIO_IN_TT_PROJECT0),
    .UIO_IN_TT_PROJECT1(Tile_X5Y8_UIO_IN_TT_PROJECT1),
    .UIO_IN_TT_PROJECT2(Tile_X5Y8_UIO_IN_TT_PROJECT2),
    .UIO_IN_TT_PROJECT3(Tile_X5Y8_UIO_IN_TT_PROJECT3),
    .UIO_IN_TT_PROJECT4(Tile_X5Y8_UIO_IN_TT_PROJECT4),
    .UIO_IN_TT_PROJECT5(Tile_X5Y8_UIO_IN_TT_PROJECT5),
    .UIO_IN_TT_PROJECT6(Tile_X5Y8_UIO_IN_TT_PROJECT6),
    .UIO_IN_TT_PROJECT7(Tile_X5Y8_UIO_IN_TT_PROJECT7),
    .ENA_TT_PROJECT(Tile_X5Y8_ENA_TT_PROJECT),
    .CLK_TT_PROJECT(Tile_X5Y8_CLK_TT_PROJECT),
    .RST_N_TT_PROJECT(Tile_X5Y8_RST_N_TT_PROJECT),
    .UserCLK(Tile_X5Y9_UserCLKo),
    .UserCLKo(Tile_X5Y8_UserCLKo),
    .FrameData(Tile_X4Y8_FrameData_O),
    .FrameData_O(Tile_X5Y8_FrameData_O),
    .FrameStrobe(Tile_X5Y9_FrameStrobe_O),
    .FrameStrobe_O(Tile_X5Y8_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
SW_term Tile_X0Y9_SW_term (
    .S1END(Tile_X0Y8_S1BEG),
    .S2MID(Tile_X0Y8_S2BEG),
    .S2END(Tile_X0Y8_S2BEGb),
    .S4END(Tile_X0Y8_S4BEG),
    .N1BEG(Tile_X0Y9_N1BEG),
    .N2BEG(Tile_X0Y9_N2BEG),
    .N2BEGb(Tile_X0Y9_N2BEGb),
    .N4BEG(Tile_X0Y9_N4BEG),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X0Y9_UserCLKo),
    .FrameData(Row_Y9_FrameData),
    .FrameData_O(Tile_X0Y9_FrameData_O),
    .FrameStrobe(Column_X0_FrameStrobe),
    .FrameStrobe_O(Tile_X0Y9_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_IO4 Tile_X1Y9_S_IO4 (
    .S1END(Tile_X1Y8_S1BEG),
    .S2MID(Tile_X1Y8_S2BEG),
    .S2END(Tile_X1Y8_S2BEGb),
    .S4END(Tile_X1Y8_S4BEG),
    .SS4END(Tile_X1Y8_SS4BEG),
    .N1BEG(Tile_X1Y9_N1BEG),
    .N2BEG(Tile_X1Y9_N2BEG),
    .N2BEGb(Tile_X1Y9_N2BEGb),
    .N4BEG(Tile_X1Y9_N4BEG),
    .NN4BEG(Tile_X1Y9_NN4BEG),
    .Co(Tile_X1Y9_Co),
    .A_O_top(Tile_X1Y9_A_O_top),
    .A_I_top(Tile_X1Y9_A_I_top),
    .A_T_top(Tile_X1Y9_A_T_top),
    .B_O_top(Tile_X1Y9_B_O_top),
    .B_I_top(Tile_X1Y9_B_I_top),
    .B_T_top(Tile_X1Y9_B_T_top),
    .C_O_top(Tile_X1Y9_C_O_top),
    .C_I_top(Tile_X1Y9_C_I_top),
    .C_T_top(Tile_X1Y9_C_T_top),
    .D_O_top(Tile_X1Y9_D_O_top),
    .D_I_top(Tile_X1Y9_D_I_top),
    .D_T_top(Tile_X1Y9_D_T_top),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X1Y9_UserCLKo),
    .FrameData(Tile_X0Y9_FrameData_O),
    .FrameData_O(Tile_X1Y9_FrameData_O),
    .FrameStrobe(Column_X1_FrameStrobe),
    .FrameStrobe_O(Tile_X1Y9_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_IO4 Tile_X2Y9_S_IO4 (
    .S1END(Tile_X2Y8_S1BEG),
    .S2MID(Tile_X2Y8_S2BEG),
    .S2END(Tile_X2Y8_S2BEGb),
    .S4END(Tile_X2Y8_S4BEG),
    .SS4END(Tile_X2Y8_SS4BEG),
    .N1BEG(Tile_X2Y9_N1BEG),
    .N2BEG(Tile_X2Y9_N2BEG),
    .N2BEGb(Tile_X2Y9_N2BEGb),
    .N4BEG(Tile_X2Y9_N4BEG),
    .NN4BEG(Tile_X2Y9_NN4BEG),
    .Co(Tile_X2Y9_Co),
    .A_O_top(Tile_X2Y9_A_O_top),
    .A_I_top(Tile_X2Y9_A_I_top),
    .A_T_top(Tile_X2Y9_A_T_top),
    .B_O_top(Tile_X2Y9_B_O_top),
    .B_I_top(Tile_X2Y9_B_I_top),
    .B_T_top(Tile_X2Y9_B_T_top),
    .C_O_top(Tile_X2Y9_C_O_top),
    .C_I_top(Tile_X2Y9_C_I_top),
    .C_T_top(Tile_X2Y9_C_T_top),
    .D_O_top(Tile_X2Y9_D_O_top),
    .D_I_top(Tile_X2Y9_D_I_top),
    .D_T_top(Tile_X2Y9_D_T_top),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X2Y9_UserCLKo),
    .FrameData(Tile_X1Y9_FrameData_O),
    .FrameData_O(Tile_X2Y9_FrameData_O),
    .FrameStrobe(Column_X2_FrameStrobe),
    .FrameStrobe_O(Tile_X2Y9_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_IO4 Tile_X3Y9_S_IO4 (
    .S1END(Tile_X3Y8_S1BEG),
    .S2MID(Tile_X3Y8_S2BEG),
    .S2END(Tile_X3Y8_S2BEGb),
    .S4END(Tile_X3Y8_S4BEG),
    .SS4END(Tile_X3Y8_SS4BEG),
    .N1BEG(Tile_X3Y9_N1BEG),
    .N2BEG(Tile_X3Y9_N2BEG),
    .N2BEGb(Tile_X3Y9_N2BEGb),
    .N4BEG(Tile_X3Y9_N4BEG),
    .NN4BEG(Tile_X3Y9_NN4BEG),
    .Co(Tile_X3Y9_Co),
    .A_O_top(Tile_X3Y9_A_O_top),
    .A_I_top(Tile_X3Y9_A_I_top),
    .A_T_top(Tile_X3Y9_A_T_top),
    .B_O_top(Tile_X3Y9_B_O_top),
    .B_I_top(Tile_X3Y9_B_I_top),
    .B_T_top(Tile_X3Y9_B_T_top),
    .C_O_top(Tile_X3Y9_C_O_top),
    .C_I_top(Tile_X3Y9_C_I_top),
    .C_T_top(Tile_X3Y9_C_T_top),
    .D_O_top(Tile_X3Y9_D_O_top),
    .D_I_top(Tile_X3Y9_D_I_top),
    .D_T_top(Tile_X3Y9_D_T_top),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X3Y9_UserCLKo),
    .FrameData(Tile_X2Y9_FrameData_O),
    .FrameData_O(Tile_X3Y9_FrameData_O),
    .FrameStrobe(Column_X3_FrameStrobe),
    .FrameStrobe_O(Tile_X3Y9_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
S_IO4 Tile_X4Y9_S_IO4 (
    .S1END(Tile_X4Y8_S1BEG),
    .S2MID(Tile_X4Y8_S2BEG),
    .S2END(Tile_X4Y8_S2BEGb),
    .S4END(Tile_X4Y8_S4BEG),
    .SS4END(Tile_X4Y8_SS4BEG),
    .N1BEG(Tile_X4Y9_N1BEG),
    .N2BEG(Tile_X4Y9_N2BEG),
    .N2BEGb(Tile_X4Y9_N2BEGb),
    .N4BEG(Tile_X4Y9_N4BEG),
    .NN4BEG(Tile_X4Y9_NN4BEG),
    .Co(Tile_X4Y9_Co),
    .A_O_top(Tile_X4Y9_A_O_top),
    .A_I_top(Tile_X4Y9_A_I_top),
    .A_T_top(Tile_X4Y9_A_T_top),
    .B_O_top(Tile_X4Y9_B_O_top),
    .B_I_top(Tile_X4Y9_B_I_top),
    .B_T_top(Tile_X4Y9_B_T_top),
    .C_O_top(Tile_X4Y9_C_O_top),
    .C_I_top(Tile_X4Y9_C_I_top),
    .C_T_top(Tile_X4Y9_C_T_top),
    .D_O_top(Tile_X4Y9_D_O_top),
    .D_I_top(Tile_X4Y9_D_I_top),
    .D_T_top(Tile_X4Y9_D_T_top),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X4Y9_UserCLKo),
    .FrameData(Tile_X3Y9_FrameData_O),
    .FrameData_O(Tile_X4Y9_FrameData_O),
    .FrameStrobe(Column_X4_FrameStrobe),
    .FrameStrobe_O(Tile_X4Y9_FrameStrobe_O)
);


 //tile IO port will get directly connected to top-level tile module
SE_term Tile_X5Y9_SE_term (
    .S1END(Tile_X5Y8_S1BEG),
    .S2MID(Tile_X5Y8_S2BEG),
    .S2END(Tile_X5Y8_S2BEGb),
    .S4END(Tile_X5Y8_S4BEG),
    .N1BEG(Tile_X5Y9_N1BEG),
    .N2BEG(Tile_X5Y9_N2BEG),
    .N2BEGb(Tile_X5Y9_N2BEGb),
    .N4BEG(Tile_X5Y9_N4BEG),
    .UserCLK(UserCLK),
    .UserCLKo(Tile_X5Y9_UserCLKo),
    .FrameData(Tile_X4Y9_FrameData_O),
    .FrameData_O(Tile_X5Y9_FrameData_O),
    .FrameStrobe(Column_X5_FrameStrobe),
    .FrameStrobe_O(Tile_X5Y9_FrameStrobe_O)
);

endmodule