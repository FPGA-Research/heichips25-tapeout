module W_TT_IF (CLK_TT_PROJECT,
    ENA_TT_PROJECT,
    RST_N_TT_PROJECT,
    UIO_IN_TT_PROJECT0,
    UIO_IN_TT_PROJECT1,
    UIO_IN_TT_PROJECT2,
    UIO_IN_TT_PROJECT3,
    UIO_IN_TT_PROJECT4,
    UIO_IN_TT_PROJECT5,
    UIO_IN_TT_PROJECT6,
    UIO_IN_TT_PROJECT7,
    UIO_OE_TT_PROJECT0,
    UIO_OE_TT_PROJECT1,
    UIO_OE_TT_PROJECT2,
    UIO_OE_TT_PROJECT3,
    UIO_OE_TT_PROJECT4,
    UIO_OE_TT_PROJECT5,
    UIO_OE_TT_PROJECT6,
    UIO_OE_TT_PROJECT7,
    UIO_OUT_TT_PROJECT0,
    UIO_OUT_TT_PROJECT1,
    UIO_OUT_TT_PROJECT2,
    UIO_OUT_TT_PROJECT3,
    UIO_OUT_TT_PROJECT4,
    UIO_OUT_TT_PROJECT5,
    UIO_OUT_TT_PROJECT6,
    UIO_OUT_TT_PROJECT7,
    UI_IN_TT_PROJECT0,
    UI_IN_TT_PROJECT1,
    UI_IN_TT_PROJECT2,
    UI_IN_TT_PROJECT3,
    UI_IN_TT_PROJECT4,
    UI_IN_TT_PROJECT5,
    UI_IN_TT_PROJECT6,
    UI_IN_TT_PROJECT7,
    UO_OUT_TT_PROJECT0,
    UO_OUT_TT_PROJECT1,
    UO_OUT_TT_PROJECT2,
    UO_OUT_TT_PROJECT3,
    UO_OUT_TT_PROJECT4,
    UO_OUT_TT_PROJECT5,
    UO_OUT_TT_PROJECT6,
    UO_OUT_TT_PROJECT7,
    UserCLK,
    UserCLKo,
    E1BEG,
    E2BEG,
    E2BEGb,
    E6BEG,
    EE4BEG,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N1END,
    N2BEG,
    N2BEGb,
    N2END,
    N2MID,
    N4BEG,
    N4END,
    S1BEG,
    S1END,
    S2BEG,
    S2BEGb,
    S2END,
    S2MID,
    S4BEG,
    S4END,
    W1END,
    W2END,
    W2MID,
    W6END,
    WW4END);
 output CLK_TT_PROJECT;
 output ENA_TT_PROJECT;
 output RST_N_TT_PROJECT;
 output UIO_IN_TT_PROJECT0;
 output UIO_IN_TT_PROJECT1;
 output UIO_IN_TT_PROJECT2;
 output UIO_IN_TT_PROJECT3;
 output UIO_IN_TT_PROJECT4;
 output UIO_IN_TT_PROJECT5;
 output UIO_IN_TT_PROJECT6;
 output UIO_IN_TT_PROJECT7;
 input UIO_OE_TT_PROJECT0;
 input UIO_OE_TT_PROJECT1;
 input UIO_OE_TT_PROJECT2;
 input UIO_OE_TT_PROJECT3;
 input UIO_OE_TT_PROJECT4;
 input UIO_OE_TT_PROJECT5;
 input UIO_OE_TT_PROJECT6;
 input UIO_OE_TT_PROJECT7;
 input UIO_OUT_TT_PROJECT0;
 input UIO_OUT_TT_PROJECT1;
 input UIO_OUT_TT_PROJECT2;
 input UIO_OUT_TT_PROJECT3;
 input UIO_OUT_TT_PROJECT4;
 input UIO_OUT_TT_PROJECT5;
 input UIO_OUT_TT_PROJECT6;
 input UIO_OUT_TT_PROJECT7;
 output UI_IN_TT_PROJECT0;
 output UI_IN_TT_PROJECT1;
 output UI_IN_TT_PROJECT2;
 output UI_IN_TT_PROJECT3;
 output UI_IN_TT_PROJECT4;
 output UI_IN_TT_PROJECT5;
 output UI_IN_TT_PROJECT6;
 output UI_IN_TT_PROJECT7;
 input UO_OUT_TT_PROJECT0;
 input UO_OUT_TT_PROJECT1;
 input UO_OUT_TT_PROJECT2;
 input UO_OUT_TT_PROJECT3;
 input UO_OUT_TT_PROJECT4;
 input UO_OUT_TT_PROJECT5;
 input UO_OUT_TT_PROJECT6;
 input UO_OUT_TT_PROJECT7;
 input UserCLK;
 output UserCLKo;
 output [3:0] E1BEG;
 output [7:0] E2BEG;
 output [7:0] E2BEGb;
 output [11:0] E6BEG;
 output [15:0] EE4BEG;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 input [3:0] N1END;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 input [7:0] N2END;
 input [7:0] N2MID;
 output [15:0] N4BEG;
 input [15:0] N4END;
 output [3:0] S1BEG;
 input [3:0] S1END;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 input [7:0] S2END;
 input [7:0] S2MID;
 output [15:0] S4BEG;
 input [15:0] S4END;
 input [3:0] W1END;
 input [7:0] W2END;
 input [7:0] W2MID;
 input [11:0] W6END;
 input [15:0] WW4END;

 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit0.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit1.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit2.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit3.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit4.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit5.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit6.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit7.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit10.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit11.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit12.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit13.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit14.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit15.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit16.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit17.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit18.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit19.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit20.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit21.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit22.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit23.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit24.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit25.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit26.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit27.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit28.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit29.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit30.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit31.Q ;
 wire \Inst_W_TT_IF_switch_matrix.E1BEG0 ;
 wire \Inst_W_TT_IF_switch_matrix.E1BEG1 ;
 wire \Inst_W_TT_IF_switch_matrix.E1BEG2 ;
 wire \Inst_W_TT_IF_switch_matrix.E1BEG3 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEG0 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEG1 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEG2 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEG3 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEG4 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEG5 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEG6 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEG7 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEGb0 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEGb1 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEGb2 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEGb3 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEGb4 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEGb5 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEGb6 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEGb7 ;
 wire \Inst_W_TT_IF_switch_matrix.E6BEG0 ;
 wire \Inst_W_TT_IF_switch_matrix.E6BEG1 ;
 wire \Inst_W_TT_IF_switch_matrix.E6BEG10 ;
 wire \Inst_W_TT_IF_switch_matrix.E6BEG11 ;
 wire \Inst_W_TT_IF_switch_matrix.E6BEG2 ;
 wire \Inst_W_TT_IF_switch_matrix.E6BEG3 ;
 wire \Inst_W_TT_IF_switch_matrix.E6BEG4 ;
 wire \Inst_W_TT_IF_switch_matrix.E6BEG5 ;
 wire \Inst_W_TT_IF_switch_matrix.E6BEG6 ;
 wire \Inst_W_TT_IF_switch_matrix.E6BEG7 ;
 wire \Inst_W_TT_IF_switch_matrix.E6BEG8 ;
 wire \Inst_W_TT_IF_switch_matrix.E6BEG9 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG0 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG1 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG10 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG11 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG12 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG13 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG14 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG15 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG2 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG3 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG4 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG5 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG6 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG7 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG8 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG9 ;
 wire \Inst_W_TT_IF_switch_matrix.N1BEG0 ;
 wire \Inst_W_TT_IF_switch_matrix.N1BEG1 ;
 wire \Inst_W_TT_IF_switch_matrix.N1BEG2 ;
 wire \Inst_W_TT_IF_switch_matrix.N1BEG3 ;
 wire \Inst_W_TT_IF_switch_matrix.N2BEG0 ;
 wire \Inst_W_TT_IF_switch_matrix.N2BEG1 ;
 wire \Inst_W_TT_IF_switch_matrix.N2BEG2 ;
 wire \Inst_W_TT_IF_switch_matrix.N2BEG3 ;
 wire \Inst_W_TT_IF_switch_matrix.N2BEG4 ;
 wire \Inst_W_TT_IF_switch_matrix.N2BEG5 ;
 wire \Inst_W_TT_IF_switch_matrix.N2BEG6 ;
 wire \Inst_W_TT_IF_switch_matrix.N2BEG7 ;
 wire \Inst_W_TT_IF_switch_matrix.N4BEG0 ;
 wire \Inst_W_TT_IF_switch_matrix.N4BEG1 ;
 wire \Inst_W_TT_IF_switch_matrix.N4BEG2 ;
 wire \Inst_W_TT_IF_switch_matrix.N4BEG3 ;
 wire \Inst_W_TT_IF_switch_matrix.S1BEG0 ;
 wire \Inst_W_TT_IF_switch_matrix.S1BEG1 ;
 wire \Inst_W_TT_IF_switch_matrix.S1BEG2 ;
 wire \Inst_W_TT_IF_switch_matrix.S1BEG3 ;
 wire \Inst_W_TT_IF_switch_matrix.S2BEG0 ;
 wire \Inst_W_TT_IF_switch_matrix.S2BEG1 ;
 wire \Inst_W_TT_IF_switch_matrix.S2BEG2 ;
 wire \Inst_W_TT_IF_switch_matrix.S2BEG3 ;
 wire \Inst_W_TT_IF_switch_matrix.S2BEG4 ;
 wire \Inst_W_TT_IF_switch_matrix.S2BEG5 ;
 wire \Inst_W_TT_IF_switch_matrix.S2BEG6 ;
 wire \Inst_W_TT_IF_switch_matrix.S2BEG7 ;
 wire \Inst_W_TT_IF_switch_matrix.S4BEG0 ;
 wire \Inst_W_TT_IF_switch_matrix.S4BEG1 ;
 wire \Inst_W_TT_IF_switch_matrix.S4BEG2 ;
 wire \Inst_W_TT_IF_switch_matrix.S4BEG3 ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire clknet_0_UserCLK;
 wire clknet_1_0__leaf_UserCLK;
 wire clknet_1_1__leaf_UserCLK;

 sg13g2_inv_1 _209_ (.Y(_000_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit5.Q ));
 sg13g2_inv_1 _210_ (.Y(_001_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit6.Q ));
 sg13g2_inv_1 _211_ (.Y(_002_),
    .A(S1END[3]));
 sg13g2_inv_1 _212_ (.Y(_003_),
    .A(S1END[2]));
 sg13g2_inv_1 _213_ (.Y(_004_),
    .A(S1END[1]));
 sg13g2_inv_1 _214_ (.Y(_005_),
    .A(S1END[0]));
 sg13g2_inv_1 _215_ (.Y(_006_),
    .A(WW4END[1]));
 sg13g2_inv_1 _216_ (.Y(_007_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit10.Q ));
 sg13g2_inv_1 _217_ (.Y(_008_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit18.Q ));
 sg13g2_inv_1 _218_ (.Y(_009_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit15.Q ));
 sg13g2_inv_1 _219_ (.Y(_010_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit16.Q ));
 sg13g2_inv_1 _220_ (.Y(_011_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit6.Q ));
 sg13g2_inv_1 _221_ (.Y(_012_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit7.Q ));
 sg13g2_inv_1 _222_ (.Y(_013_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit12.Q ));
 sg13g2_inv_1 _223_ (.Y(_014_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit13.Q ));
 sg13g2_inv_1 _224_ (.Y(_015_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit5.Q ));
 sg13g2_inv_1 _225_ (.Y(_016_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit6.Q ));
 sg13g2_inv_1 _226_ (.Y(_017_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit7.Q ));
 sg13g2_inv_1 _227_ (.Y(_018_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit2.Q ));
 sg13g2_inv_1 _228_ (.Y(_019_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit3.Q ));
 sg13g2_mux2_1 _229_ (.A0(W2END[1]),
    .A1(W2END[2]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_020_));
 sg13g2_nand2_1 _230_ (.Y(_021_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit5.Q ),
    .B(_020_));
 sg13g2_mux2_1 _231_ (.A0(W2MID[3]),
    .A1(W2MID[6]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_022_));
 sg13g2_a21oi_1 _232_ (.A1(_000_),
    .A2(_022_),
    .Y(_023_),
    .B1(_001_));
 sg13g2_mux2_1 _233_ (.A0(N2MID[6]),
    .A1(N2END[2]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_024_));
 sg13g2_nand2b_1 _234_ (.Y(_025_),
    .B(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit4.Q ),
    .A_N(W2MID[0]));
 sg13g2_o21ai_1 _235_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit5.Q ),
    .Y(_026_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit4.Q ),
    .A2(N2END[3]));
 sg13g2_nand2b_1 _236_ (.Y(_027_),
    .B(_025_),
    .A_N(_026_));
 sg13g2_a21oi_1 _237_ (.A1(_000_),
    .A2(_024_),
    .Y(_028_),
    .B1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit6.Q ));
 sg13g2_a221oi_1 _238_ (.B2(_028_),
    .C1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit7.Q ),
    .B1(_027_),
    .A1(_021_),
    .Y(_029_),
    .A2(_023_));
 sg13g2_nor2_1 _239_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit5.Q ),
    .B(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit6.Q ),
    .Y(_030_));
 sg13g2_nor2b_1 _240_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit6.Q ),
    .B_N(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit5.Q ),
    .Y(_031_));
 sg13g2_nor2b_1 _241_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit5.Q ),
    .B_N(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit6.Q ),
    .Y(_032_));
 sg13g2_a22oi_1 _242_ (.Y(_033_),
    .B1(_032_),
    .B2(S2END[2]),
    .A2(_030_),
    .A1(W2END[3]));
 sg13g2_a21oi_1 _243_ (.A1(W2END[5]),
    .A2(_031_),
    .Y(_034_),
    .B1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit4.Q ));
 sg13g2_o21ai_1 _244_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit6.Q ),
    .Y(_035_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit5.Q ),
    .A2(S2END[3]));
 sg13g2_a22oi_1 _245_ (.Y(_036_),
    .B1(_030_),
    .B2(W2END[4]),
    .A2(S2MID[0]),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit5.Q ));
 sg13g2_and2_1 _246_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit4.Q ),
    .B(_035_),
    .X(_037_));
 sg13g2_a22oi_1 _247_ (.Y(_038_),
    .B1(_036_),
    .B2(_037_),
    .A2(_034_),
    .A1(_033_));
 sg13g2_a21o_1 _248_ (.A2(_038_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit7.Q ),
    .B1(_029_),
    .X(RST_N_TT_PROJECT));
 sg13g2_mux4_1 _249_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit22.Q ),
    .A0(N2MID[7]),
    .A1(N2END[7]),
    .A2(S2MID[7]),
    .A3(S2END[7]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit23.Q ),
    .X(_039_));
 sg13g2_inv_1 _250_ (.Y(_040_),
    .A(_039_));
 sg13g2_mux4_1 _251_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit6.Q ),
    .A0(N1END[3]),
    .A1(N4END[3]),
    .A2(S1END[3]),
    .A3(S4END[3]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit7.Q ),
    .X(_041_));
 sg13g2_nor2b_1 _252_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit31.Q ),
    .B_N(WW4END[15]),
    .Y(_042_));
 sg13g2_a21oi_1 _253_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit31.Q ),
    .A2(_041_),
    .Y(_043_),
    .B1(_042_));
 sg13g2_nand3b_1 _254_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit0.Q ),
    .C(_039_),
    .Y(_044_),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit31.Q ));
 sg13g2_o21ai_1 _255_ (.B1(_044_),
    .Y(_045_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit0.Q ),
    .A2(_043_));
 sg13g2_mux4_1 _256_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit31.Q ),
    .A0(W1END[3]),
    .A1(W2MID[7]),
    .A2(W2END[7]),
    .A3(WW4END[7]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit0.Q ),
    .X(_046_));
 sg13g2_mux2_1 _257_ (.A0(_046_),
    .A1(_045_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit1.Q ),
    .X(UIO_IN_TT_PROJECT7));
 sg13g2_mux4_1 _258_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit20.Q ),
    .A0(N2MID[6]),
    .A1(N2END[6]),
    .A2(S2MID[6]),
    .A3(S2END[6]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit21.Q ),
    .X(_047_));
 sg13g2_mux4_1 _259_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit4.Q ),
    .A0(N1END[2]),
    .A1(N4END[2]),
    .A2(S1END[2]),
    .A3(S4END[2]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit5.Q ),
    .X(_048_));
 sg13g2_nor2b_1 _260_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit28.Q ),
    .B_N(WW4END[14]),
    .Y(_049_));
 sg13g2_a21oi_1 _261_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit28.Q ),
    .A2(_048_),
    .Y(_050_),
    .B1(_049_));
 sg13g2_nand3b_1 _262_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit29.Q ),
    .C(_047_),
    .Y(_051_),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit28.Q ));
 sg13g2_o21ai_1 _263_ (.B1(_051_),
    .Y(_052_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit29.Q ),
    .A2(_050_));
 sg13g2_mux4_1 _264_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit29.Q ),
    .A0(W1END[2]),
    .A1(W2END[6]),
    .A2(W2MID[6]),
    .A3(WW4END[6]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit28.Q ),
    .X(_053_));
 sg13g2_mux2_1 _265_ (.A0(_053_),
    .A1(_052_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit30.Q ),
    .X(UIO_IN_TT_PROJECT6));
 sg13g2_mux4_1 _266_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit2.Q ),
    .A0(N1END[1]),
    .A1(N4END[1]),
    .A2(S1END[1]),
    .A3(S4END[1]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit3.Q ),
    .X(_054_));
 sg13g2_mux4_1 _267_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit18.Q ),
    .A0(N2MID[5]),
    .A1(N2END[5]),
    .A2(S2MID[5]),
    .A3(S2END[5]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit19.Q ),
    .X(_055_));
 sg13g2_mux4_1 _268_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit25.Q ),
    .A0(W1END[1]),
    .A1(W2MID[5]),
    .A2(W2END[5]),
    .A3(WW4END[5]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit26.Q ),
    .X(_056_));
 sg13g2_nand3b_1 _269_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit26.Q ),
    .C(_055_),
    .Y(_057_),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit25.Q ));
 sg13g2_nor2b_1 _270_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit25.Q ),
    .B_N(WW4END[13]),
    .Y(_058_));
 sg13g2_a21oi_1 _271_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit25.Q ),
    .A2(_054_),
    .Y(_059_),
    .B1(_058_));
 sg13g2_o21ai_1 _272_ (.B1(_057_),
    .Y(_060_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit26.Q ),
    .A2(_059_));
 sg13g2_mux2_1 _273_ (.A0(_056_),
    .A1(_060_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit27.Q ),
    .X(UIO_IN_TT_PROJECT5));
 sg13g2_mux4_1 _274_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit0.Q ),
    .A0(N1END[0]),
    .A1(N4END[0]),
    .A2(S1END[0]),
    .A3(S4END[0]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit1.Q ),
    .X(_061_));
 sg13g2_mux4_1 _275_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit16.Q ),
    .A0(N2MID[4]),
    .A1(N2END[4]),
    .A2(S2MID[4]),
    .A3(S2END[4]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit17.Q ),
    .X(_062_));
 sg13g2_inv_1 _276_ (.Y(_063_),
    .A(_062_));
 sg13g2_nor2b_1 _277_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit22.Q ),
    .B_N(WW4END[12]),
    .Y(_064_));
 sg13g2_a21oi_1 _278_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit22.Q ),
    .A2(_061_),
    .Y(_065_),
    .B1(_064_));
 sg13g2_nand3b_1 _279_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit23.Q ),
    .C(_062_),
    .Y(_066_),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit22.Q ));
 sg13g2_o21ai_1 _280_ (.B1(_066_),
    .Y(_067_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit23.Q ),
    .A2(_065_));
 sg13g2_mux4_1 _281_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit22.Q ),
    .A0(W1END[0]),
    .A1(W2MID[4]),
    .A2(W2END[4]),
    .A3(WW4END[4]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit23.Q ),
    .X(_068_));
 sg13g2_mux2_1 _282_ (.A0(_068_),
    .A1(_067_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit24.Q ),
    .X(UIO_IN_TT_PROJECT4));
 sg13g2_mux4_1 _283_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit30.Q ),
    .A0(N1END[3]),
    .A1(N4END[3]),
    .A2(S1END[3]),
    .A3(S4END[3]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit31.Q ),
    .X(_069_));
 sg13g2_mux4_1 _284_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit15.Q ),
    .A0(N2MID[3]),
    .A1(S2MID[3]),
    .A2(N2END[3]),
    .A3(S2END[3]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit14.Q ),
    .X(_070_));
 sg13g2_nand3b_1 _285_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit20.Q ),
    .C(_070_),
    .Y(_071_),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit19.Q ));
 sg13g2_nor2b_1 _286_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit19.Q ),
    .B_N(W6END[11]),
    .Y(_072_));
 sg13g2_a21oi_1 _287_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit19.Q ),
    .A2(_069_),
    .Y(_073_),
    .B1(_072_));
 sg13g2_o21ai_1 _288_ (.B1(_071_),
    .Y(_074_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit20.Q ),
    .A2(_073_));
 sg13g2_mux4_1 _289_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit19.Q ),
    .A0(W2MID[3]),
    .A1(W2END[3]),
    .A2(WW4END[3]),
    .A3(WW4END[11]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit20.Q ),
    .X(_075_));
 sg13g2_mux2_1 _290_ (.A0(_075_),
    .A1(_074_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit21.Q ),
    .X(UIO_IN_TT_PROJECT3));
 sg13g2_mux4_1 _291_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit28.Q ),
    .A0(N1END[2]),
    .A1(N4END[2]),
    .A2(S1END[2]),
    .A3(S4END[2]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit29.Q ),
    .X(_076_));
 sg13g2_mux4_1 _292_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit13.Q ),
    .A0(N2MID[2]),
    .A1(S2MID[2]),
    .A2(N2END[2]),
    .A3(S2END[2]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit12.Q ),
    .X(_077_));
 sg13g2_mux4_1 _293_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit17.Q ),
    .A0(W2MID[2]),
    .A1(WW4END[2]),
    .A2(W2END[2]),
    .A3(WW4END[10]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit16.Q ),
    .X(_078_));
 sg13g2_nand3b_1 _294_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit17.Q ),
    .C(_077_),
    .Y(_079_),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit16.Q ));
 sg13g2_nor2b_1 _295_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit16.Q ),
    .B_N(W6END[10]),
    .Y(_080_));
 sg13g2_a21oi_1 _296_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit16.Q ),
    .A2(_076_),
    .Y(_081_),
    .B1(_080_));
 sg13g2_o21ai_1 _297_ (.B1(_079_),
    .Y(_082_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit17.Q ),
    .A2(_081_));
 sg13g2_mux2_1 _298_ (.A0(_078_),
    .A1(_082_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit18.Q ),
    .X(UIO_IN_TT_PROJECT2));
 sg13g2_mux4_1 _299_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit26.Q ),
    .A0(N1END[1]),
    .A1(N4END[1]),
    .A2(S1END[1]),
    .A3(S4END[1]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit27.Q ),
    .X(_083_));
 sg13g2_mux4_1 _300_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit10.Q ),
    .A0(N2MID[1]),
    .A1(N2END[1]),
    .A2(S2MID[1]),
    .A3(S2END[1]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit11.Q ),
    .X(_084_));
 sg13g2_nor2b_1 _301_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit13.Q ),
    .B_N(W6END[9]),
    .Y(_085_));
 sg13g2_a21oi_1 _302_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit13.Q ),
    .A2(_083_),
    .Y(_086_),
    .B1(_085_));
 sg13g2_nand3b_1 _303_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit14.Q ),
    .C(_084_),
    .Y(_087_),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit13.Q ));
 sg13g2_o21ai_1 _304_ (.B1(_087_),
    .Y(_088_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit14.Q ),
    .A2(_086_));
 sg13g2_mux4_1 _305_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit14.Q ),
    .A0(W2MID[1]),
    .A1(WW4END[1]),
    .A2(W2END[1]),
    .A3(WW4END[9]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit13.Q ),
    .X(_089_));
 sg13g2_mux2_1 _306_ (.A0(_089_),
    .A1(_088_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit15.Q ),
    .X(UIO_IN_TT_PROJECT1));
 sg13g2_mux4_1 _307_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit8.Q ),
    .A0(N2MID[0]),
    .A1(N2END[0]),
    .A2(S2MID[0]),
    .A3(S2END[0]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit9.Q ),
    .X(_090_));
 sg13g2_inv_1 _308_ (.Y(_091_),
    .A(_090_));
 sg13g2_mux4_1 _309_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit24.Q ),
    .A0(N1END[0]),
    .A1(N4END[0]),
    .A2(S1END[0]),
    .A3(S4END[0]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit25.Q ),
    .X(_092_));
 sg13g2_inv_1 _310_ (.Y(_093_),
    .A(_092_));
 sg13g2_nand3_1 _311_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit11.Q ),
    .C(_090_),
    .A(_007_),
    .Y(_094_));
 sg13g2_or2_1 _312_ (.X(_095_),
    .B(W6END[8]),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit10.Q ));
 sg13g2_o21ai_1 _313_ (.B1(_095_),
    .Y(_096_),
    .A1(_007_),
    .A2(_092_));
 sg13g2_o21ai_1 _314_ (.B1(_094_),
    .Y(_097_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit11.Q ),
    .A2(_096_));
 sg13g2_mux4_1 _315_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit10.Q ),
    .A0(W2MID[0]),
    .A1(W2END[0]),
    .A2(WW4END[0]),
    .A3(WW4END[8]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit11.Q ),
    .X(_098_));
 sg13g2_mux2_1 _316_ (.A0(_098_),
    .A1(_097_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit12.Q ),
    .X(UIO_IN_TT_PROJECT0));
 sg13g2_mux4_1 _317_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit22.Q ),
    .A0(N1END[3]),
    .A1(N4END[3]),
    .A2(S1END[3]),
    .A3(S4END[3]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit23.Q ),
    .X(_099_));
 sg13g2_mux4_1 _318_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit7.Q ),
    .A0(W2MID[7]),
    .A1(W2END[7]),
    .A2(WW4END[7]),
    .A3(WW4END[15]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit8.Q ),
    .X(_100_));
 sg13g2_nand3b_1 _319_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit8.Q ),
    .C(_039_),
    .Y(_101_),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit7.Q ));
 sg13g2_nor2b_1 _320_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit7.Q ),
    .B_N(W6END[7]),
    .Y(_102_));
 sg13g2_a21oi_1 _321_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit7.Q ),
    .A2(_099_),
    .Y(_103_),
    .B1(_102_));
 sg13g2_o21ai_1 _322_ (.B1(_101_),
    .Y(_104_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit8.Q ),
    .A2(_103_));
 sg13g2_mux2_1 _323_ (.A0(_100_),
    .A1(_104_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit9.Q ),
    .X(UI_IN_TT_PROJECT7));
 sg13g2_mux4_1 _324_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit20.Q ),
    .A0(N1END[2]),
    .A1(N4END[2]),
    .A2(S1END[2]),
    .A3(S4END[2]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit21.Q ),
    .X(_105_));
 sg13g2_mux4_1 _325_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit4.Q ),
    .A0(W2MID[6]),
    .A1(W2END[6]),
    .A2(WW4END[6]),
    .A3(WW4END[14]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit5.Q ),
    .X(_106_));
 sg13g2_nand3b_1 _326_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit5.Q ),
    .C(_047_),
    .Y(_107_),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit4.Q ));
 sg13g2_nor2b_1 _327_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit4.Q ),
    .B_N(W6END[6]),
    .Y(_108_));
 sg13g2_a21oi_1 _328_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit4.Q ),
    .A2(_105_),
    .Y(_109_),
    .B1(_108_));
 sg13g2_o21ai_1 _329_ (.B1(_107_),
    .Y(_110_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit5.Q ),
    .A2(_109_));
 sg13g2_mux2_1 _330_ (.A0(_106_),
    .A1(_110_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit6.Q ),
    .X(UI_IN_TT_PROJECT6));
 sg13g2_mux4_1 _331_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit18.Q ),
    .A0(N1END[1]),
    .A1(N4END[1]),
    .A2(S1END[1]),
    .A3(S4END[1]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit19.Q ),
    .X(_111_));
 sg13g2_nor2b_1 _332_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit1.Q ),
    .B_N(W6END[5]),
    .Y(_112_));
 sg13g2_a21oi_1 _333_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit1.Q ),
    .A2(_111_),
    .Y(_113_),
    .B1(_112_));
 sg13g2_nand3b_1 _334_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit2.Q ),
    .C(_055_),
    .Y(_114_),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit1.Q ));
 sg13g2_o21ai_1 _335_ (.B1(_114_),
    .Y(_115_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit2.Q ),
    .A2(_113_));
 sg13g2_mux4_1 _336_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit2.Q ),
    .A0(W2MID[5]),
    .A1(WW4END[5]),
    .A2(W2END[5]),
    .A3(WW4END[13]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit1.Q ),
    .X(_116_));
 sg13g2_mux2_1 _337_ (.A0(_116_),
    .A1(_115_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit3.Q ),
    .X(UI_IN_TT_PROJECT5));
 sg13g2_mux4_1 _338_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit16.Q ),
    .A0(N1END[0]),
    .A1(N4END[0]),
    .A2(S1END[0]),
    .A3(S4END[0]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit17.Q ),
    .X(_117_));
 sg13g2_nor2b_1 _339_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit30.Q ),
    .B_N(W6END[4]),
    .Y(_118_));
 sg13g2_a21oi_1 _340_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit30.Q ),
    .A2(_117_),
    .Y(_119_),
    .B1(_118_));
 sg13g2_nand3b_1 _341_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit31.Q ),
    .C(_062_),
    .Y(_120_),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit30.Q ));
 sg13g2_o21ai_1 _342_ (.B1(_120_),
    .Y(_121_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit31.Q ),
    .A2(_119_));
 sg13g2_mux4_1 _343_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit31.Q ),
    .A0(W2MID[4]),
    .A1(WW4END[4]),
    .A2(W2END[4]),
    .A3(WW4END[12]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit30.Q ),
    .X(_122_));
 sg13g2_mux2_1 _344_ (.A0(_122_),
    .A1(_121_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit0.Q ),
    .X(UI_IN_TT_PROJECT4));
 sg13g2_mux4_1 _345_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit14.Q ),
    .A0(N1END[3]),
    .A1(N4END[3]),
    .A2(S1END[3]),
    .A3(S4END[3]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit15.Q ),
    .X(_123_));
 sg13g2_mux4_1 _346_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit27.Q ),
    .A0(W2MID[3]),
    .A1(W2END[3]),
    .A2(WW4END[3]),
    .A3(WW4END[11]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit28.Q ),
    .X(_124_));
 sg13g2_nand3b_1 _347_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit28.Q ),
    .C(_070_),
    .Y(_125_),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit27.Q ));
 sg13g2_nor2b_1 _348_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit27.Q ),
    .B_N(W6END[3]),
    .Y(_126_));
 sg13g2_a21oi_1 _349_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit27.Q ),
    .A2(_123_),
    .Y(_127_),
    .B1(_126_));
 sg13g2_o21ai_1 _350_ (.B1(_125_),
    .Y(_128_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit28.Q ),
    .A2(_127_));
 sg13g2_mux2_1 _351_ (.A0(_124_),
    .A1(_128_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit29.Q ),
    .X(UI_IN_TT_PROJECT3));
 sg13g2_mux4_1 _352_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit12.Q ),
    .A0(N1END[2]),
    .A1(N4END[2]),
    .A2(S1END[2]),
    .A3(S4END[2]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_129_));
 sg13g2_mux4_1 _353_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit25.Q ),
    .A0(W2MID[2]),
    .A1(WW4END[2]),
    .A2(W2END[2]),
    .A3(WW4END[10]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit24.Q ),
    .X(_130_));
 sg13g2_nand3b_1 _354_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit25.Q ),
    .C(_077_),
    .Y(_131_),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit24.Q ));
 sg13g2_nor2b_1 _355_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit24.Q ),
    .B_N(W6END[2]),
    .Y(_132_));
 sg13g2_a21oi_1 _356_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit24.Q ),
    .A2(_129_),
    .Y(_133_),
    .B1(_132_));
 sg13g2_o21ai_1 _357_ (.B1(_131_),
    .Y(_134_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit25.Q ),
    .A2(_133_));
 sg13g2_mux2_1 _358_ (.A0(_130_),
    .A1(_134_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit26.Q ),
    .X(UI_IN_TT_PROJECT2));
 sg13g2_mux4_1 _359_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit10.Q ),
    .A0(N1END[1]),
    .A1(N4END[1]),
    .A2(S1END[1]),
    .A3(S4END[1]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit11.Q ),
    .X(_135_));
 sg13g2_nor2b_1 _360_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit21.Q ),
    .B_N(W6END[1]),
    .Y(_136_));
 sg13g2_a21oi_1 _361_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit21.Q ),
    .A2(_135_),
    .Y(_137_),
    .B1(_136_));
 sg13g2_nand3b_1 _362_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit22.Q ),
    .C(_084_),
    .Y(_138_),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit21.Q ));
 sg13g2_o21ai_1 _363_ (.B1(_138_),
    .Y(_139_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit22.Q ),
    .A2(_137_));
 sg13g2_mux4_1 _364_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit22.Q ),
    .A0(W2MID[1]),
    .A1(WW4END[1]),
    .A2(W2END[1]),
    .A3(WW4END[9]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit21.Q ),
    .X(_140_));
 sg13g2_mux2_1 _365_ (.A0(_140_),
    .A1(_139_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit23.Q ),
    .X(UI_IN_TT_PROJECT1));
 sg13g2_mux4_1 _366_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit8.Q ),
    .A0(N1END[0]),
    .A1(N4END[0]),
    .A2(S1END[0]),
    .A3(S4END[0]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_141_));
 sg13g2_nand3_1 _367_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit19.Q ),
    .C(_090_),
    .A(_008_),
    .Y(_142_));
 sg13g2_or2_1 _368_ (.X(_143_),
    .B(W6END[0]),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit18.Q ));
 sg13g2_o21ai_1 _369_ (.B1(_143_),
    .Y(_144_),
    .A1(_008_),
    .A2(_141_));
 sg13g2_o21ai_1 _370_ (.B1(_142_),
    .Y(_145_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit19.Q ),
    .A2(_144_));
 sg13g2_mux4_1 _371_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit18.Q ),
    .A0(W2MID[0]),
    .A1(W2END[0]),
    .A2(WW4END[0]),
    .A3(WW4END[8]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit19.Q ),
    .X(_146_));
 sg13g2_mux2_1 _372_ (.A0(_146_),
    .A1(_145_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit20.Q ),
    .X(UI_IN_TT_PROJECT0));
 sg13g2_o21ai_1 _373_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit15.Q ),
    .Y(_147_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit17.Q ),
    .A2(_123_));
 sg13g2_a21o_1 _374_ (.A2(_040_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit17.Q ),
    .B1(_147_),
    .X(_148_));
 sg13g2_mux2_1 _375_ (.A0(W6END[7]),
    .A1(_041_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit17.Q ),
    .X(_149_));
 sg13g2_a21oi_1 _376_ (.A1(_009_),
    .A2(_149_),
    .Y(_150_),
    .B1(_010_));
 sg13g2_mux4_1 _377_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit15.Q ),
    .A0(W1END[3]),
    .A1(WW4END[15]),
    .A2(_099_),
    .A3(_069_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit17.Q ),
    .X(_151_));
 sg13g2_nor2_1 _378_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit16.Q ),
    .B(_151_),
    .Y(_152_));
 sg13g2_a21oi_1 _379_ (.A1(_148_),
    .A2(_150_),
    .Y(\Inst_W_TT_IF_switch_matrix.S4BEG3 ),
    .B1(_152_));
 sg13g2_mux4_1 _380_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit12.Q ),
    .A0(W1END[2]),
    .A1(WW4END[14]),
    .A2(W6END[6]),
    .A3(_129_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit13.Q ),
    .X(_153_));
 sg13g2_mux4_1 _381_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit12.Q ),
    .A0(_105_),
    .A1(_076_),
    .A2(_048_),
    .A3(_047_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit13.Q ),
    .X(_154_));
 sg13g2_mux2_1 _382_ (.A0(_153_),
    .A1(_154_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit14.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.S4BEG2 ));
 sg13g2_mux4_1 _383_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit9.Q ),
    .A0(W1END[1]),
    .A1(WW4END[13]),
    .A2(W6END[5]),
    .A3(_135_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit10.Q ),
    .X(_155_));
 sg13g2_nand2b_1 _384_ (.Y(_156_),
    .B(_155_),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit11.Q ));
 sg13g2_mux2_1 _385_ (.A0(_111_),
    .A1(_083_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit9.Q ),
    .X(_157_));
 sg13g2_nand2b_1 _386_ (.Y(_158_),
    .B(_054_),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit9.Q ));
 sg13g2_nand2_1 _387_ (.Y(_159_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit9.Q ),
    .B(_055_));
 sg13g2_and3_1 _388_ (.X(_160_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit10.Q ),
    .B(_158_),
    .C(_159_));
 sg13g2_o21ai_1 _389_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit11.Q ),
    .Y(_161_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit10.Q ),
    .A2(_157_));
 sg13g2_o21ai_1 _390_ (.B1(_156_),
    .Y(\Inst_W_TT_IF_switch_matrix.S4BEG1 ),
    .A1(_160_),
    .A2(_161_));
 sg13g2_o21ai_1 _391_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit6.Q ),
    .Y(_162_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit8.Q ),
    .A2(_141_));
 sg13g2_a21o_1 _392_ (.A2(_063_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit8.Q ),
    .B1(_162_),
    .X(_163_));
 sg13g2_mux2_1 _393_ (.A0(W6END[4]),
    .A1(_061_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit8.Q ),
    .X(_164_));
 sg13g2_a21oi_1 _394_ (.A1(_011_),
    .A2(_164_),
    .Y(_165_),
    .B1(_012_));
 sg13g2_o21ai_1 _395_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit6.Q ),
    .Y(_166_),
    .A1(WW4END[12]),
    .A2(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit8.Q ));
 sg13g2_a21o_1 _396_ (.A2(_093_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit8.Q ),
    .B1(_166_),
    .X(_167_));
 sg13g2_mux2_1 _397_ (.A0(W1END[0]),
    .A1(_117_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit8.Q ),
    .X(_168_));
 sg13g2_a21oi_1 _398_ (.A1(_011_),
    .A2(_168_),
    .Y(_169_),
    .B1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit7.Q ));
 sg13g2_a22oi_1 _399_ (.Y(\Inst_W_TT_IF_switch_matrix.S4BEG0 ),
    .B1(_167_),
    .B2(_169_),
    .A2(_165_),
    .A1(_163_));
 sg13g2_mux4_1 _400_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit11.Q ),
    .A0(W1END[3]),
    .A1(WW4END[3]),
    .A2(W6END[11]),
    .A3(_123_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit12.Q ),
    .X(_170_));
 sg13g2_nand2b_1 _401_ (.Y(_171_),
    .B(_099_),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit11.Q ));
 sg13g2_a21oi_1 _402_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit11.Q ),
    .A2(_069_),
    .Y(_172_),
    .B1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit12.Q ));
 sg13g2_nand2b_1 _403_ (.Y(_173_),
    .B(_041_),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit11.Q ));
 sg13g2_a21oi_1 _404_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit11.Q ),
    .A2(_070_),
    .Y(_174_),
    .B1(_013_));
 sg13g2_a221oi_1 _405_ (.B2(_174_),
    .C1(_014_),
    .B1(_173_),
    .A1(_171_),
    .Y(_175_),
    .A2(_172_));
 sg13g2_a21o_1 _406_ (.A2(_170_),
    .A1(_014_),
    .B1(_175_),
    .X(\Inst_W_TT_IF_switch_matrix.N4BEG3 ));
 sg13g2_mux4_1 _407_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit8.Q ),
    .A0(W1END[2]),
    .A1(WW4END[2]),
    .A2(W6END[10]),
    .A3(_129_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit9.Q ),
    .X(_176_));
 sg13g2_mux4_1 _408_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit8.Q ),
    .A0(_105_),
    .A1(_076_),
    .A2(_048_),
    .A3(_077_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit9.Q ),
    .X(_177_));
 sg13g2_mux2_1 _409_ (.A0(_176_),
    .A1(_177_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit10.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.N4BEG2 ));
 sg13g2_nor2_1 _410_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit7.Q ),
    .B(_135_),
    .Y(_178_));
 sg13g2_o21ai_1 _411_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit5.Q ),
    .Y(_179_),
    .A1(_017_),
    .A2(_084_));
 sg13g2_or2_1 _412_ (.X(_180_),
    .B(_179_),
    .A(_178_));
 sg13g2_mux2_1 _413_ (.A0(W6END[9]),
    .A1(_054_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit7.Q ),
    .X(_181_));
 sg13g2_a21oi_1 _414_ (.A1(_015_),
    .A2(_181_),
    .Y(_182_),
    .B1(_016_));
 sg13g2_a21oi_1 _415_ (.A1(_006_),
    .A2(_017_),
    .Y(_183_),
    .B1(_015_));
 sg13g2_o21ai_1 _416_ (.B1(_183_),
    .Y(_184_),
    .A1(_017_),
    .A2(_083_));
 sg13g2_mux2_1 _417_ (.A0(W1END[1]),
    .A1(_111_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit7.Q ),
    .X(_185_));
 sg13g2_a21oi_1 _418_ (.A1(_015_),
    .A2(_185_),
    .Y(_186_),
    .B1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit6.Q ));
 sg13g2_a22oi_1 _419_ (.Y(\Inst_W_TT_IF_switch_matrix.N4BEG1 ),
    .B1(_184_),
    .B2(_186_),
    .A2(_182_),
    .A1(_180_));
 sg13g2_o21ai_1 _420_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit2.Q ),
    .Y(_187_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit4.Q ),
    .A2(_141_));
 sg13g2_a21o_1 _421_ (.A2(_091_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit4.Q ),
    .B1(_187_),
    .X(_188_));
 sg13g2_mux2_1 _422_ (.A0(W6END[8]),
    .A1(_061_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit4.Q ),
    .X(_189_));
 sg13g2_a21oi_1 _423_ (.A1(_018_),
    .A2(_189_),
    .Y(_190_),
    .B1(_019_));
 sg13g2_mux2_1 _424_ (.A0(W1END[0]),
    .A1(_117_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit4.Q ),
    .X(_191_));
 sg13g2_o21ai_1 _425_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit2.Q ),
    .Y(_192_),
    .A1(WW4END[0]),
    .A2(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit4.Q ));
 sg13g2_a21o_1 _426_ (.A2(_093_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit4.Q ),
    .B1(_192_),
    .X(_193_));
 sg13g2_a21oi_1 _427_ (.A1(_018_),
    .A2(_191_),
    .Y(_194_),
    .B1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit3.Q ));
 sg13g2_a22oi_1 _428_ (.Y(\Inst_W_TT_IF_switch_matrix.N4BEG0 ),
    .B1(_193_),
    .B2(_194_),
    .A2(_190_),
    .A1(_188_));
 sg13g2_o21ai_1 _429_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit2.Q ),
    .Y(_195_),
    .A1(W2MID[6]),
    .A2(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit3.Q ));
 sg13g2_nand2b_1 _430_ (.Y(_196_),
    .B(N2MID[6]),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit2.Q ));
 sg13g2_o21ai_1 _431_ (.B1(_195_),
    .Y(ENA_TT_PROJECT),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit3.Q ),
    .A2(_196_));
 sg13g2_mux4_1 _432_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit17.Q ),
    .A0(UIO_OUT_TT_PROJECT3),
    .A1(_117_),
    .A2(_141_),
    .A3(_039_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit16.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E6BEG11 ));
 sg13g2_mux4_1 _433_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit15.Q ),
    .A0(UIO_OUT_TT_PROJECT2),
    .A1(_111_),
    .A2(_135_),
    .A3(_047_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit14.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E6BEG10 ));
 sg13g2_mux4_1 _434_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit13.Q ),
    .A0(UIO_OUT_TT_PROJECT1),
    .A1(_105_),
    .A2(_129_),
    .A3(_055_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit12.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E6BEG9 ));
 sg13g2_mux4_1 _435_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit11.Q ),
    .A0(UIO_OUT_TT_PROJECT0),
    .A1(_099_),
    .A2(_123_),
    .A3(_062_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit10.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E6BEG8 ));
 sg13g2_mux4_1 _436_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit9.Q ),
    .A0(UIO_OUT_TT_PROJECT7),
    .A1(_092_),
    .A2(_117_),
    .A3(_070_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit8.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E6BEG7 ));
 sg13g2_mux4_1 _437_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit7.Q ),
    .A0(UIO_OUT_TT_PROJECT6),
    .A1(_083_),
    .A2(_111_),
    .A3(_077_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit6.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E6BEG6 ));
 sg13g2_mux4_1 _438_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit5.Q ),
    .A0(UIO_OUT_TT_PROJECT5),
    .A1(_076_),
    .A2(_105_),
    .A3(_084_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit4.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E6BEG5 ));
 sg13g2_mux4_1 _439_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit3.Q ),
    .A0(UIO_OUT_TT_PROJECT4),
    .A1(_069_),
    .A2(_099_),
    .A3(_090_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit2.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E6BEG4 ));
 sg13g2_mux4_1 _440_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit0.Q ),
    .A0(N4END[3]),
    .A1(S4END[3]),
    .A2(_092_),
    .A3(_061_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit1.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E6BEG3 ));
 sg13g2_mux4_1 _441_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit30.Q ),
    .A0(N4END[2]),
    .A1(S4END[2]),
    .A2(_083_),
    .A3(_054_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit31.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E6BEG2 ));
 sg13g2_mux4_1 _442_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit28.Q ),
    .A0(N4END[1]),
    .A1(S4END[1]),
    .A2(_076_),
    .A3(_048_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit29.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E6BEG1 ));
 sg13g2_mux4_1 _443_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit26.Q ),
    .A0(N4END[0]),
    .A1(S4END[0]),
    .A2(_069_),
    .A3(_041_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit27.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E6BEG0 ));
 sg13g2_mux4_1 _444_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit25.Q ),
    .A0(UO_OUT_TT_PROJECT3),
    .A1(_141_),
    .A2(UIO_OUT_TT_PROJECT7),
    .A3(_090_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit24.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG15 ));
 sg13g2_mux4_1 _445_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit23.Q ),
    .A0(UO_OUT_TT_PROJECT2),
    .A1(_135_),
    .A2(UIO_OUT_TT_PROJECT6),
    .A3(_084_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit22.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG14 ));
 sg13g2_mux4_1 _446_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit21.Q ),
    .A0(UO_OUT_TT_PROJECT1),
    .A1(_129_),
    .A2(UIO_OUT_TT_PROJECT5),
    .A3(_077_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit20.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG13 ));
 sg13g2_mux4_1 _447_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit19.Q ),
    .A0(UO_OUT_TT_PROJECT0),
    .A1(_123_),
    .A2(UIO_OUT_TT_PROJECT4),
    .A3(_070_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit18.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG12 ));
 sg13g2_mux4_1 _448_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit17.Q ),
    .A0(UO_OUT_TT_PROJECT7),
    .A1(_117_),
    .A2(UIO_OUT_TT_PROJECT3),
    .A3(_062_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit16.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG11 ));
 sg13g2_mux4_1 _449_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit15.Q ),
    .A0(UO_OUT_TT_PROJECT6),
    .A1(_111_),
    .A2(UIO_OUT_TT_PROJECT2),
    .A3(_055_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit14.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG10 ));
 sg13g2_mux4_1 _450_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit13.Q ),
    .A0(UO_OUT_TT_PROJECT5),
    .A1(_105_),
    .A2(UIO_OUT_TT_PROJECT1),
    .A3(_047_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit12.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG9 ));
 sg13g2_mux4_1 _451_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit11.Q ),
    .A0(UO_OUT_TT_PROJECT4),
    .A1(_099_),
    .A2(UIO_OUT_TT_PROJECT0),
    .A3(_039_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit10.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG8 ));
 sg13g2_mux4_1 _452_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit8.Q ),
    .A0(UO_OUT_TT_PROJECT7),
    .A1(UIO_OE_TT_PROJECT3),
    .A2(_092_),
    .A3(_090_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit9.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG7 ));
 sg13g2_mux4_1 _453_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit6.Q ),
    .A0(UO_OUT_TT_PROJECT6),
    .A1(UIO_OE_TT_PROJECT2),
    .A2(_083_),
    .A3(_084_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit7.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG6 ));
 sg13g2_mux4_1 _454_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit4.Q ),
    .A0(UO_OUT_TT_PROJECT5),
    .A1(UIO_OE_TT_PROJECT1),
    .A2(_076_),
    .A3(_077_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit5.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG5 ));
 sg13g2_mux4_1 _455_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit2.Q ),
    .A0(UO_OUT_TT_PROJECT4),
    .A1(UIO_OE_TT_PROJECT0),
    .A2(_069_),
    .A3(_070_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit3.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG4 ));
 sg13g2_mux4_1 _456_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit0.Q ),
    .A0(UO_OUT_TT_PROJECT3),
    .A1(UIO_OE_TT_PROJECT7),
    .A2(_061_),
    .A3(_062_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit1.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG3 ));
 sg13g2_mux4_1 _457_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit30.Q ),
    .A0(UO_OUT_TT_PROJECT2),
    .A1(UIO_OE_TT_PROJECT6),
    .A2(_054_),
    .A3(_055_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit31.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG2 ));
 sg13g2_mux4_1 _458_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit28.Q ),
    .A0(UO_OUT_TT_PROJECT1),
    .A1(UIO_OE_TT_PROJECT5),
    .A2(_048_),
    .A3(_047_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit29.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG1 ));
 sg13g2_mux4_1 _459_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit26.Q ),
    .A0(UO_OUT_TT_PROJECT0),
    .A1(UIO_OE_TT_PROJECT4),
    .A2(_041_),
    .A3(_039_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit27.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG0 ));
 sg13g2_mux4_1 _460_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit24.Q ),
    .A0(UIO_OUT_TT_PROJECT7),
    .A1(UIO_OE_TT_PROJECT7),
    .A2(_090_),
    .A3(_039_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit25.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E2BEGb7 ));
 sg13g2_mux4_1 _461_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit22.Q ),
    .A0(UIO_OUT_TT_PROJECT6),
    .A1(UIO_OE_TT_PROJECT6),
    .A2(_084_),
    .A3(_047_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit23.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E2BEGb6 ));
 sg13g2_mux4_1 _462_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit20.Q ),
    .A0(UIO_OUT_TT_PROJECT5),
    .A1(UIO_OE_TT_PROJECT5),
    .A2(_077_),
    .A3(_055_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit21.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E2BEGb5 ));
 sg13g2_mux4_1 _463_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit18.Q ),
    .A0(UIO_OUT_TT_PROJECT4),
    .A1(UIO_OE_TT_PROJECT4),
    .A2(_070_),
    .A3(_062_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit19.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E2BEGb4 ));
 sg13g2_mux4_1 _464_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit16.Q ),
    .A0(UIO_OUT_TT_PROJECT3),
    .A1(UIO_OE_TT_PROJECT3),
    .A2(_070_),
    .A3(_062_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit17.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E2BEGb3 ));
 sg13g2_mux4_1 _465_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit14.Q ),
    .A0(UIO_OUT_TT_PROJECT2),
    .A1(UIO_OE_TT_PROJECT2),
    .A2(_077_),
    .A3(_055_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit15.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E2BEGb2 ));
 sg13g2_mux4_1 _466_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit12.Q ),
    .A0(UIO_OUT_TT_PROJECT1),
    .A1(UIO_OE_TT_PROJECT1),
    .A2(_084_),
    .A3(_047_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit13.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E2BEGb1 ));
 sg13g2_mux4_1 _467_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit10.Q ),
    .A0(UIO_OUT_TT_PROJECT0),
    .A1(UIO_OE_TT_PROJECT0),
    .A2(_090_),
    .A3(_039_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit11.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E2BEGb0 ));
 sg13g2_mux4_1 _468_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit9.Q ),
    .A0(UO_OUT_TT_PROJECT7),
    .A1(_090_),
    .A2(UIO_OUT_TT_PROJECT7),
    .A3(_039_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit8.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E2BEG7 ));
 sg13g2_mux4_1 _469_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit7.Q ),
    .A0(UO_OUT_TT_PROJECT6),
    .A1(_084_),
    .A2(UIO_OUT_TT_PROJECT6),
    .A3(_047_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit6.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E2BEG6 ));
 sg13g2_mux4_1 _470_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit5.Q ),
    .A0(UO_OUT_TT_PROJECT5),
    .A1(_077_),
    .A2(UIO_OUT_TT_PROJECT5),
    .A3(_055_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit4.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E2BEG5 ));
 sg13g2_mux4_1 _471_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit3.Q ),
    .A0(UO_OUT_TT_PROJECT4),
    .A1(_070_),
    .A2(UIO_OUT_TT_PROJECT4),
    .A3(_062_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit2.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E2BEG4 ));
 sg13g2_mux4_1 _472_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit1.Q ),
    .A0(UO_OUT_TT_PROJECT3),
    .A1(_070_),
    .A2(UIO_OUT_TT_PROJECT3),
    .A3(_062_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit0.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E2BEG3 ));
 sg13g2_mux4_1 _473_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit31.Q ),
    .A0(UO_OUT_TT_PROJECT2),
    .A1(_077_),
    .A2(UIO_OUT_TT_PROJECT2),
    .A3(_055_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit30.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E2BEG2 ));
 sg13g2_mux4_1 _474_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit29.Q ),
    .A0(UO_OUT_TT_PROJECT1),
    .A1(_084_),
    .A2(UIO_OUT_TT_PROJECT1),
    .A3(_047_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit28.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E2BEG1 ));
 sg13g2_mux4_1 _475_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit27.Q ),
    .A0(UO_OUT_TT_PROJECT0),
    .A1(_090_),
    .A2(UIO_OUT_TT_PROJECT0),
    .A3(_039_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit26.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E2BEG0 ));
 sg13g2_mux4_1 _476_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit24.Q ),
    .A0(N1END[3]),
    .A1(S1END[3]),
    .A2(UO_OUT_TT_PROJECT1),
    .A3(UO_OUT_TT_PROJECT4),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit25.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E1BEG3 ));
 sg13g2_mux4_1 _477_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit22.Q ),
    .A0(N1END[2]),
    .A1(S1END[2]),
    .A2(UO_OUT_TT_PROJECT0),
    .A3(UO_OUT_TT_PROJECT5),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit23.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E1BEG2 ));
 sg13g2_mux4_1 _478_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit20.Q ),
    .A0(N1END[1]),
    .A1(S1END[1]),
    .A2(UO_OUT_TT_PROJECT3),
    .A3(UO_OUT_TT_PROJECT6),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit21.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E1BEG1 ));
 sg13g2_mux4_1 _479_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit18.Q ),
    .A0(N1END[0]),
    .A1(S1END[0]),
    .A2(UO_OUT_TT_PROJECT2),
    .A3(UO_OUT_TT_PROJECT7),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit19.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E1BEG0 ));
 sg13g2_mux4_1 _480_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit5.Q ),
    .A0(W1END[3]),
    .A1(W2END[0]),
    .A2(W2MID[0]),
    .A3(_039_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit4.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.S2BEG7 ));
 sg13g2_mux4_1 _481_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit2.Q ),
    .A0(W1END[2]),
    .A1(W2MID[1]),
    .A2(W2END[1]),
    .A3(_047_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit3.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.S2BEG6 ));
 sg13g2_mux4_1 _482_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit0.Q ),
    .A0(W1END[1]),
    .A1(W2MID[2]),
    .A2(W2END[2]),
    .A3(_055_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit1.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.S2BEG5 ));
 sg13g2_mux4_1 _483_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit31.Q ),
    .A0(W1END[0]),
    .A1(W2END[3]),
    .A2(W2MID[3]),
    .A3(_062_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit30.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.S2BEG4 ));
 sg13g2_mux4_1 _484_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit29.Q ),
    .A0(W2MID[4]),
    .A1(W6END[11]),
    .A2(W2END[4]),
    .A3(_070_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit28.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.S2BEG3 ));
 sg13g2_mux4_1 _485_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit27.Q ),
    .A0(W2MID[5]),
    .A1(W6END[10]),
    .A2(W2END[5]),
    .A3(_077_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit26.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.S2BEG2 ));
 sg13g2_mux4_1 _486_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit24.Q ),
    .A0(W2MID[6]),
    .A1(W2END[6]),
    .A2(W6END[9]),
    .A3(_084_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit25.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.S2BEG1 ));
 sg13g2_mux4_1 _487_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit22.Q ),
    .A0(W2MID[7]),
    .A1(W2END[7]),
    .A2(W6END[8]),
    .A3(_090_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit23.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.S2BEG0 ));
 sg13g2_nor3_1 _488_ (.A(N1END[3]),
    .B(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit30.Q ),
    .C(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit31.Q ),
    .Y(_197_));
 sg13g2_nand2b_1 _489_ (.Y(_198_),
    .B(W6END[3]),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit31.Q ));
 sg13g2_a221oi_1 _490_ (.B2(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit30.Q ),
    .C1(_197_),
    .B1(_198_),
    .A1(_002_),
    .Y(_199_),
    .A2(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit31.Q ));
 sg13g2_mux4_1 _491_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit20.Q ),
    .A0(W1END[3]),
    .A1(W6END[11]),
    .A2(_041_),
    .A3(_199_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit21.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.S1BEG3 ));
 sg13g2_nor3_1 _492_ (.A(N1END[2]),
    .B(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit28.Q ),
    .C(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit29.Q ),
    .Y(_200_));
 sg13g2_nand2b_1 _493_ (.Y(_201_),
    .B(W6END[2]),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit29.Q ));
 sg13g2_a221oi_1 _494_ (.B2(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit28.Q ),
    .C1(_200_),
    .B1(_201_),
    .A1(_003_),
    .Y(_202_),
    .A2(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit29.Q ));
 sg13g2_mux4_1 _495_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit18.Q ),
    .A0(W1END[2]),
    .A1(W6END[10]),
    .A2(_048_),
    .A3(_202_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit19.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.S1BEG2 ));
 sg13g2_nor3_1 _496_ (.A(N1END[1]),
    .B(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit26.Q ),
    .C(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit27.Q ),
    .Y(_203_));
 sg13g2_nand2b_1 _497_ (.Y(_204_),
    .B(W6END[1]),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit27.Q ));
 sg13g2_a221oi_1 _498_ (.B2(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit26.Q ),
    .C1(_203_),
    .B1(_204_),
    .A1(_004_),
    .Y(_205_),
    .A2(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit27.Q ));
 sg13g2_mux4_1 _499_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit16.Q ),
    .A0(W1END[1]),
    .A1(W6END[9]),
    .A2(_054_),
    .A3(_205_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit17.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.S1BEG1 ));
 sg13g2_nor3_1 _500_ (.A(N1END[0]),
    .B(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit24.Q ),
    .C(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit25.Q ),
    .Y(_206_));
 sg13g2_nand2b_1 _501_ (.Y(_207_),
    .B(W6END[0]),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit25.Q ));
 sg13g2_a221oi_1 _502_ (.B2(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit24.Q ),
    .C1(_206_),
    .B1(_207_),
    .A1(_005_),
    .Y(_208_),
    .A2(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit25.Q ));
 sg13g2_mux4_1 _503_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit14.Q ),
    .A0(W1END[0]),
    .A1(W6END[8]),
    .A2(_061_),
    .A3(_208_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit15.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.S1BEG0 ));
 sg13g2_mux4_1 _504_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit0.Q ),
    .A0(W2MID[0]),
    .A1(W2END[0]),
    .A2(W6END[0]),
    .A3(_039_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit1.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.N2BEG7 ));
 sg13g2_mux4_1 _505_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit31.Q ),
    .A0(W2MID[1]),
    .A1(W6END[1]),
    .A2(W2END[1]),
    .A3(_047_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit30.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.N2BEG6 ));
 sg13g2_mux4_1 _506_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit29.Q ),
    .A0(W2MID[2]),
    .A1(W6END[2]),
    .A2(W2END[2]),
    .A3(_055_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit28.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.N2BEG5 ));
 sg13g2_mux4_1 _507_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit26.Q ),
    .A0(W2MID[3]),
    .A1(W2END[3]),
    .A2(W6END[3]),
    .A3(_062_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit27.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.N2BEG4 ));
 sg13g2_mux4_1 _508_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit25.Q ),
    .A0(W2MID[4]),
    .A1(W6END[4]),
    .A2(W2END[4]),
    .A3(_070_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit24.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.N2BEG3 ));
 sg13g2_mux4_1 _509_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit23.Q ),
    .A0(W2MID[5]),
    .A1(W6END[5]),
    .A2(W2END[5]),
    .A3(_077_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit22.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.N2BEG2 ));
 sg13g2_mux4_1 _510_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit20.Q ),
    .A0(W2MID[6]),
    .A1(W2END[6]),
    .A2(W6END[6]),
    .A3(_084_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit21.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.N2BEG1 ));
 sg13g2_mux4_1 _511_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit18.Q ),
    .A0(W2MID[7]),
    .A1(W2END[7]),
    .A2(W6END[7]),
    .A3(_090_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit19.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.N2BEG0 ));
 sg13g2_mux4_1 _512_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit16.Q ),
    .A0(W1END[3]),
    .A1(W6END[7]),
    .A2(_041_),
    .A3(_199_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit17.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.N1BEG3 ));
 sg13g2_mux4_1 _513_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit14.Q ),
    .A0(W1END[2]),
    .A1(W6END[6]),
    .A2(_048_),
    .A3(_202_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit15.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.N1BEG2 ));
 sg13g2_mux4_1 _514_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit12.Q ),
    .A0(W1END[1]),
    .A1(W6END[5]),
    .A2(_054_),
    .A3(_205_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit13.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.N1BEG1 ));
 sg13g2_mux4_1 _515_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit10.Q ),
    .A0(W1END[0]),
    .A1(W6END[4]),
    .A2(_061_),
    .A3(_208_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit11.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.N1BEG0 ));
 sg13g2_dlhq_1 _516_ (.D(FrameData[10]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit10.Q ));
 sg13g2_dlhq_1 _517_ (.D(FrameData[11]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit11.Q ));
 sg13g2_dlhq_1 _518_ (.D(FrameData[12]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit12.Q ));
 sg13g2_dlhq_1 _519_ (.D(FrameData[13]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit13.Q ));
 sg13g2_dlhq_1 _520_ (.D(FrameData[14]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit14.Q ));
 sg13g2_dlhq_1 _521_ (.D(FrameData[15]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit15.Q ));
 sg13g2_dlhq_1 _522_ (.D(FrameData[16]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit16.Q ));
 sg13g2_dlhq_1 _523_ (.D(FrameData[17]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit17.Q ));
 sg13g2_dlhq_1 _524_ (.D(FrameData[18]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit18.Q ));
 sg13g2_dlhq_1 _525_ (.D(FrameData[19]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit19.Q ));
 sg13g2_dlhq_1 _526_ (.D(FrameData[20]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit20.Q ));
 sg13g2_dlhq_1 _527_ (.D(FrameData[21]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit21.Q ));
 sg13g2_dlhq_1 _528_ (.D(FrameData[22]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit22.Q ));
 sg13g2_dlhq_1 _529_ (.D(FrameData[23]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit23.Q ));
 sg13g2_dlhq_1 _530_ (.D(FrameData[24]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit24.Q ));
 sg13g2_dlhq_1 _531_ (.D(FrameData[25]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit25.Q ));
 sg13g2_dlhq_1 _532_ (.D(FrameData[26]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit26.Q ));
 sg13g2_dlhq_1 _533_ (.D(FrameData[27]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit27.Q ));
 sg13g2_dlhq_1 _534_ (.D(FrameData[28]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit28.Q ));
 sg13g2_dlhq_1 _535_ (.D(FrameData[29]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit29.Q ));
 sg13g2_dlhq_1 _536_ (.D(FrameData[30]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit30.Q ));
 sg13g2_dlhq_1 _537_ (.D(FrameData[31]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit31.Q ));
 sg13g2_dlhq_1 _538_ (.D(FrameData[0]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit0.Q ));
 sg13g2_dlhq_1 _539_ (.D(FrameData[1]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit1.Q ));
 sg13g2_dlhq_1 _540_ (.D(FrameData[2]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit2.Q ));
 sg13g2_dlhq_1 _541_ (.D(FrameData[3]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit3.Q ));
 sg13g2_dlhq_1 _542_ (.D(FrameData[4]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit4.Q ));
 sg13g2_dlhq_1 _543_ (.D(FrameData[5]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit5.Q ));
 sg13g2_dlhq_1 _544_ (.D(FrameData[6]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit6.Q ));
 sg13g2_dlhq_1 _545_ (.D(FrameData[7]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit7.Q ));
 sg13g2_dlhq_1 _546_ (.D(FrameData[8]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit8.Q ));
 sg13g2_dlhq_1 _547_ (.D(FrameData[9]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit9.Q ));
 sg13g2_dlhq_1 _548_ (.D(FrameData[10]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit10.Q ));
 sg13g2_dlhq_1 _549_ (.D(FrameData[11]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit11.Q ));
 sg13g2_dlhq_1 _550_ (.D(FrameData[12]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit12.Q ));
 sg13g2_dlhq_1 _551_ (.D(FrameData[13]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit13.Q ));
 sg13g2_dlhq_1 _552_ (.D(FrameData[14]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit14.Q ));
 sg13g2_dlhq_1 _553_ (.D(FrameData[15]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit15.Q ));
 sg13g2_dlhq_1 _554_ (.D(FrameData[16]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit16.Q ));
 sg13g2_dlhq_1 _555_ (.D(FrameData[17]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit17.Q ));
 sg13g2_dlhq_1 _556_ (.D(FrameData[18]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit18.Q ));
 sg13g2_dlhq_1 _557_ (.D(FrameData[19]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit19.Q ));
 sg13g2_dlhq_1 _558_ (.D(FrameData[20]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit20.Q ));
 sg13g2_dlhq_1 _559_ (.D(FrameData[21]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit21.Q ));
 sg13g2_dlhq_1 _560_ (.D(FrameData[22]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit22.Q ));
 sg13g2_dlhq_1 _561_ (.D(FrameData[23]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit23.Q ));
 sg13g2_dlhq_1 _562_ (.D(FrameData[24]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit24.Q ));
 sg13g2_dlhq_1 _563_ (.D(FrameData[25]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit25.Q ));
 sg13g2_dlhq_1 _564_ (.D(FrameData[26]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit26.Q ));
 sg13g2_dlhq_1 _565_ (.D(FrameData[27]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit27.Q ));
 sg13g2_dlhq_1 _566_ (.D(FrameData[28]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit28.Q ));
 sg13g2_dlhq_1 _567_ (.D(FrameData[29]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit29.Q ));
 sg13g2_dlhq_1 _568_ (.D(FrameData[30]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit30.Q ));
 sg13g2_dlhq_1 _569_ (.D(FrameData[31]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit31.Q ));
 sg13g2_dlhq_1 _570_ (.D(FrameData[0]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit0.Q ));
 sg13g2_dlhq_1 _571_ (.D(FrameData[1]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit1.Q ));
 sg13g2_dlhq_1 _572_ (.D(FrameData[2]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit2.Q ));
 sg13g2_dlhq_1 _573_ (.D(FrameData[3]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit3.Q ));
 sg13g2_dlhq_1 _574_ (.D(FrameData[4]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit4.Q ));
 sg13g2_dlhq_1 _575_ (.D(FrameData[5]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit5.Q ));
 sg13g2_dlhq_1 _576_ (.D(FrameData[6]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit6.Q ));
 sg13g2_dlhq_1 _577_ (.D(FrameData[7]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit7.Q ));
 sg13g2_dlhq_1 _578_ (.D(FrameData[8]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit8.Q ));
 sg13g2_dlhq_1 _579_ (.D(FrameData[9]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit9.Q ));
 sg13g2_dlhq_1 _580_ (.D(FrameData[10]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit10.Q ));
 sg13g2_dlhq_1 _581_ (.D(FrameData[11]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit11.Q ));
 sg13g2_dlhq_1 _582_ (.D(FrameData[12]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit12.Q ));
 sg13g2_dlhq_1 _583_ (.D(FrameData[13]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit13.Q ));
 sg13g2_dlhq_1 _584_ (.D(FrameData[14]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit14.Q ));
 sg13g2_dlhq_1 _585_ (.D(FrameData[15]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit15.Q ));
 sg13g2_dlhq_1 _586_ (.D(FrameData[16]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit16.Q ));
 sg13g2_dlhq_1 _587_ (.D(FrameData[17]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit17.Q ));
 sg13g2_dlhq_1 _588_ (.D(FrameData[18]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit18.Q ));
 sg13g2_dlhq_1 _589_ (.D(FrameData[19]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit19.Q ));
 sg13g2_dlhq_1 _590_ (.D(FrameData[20]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit20.Q ));
 sg13g2_dlhq_1 _591_ (.D(FrameData[21]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit21.Q ));
 sg13g2_dlhq_1 _592_ (.D(FrameData[22]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit22.Q ));
 sg13g2_dlhq_1 _593_ (.D(FrameData[23]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit23.Q ));
 sg13g2_dlhq_1 _594_ (.D(FrameData[24]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit24.Q ));
 sg13g2_dlhq_1 _595_ (.D(FrameData[25]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit25.Q ));
 sg13g2_dlhq_1 _596_ (.D(FrameData[26]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit26.Q ));
 sg13g2_dlhq_1 _597_ (.D(FrameData[27]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit27.Q ));
 sg13g2_dlhq_1 _598_ (.D(FrameData[28]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit28.Q ));
 sg13g2_dlhq_1 _599_ (.D(FrameData[29]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit29.Q ));
 sg13g2_dlhq_1 _600_ (.D(FrameData[30]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit30.Q ));
 sg13g2_dlhq_1 _601_ (.D(FrameData[31]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit31.Q ));
 sg13g2_dlhq_1 _602_ (.D(FrameData[0]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit0.Q ));
 sg13g2_dlhq_1 _603_ (.D(FrameData[1]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit1.Q ));
 sg13g2_dlhq_1 _604_ (.D(FrameData[2]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit2.Q ));
 sg13g2_dlhq_1 _605_ (.D(FrameData[3]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit3.Q ));
 sg13g2_dlhq_1 _606_ (.D(FrameData[4]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit4.Q ));
 sg13g2_dlhq_1 _607_ (.D(FrameData[5]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit5.Q ));
 sg13g2_dlhq_1 _608_ (.D(FrameData[6]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit6.Q ));
 sg13g2_dlhq_1 _609_ (.D(FrameData[7]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit7.Q ));
 sg13g2_dlhq_1 _610_ (.D(FrameData[8]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit8.Q ));
 sg13g2_dlhq_1 _611_ (.D(FrameData[9]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit9.Q ));
 sg13g2_dlhq_1 _612_ (.D(FrameData[10]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit10.Q ));
 sg13g2_dlhq_1 _613_ (.D(FrameData[11]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit11.Q ));
 sg13g2_dlhq_1 _614_ (.D(FrameData[12]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit12.Q ));
 sg13g2_dlhq_1 _615_ (.D(FrameData[13]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit13.Q ));
 sg13g2_dlhq_1 _616_ (.D(FrameData[14]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit14.Q ));
 sg13g2_dlhq_1 _617_ (.D(FrameData[15]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit15.Q ));
 sg13g2_dlhq_1 _618_ (.D(FrameData[16]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit16.Q ));
 sg13g2_dlhq_1 _619_ (.D(FrameData[17]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit17.Q ));
 sg13g2_dlhq_1 _620_ (.D(FrameData[18]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit18.Q ));
 sg13g2_dlhq_1 _621_ (.D(FrameData[19]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit19.Q ));
 sg13g2_dlhq_1 _622_ (.D(FrameData[20]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit20.Q ));
 sg13g2_dlhq_1 _623_ (.D(FrameData[21]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit21.Q ));
 sg13g2_dlhq_1 _624_ (.D(FrameData[22]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit22.Q ));
 sg13g2_dlhq_1 _625_ (.D(FrameData[23]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit23.Q ));
 sg13g2_dlhq_1 _626_ (.D(FrameData[24]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit24.Q ));
 sg13g2_dlhq_1 _627_ (.D(FrameData[25]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit25.Q ));
 sg13g2_dlhq_1 _628_ (.D(FrameData[26]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit26.Q ));
 sg13g2_dlhq_1 _629_ (.D(FrameData[27]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit27.Q ));
 sg13g2_dlhq_1 _630_ (.D(FrameData[28]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit28.Q ));
 sg13g2_dlhq_1 _631_ (.D(FrameData[29]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit29.Q ));
 sg13g2_dlhq_1 _632_ (.D(FrameData[30]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit30.Q ));
 sg13g2_dlhq_1 _633_ (.D(FrameData[31]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit31.Q ));
 sg13g2_dlhq_1 _634_ (.D(FrameData[0]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit0.Q ));
 sg13g2_dlhq_1 _635_ (.D(FrameData[1]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit1.Q ));
 sg13g2_dlhq_1 _636_ (.D(FrameData[2]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit2.Q ));
 sg13g2_dlhq_1 _637_ (.D(FrameData[3]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit3.Q ));
 sg13g2_dlhq_1 _638_ (.D(FrameData[4]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit4.Q ));
 sg13g2_dlhq_1 _639_ (.D(FrameData[5]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit5.Q ));
 sg13g2_dlhq_1 _640_ (.D(FrameData[6]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit6.Q ));
 sg13g2_dlhq_1 _641_ (.D(FrameData[7]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit7.Q ));
 sg13g2_dlhq_1 _642_ (.D(FrameData[8]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit8.Q ));
 sg13g2_dlhq_1 _643_ (.D(FrameData[9]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit9.Q ));
 sg13g2_dlhq_1 _644_ (.D(FrameData[10]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit10.Q ));
 sg13g2_dlhq_1 _645_ (.D(FrameData[11]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit11.Q ));
 sg13g2_dlhq_1 _646_ (.D(FrameData[12]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit12.Q ));
 sg13g2_dlhq_1 _647_ (.D(FrameData[13]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit13.Q ));
 sg13g2_dlhq_1 _648_ (.D(FrameData[14]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit14.Q ));
 sg13g2_dlhq_1 _649_ (.D(FrameData[15]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit15.Q ));
 sg13g2_dlhq_1 _650_ (.D(FrameData[16]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit16.Q ));
 sg13g2_dlhq_1 _651_ (.D(FrameData[17]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit17.Q ));
 sg13g2_dlhq_1 _652_ (.D(FrameData[18]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit18.Q ));
 sg13g2_dlhq_1 _653_ (.D(FrameData[19]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit19.Q ));
 sg13g2_dlhq_1 _654_ (.D(FrameData[20]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit20.Q ));
 sg13g2_dlhq_1 _655_ (.D(FrameData[21]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit21.Q ));
 sg13g2_dlhq_1 _656_ (.D(FrameData[22]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit22.Q ));
 sg13g2_dlhq_1 _657_ (.D(FrameData[23]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit23.Q ));
 sg13g2_dlhq_1 _658_ (.D(FrameData[24]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit24.Q ));
 sg13g2_dlhq_1 _659_ (.D(FrameData[25]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit25.Q ));
 sg13g2_dlhq_1 _660_ (.D(FrameData[26]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit26.Q ));
 sg13g2_dlhq_1 _661_ (.D(FrameData[27]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit27.Q ));
 sg13g2_dlhq_1 _662_ (.D(FrameData[28]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit28.Q ));
 sg13g2_dlhq_1 _663_ (.D(FrameData[29]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit29.Q ));
 sg13g2_dlhq_1 _664_ (.D(FrameData[30]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit30.Q ));
 sg13g2_dlhq_1 _665_ (.D(FrameData[31]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit31.Q ));
 sg13g2_dlhq_1 _666_ (.D(FrameData[0]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit0.Q ));
 sg13g2_dlhq_1 _667_ (.D(FrameData[1]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit1.Q ));
 sg13g2_dlhq_1 _668_ (.D(FrameData[2]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit2.Q ));
 sg13g2_dlhq_1 _669_ (.D(FrameData[3]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit3.Q ));
 sg13g2_dlhq_1 _670_ (.D(FrameData[4]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit4.Q ));
 sg13g2_dlhq_1 _671_ (.D(FrameData[5]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit5.Q ));
 sg13g2_dlhq_1 _672_ (.D(FrameData[6]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit6.Q ));
 sg13g2_dlhq_1 _673_ (.D(FrameData[7]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit7.Q ));
 sg13g2_dlhq_1 _674_ (.D(FrameData[8]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit8.Q ));
 sg13g2_dlhq_1 _675_ (.D(FrameData[9]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit9.Q ));
 sg13g2_dlhq_1 _676_ (.D(FrameData[10]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit10.Q ));
 sg13g2_dlhq_1 _677_ (.D(FrameData[11]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit11.Q ));
 sg13g2_dlhq_1 _678_ (.D(FrameData[12]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit12.Q ));
 sg13g2_dlhq_1 _679_ (.D(FrameData[13]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit13.Q ));
 sg13g2_dlhq_1 _680_ (.D(FrameData[14]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit14.Q ));
 sg13g2_dlhq_1 _681_ (.D(FrameData[15]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit15.Q ));
 sg13g2_dlhq_1 _682_ (.D(FrameData[16]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit16.Q ));
 sg13g2_dlhq_1 _683_ (.D(FrameData[17]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit17.Q ));
 sg13g2_dlhq_1 _684_ (.D(FrameData[18]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit18.Q ));
 sg13g2_dlhq_1 _685_ (.D(FrameData[19]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit19.Q ));
 sg13g2_dlhq_1 _686_ (.D(FrameData[20]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit20.Q ));
 sg13g2_dlhq_1 _687_ (.D(FrameData[21]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit21.Q ));
 sg13g2_dlhq_1 _688_ (.D(FrameData[22]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit22.Q ));
 sg13g2_dlhq_1 _689_ (.D(FrameData[23]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit23.Q ));
 sg13g2_dlhq_1 _690_ (.D(FrameData[24]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit24.Q ));
 sg13g2_dlhq_1 _691_ (.D(FrameData[25]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit25.Q ));
 sg13g2_dlhq_1 _692_ (.D(FrameData[26]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit26.Q ));
 sg13g2_dlhq_1 _693_ (.D(FrameData[27]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit27.Q ));
 sg13g2_dlhq_1 _694_ (.D(FrameData[28]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit28.Q ));
 sg13g2_dlhq_1 _695_ (.D(FrameData[29]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit29.Q ));
 sg13g2_dlhq_1 _696_ (.D(FrameData[30]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit30.Q ));
 sg13g2_dlhq_1 _697_ (.D(FrameData[31]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit31.Q ));
 sg13g2_dlhq_1 _698_ (.D(FrameData[0]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit0.Q ));
 sg13g2_dlhq_1 _699_ (.D(FrameData[1]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit1.Q ));
 sg13g2_dlhq_1 _700_ (.D(FrameData[2]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit2.Q ));
 sg13g2_dlhq_1 _701_ (.D(FrameData[3]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit3.Q ));
 sg13g2_dlhq_1 _702_ (.D(FrameData[4]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit4.Q ));
 sg13g2_dlhq_1 _703_ (.D(FrameData[5]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit5.Q ));
 sg13g2_dlhq_1 _704_ (.D(FrameData[6]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit6.Q ));
 sg13g2_dlhq_1 _705_ (.D(FrameData[7]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit7.Q ));
 sg13g2_dlhq_1 _706_ (.D(FrameData[8]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit8.Q ));
 sg13g2_dlhq_1 _707_ (.D(FrameData[9]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit9.Q ));
 sg13g2_dlhq_1 _708_ (.D(FrameData[10]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit10.Q ));
 sg13g2_dlhq_1 _709_ (.D(FrameData[11]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit11.Q ));
 sg13g2_dlhq_1 _710_ (.D(FrameData[12]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit12.Q ));
 sg13g2_dlhq_1 _711_ (.D(FrameData[13]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit13.Q ));
 sg13g2_dlhq_1 _712_ (.D(FrameData[14]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit14.Q ));
 sg13g2_dlhq_1 _713_ (.D(FrameData[15]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit15.Q ));
 sg13g2_dlhq_1 _714_ (.D(FrameData[16]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit16.Q ));
 sg13g2_dlhq_1 _715_ (.D(FrameData[17]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit17.Q ));
 sg13g2_dlhq_1 _716_ (.D(FrameData[18]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit18.Q ));
 sg13g2_dlhq_1 _717_ (.D(FrameData[19]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit19.Q ));
 sg13g2_dlhq_1 _718_ (.D(FrameData[20]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit20.Q ));
 sg13g2_dlhq_1 _719_ (.D(FrameData[21]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit21.Q ));
 sg13g2_dlhq_1 _720_ (.D(FrameData[22]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit22.Q ));
 sg13g2_dlhq_1 _721_ (.D(FrameData[23]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit23.Q ));
 sg13g2_dlhq_1 _722_ (.D(FrameData[24]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit24.Q ));
 sg13g2_dlhq_1 _723_ (.D(FrameData[25]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit25.Q ));
 sg13g2_dlhq_1 _724_ (.D(FrameData[26]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit26.Q ));
 sg13g2_dlhq_1 _725_ (.D(FrameData[27]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit27.Q ));
 sg13g2_dlhq_1 _726_ (.D(FrameData[28]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit28.Q ));
 sg13g2_dlhq_1 _727_ (.D(FrameData[29]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit29.Q ));
 sg13g2_dlhq_1 _728_ (.D(FrameData[30]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit30.Q ));
 sg13g2_dlhq_1 _729_ (.D(FrameData[31]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit31.Q ));
 sg13g2_dlhq_1 _730_ (.D(FrameData[0]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit0.Q ));
 sg13g2_dlhq_1 _731_ (.D(FrameData[1]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit1.Q ));
 sg13g2_dlhq_1 _732_ (.D(FrameData[2]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit2.Q ));
 sg13g2_dlhq_1 _733_ (.D(FrameData[3]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit3.Q ));
 sg13g2_dlhq_1 _734_ (.D(FrameData[4]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit4.Q ));
 sg13g2_dlhq_1 _735_ (.D(FrameData[5]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit5.Q ));
 sg13g2_dlhq_1 _736_ (.D(FrameData[6]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit6.Q ));
 sg13g2_dlhq_1 _737_ (.D(FrameData[7]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit7.Q ));
 sg13g2_dlhq_1 _738_ (.D(FrameData[8]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit8.Q ));
 sg13g2_dlhq_1 _739_ (.D(FrameData[9]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit9.Q ));
 sg13g2_dlhq_1 _740_ (.D(FrameData[10]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit10.Q ));
 sg13g2_dlhq_1 _741_ (.D(FrameData[11]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit11.Q ));
 sg13g2_dlhq_1 _742_ (.D(FrameData[12]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit12.Q ));
 sg13g2_dlhq_1 _743_ (.D(FrameData[13]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit13.Q ));
 sg13g2_dlhq_1 _744_ (.D(FrameData[14]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit14.Q ));
 sg13g2_dlhq_1 _745_ (.D(FrameData[15]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit15.Q ));
 sg13g2_dlhq_1 _746_ (.D(FrameData[16]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit16.Q ));
 sg13g2_dlhq_1 _747_ (.D(FrameData[17]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit17.Q ));
 sg13g2_dlhq_1 _748_ (.D(FrameData[18]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit18.Q ));
 sg13g2_dlhq_1 _749_ (.D(FrameData[19]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit19.Q ));
 sg13g2_dlhq_1 _750_ (.D(FrameData[20]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit20.Q ));
 sg13g2_dlhq_1 _751_ (.D(FrameData[21]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit21.Q ));
 sg13g2_dlhq_1 _752_ (.D(FrameData[22]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit22.Q ));
 sg13g2_dlhq_1 _753_ (.D(FrameData[23]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit23.Q ));
 sg13g2_dlhq_1 _754_ (.D(FrameData[24]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit24.Q ));
 sg13g2_dlhq_1 _755_ (.D(FrameData[25]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit25.Q ));
 sg13g2_dlhq_1 _756_ (.D(FrameData[26]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit26.Q ));
 sg13g2_dlhq_1 _757_ (.D(FrameData[27]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit27.Q ));
 sg13g2_dlhq_1 _758_ (.D(FrameData[28]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit28.Q ));
 sg13g2_dlhq_1 _759_ (.D(FrameData[29]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit29.Q ));
 sg13g2_dlhq_1 _760_ (.D(FrameData[30]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit30.Q ));
 sg13g2_dlhq_1 _761_ (.D(FrameData[31]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit31.Q ));
 sg13g2_dlhq_1 _762_ (.D(FrameData[0]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit0.Q ));
 sg13g2_dlhq_1 _763_ (.D(FrameData[1]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit1.Q ));
 sg13g2_dlhq_1 _764_ (.D(FrameData[2]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit2.Q ));
 sg13g2_dlhq_1 _765_ (.D(FrameData[3]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit3.Q ));
 sg13g2_dlhq_1 _766_ (.D(FrameData[4]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit4.Q ));
 sg13g2_dlhq_1 _767_ (.D(FrameData[5]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit5.Q ));
 sg13g2_dlhq_1 _768_ (.D(FrameData[6]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit6.Q ));
 sg13g2_dlhq_1 _769_ (.D(FrameData[7]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit7.Q ));
 sg13g2_dlhq_1 _770_ (.D(FrameData[8]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit8.Q ));
 sg13g2_dlhq_1 _771_ (.D(FrameData[9]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit9.Q ));
 sg13g2_dlhq_1 _772_ (.D(FrameData[10]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit10.Q ));
 sg13g2_dlhq_1 _773_ (.D(FrameData[11]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit11.Q ));
 sg13g2_dlhq_1 _774_ (.D(FrameData[12]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit12.Q ));
 sg13g2_dlhq_1 _775_ (.D(FrameData[13]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit13.Q ));
 sg13g2_dlhq_1 _776_ (.D(FrameData[14]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit14.Q ));
 sg13g2_dlhq_1 _777_ (.D(FrameData[15]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit15.Q ));
 sg13g2_dlhq_1 _778_ (.D(FrameData[16]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit16.Q ));
 sg13g2_dlhq_1 _779_ (.D(FrameData[17]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit17.Q ));
 sg13g2_dlhq_1 _780_ (.D(FrameData[18]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit18.Q ));
 sg13g2_dlhq_1 _781_ (.D(FrameData[19]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit19.Q ));
 sg13g2_dlhq_1 _782_ (.D(FrameData[20]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit20.Q ));
 sg13g2_dlhq_1 _783_ (.D(FrameData[21]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit21.Q ));
 sg13g2_dlhq_1 _784_ (.D(FrameData[22]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit22.Q ));
 sg13g2_dlhq_1 _785_ (.D(FrameData[23]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit23.Q ));
 sg13g2_dlhq_1 _786_ (.D(FrameData[24]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_dlhq_1 _787_ (.D(FrameData[25]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit25.Q ));
 sg13g2_dlhq_1 _788_ (.D(FrameData[26]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_dlhq_1 _789_ (.D(FrameData[27]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit27.Q ));
 sg13g2_dlhq_1 _790_ (.D(FrameData[28]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit28.Q ));
 sg13g2_dlhq_1 _791_ (.D(FrameData[29]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit29.Q ));
 sg13g2_dlhq_1 _792_ (.D(FrameData[30]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_dlhq_1 _793_ (.D(FrameData[31]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit31.Q ));
 sg13g2_buf_1 _794_ (.A(clknet_1_0__leaf_UserCLK),
    .X(CLK_TT_PROJECT));
 sg13g2_buf_1 _795_ (.A(\Inst_W_TT_IF_switch_matrix.E1BEG0 ),
    .X(E1BEG[0]));
 sg13g2_buf_1 _796_ (.A(\Inst_W_TT_IF_switch_matrix.E1BEG1 ),
    .X(E1BEG[1]));
 sg13g2_buf_1 _797_ (.A(\Inst_W_TT_IF_switch_matrix.E1BEG2 ),
    .X(E1BEG[2]));
 sg13g2_buf_1 _798_ (.A(\Inst_W_TT_IF_switch_matrix.E1BEG3 ),
    .X(E1BEG[3]));
 sg13g2_buf_1 _799_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEG0 ),
    .X(E2BEG[0]));
 sg13g2_buf_1 _800_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEG1 ),
    .X(E2BEG[1]));
 sg13g2_buf_1 _801_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEG2 ),
    .X(E2BEG[2]));
 sg13g2_buf_1 _802_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEG3 ),
    .X(E2BEG[3]));
 sg13g2_buf_1 _803_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEG4 ),
    .X(E2BEG[4]));
 sg13g2_buf_1 _804_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEG5 ),
    .X(E2BEG[5]));
 sg13g2_buf_1 _805_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEG6 ),
    .X(E2BEG[6]));
 sg13g2_buf_1 _806_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEG7 ),
    .X(E2BEG[7]));
 sg13g2_buf_1 _807_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEGb0 ),
    .X(E2BEGb[0]));
 sg13g2_buf_1 _808_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEGb1 ),
    .X(E2BEGb[1]));
 sg13g2_buf_1 _809_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEGb2 ),
    .X(E2BEGb[2]));
 sg13g2_buf_1 _810_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEGb3 ),
    .X(E2BEGb[3]));
 sg13g2_buf_1 _811_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEGb4 ),
    .X(E2BEGb[4]));
 sg13g2_buf_1 _812_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEGb5 ),
    .X(E2BEGb[5]));
 sg13g2_buf_1 _813_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEGb6 ),
    .X(E2BEGb[6]));
 sg13g2_buf_1 _814_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEGb7 ),
    .X(E2BEGb[7]));
 sg13g2_buf_1 _815_ (.A(\Inst_W_TT_IF_switch_matrix.E6BEG0 ),
    .X(E6BEG[0]));
 sg13g2_buf_1 _816_ (.A(\Inst_W_TT_IF_switch_matrix.E6BEG1 ),
    .X(E6BEG[1]));
 sg13g2_buf_1 _817_ (.A(\Inst_W_TT_IF_switch_matrix.E6BEG2 ),
    .X(E6BEG[2]));
 sg13g2_buf_1 _818_ (.A(\Inst_W_TT_IF_switch_matrix.E6BEG3 ),
    .X(E6BEG[3]));
 sg13g2_buf_1 _819_ (.A(\Inst_W_TT_IF_switch_matrix.E6BEG4 ),
    .X(E6BEG[4]));
 sg13g2_buf_1 _820_ (.A(\Inst_W_TT_IF_switch_matrix.E6BEG5 ),
    .X(E6BEG[5]));
 sg13g2_buf_1 _821_ (.A(\Inst_W_TT_IF_switch_matrix.E6BEG6 ),
    .X(E6BEG[6]));
 sg13g2_buf_1 _822_ (.A(\Inst_W_TT_IF_switch_matrix.E6BEG7 ),
    .X(E6BEG[7]));
 sg13g2_buf_1 _823_ (.A(\Inst_W_TT_IF_switch_matrix.E6BEG8 ),
    .X(E6BEG[8]));
 sg13g2_buf_1 _824_ (.A(\Inst_W_TT_IF_switch_matrix.E6BEG9 ),
    .X(E6BEG[9]));
 sg13g2_buf_1 _825_ (.A(\Inst_W_TT_IF_switch_matrix.E6BEG10 ),
    .X(E6BEG[10]));
 sg13g2_buf_1 _826_ (.A(\Inst_W_TT_IF_switch_matrix.E6BEG11 ),
    .X(E6BEG[11]));
 sg13g2_buf_1 _827_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG0 ),
    .X(EE4BEG[0]));
 sg13g2_buf_1 _828_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG1 ),
    .X(EE4BEG[1]));
 sg13g2_buf_1 _829_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG2 ),
    .X(EE4BEG[2]));
 sg13g2_buf_1 _830_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG3 ),
    .X(EE4BEG[3]));
 sg13g2_buf_1 _831_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG4 ),
    .X(EE4BEG[4]));
 sg13g2_buf_1 _832_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG5 ),
    .X(EE4BEG[5]));
 sg13g2_buf_1 _833_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG6 ),
    .X(EE4BEG[6]));
 sg13g2_buf_1 _834_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG7 ),
    .X(EE4BEG[7]));
 sg13g2_buf_1 _835_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG8 ),
    .X(EE4BEG[8]));
 sg13g2_buf_1 _836_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG9 ),
    .X(EE4BEG[9]));
 sg13g2_buf_1 _837_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG10 ),
    .X(EE4BEG[10]));
 sg13g2_buf_1 _838_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG11 ),
    .X(EE4BEG[11]));
 sg13g2_buf_1 _839_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG12 ),
    .X(EE4BEG[12]));
 sg13g2_buf_1 _840_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG13 ),
    .X(EE4BEG[13]));
 sg13g2_buf_1 _841_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG14 ),
    .X(EE4BEG[14]));
 sg13g2_buf_1 _842_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG15 ),
    .X(EE4BEG[15]));
 sg13g2_buf_1 _843_ (.A(FrameData[0]),
    .X(FrameData_O[0]));
 sg13g2_buf_1 _844_ (.A(FrameData[1]),
    .X(FrameData_O[1]));
 sg13g2_buf_1 _845_ (.A(FrameData[2]),
    .X(FrameData_O[2]));
 sg13g2_buf_1 _846_ (.A(FrameData[3]),
    .X(FrameData_O[3]));
 sg13g2_buf_1 _847_ (.A(FrameData[4]),
    .X(FrameData_O[4]));
 sg13g2_buf_1 _848_ (.A(FrameData[5]),
    .X(FrameData_O[5]));
 sg13g2_buf_1 _849_ (.A(FrameData[6]),
    .X(FrameData_O[6]));
 sg13g2_buf_1 _850_ (.A(FrameData[7]),
    .X(FrameData_O[7]));
 sg13g2_buf_1 _851_ (.A(FrameData[8]),
    .X(FrameData_O[8]));
 sg13g2_buf_1 _852_ (.A(FrameData[9]),
    .X(FrameData_O[9]));
 sg13g2_buf_1 _853_ (.A(FrameData[10]),
    .X(FrameData_O[10]));
 sg13g2_buf_1 _854_ (.A(FrameData[11]),
    .X(FrameData_O[11]));
 sg13g2_buf_1 _855_ (.A(FrameData[12]),
    .X(FrameData_O[12]));
 sg13g2_buf_1 _856_ (.A(FrameData[13]),
    .X(FrameData_O[13]));
 sg13g2_buf_1 _857_ (.A(FrameData[14]),
    .X(FrameData_O[14]));
 sg13g2_buf_1 _858_ (.A(FrameData[15]),
    .X(FrameData_O[15]));
 sg13g2_buf_1 _859_ (.A(FrameData[16]),
    .X(FrameData_O[16]));
 sg13g2_buf_1 _860_ (.A(FrameData[17]),
    .X(FrameData_O[17]));
 sg13g2_buf_1 _861_ (.A(FrameData[18]),
    .X(FrameData_O[18]));
 sg13g2_buf_1 _862_ (.A(FrameData[19]),
    .X(FrameData_O[19]));
 sg13g2_buf_1 _863_ (.A(FrameData[20]),
    .X(FrameData_O[20]));
 sg13g2_buf_1 _864_ (.A(FrameData[21]),
    .X(FrameData_O[21]));
 sg13g2_buf_1 _865_ (.A(FrameData[22]),
    .X(FrameData_O[22]));
 sg13g2_buf_1 _866_ (.A(FrameData[23]),
    .X(FrameData_O[23]));
 sg13g2_buf_1 _867_ (.A(FrameData[24]),
    .X(FrameData_O[24]));
 sg13g2_buf_1 _868_ (.A(FrameData[25]),
    .X(FrameData_O[25]));
 sg13g2_buf_1 _869_ (.A(FrameData[26]),
    .X(FrameData_O[26]));
 sg13g2_buf_1 _870_ (.A(FrameData[27]),
    .X(FrameData_O[27]));
 sg13g2_buf_1 _871_ (.A(FrameData[28]),
    .X(FrameData_O[28]));
 sg13g2_buf_1 _872_ (.A(FrameData[29]),
    .X(FrameData_O[29]));
 sg13g2_buf_1 _873_ (.A(FrameData[30]),
    .X(FrameData_O[30]));
 sg13g2_buf_1 _874_ (.A(FrameData[31]),
    .X(FrameData_O[31]));
 sg13g2_buf_1 _875_ (.A(FrameStrobe[0]),
    .X(FrameStrobe_O[0]));
 sg13g2_buf_1 _876_ (.A(FrameStrobe[1]),
    .X(FrameStrobe_O[1]));
 sg13g2_buf_1 _877_ (.A(FrameStrobe[2]),
    .X(FrameStrobe_O[2]));
 sg13g2_buf_1 _878_ (.A(FrameStrobe[3]),
    .X(FrameStrobe_O[3]));
 sg13g2_buf_1 _879_ (.A(FrameStrobe[4]),
    .X(FrameStrobe_O[4]));
 sg13g2_buf_1 _880_ (.A(FrameStrobe[5]),
    .X(FrameStrobe_O[5]));
 sg13g2_buf_1 _881_ (.A(FrameStrobe[6]),
    .X(FrameStrobe_O[6]));
 sg13g2_buf_1 _882_ (.A(FrameStrobe[7]),
    .X(FrameStrobe_O[7]));
 sg13g2_buf_1 _883_ (.A(FrameStrobe[8]),
    .X(FrameStrobe_O[8]));
 sg13g2_buf_1 _884_ (.A(FrameStrobe[9]),
    .X(FrameStrobe_O[9]));
 sg13g2_buf_1 _885_ (.A(FrameStrobe[10]),
    .X(FrameStrobe_O[10]));
 sg13g2_buf_1 _886_ (.A(FrameStrobe[11]),
    .X(FrameStrobe_O[11]));
 sg13g2_buf_1 _887_ (.A(FrameStrobe[12]),
    .X(FrameStrobe_O[12]));
 sg13g2_buf_1 _888_ (.A(FrameStrobe[13]),
    .X(FrameStrobe_O[13]));
 sg13g2_buf_1 _889_ (.A(FrameStrobe[14]),
    .X(FrameStrobe_O[14]));
 sg13g2_buf_1 _890_ (.A(FrameStrobe[15]),
    .X(FrameStrobe_O[15]));
 sg13g2_buf_1 _891_ (.A(FrameStrobe[16]),
    .X(FrameStrobe_O[16]));
 sg13g2_buf_1 _892_ (.A(FrameStrobe[17]),
    .X(FrameStrobe_O[17]));
 sg13g2_buf_1 _893_ (.A(FrameStrobe[18]),
    .X(FrameStrobe_O[18]));
 sg13g2_buf_1 _894_ (.A(FrameStrobe[19]),
    .X(FrameStrobe_O[19]));
 sg13g2_buf_1 _895_ (.A(\Inst_W_TT_IF_switch_matrix.N1BEG0 ),
    .X(N1BEG[0]));
 sg13g2_buf_1 _896_ (.A(\Inst_W_TT_IF_switch_matrix.N1BEG1 ),
    .X(N1BEG[1]));
 sg13g2_buf_1 _897_ (.A(\Inst_W_TT_IF_switch_matrix.N1BEG2 ),
    .X(N1BEG[2]));
 sg13g2_buf_1 _898_ (.A(\Inst_W_TT_IF_switch_matrix.N1BEG3 ),
    .X(N1BEG[3]));
 sg13g2_buf_1 _899_ (.A(\Inst_W_TT_IF_switch_matrix.N2BEG0 ),
    .X(N2BEG[0]));
 sg13g2_buf_1 _900_ (.A(\Inst_W_TT_IF_switch_matrix.N2BEG1 ),
    .X(N2BEG[1]));
 sg13g2_buf_1 _901_ (.A(\Inst_W_TT_IF_switch_matrix.N2BEG2 ),
    .X(N2BEG[2]));
 sg13g2_buf_1 _902_ (.A(\Inst_W_TT_IF_switch_matrix.N2BEG3 ),
    .X(N2BEG[3]));
 sg13g2_buf_1 _903_ (.A(\Inst_W_TT_IF_switch_matrix.N2BEG4 ),
    .X(N2BEG[4]));
 sg13g2_buf_1 _904_ (.A(\Inst_W_TT_IF_switch_matrix.N2BEG5 ),
    .X(N2BEG[5]));
 sg13g2_buf_1 _905_ (.A(\Inst_W_TT_IF_switch_matrix.N2BEG6 ),
    .X(N2BEG[6]));
 sg13g2_buf_1 _906_ (.A(\Inst_W_TT_IF_switch_matrix.N2BEG7 ),
    .X(N2BEG[7]));
 sg13g2_buf_1 _907_ (.A(N2MID[0]),
    .X(N2BEGb[0]));
 sg13g2_buf_1 _908_ (.A(N2MID[1]),
    .X(N2BEGb[1]));
 sg13g2_buf_1 _909_ (.A(N2MID[2]),
    .X(N2BEGb[2]));
 sg13g2_buf_1 _910_ (.A(N2MID[3]),
    .X(N2BEGb[3]));
 sg13g2_buf_1 _911_ (.A(N2MID[4]),
    .X(N2BEGb[4]));
 sg13g2_buf_1 _912_ (.A(N2MID[5]),
    .X(N2BEGb[5]));
 sg13g2_buf_1 _913_ (.A(N2MID[6]),
    .X(N2BEGb[6]));
 sg13g2_buf_1 _914_ (.A(N2MID[7]),
    .X(N2BEGb[7]));
 sg13g2_buf_1 _915_ (.A(N4END[4]),
    .X(N4BEG[0]));
 sg13g2_buf_1 _916_ (.A(N4END[5]),
    .X(N4BEG[1]));
 sg13g2_buf_1 _917_ (.A(N4END[6]),
    .X(N4BEG[2]));
 sg13g2_buf_1 _918_ (.A(N4END[7]),
    .X(N4BEG[3]));
 sg13g2_buf_1 _919_ (.A(N4END[8]),
    .X(N4BEG[4]));
 sg13g2_buf_1 _920_ (.A(N4END[9]),
    .X(N4BEG[5]));
 sg13g2_buf_1 _921_ (.A(N4END[10]),
    .X(N4BEG[6]));
 sg13g2_buf_1 _922_ (.A(N4END[11]),
    .X(N4BEG[7]));
 sg13g2_buf_1 _923_ (.A(N4END[12]),
    .X(N4BEG[8]));
 sg13g2_buf_1 _924_ (.A(N4END[13]),
    .X(N4BEG[9]));
 sg13g2_buf_1 _925_ (.A(N4END[14]),
    .X(N4BEG[10]));
 sg13g2_buf_1 _926_ (.A(N4END[15]),
    .X(N4BEG[11]));
 sg13g2_buf_1 _927_ (.A(\Inst_W_TT_IF_switch_matrix.N4BEG0 ),
    .X(N4BEG[12]));
 sg13g2_buf_1 _928_ (.A(\Inst_W_TT_IF_switch_matrix.N4BEG1 ),
    .X(N4BEG[13]));
 sg13g2_buf_1 _929_ (.A(\Inst_W_TT_IF_switch_matrix.N4BEG2 ),
    .X(N4BEG[14]));
 sg13g2_buf_1 _930_ (.A(\Inst_W_TT_IF_switch_matrix.N4BEG3 ),
    .X(N4BEG[15]));
 sg13g2_buf_1 _931_ (.A(\Inst_W_TT_IF_switch_matrix.S1BEG0 ),
    .X(S1BEG[0]));
 sg13g2_buf_1 _932_ (.A(\Inst_W_TT_IF_switch_matrix.S1BEG1 ),
    .X(S1BEG[1]));
 sg13g2_buf_1 _933_ (.A(\Inst_W_TT_IF_switch_matrix.S1BEG2 ),
    .X(S1BEG[2]));
 sg13g2_buf_1 _934_ (.A(\Inst_W_TT_IF_switch_matrix.S1BEG3 ),
    .X(S1BEG[3]));
 sg13g2_buf_1 _935_ (.A(\Inst_W_TT_IF_switch_matrix.S2BEG0 ),
    .X(S2BEG[0]));
 sg13g2_buf_1 _936_ (.A(\Inst_W_TT_IF_switch_matrix.S2BEG1 ),
    .X(S2BEG[1]));
 sg13g2_buf_1 _937_ (.A(\Inst_W_TT_IF_switch_matrix.S2BEG2 ),
    .X(S2BEG[2]));
 sg13g2_buf_1 _938_ (.A(\Inst_W_TT_IF_switch_matrix.S2BEG3 ),
    .X(S2BEG[3]));
 sg13g2_buf_1 _939_ (.A(\Inst_W_TT_IF_switch_matrix.S2BEG4 ),
    .X(S2BEG[4]));
 sg13g2_buf_1 _940_ (.A(\Inst_W_TT_IF_switch_matrix.S2BEG5 ),
    .X(S2BEG[5]));
 sg13g2_buf_1 _941_ (.A(\Inst_W_TT_IF_switch_matrix.S2BEG6 ),
    .X(S2BEG[6]));
 sg13g2_buf_1 _942_ (.A(\Inst_W_TT_IF_switch_matrix.S2BEG7 ),
    .X(S2BEG[7]));
 sg13g2_buf_1 _943_ (.A(S2MID[0]),
    .X(S2BEGb[0]));
 sg13g2_buf_1 _944_ (.A(S2MID[1]),
    .X(S2BEGb[1]));
 sg13g2_buf_1 _945_ (.A(S2MID[2]),
    .X(S2BEGb[2]));
 sg13g2_buf_1 _946_ (.A(S2MID[3]),
    .X(S2BEGb[3]));
 sg13g2_buf_1 _947_ (.A(S2MID[4]),
    .X(S2BEGb[4]));
 sg13g2_buf_1 _948_ (.A(S2MID[5]),
    .X(S2BEGb[5]));
 sg13g2_buf_1 _949_ (.A(S2MID[6]),
    .X(S2BEGb[6]));
 sg13g2_buf_1 _950_ (.A(S2MID[7]),
    .X(S2BEGb[7]));
 sg13g2_buf_1 _951_ (.A(S4END[4]),
    .X(S4BEG[0]));
 sg13g2_buf_1 _952_ (.A(S4END[5]),
    .X(S4BEG[1]));
 sg13g2_buf_1 _953_ (.A(S4END[6]),
    .X(S4BEG[2]));
 sg13g2_buf_1 _954_ (.A(S4END[7]),
    .X(S4BEG[3]));
 sg13g2_buf_1 _955_ (.A(S4END[8]),
    .X(S4BEG[4]));
 sg13g2_buf_1 _956_ (.A(S4END[9]),
    .X(S4BEG[5]));
 sg13g2_buf_1 _957_ (.A(S4END[10]),
    .X(S4BEG[6]));
 sg13g2_buf_1 _958_ (.A(S4END[11]),
    .X(S4BEG[7]));
 sg13g2_buf_1 _959_ (.A(S4END[12]),
    .X(S4BEG[8]));
 sg13g2_buf_1 _960_ (.A(S4END[13]),
    .X(S4BEG[9]));
 sg13g2_buf_1 _961_ (.A(S4END[14]),
    .X(S4BEG[10]));
 sg13g2_buf_1 _962_ (.A(S4END[15]),
    .X(S4BEG[11]));
 sg13g2_buf_1 _963_ (.A(\Inst_W_TT_IF_switch_matrix.S4BEG0 ),
    .X(S4BEG[12]));
 sg13g2_buf_1 _964_ (.A(\Inst_W_TT_IF_switch_matrix.S4BEG1 ),
    .X(S4BEG[13]));
 sg13g2_buf_1 _965_ (.A(\Inst_W_TT_IF_switch_matrix.S4BEG2 ),
    .X(S4BEG[14]));
 sg13g2_buf_1 _966_ (.A(\Inst_W_TT_IF_switch_matrix.S4BEG3 ),
    .X(S4BEG[15]));
 sg13g2_buf_1 _967_ (.A(clknet_1_1__leaf_UserCLK),
    .X(UserCLKo));
 sg13g2_buf_8 clkbuf_0_UserCLK (.A(UserCLK),
    .X(clknet_0_UserCLK));
 sg13g2_buf_8 clkbuf_1_0__f_UserCLK (.A(clknet_0_UserCLK),
    .X(clknet_1_0__leaf_UserCLK));
 sg13g2_buf_8 clkbuf_1_1__f_UserCLK (.A(clknet_0_UserCLK),
    .X(clknet_1_1__leaf_UserCLK));
 sg13g2_antennanp ANTENNA_1 (.A(FrameStrobe[12]));
 sg13g2_antennanp ANTENNA_2 (.A(FrameStrobe[15]));
 sg13g2_antennanp ANTENNA_3 (.A(FrameStrobe[16]));
 sg13g2_antennanp ANTENNA_4 (.A(FrameStrobe[9]));
 sg13g2_antennanp ANTENNA_5 (.A(N2END[6]));
 sg13g2_antennanp ANTENNA_6 (.A(N2END[7]));
 sg13g2_antennanp ANTENNA_7 (.A(N2MID[3]));
 sg13g2_antennanp ANTENNA_8 (.A(N2MID[3]));
 sg13g2_antennanp ANTENNA_9 (.A(N2MID[3]));
 sg13g2_antennanp ANTENNA_10 (.A(N2MID[4]));
 sg13g2_antennanp ANTENNA_11 (.A(N2MID[4]));
 sg13g2_antennanp ANTENNA_12 (.A(N2MID[4]));
 sg13g2_antennanp ANTENNA_13 (.A(N4END[8]));
 sg13g2_antennanp ANTENNA_14 (.A(FrameStrobe[11]));
 sg13g2_antennanp ANTENNA_15 (.A(FrameStrobe[13]));
 sg13g2_antennanp ANTENNA_16 (.A(FrameStrobe[17]));
 sg13g2_antennanp ANTENNA_17 (.A(FrameStrobe[18]));
 sg13g2_antennanp ANTENNA_18 (.A(N4END[12]));
 sg13g2_antennanp ANTENNA_19 (.A(N4END[13]));
 sg13g2_antennanp ANTENNA_20 (.A(N4END[15]));
 sg13g2_antennanp ANTENNA_21 (.A(N4END[4]));
 sg13g2_antennanp ANTENNA_22 (.A(N4END[5]));
 sg13g2_antennanp ANTENNA_23 (.A(N4END[7]));
 sg13g2_antennanp ANTENNA_24 (.A(S2MID[1]));
 sg13g2_antennanp ANTENNA_25 (.A(S2MID[1]));
 sg13g2_antennanp ANTENNA_26 (.A(S2MID[1]));
 sg13g2_antennanp ANTENNA_27 (.A(S2MID[1]));
 sg13g2_antennanp ANTENNA_28 (.A(FrameStrobe[14]));
 sg13g2_antennanp ANTENNA_29 (.A(N4END[11]));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_4 FILLER_0_7 ();
 sg13g2_fill_1 FILLER_0_11 ();
 sg13g2_fill_2 FILLER_0_60 ();
 sg13g2_fill_1 FILLER_0_86 ();
 sg13g2_fill_1 FILLER_0_103 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_4 FILLER_0_119 ();
 sg13g2_fill_2 FILLER_0_123 ();
 sg13g2_fill_1 FILLER_0_146 ();
 sg13g2_fill_2 FILLER_0_174 ();
 sg13g2_decap_8 FILLER_0_193 ();
 sg13g2_fill_1 FILLER_1_0 ();
 sg13g2_fill_2 FILLER_1_65 ();
 sg13g2_fill_1 FILLER_1_82 ();
 sg13g2_fill_2 FILLER_1_87 ();
 sg13g2_fill_1 FILLER_1_94 ();
 sg13g2_fill_1 FILLER_1_145 ();
 sg13g2_fill_1 FILLER_1_178 ();
 sg13g2_decap_4 FILLER_1_196 ();
 sg13g2_decap_4 FILLER_2_0 ();
 sg13g2_fill_2 FILLER_2_25 ();
 sg13g2_fill_1 FILLER_2_66 ();
 sg13g2_fill_1 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_121 ();
 sg13g2_fill_2 FILLER_2_128 ();
 sg13g2_fill_1 FILLER_2_130 ();
 sg13g2_fill_2 FILLER_2_139 ();
 sg13g2_fill_2 FILLER_2_178 ();
 sg13g2_fill_2 FILLER_2_197 ();
 sg13g2_fill_1 FILLER_2_199 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_4 FILLER_3_7 ();
 sg13g2_fill_2 FILLER_3_11 ();
 sg13g2_fill_1 FILLER_3_34 ();
 sg13g2_fill_1 FILLER_3_59 ();
 sg13g2_decap_4 FILLER_3_100 ();
 sg13g2_decap_8 FILLER_3_121 ();
 sg13g2_decap_8 FILLER_3_128 ();
 sg13g2_fill_2 FILLER_3_174 ();
 sg13g2_fill_2 FILLER_3_198 ();
 sg13g2_fill_1 FILLER_4_80 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_143 ();
 sg13g2_decap_8 FILLER_4_150 ();
 sg13g2_decap_4 FILLER_4_173 ();
 sg13g2_fill_2 FILLER_4_177 ();
 sg13g2_fill_2 FILLER_5_39 ();
 sg13g2_fill_1 FILLER_5_41 ();
 sg13g2_fill_1 FILLER_5_59 ();
 sg13g2_decap_8 FILLER_5_81 ();
 sg13g2_fill_1 FILLER_5_88 ();
 sg13g2_decap_4 FILLER_5_174 ();
 sg13g2_fill_2 FILLER_5_183 ();
 sg13g2_fill_1 FILLER_5_185 ();
 sg13g2_decap_4 FILLER_5_196 ();
 sg13g2_fill_2 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_2 ();
 sg13g2_fill_2 FILLER_6_58 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_fill_1 FILLER_6_105 ();
 sg13g2_fill_2 FILLER_6_123 ();
 sg13g2_fill_1 FILLER_6_142 ();
 sg13g2_fill_2 FILLER_6_176 ();
 sg13g2_fill_1 FILLER_7_17 ();
 sg13g2_decap_8 FILLER_7_64 ();
 sg13g2_decap_4 FILLER_7_71 ();
 sg13g2_fill_2 FILLER_7_75 ();
 sg13g2_decap_4 FILLER_7_98 ();
 sg13g2_fill_2 FILLER_7_102 ();
 sg13g2_decap_8 FILLER_7_142 ();
 sg13g2_fill_2 FILLER_7_149 ();
 sg13g2_fill_2 FILLER_7_168 ();
 sg13g2_fill_2 FILLER_7_198 ();
 sg13g2_decap_8 FILLER_8_39 ();
 sg13g2_decap_8 FILLER_8_46 ();
 sg13g2_fill_1 FILLER_8_53 ();
 sg13g2_fill_2 FILLER_8_71 ();
 sg13g2_fill_1 FILLER_8_73 ();
 sg13g2_decap_8 FILLER_8_129 ();
 sg13g2_decap_4 FILLER_8_195 ();
 sg13g2_fill_1 FILLER_8_199 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_35 ();
 sg13g2_fill_1 FILLER_9_74 ();
 sg13g2_decap_4 FILLER_9_126 ();
 sg13g2_fill_2 FILLER_9_130 ();
 sg13g2_decap_8 FILLER_9_166 ();
 sg13g2_fill_2 FILLER_9_173 ();
 sg13g2_fill_2 FILLER_9_183 ();
 sg13g2_fill_1 FILLER_9_185 ();
 sg13g2_decap_4 FILLER_9_196 ();
 sg13g2_fill_2 FILLER_10_17 ();
 sg13g2_decap_8 FILLER_10_39 ();
 sg13g2_fill_1 FILLER_10_46 ();
 sg13g2_decap_8 FILLER_10_64 ();
 sg13g2_fill_2 FILLER_10_71 ();
 sg13g2_fill_1 FILLER_10_73 ();
 sg13g2_decap_8 FILLER_10_112 ();
 sg13g2_decap_4 FILLER_10_119 ();
 sg13g2_fill_1 FILLER_10_140 ();
 sg13g2_fill_2 FILLER_10_154 ();
 sg13g2_fill_1 FILLER_10_199 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_2 ();
 sg13g2_fill_1 FILLER_11_20 ();
 sg13g2_fill_2 FILLER_11_28 ();
 sg13g2_fill_2 FILLER_11_85 ();
 sg13g2_fill_1 FILLER_11_87 ();
 sg13g2_decap_4 FILLER_11_100 ();
 sg13g2_fill_2 FILLER_11_162 ();
 sg13g2_decap_8 FILLER_12_38 ();
 sg13g2_decap_8 FILLER_12_45 ();
 sg13g2_decap_8 FILLER_12_52 ();
 sg13g2_decap_4 FILLER_12_59 ();
 sg13g2_fill_2 FILLER_12_63 ();
 sg13g2_fill_2 FILLER_12_103 ();
 sg13g2_fill_1 FILLER_12_105 ();
 sg13g2_fill_2 FILLER_12_123 ();
 sg13g2_decap_4 FILLER_12_163 ();
 sg13g2_fill_2 FILLER_12_167 ();
 sg13g2_decap_4 FILLER_12_196 ();
 sg13g2_fill_2 FILLER_13_17 ();
 sg13g2_decap_4 FILLER_13_29 ();
 sg13g2_decap_4 FILLER_13_43 ();
 sg13g2_fill_1 FILLER_13_47 ();
 sg13g2_fill_2 FILLER_13_65 ();
 sg13g2_fill_1 FILLER_13_67 ();
 sg13g2_fill_2 FILLER_13_94 ();
 sg13g2_fill_1 FILLER_13_96 ();
 sg13g2_fill_2 FILLER_13_114 ();
 sg13g2_fill_1 FILLER_13_116 ();
 sg13g2_decap_8 FILLER_13_132 ();
 sg13g2_decap_8 FILLER_13_139 ();
 sg13g2_decap_8 FILLER_13_146 ();
 sg13g2_decap_8 FILLER_13_153 ();
 sg13g2_decap_8 FILLER_13_160 ();
 sg13g2_decap_4 FILLER_13_167 ();
 sg13g2_fill_1 FILLER_13_171 ();
 sg13g2_fill_2 FILLER_13_198 ();
 sg13g2_decap_8 FILLER_14_17 ();
 sg13g2_decap_8 FILLER_14_29 ();
 sg13g2_decap_8 FILLER_14_36 ();
 sg13g2_fill_1 FILLER_14_43 ();
 sg13g2_fill_2 FILLER_14_141 ();
 sg13g2_fill_1 FILLER_14_143 ();
 sg13g2_fill_2 FILLER_14_161 ();
 sg13g2_fill_1 FILLER_14_185 ();
 sg13g2_fill_1 FILLER_14_199 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_4 FILLER_15_7 ();
 sg13g2_fill_1 FILLER_15_66 ();
 sg13g2_decap_4 FILLER_15_94 ();
 sg13g2_fill_2 FILLER_15_98 ();
 sg13g2_decap_4 FILLER_15_117 ();
 sg13g2_fill_2 FILLER_15_128 ();
 sg13g2_fill_1 FILLER_15_130 ();
 sg13g2_fill_1 FILLER_15_148 ();
 sg13g2_decap_4 FILLER_15_196 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_4 FILLER_16_42 ();
 sg13g2_fill_1 FILLER_16_139 ();
 sg13g2_fill_2 FILLER_16_171 ();
 sg13g2_decap_4 FILLER_16_195 ();
 sg13g2_fill_1 FILLER_16_199 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_fill_1 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_36 ();
 sg13g2_decap_4 FILLER_17_43 ();
 sg13g2_fill_1 FILLER_17_47 ();
 sg13g2_decap_4 FILLER_17_69 ();
 sg13g2_fill_2 FILLER_17_73 ();
 sg13g2_decap_8 FILLER_17_90 ();
 sg13g2_decap_4 FILLER_17_97 ();
 sg13g2_fill_1 FILLER_17_101 ();
 sg13g2_fill_2 FILLER_17_119 ();
 sg13g2_decap_8 FILLER_17_170 ();
 sg13g2_fill_1 FILLER_17_199 ();
 sg13g2_fill_1 FILLER_18_32 ();
 sg13g2_fill_2 FILLER_18_50 ();
 sg13g2_fill_1 FILLER_18_69 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_fill_1 FILLER_18_98 ();
 sg13g2_fill_2 FILLER_18_116 ();
 sg13g2_fill_1 FILLER_18_118 ();
 sg13g2_fill_1 FILLER_18_146 ();
 sg13g2_decap_8 FILLER_18_164 ();
 sg13g2_fill_1 FILLER_19_17 ();
 sg13g2_decap_8 FILLER_19_90 ();
 sg13g2_fill_2 FILLER_19_97 ();
 sg13g2_fill_1 FILLER_19_137 ();
 sg13g2_fill_2 FILLER_19_176 ();
 sg13g2_fill_1 FILLER_19_178 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_19 ();
 sg13g2_fill_2 FILLER_20_67 ();
 sg13g2_decap_8 FILLER_20_103 ();
 sg13g2_fill_1 FILLER_20_110 ();
 sg13g2_decap_8 FILLER_20_128 ();
 sg13g2_decap_8 FILLER_20_135 ();
 sg13g2_decap_4 FILLER_20_142 ();
 sg13g2_fill_2 FILLER_20_146 ();
 sg13g2_fill_2 FILLER_20_175 ();
 sg13g2_fill_1 FILLER_20_199 ();
 sg13g2_fill_2 FILLER_21_17 ();
 sg13g2_fill_1 FILLER_21_41 ();
 sg13g2_fill_1 FILLER_21_64 ();
 sg13g2_decap_8 FILLER_21_82 ();
 sg13g2_fill_2 FILLER_21_89 ();
 sg13g2_fill_1 FILLER_21_129 ();
 sg13g2_fill_1 FILLER_21_152 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_31 ();
 sg13g2_decap_4 FILLER_22_38 ();
 sg13g2_fill_2 FILLER_22_59 ();
 sg13g2_decap_8 FILLER_22_103 ();
 sg13g2_decap_8 FILLER_22_110 ();
 sg13g2_decap_8 FILLER_22_117 ();
 sg13g2_decap_4 FILLER_22_124 ();
 sg13g2_fill_2 FILLER_22_128 ();
 sg13g2_decap_8 FILLER_22_159 ();
 sg13g2_fill_1 FILLER_22_166 ();
 sg13g2_fill_2 FILLER_22_184 ();
 sg13g2_decap_4 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_4 FILLER_23_7 ();
 sg13g2_fill_1 FILLER_23_11 ();
 sg13g2_decap_8 FILLER_23_33 ();
 sg13g2_fill_2 FILLER_23_40 ();
 sg13g2_fill_1 FILLER_23_42 ();
 sg13g2_decap_4 FILLER_23_67 ();
 sg13g2_fill_2 FILLER_23_71 ();
 sg13g2_fill_1 FILLER_23_153 ();
 sg13g2_decap_8 FILLER_24_17 ();
 sg13g2_fill_1 FILLER_24_24 ();
 sg13g2_decap_8 FILLER_24_47 ();
 sg13g2_decap_8 FILLER_24_54 ();
 sg13g2_fill_2 FILLER_24_61 ();
 sg13g2_decap_8 FILLER_24_97 ();
 sg13g2_decap_4 FILLER_24_104 ();
 sg13g2_fill_1 FILLER_24_130 ();
 sg13g2_fill_1 FILLER_24_184 ();
 sg13g2_fill_2 FILLER_24_197 ();
 sg13g2_fill_1 FILLER_24_199 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_2 ();
 sg13g2_fill_1 FILLER_25_20 ();
 sg13g2_decap_4 FILLER_25_38 ();
 sg13g2_fill_1 FILLER_25_42 ();
 sg13g2_fill_1 FILLER_25_98 ();
 sg13g2_decap_4 FILLER_25_124 ();
 sg13g2_fill_2 FILLER_25_150 ();
 sg13g2_decap_8 FILLER_25_169 ();
 sg13g2_fill_1 FILLER_25_176 ();
 sg13g2_fill_2 FILLER_25_198 ();
 sg13g2_decap_4 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_21 ();
 sg13g2_decap_4 FILLER_26_44 ();
 sg13g2_fill_2 FILLER_26_48 ();
 sg13g2_decap_8 FILLER_26_88 ();
 sg13g2_decap_8 FILLER_26_95 ();
 sg13g2_decap_8 FILLER_26_162 ();
 sg13g2_fill_2 FILLER_26_198 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_4 FILLER_27_14 ();
 sg13g2_fill_1 FILLER_27_28 ();
 sg13g2_fill_1 FILLER_27_63 ();
 sg13g2_decap_4 FILLER_27_85 ();
 sg13g2_fill_1 FILLER_27_89 ();
 sg13g2_decap_8 FILLER_27_107 ();
 sg13g2_fill_2 FILLER_27_114 ();
 sg13g2_fill_1 FILLER_27_116 ();
 sg13g2_fill_1 FILLER_27_141 ();
 sg13g2_decap_4 FILLER_27_159 ();
 sg13g2_fill_1 FILLER_27_184 ();
 sg13g2_decap_8 FILLER_27_193 ();
 sg13g2_fill_2 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_46 ();
 sg13g2_decap_8 FILLER_28_53 ();
 sg13g2_fill_1 FILLER_28_72 ();
 sg13g2_fill_1 FILLER_28_145 ();
 sg13g2_fill_2 FILLER_28_163 ();
 sg13g2_fill_1 FILLER_28_165 ();
 sg13g2_fill_2 FILLER_28_183 ();
 sg13g2_fill_2 FILLER_28_197 ();
 sg13g2_fill_1 FILLER_28_199 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_19 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_fill_1 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_147 ();
 sg13g2_decap_8 FILLER_29_154 ();
 sg13g2_decap_8 FILLER_29_161 ();
 sg13g2_decap_8 FILLER_29_168 ();
 sg13g2_fill_2 FILLER_29_175 ();
 sg13g2_fill_1 FILLER_29_177 ();
 sg13g2_fill_1 FILLER_29_199 ();
 sg13g2_fill_2 FILLER_30_31 ();
 sg13g2_fill_1 FILLER_30_45 ();
 sg13g2_fill_1 FILLER_30_80 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_4 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_193 ();
 sg13g2_fill_2 FILLER_31_22 ();
 sg13g2_fill_1 FILLER_31_24 ();
 sg13g2_fill_2 FILLER_31_59 ();
 sg13g2_fill_2 FILLER_31_71 ();
 sg13g2_decap_8 FILLER_31_111 ();
 sg13g2_decap_8 FILLER_31_118 ();
 sg13g2_decap_8 FILLER_31_125 ();
 sg13g2_decap_8 FILLER_31_149 ();
 sg13g2_fill_2 FILLER_31_156 ();
 sg13g2_fill_2 FILLER_31_179 ();
 sg13g2_fill_2 FILLER_31_197 ();
 sg13g2_fill_1 FILLER_31_199 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_4 ();
 sg13g2_fill_2 FILLER_32_22 ();
 sg13g2_fill_1 FILLER_32_24 ();
 sg13g2_decap_8 FILLER_32_46 ();
 sg13g2_decap_8 FILLER_32_53 ();
 sg13g2_fill_1 FILLER_32_81 ();
 sg13g2_decap_8 FILLER_32_120 ();
 sg13g2_fill_2 FILLER_32_127 ();
 sg13g2_decap_8 FILLER_32_150 ();
 sg13g2_fill_1 FILLER_32_157 ();
 sg13g2_decap_4 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_42 ();
 sg13g2_decap_4 FILLER_33_78 ();
 sg13g2_fill_1 FILLER_33_82 ();
 sg13g2_decap_8 FILLER_33_134 ();
 sg13g2_fill_1 FILLER_33_141 ();
 sg13g2_decap_8 FILLER_33_159 ();
 sg13g2_fill_2 FILLER_33_166 ();
 sg13g2_fill_2 FILLER_33_197 ();
 sg13g2_fill_1 FILLER_33_199 ();
 sg13g2_decap_8 FILLER_34_68 ();
 sg13g2_decap_4 FILLER_34_75 ();
 sg13g2_fill_1 FILLER_34_79 ();
 sg13g2_fill_2 FILLER_34_97 ();
 sg13g2_fill_1 FILLER_34_99 ();
 sg13g2_decap_8 FILLER_34_117 ();
 sg13g2_decap_4 FILLER_34_124 ();
 sg13g2_fill_1 FILLER_34_128 ();
 sg13g2_decap_8 FILLER_34_146 ();
 sg13g2_decap_4 FILLER_34_153 ();
 sg13g2_fill_2 FILLER_34_157 ();
 sg13g2_fill_2 FILLER_34_197 ();
 sg13g2_fill_1 FILLER_34_199 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_4 FILLER_35_7 ();
 sg13g2_fill_1 FILLER_35_11 ();
 sg13g2_decap_8 FILLER_35_33 ();
 sg13g2_decap_4 FILLER_35_40 ();
 sg13g2_decap_8 FILLER_35_86 ();
 sg13g2_fill_2 FILLER_35_93 ();
 sg13g2_decap_8 FILLER_35_116 ();
 sg13g2_fill_1 FILLER_35_199 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_4 FILLER_36_45 ();
 sg13g2_fill_2 FILLER_36_66 ();
 sg13g2_decap_8 FILLER_36_85 ();
 sg13g2_decap_8 FILLER_36_113 ();
 sg13g2_decap_4 FILLER_36_120 ();
 sg13g2_fill_1 FILLER_36_124 ();
 sg13g2_fill_2 FILLER_36_163 ();
 sg13g2_fill_2 FILLER_36_198 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_2 ();
 sg13g2_decap_8 FILLER_37_20 ();
 sg13g2_decap_8 FILLER_37_44 ();
 sg13g2_decap_8 FILLER_37_51 ();
 sg13g2_fill_2 FILLER_37_58 ();
 sg13g2_fill_1 FILLER_37_77 ();
 sg13g2_fill_2 FILLER_37_197 ();
 sg13g2_fill_1 FILLER_37_199 ();
 sg13g2_decap_8 FILLER_38_30 ();
 sg13g2_decap_4 FILLER_38_37 ();
 sg13g2_fill_2 FILLER_38_92 ();
 sg13g2_fill_1 FILLER_38_94 ();
 sg13g2_decap_8 FILLER_38_116 ();
 sg13g2_decap_8 FILLER_38_123 ();
 sg13g2_fill_1 FILLER_38_130 ();
 sg13g2_fill_2 FILLER_38_152 ();
 sg13g2_fill_1 FILLER_38_154 ();
 sg13g2_fill_2 FILLER_38_163 ();
 sg13g2_fill_2 FILLER_38_186 ();
 sg13g2_fill_1 FILLER_38_188 ();
 sg13g2_fill_2 FILLER_38_197 ();
 sg13g2_fill_1 FILLER_38_199 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_fill_2 FILLER_39_7 ();
 sg13g2_fill_1 FILLER_39_9 ();
 sg13g2_fill_2 FILLER_39_58 ();
 sg13g2_decap_8 FILLER_39_67 ();
 sg13g2_decap_4 FILLER_39_74 ();
 sg13g2_fill_2 FILLER_39_78 ();
 sg13g2_fill_2 FILLER_39_97 ();
 sg13g2_fill_1 FILLER_39_99 ();
 sg13g2_fill_2 FILLER_39_168 ();
 sg13g2_fill_1 FILLER_39_170 ();
 sg13g2_fill_2 FILLER_40_17 ();
 sg13g2_decap_8 FILLER_40_22 ();
 sg13g2_fill_1 FILLER_40_29 ();
 sg13g2_fill_2 FILLER_40_88 ();
 sg13g2_fill_1 FILLER_40_90 ();
 sg13g2_decap_4 FILLER_40_112 ();
 sg13g2_fill_2 FILLER_40_116 ();
 sg13g2_decap_8 FILLER_40_135 ();
 sg13g2_fill_2 FILLER_40_176 ();
 sg13g2_fill_1 FILLER_40_178 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_fill_2 FILLER_41_14 ();
 sg13g2_fill_2 FILLER_41_64 ();
 sg13g2_fill_1 FILLER_41_76 ();
 sg13g2_decap_4 FILLER_41_94 ();
 sg13g2_fill_1 FILLER_41_98 ();
 sg13g2_fill_2 FILLER_41_137 ();
 sg13g2_fill_1 FILLER_41_139 ();
 sg13g2_fill_2 FILLER_41_186 ();
 sg13g2_fill_1 FILLER_41_188 ();
 sg13g2_fill_2 FILLER_41_197 ();
 sg13g2_fill_1 FILLER_41_199 ();
 sg13g2_fill_1 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_9 ();
 sg13g2_fill_1 FILLER_42_28 ();
 sg13g2_fill_2 FILLER_42_46 ();
 sg13g2_decap_4 FILLER_42_88 ();
 sg13g2_fill_1 FILLER_42_92 ();
 sg13g2_fill_2 FILLER_42_123 ();
 sg13g2_fill_1 FILLER_42_125 ();
 sg13g2_decap_4 FILLER_42_143 ();
 sg13g2_fill_1 FILLER_42_147 ();
 sg13g2_fill_2 FILLER_42_186 ();
 sg13g2_fill_1 FILLER_42_188 ();
 sg13g2_fill_2 FILLER_42_197 ();
 sg13g2_fill_1 FILLER_42_199 ();
 sg13g2_fill_2 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_30 ();
 sg13g2_fill_2 FILLER_43_71 ();
 sg13g2_decap_4 FILLER_43_111 ();
 sg13g2_fill_1 FILLER_43_115 ();
 sg13g2_decap_8 FILLER_43_137 ();
 sg13g2_fill_2 FILLER_43_144 ();
 sg13g2_fill_2 FILLER_43_174 ();
 sg13g2_fill_1 FILLER_43_176 ();
 sg13g2_fill_2 FILLER_43_197 ();
 sg13g2_fill_1 FILLER_43_199 ();
 sg13g2_fill_1 FILLER_44_17 ();
 sg13g2_fill_1 FILLER_44_30 ();
 sg13g2_fill_1 FILLER_44_48 ();
 sg13g2_decap_8 FILLER_44_90 ();
 sg13g2_decap_4 FILLER_44_97 ();
 sg13g2_fill_1 FILLER_44_101 ();
 sg13g2_decap_4 FILLER_44_119 ();
 sg13g2_fill_2 FILLER_44_123 ();
 sg13g2_fill_1 FILLER_44_180 ();
 sg13g2_fill_2 FILLER_44_197 ();
 sg13g2_fill_1 FILLER_44_199 ();
 sg13g2_fill_2 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_48 ();
 sg13g2_fill_1 FILLER_45_50 ();
 sg13g2_fill_2 FILLER_45_198 ();
 sg13g2_fill_1 FILLER_46_0 ();
 sg13g2_decap_4 FILLER_46_5 ();
 sg13g2_fill_1 FILLER_46_9 ();
 sg13g2_decap_8 FILLER_46_13 ();
 sg13g2_fill_2 FILLER_46_20 ();
 sg13g2_fill_1 FILLER_46_22 ();
 sg13g2_fill_2 FILLER_46_31 ();
 sg13g2_fill_1 FILLER_46_33 ();
 sg13g2_decap_8 FILLER_46_75 ();
 sg13g2_fill_2 FILLER_46_82 ();
 sg13g2_fill_1 FILLER_46_84 ();
 sg13g2_fill_1 FILLER_46_199 ();
 sg13g2_fill_1 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_9 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_4 FILLER_47_21 ();
 sg13g2_fill_2 FILLER_47_25 ();
 sg13g2_fill_1 FILLER_47_30 ();
 sg13g2_fill_1 FILLER_47_38 ();
 sg13g2_fill_2 FILLER_47_63 ();
 sg13g2_fill_1 FILLER_47_137 ();
 sg13g2_fill_1 FILLER_47_184 ();
 sg13g2_fill_2 FILLER_47_197 ();
 sg13g2_fill_1 FILLER_47_199 ();
 sg13g2_fill_1 FILLER_48_11 ();
 sg13g2_fill_1 FILLER_48_33 ();
 sg13g2_fill_2 FILLER_48_104 ();
 sg13g2_fill_1 FILLER_48_106 ();
 sg13g2_fill_2 FILLER_48_124 ();
 sg13g2_fill_2 FILLER_48_143 ();
 sg13g2_fill_1 FILLER_48_145 ();
 sg13g2_fill_2 FILLER_49_33 ();
 sg13g2_fill_1 FILLER_49_35 ();
 sg13g2_fill_2 FILLER_49_57 ();
 sg13g2_fill_2 FILLER_49_67 ();
 sg13g2_fill_1 FILLER_49_86 ();
 sg13g2_fill_2 FILLER_49_111 ();
 sg13g2_fill_1 FILLER_49_184 ();
 sg13g2_fill_1 FILLER_50_0 ();
 sg13g2_decap_4 FILLER_50_25 ();
 sg13g2_fill_2 FILLER_50_29 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_4 FILLER_50_42 ();
 sg13g2_fill_1 FILLER_50_46 ();
 sg13g2_decap_4 FILLER_50_89 ();
 sg13g2_fill_1 FILLER_50_93 ();
 sg13g2_fill_2 FILLER_50_111 ();
 sg13g2_fill_1 FILLER_50_117 ();
 sg13g2_fill_2 FILLER_50_135 ();
 sg13g2_fill_1 FILLER_50_137 ();
 sg13g2_fill_2 FILLER_50_175 ();
 sg13g2_fill_1 FILLER_50_184 ();
 sg13g2_fill_1 FILLER_51_4 ();
 sg13g2_decap_4 FILLER_51_29 ();
 sg13g2_decap_8 FILLER_51_53 ();
 sg13g2_fill_2 FILLER_51_143 ();
 sg13g2_fill_1 FILLER_51_145 ();
 sg13g2_fill_2 FILLER_52_7 ();
 sg13g2_fill_2 FILLER_52_47 ();
 sg13g2_fill_1 FILLER_52_49 ();
 sg13g2_fill_1 FILLER_52_71 ();
 sg13g2_fill_1 FILLER_52_166 ();
 sg13g2_fill_2 FILLER_52_198 ();
 sg13g2_fill_2 FILLER_53_3 ();
 sg13g2_fill_1 FILLER_53_5 ();
 sg13g2_decap_8 FILLER_53_40 ();
 sg13g2_decap_4 FILLER_53_47 ();
 sg13g2_fill_2 FILLER_53_68 ();
 sg13g2_fill_1 FILLER_53_70 ();
 sg13g2_fill_2 FILLER_53_75 ();
 sg13g2_fill_1 FILLER_53_77 ();
 sg13g2_fill_2 FILLER_53_158 ();
 sg13g2_fill_1 FILLER_53_160 ();
 sg13g2_fill_2 FILLER_53_197 ();
 sg13g2_fill_1 FILLER_53_199 ();
endmodule
