* NGSPICE file created from N_IO.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlhq_1 abstract view
.subckt sg13g2_dlhq_1 D GATE Q VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux4_1 abstract view
.subckt sg13g2_mux4_1 S0 A0 A1 A2 A3 S1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

.subckt N_IO A_I_top A_O_top A_T_top A_config_C_bit0 A_config_C_bit1 A_config_C_bit2
+ A_config_C_bit3 B_I_top B_O_top B_T_top B_config_C_bit0 B_config_C_bit1 B_config_C_bit2
+ B_config_C_bit3 Ci FrameData[0] FrameData[10] FrameData[11] FrameData[12] FrameData[13]
+ FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18] FrameData[19]
+ FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23] FrameData[24]
+ FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29] FrameData[2]
+ FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5] FrameData[6]
+ FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10] FrameData_O[11]
+ FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15] FrameData_O[16]
+ FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20] FrameData_O[21]
+ FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25] FrameData_O[26]
+ FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30] FrameData_O[31]
+ FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7] FrameData_O[8]
+ FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12] FrameStrobe[13]
+ FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17] FrameStrobe[18]
+ FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4] FrameStrobe[5]
+ FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10]
+ FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15]
+ FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1]
+ FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6]
+ FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1END[0] N1END[1] N1END[2] N1END[3]
+ N2END[0] N2END[1] N2END[2] N2END[3] N2END[4] N2END[5] N2END[6] N2END[7] N2MID[0]
+ N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5] N2MID[6] N2MID[7] N4END[0] N4END[10]
+ N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2] N4END[3] N4END[4]
+ N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] NN4END[0] NN4END[10] NN4END[11] NN4END[12]
+ NN4END[13] NN4END[14] NN4END[15] NN4END[1] NN4END[2] NN4END[3] NN4END[4] NN4END[5]
+ NN4END[6] NN4END[7] NN4END[8] NN4END[9] S1BEG[0] S1BEG[1] S1BEG[2] S1BEG[3] S2BEG[0]
+ S2BEG[1] S2BEG[2] S2BEG[3] S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7] S2BEGb[0] S2BEGb[1]
+ S2BEGb[2] S2BEGb[3] S2BEGb[4] S2BEGb[5] S2BEGb[6] S2BEGb[7] S4BEG[0] S4BEG[10] S4BEG[11]
+ S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1] S4BEG[2] S4BEG[3] S4BEG[4] S4BEG[5]
+ S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] SS4BEG[0] SS4BEG[10] SS4BEG[11] SS4BEG[12] SS4BEG[13]
+ SS4BEG[14] SS4BEG[15] SS4BEG[1] SS4BEG[2] SS4BEG[3] SS4BEG[4] SS4BEG[5] SS4BEG[6]
+ SS4BEG[7] SS4BEG[8] SS4BEG[9] UserCLK UserCLKo VGND VPWR
XFILLER_9_148 VPWR VGND sg13g2_decap_8
X_294_ FrameData[20] FrameData_O[20] VPWR VGND sg13g2_buf_1
X_363_ Inst_N_IO_switch_matrix.SS4BEG1 SS4BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_8_181 VPWR VGND sg13g2_decap_4
X_346_ Inst_N_IO_switch_matrix.S4BEG0 S4BEG[0] VPWR VGND sg13g2_buf_1
X_277_ FrameData[3] FrameData_O[3] VPWR VGND sg13g2_buf_1
XFILLER_11_423 VPWR VGND sg13g2_fill_1
X_200_ FrameData[26] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit26.Q VPWR VGND
+ sg13g2_dlhq_1
X_062_ Inst_N_IO_ConfigMem.Inst_frame3_bit20.Q N2MID[6] N4END[6] NN4END[6] NN4END[14]
+ Inst_N_IO_ConfigMem.Inst_frame3_bit21.Q Inst_N_IO_switch_matrix.S2BEG1 VPWR VGND
+ sg13g2_mux4_1
X_131_ Inst_N_IO_ConfigMem.Inst_frame1_bit20.Q N4END[6] N4END[8] N4END[10] B_O_top
+ Inst_N_IO_ConfigMem.Inst_frame1_bit21.Q Inst_N_IO_switch_matrix.SS4BEG1 VPWR VGND
+ sg13g2_mux4_1
XFILLER_9_66 VPWR VGND sg13g2_fill_2
X_329_ Inst_N_IO_switch_matrix.S1BEG3 S1BEG[3] VPWR VGND sg13g2_buf_1
XFILLER_2_121 VPWR VGND sg13g2_decap_8
XFILLER_11_275 VPWR VGND sg13g2_fill_1
XFILLER_11_264 VPWR VGND sg13g2_decap_8
X_114_ _028_ _029_ Inst_N_IO_ConfigMem.Inst_frame0_bit20.Q _030_ VPWR VGND sg13g2_mux2_1
XFILLER_4_205 VPWR VGND sg13g2_fill_1
XFILLER_1_219 VPWR VGND sg13g2_fill_2
XFILLER_0_230 VPWR VGND sg13g2_fill_2
XFILLER_11_0 VPWR VGND sg13g2_fill_2
X_293_ FrameData[19] FrameData_O[19] VPWR VGND sg13g2_buf_1
X_362_ Inst_N_IO_switch_matrix.SS4BEG0 SS4BEG[0] VPWR VGND sg13g2_buf_1
XFILLER_2_325 VPWR VGND sg13g2_fill_1
XFILLER_2_347 VPWR VGND sg13g2_decap_8
XFILLER_6_119 VPWR VGND sg13g2_decap_4
X_276_ FrameData[2] FrameData_O[2] VPWR VGND sg13g2_buf_1
X_345_ Inst_N_IO_switch_matrix.S2BEGb7 S2BEGb[7] VPWR VGND sg13g2_buf_1
XFILLER_5_152 VPWR VGND sg13g2_decap_8
X_130_ Inst_N_IO_ConfigMem.Inst_frame1_bit22.Q N4END[1] N4END[3] N4END[5] Inst_A_IO_1_bidirectional_frame_config_pass.Q
+ Inst_N_IO_ConfigMem.Inst_frame1_bit23.Q Inst_N_IO_switch_matrix.SS4BEG2 VPWR VGND
+ sg13g2_mux4_1
XFILLER_7_417 VPWR VGND sg13g2_decap_8
X_061_ Inst_N_IO_ConfigMem.Inst_frame3_bit22.Q N2MID[5] N4END[5] NN4END[5] NN4END[13]
+ Inst_N_IO_ConfigMem.Inst_frame3_bit23.Q Inst_N_IO_switch_matrix.S2BEG2 VPWR VGND
+ sg13g2_mux4_1
X_328_ Inst_N_IO_switch_matrix.S1BEG2 S1BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_0_69 VPWR VGND sg13g2_decap_8
XFILLER_0_36 VPWR VGND sg13g2_decap_4
X_259_ FrameData[21] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit21.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_7_258 VPWR VGND sg13g2_fill_1
XFILLER_7_236 VPWR VGND sg13g2_decap_4
X_113_ Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q N2MID[4] N2MID[5] N2MID[6] N2MID[7]
+ Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q _029_ VPWR VGND sg13g2_mux4_1
XFILLER_0_423 VPWR VGND sg13g2_fill_1
XFILLER_0_253 VPWR VGND sg13g2_fill_1
XFILLER_0_220 VPWR VGND sg13g2_decap_4
X_361_ Inst_N_IO_switch_matrix.S4BEG15 S4BEG[15] VPWR VGND sg13g2_buf_1
XFILLER_5_378 VPWR VGND sg13g2_decap_8
X_292_ FrameData[18] FrameData_O[18] VPWR VGND sg13g2_buf_1
XFILLER_10_116 VPWR VGND sg13g2_fill_1
XFILLER_10_105 VPWR VGND sg13g2_decap_8
X_275_ FrameData[1] FrameData_O[1] VPWR VGND sg13g2_buf_1
X_344_ Inst_N_IO_switch_matrix.S2BEGb6 S2BEGb[6] VPWR VGND sg13g2_buf_1
XFILLER_5_120 VPWR VGND sg13g2_decap_8
X_060_ Inst_N_IO_ConfigMem.Inst_frame3_bit24.Q N2MID[4] N4END[4] NN4END[4] NN4END[12]
+ Inst_N_IO_ConfigMem.Inst_frame3_bit25.Q Inst_N_IO_switch_matrix.S2BEG3 VPWR VGND
+ sg13g2_mux4_1
XFILLER_9_79 VPWR VGND sg13g2_fill_1
XFILLER_9_68 VPWR VGND sg13g2_fill_1
XFILLER_9_46 VPWR VGND sg13g2_fill_2
X_327_ Inst_N_IO_switch_matrix.S1BEG1 S1BEG[1] VPWR VGND sg13g2_buf_1
X_258_ FrameData[20] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit20.Q VPWR VGND
+ sg13g2_dlhq_1
X_189_ FrameData[15] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit15.Q VPWR VGND
+ sg13g2_dlhq_1
X_112_ Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q N2MID[0] N2MID[1] N2MID[2] N2MID[3]
+ Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q _028_ VPWR VGND sg13g2_mux4_1
XFILLER_1_0 VPWR VGND sg13g2_decap_8
XFILLER_3_421 VPWR VGND sg13g2_fill_2
XFILLER_11_2 VPWR VGND sg13g2_fill_1
X_360_ Inst_N_IO_switch_matrix.S4BEG14 S4BEG[14] VPWR VGND sg13g2_buf_1
X_291_ FrameData[17] FrameData_O[17] VPWR VGND sg13g2_buf_1
XFILLER_8_151 VPWR VGND sg13g2_decap_4
X_274_ FrameData[0] FrameData_O[0] VPWR VGND sg13g2_buf_1
X_343_ Inst_N_IO_switch_matrix.S2BEGb5 S2BEGb[5] VPWR VGND sg13g2_buf_1
XFILLER_1_382 VPWR VGND sg13g2_fill_2
XFILLER_7_408 VPWR VGND sg13g2_fill_1
X_326_ Inst_N_IO_switch_matrix.S1BEG0 S1BEG[0] VPWR VGND sg13g2_buf_1
X_188_ FrameData[14] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit14.Q VPWR VGND
+ sg13g2_dlhq_1
X_257_ FrameData[19] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_11_212 VPWR VGND sg13g2_decap_8
XFILLER_11_201 VPWR VGND sg13g2_decap_8
X_309_ FrameStrobe[3] FrameStrobe_O[3] VPWR VGND sg13g2_buf_1
X_111_ Inst_N_IO_ConfigMem.Inst_frame0_bit21.Q VPWR _027_ VGND _023_ _026_ sg13g2_o21ai_1
XFILLER_6_271 VPWR VGND sg13g2_fill_2
XFILLER_3_274 VPWR VGND sg13g2_decap_4
XFILLER_0_288 VPWR VGND sg13g2_fill_2
XFILLER_5_314 VPWR VGND sg13g2_decap_4
X_290_ FrameData[16] FrameData_O[16] VPWR VGND sg13g2_buf_1
XFILLER_8_185 VPWR VGND sg13g2_fill_2
XFILLER_8_174 VPWR VGND sg13g2_decap_8
X_273_ VPWR VGND _046_ sg13g2_tiehi
X_342_ Inst_N_IO_switch_matrix.S2BEGb4 S2BEGb[4] VPWR VGND sg13g2_buf_1
XFILLER_1_350 VPWR VGND sg13g2_decap_4
XFILLER_11_405 VPWR VGND sg13g2_decap_4
XFILLER_4_70 VPWR VGND sg13g2_fill_1
X_325_ FrameStrobe[19] FrameStrobe_O[19] VPWR VGND sg13g2_buf_1
XFILLER_9_48 VPWR VGND sg13g2_fill_1
X_187_ FrameData[13] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit13.Q VPWR VGND
+ sg13g2_dlhq_1
X_256_ FrameData[18] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_11_257 VPWR VGND sg13g2_decap_8
X_110_ Inst_N_IO_ConfigMem.Inst_frame0_bit20.Q VPWR _026_ VGND _024_ _025_ sg13g2_o21ai_1
XFILLER_3_423 VPWR VGND sg13g2_fill_1
X_308_ FrameStrobe[2] FrameStrobe_O[2] VPWR VGND sg13g2_buf_1
X_239_ FrameData[1] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit1.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_3_297 VPWR VGND sg13g2_fill_2
XFILLER_8_334 VPWR VGND sg13g2_fill_1
XFILLER_0_278 VPWR VGND sg13g2_decap_4
X_272_ VPWR VGND _045_ sg13g2_tiehi
X_341_ Inst_N_IO_switch_matrix.S2BEGb3 S2BEGb[3] VPWR VGND sg13g2_buf_1
XFILLER_1_384 VPWR VGND sg13g2_fill_1
XFILLER_5_101 VPWR VGND sg13g2_fill_2
X_324_ FrameStrobe[18] FrameStrobe_O[18] VPWR VGND sg13g2_buf_1
XFILLER_0_18 VPWR VGND sg13g2_fill_1
X_255_ FrameData[17] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit17.Q VPWR VGND
+ sg13g2_dlhq_1
X_186_ FrameData[12] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit12.Q VPWR VGND
+ sg13g2_dlhq_1
X_169_ FrameData[27] FrameStrobe[3] Inst_N_IO_ConfigMem.Inst_frame3_bit27.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_10_291 VPWR VGND sg13g2_fill_1
X_307_ FrameStrobe[1] FrameStrobe_O[1] VPWR VGND sg13g2_buf_1
X_238_ FrameData[0] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit0.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_6_273 VPWR VGND sg13g2_fill_1
XFILLER_6_28 VPWR VGND sg13g2_fill_2
XFILLER_0_224 VPWR VGND sg13g2_fill_2
XFILLER_0_202 VPWR VGND sg13g2_fill_1
X_271_ _046_ VGND VPWR B_O_top Inst_B_IO_1_bidirectional_frame_config_pass.Q clknet_1_0__leaf_UserCLK_regs
+ sg13g2_dfrbpq_1
X_340_ Inst_N_IO_switch_matrix.S2BEGb2 S2BEGb[2] VPWR VGND sg13g2_buf_1
X_185_ FrameData[11] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit11.Q VPWR VGND
+ sg13g2_dlhq_1
X_323_ FrameStrobe[17] FrameStrobe_O[17] VPWR VGND sg13g2_buf_1
X_254_ FrameData[16] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit16.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_9_282 VPWR VGND sg13g2_fill_2
XFILLER_1_193 VPWR VGND sg13g2_fill_1
X_306_ FrameStrobe[0] FrameStrobe_O[0] VPWR VGND sg13g2_buf_1
X_168_ FrameData[26] FrameStrobe[3] Inst_N_IO_ConfigMem.Inst_frame3_bit26.Q VPWR VGND
+ sg13g2_dlhq_1
X_099_ _016_ _015_ Inst_N_IO_ConfigMem.Inst_frame0_bit28.Q VPWR VGND sg13g2_nand2b_1
X_237_ FrameData[31] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit31.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_6_263 VPWR VGND sg13g2_decap_4
XFILLER_3_299 VPWR VGND sg13g2_fill_1
XFILLER_7_83 VPWR VGND sg13g2_decap_8
XFILLER_8_155 VPWR VGND sg13g2_fill_2
XFILLER_8_100 VPWR VGND sg13g2_decap_4
X_270_ _045_ VGND VPWR A_O_top Inst_A_IO_1_bidirectional_frame_config_pass.Q clknet_1_1__leaf_UserCLK_regs
+ sg13g2_dfrbpq_1
XFILLER_1_375 VPWR VGND sg13g2_fill_2
XFILLER_4_95 VPWR VGND sg13g2_fill_1
X_322_ FrameStrobe[16] FrameStrobe_O[16] VPWR VGND sg13g2_buf_1
XFILLER_2_128 VPWR VGND sg13g2_fill_2
X_184_ FrameData[10] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit10.Q VPWR VGND
+ sg13g2_dlhq_1
X_253_ FrameData[15] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit15.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_11_238 VPWR VGND sg13g2_fill_2
X_305_ FrameData[31] FrameData_O[31] VPWR VGND sg13g2_buf_1
X_167_ FrameData[25] FrameStrobe[3] Inst_N_IO_ConfigMem.Inst_frame3_bit25.Q VPWR VGND
+ sg13g2_dlhq_1
X_098_ _014_ _013_ Inst_N_IO_ConfigMem.Inst_frame0_bit27.Q _015_ VPWR VGND sg13g2_mux2_1
X_236_ FrameData[30] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit30.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_1_96 VPWR VGND sg13g2_fill_2
XFILLER_3_267 VPWR VGND sg13g2_decap_8
XFILLER_3_278 VPWR VGND sg13g2_fill_2
X_219_ FrameData[13] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit13.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_5_307 VPWR VGND sg13g2_decap_8
XFILLER_5_318 VPWR VGND sg13g2_fill_1
XFILLER_4_373 VPWR VGND sg13g2_fill_2
XFILLER_5_159 VPWR VGND sg13g2_fill_2
XFILLER_9_421 VPWR VGND sg13g2_fill_2
X_321_ FrameStrobe[15] FrameStrobe_O[15] VPWR VGND sg13g2_buf_1
X_183_ FrameData[9] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit9.Q VPWR VGND
+ sg13g2_dlhq_1
X_252_ FrameData[14] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit14.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_9_284 VPWR VGND sg13g2_fill_1
X_304_ FrameData[30] FrameData_O[30] VPWR VGND sg13g2_buf_1
XFILLER_10_250 VPWR VGND sg13g2_fill_1
X_235_ FrameData[29] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit29.Q VPWR VGND
+ sg13g2_dlhq_1
X_166_ FrameData[24] FrameStrobe[3] Inst_N_IO_ConfigMem.Inst_frame3_bit24.Q VPWR VGND
+ sg13g2_dlhq_1
X_097_ Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q N2MID[0] N2MID[1] N2MID[2] N2MID[3]
+ Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q _014_ VPWR VGND sg13g2_mux4_1
X_149_ FrameData[7] FrameStrobe[3] A_config_C_bit1 VPWR VGND sg13g2_dlhq_1
X_218_ FrameData[12] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit12.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_0_249 VPWR VGND sg13g2_decap_4
XFILLER_8_316 VPWR VGND sg13g2_fill_1
XFILLER_5_127 VPWR VGND sg13g2_decap_4
XFILLER_9_400 VPWR VGND sg13g2_decap_8
XFILLER_1_377 VPWR VGND sg13g2_fill_1
XFILLER_4_20 VPWR VGND sg13g2_fill_2
XFILLER_4_160 VPWR VGND sg13g2_decap_8
X_182_ FrameData[8] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit8.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_10_421 VPWR VGND sg13g2_fill_2
XFILLER_10_410 VPWR VGND sg13g2_fill_2
X_320_ FrameStrobe[14] FrameStrobe_O[14] VPWR VGND sg13g2_buf_1
XFILLER_8_0 VPWR VGND sg13g2_decap_8
X_251_ FrameData[13] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit13.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_6_403 VPWR VGND sg13g2_decap_4
XFILLER_1_7 VPWR VGND sg13g2_fill_2
X_303_ FrameData[29] FrameData_O[29] VPWR VGND sg13g2_buf_1
X_234_ FrameData[28] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit28.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_1_65 VPWR VGND sg13g2_fill_2
X_096_ Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q N2MID[4] N2MID[5] N2MID[6] N2MID[7]
+ Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q _013_ VPWR VGND sg13g2_mux4_1
X_165_ FrameData[23] FrameStrobe[3] Inst_N_IO_ConfigMem.Inst_frame3_bit23.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_6_299 VPWR VGND sg13g2_fill_2
X_148_ FrameData[6] FrameStrobe[3] A_config_C_bit0 VPWR VGND sg13g2_dlhq_1
X_217_ FrameData[11] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit11.Q VPWR VGND
+ sg13g2_dlhq_1
X_079_ Inst_N_IO_ConfigMem.Inst_frame0_bit29.Q VPWR _042_ VGND N2END[6] Inst_N_IO_ConfigMem.Inst_frame0_bit30.Q
+ sg13g2_o21ai_1
XFILLER_7_350 VPWR VGND sg13g2_decap_8
XFILLER_8_125 VPWR VGND sg13g2_decap_4
XFILLER_9_423 VPWR VGND sg13g2_fill_1
XFILLER_4_43 VPWR VGND sg13g2_fill_2
X_250_ FrameData[12] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit12.Q VPWR VGND
+ sg13g2_dlhq_1
X_181_ FrameData[7] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit7.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_9_275 VPWR VGND sg13g2_decap_8
XFILLER_9_242 VPWR VGND sg13g2_decap_8
XFILLER_11_219 VPWR VGND sg13g2_fill_2
X_302_ FrameData[28] FrameData_O[28] VPWR VGND sg13g2_buf_1
XFILLER_10_296 VPWR VGND sg13g2_fill_1
X_233_ FrameData[27] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit27.Q VPWR VGND
+ sg13g2_dlhq_1
X_164_ FrameData[22] FrameStrobe[3] Inst_N_IO_ConfigMem.Inst_frame3_bit22.Q VPWR VGND
+ sg13g2_dlhq_1
X_095_ Inst_N_IO_ConfigMem.Inst_frame0_bit28.Q VPWR _012_ VGND _008_ _011_ sg13g2_o21ai_1
XFILLER_6_234 VPWR VGND sg13g2_fill_1
XFILLER_6_256 VPWR VGND sg13g2_decap_8
X_078_ Inst_N_IO_ConfigMem.Inst_frame0_bit29.Q N2MID[6] N2MID[7] N2END[0] N2END[4]
+ Inst_N_IO_ConfigMem.Inst_frame0_bit30.Q _041_ VPWR VGND sg13g2_mux4_1
X_147_ Inst_N_IO_ConfigMem.Inst_frame2_bit20.Q N1END[3] N4END[14] NN4END[14] B_O_top
+ Inst_N_IO_ConfigMem.Inst_frame2_bit21.Q Inst_N_IO_switch_matrix.S4BEG1 VPWR VGND
+ sg13g2_mux4_1
X_216_ FrameData[10] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit10.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_11_391 VPWR VGND sg13g2_decap_8
XFILLER_7_65 VPWR VGND sg13g2_fill_1
Xclkbuf_1_0__f_UserCLK_regs clknet_0_UserCLK_regs clknet_1_0__leaf_UserCLK_regs VPWR
+ VGND sg13g2_buf_8
XFILLER_4_22 VPWR VGND sg13g2_fill_1
XFILLER_4_66 VPWR VGND sg13g2_decap_4
XFILLER_4_88 VPWR VGND sg13g2_decap_8
XFILLER_10_423 VPWR VGND sg13g2_fill_1
XFILLER_10_412 VPWR VGND sg13g2_fill_1
XFILLER_10_401 VPWR VGND sg13g2_fill_1
X_180_ FrameData[6] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit6.Q VPWR VGND
+ sg13g2_dlhq_1
X_378_ clknet_1_0__leaf_UserCLK UserCLKo VPWR VGND sg13g2_buf_1
XFILLER_1_165 VPWR VGND sg13g2_fill_2
XFILLER_1_9 VPWR VGND sg13g2_fill_1
X_301_ FrameData[27] FrameData_O[27] VPWR VGND sg13g2_buf_1
X_232_ FrameData[26] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit26.Q VPWR VGND
+ sg13g2_dlhq_1
X_163_ FrameData[21] FrameStrobe[3] Inst_N_IO_ConfigMem.Inst_frame3_bit21.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_6_202 VPWR VGND sg13g2_decap_8
X_094_ Inst_N_IO_ConfigMem.Inst_frame0_bit27.Q VPWR _011_ VGND _009_ _010_ sg13g2_o21ai_1
XFILLER_1_89 VPWR VGND sg13g2_decap_8
XFILLER_1_67 VPWR VGND sg13g2_fill_1
XFILLER_10_21 VPWR VGND sg13g2_fill_2
XFILLER_3_227 VPWR VGND sg13g2_fill_2
X_146_ Inst_N_IO_ConfigMem.Inst_frame2_bit23.Q N4END[11] NN4END[15] NN4END[11] A_O_top
+ Inst_N_IO_ConfigMem.Inst_frame2_bit22.Q Inst_N_IO_switch_matrix.S4BEG2 VPWR VGND
+ sg13g2_mux4_1
X_077_ _040_ N2END[5] Inst_N_IO_ConfigMem.Inst_frame0_bit30.Q VPWR VGND sg13g2_nand2b_1
X_215_ FrameData[9] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit9.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_7_22 VPWR VGND sg13g2_fill_1
X_129_ Inst_N_IO_ConfigMem.Inst_frame1_bit24.Q N4END[7] N4END[9] N4END[11] Inst_B_IO_1_bidirectional_frame_config_pass.Q
+ Inst_N_IO_ConfigMem.Inst_frame1_bit25.Q Inst_N_IO_switch_matrix.SS4BEG3 VPWR VGND
+ sg13g2_mux4_1
XFILLER_4_322 VPWR VGND sg13g2_decap_4
XFILLER_4_130 VPWR VGND sg13g2_fill_2
XFILLER_4_185 VPWR VGND sg13g2_fill_2
X_377_ Inst_N_IO_switch_matrix.SS4BEG15 SS4BEG[15] VPWR VGND sg13g2_buf_1
XFILLER_6_417 VPWR VGND sg13g2_decap_8
X_300_ FrameData[26] FrameData_O[26] VPWR VGND sg13g2_buf_1
X_231_ FrameData[25] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit25.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_10_243 VPWR VGND sg13g2_decap_8
X_162_ FrameData[20] FrameStrobe[3] Inst_N_IO_ConfigMem.Inst_frame3_bit20.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_6_0 VPWR VGND sg13g2_decap_4
X_093_ Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q VPWR _010_ VGND Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q
+ N2END[6] sg13g2_o21ai_1
X_076_ _039_ VPWR A_T_top VGND Inst_N_IO_ConfigMem.Inst_frame0_bit22.Q _035_ sg13g2_o21ai_1
XFILLER_2_250 VPWR VGND sg13g2_fill_1
X_214_ FrameData[8] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit8.Q VPWR VGND
+ sg13g2_dlhq_1
X_145_ Inst_N_IO_ConfigMem.Inst_frame2_bit25.Q N4END[10] NN4END[14] NN4END[10] B_O_top
+ Inst_N_IO_ConfigMem.Inst_frame2_bit24.Q Inst_N_IO_switch_matrix.S4BEG3 VPWR VGND
+ sg13g2_mux4_1
Xclkbuf_1_0__f_UserCLK clknet_0_UserCLK clknet_1_0__leaf_UserCLK VPWR VGND sg13g2_buf_8
XFILLER_8_309 VPWR VGND sg13g2_decap_8
X_059_ Inst_N_IO_ConfigMem.Inst_frame3_bit26.Q N2MID[3] N4END[3] NN4END[3] NN4END[11]
+ Inst_N_IO_ConfigMem.Inst_frame3_bit27.Q Inst_N_IO_switch_matrix.S2BEG4 VPWR VGND
+ sg13g2_mux4_1
X_128_ Inst_N_IO_ConfigMem.Inst_frame1_bit26.Q N2END[0] N2END[2] N2END[4] N2END[6]
+ Inst_N_IO_ConfigMem.Inst_frame1_bit27.Q Inst_N_IO_switch_matrix.SS4BEG4 VPWR VGND
+ sg13g2_mux4_1
XFILLER_7_364 VPWR VGND sg13g2_fill_2
XFILLER_7_172 VPWR VGND sg13g2_fill_1
XFILLER_4_153 VPWR VGND sg13g2_decap_8
XFILLER_1_189 VPWR VGND sg13g2_decap_4
XFILLER_1_167 VPWR VGND sg13g2_fill_1
XFILLER_6_407 VPWR VGND sg13g2_fill_2
X_376_ Inst_N_IO_switch_matrix.SS4BEG14 SS4BEG[14] VPWR VGND sg13g2_buf_1
X_230_ FrameData[24] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit24.Q VPWR VGND
+ sg13g2_dlhq_1
X_161_ FrameData[19] FrameStrobe[3] Inst_N_IO_ConfigMem.Inst_frame3_bit19.Q VPWR VGND
+ sg13g2_dlhq_1
X_359_ Inst_N_IO_switch_matrix.S4BEG13 S4BEG[13] VPWR VGND sg13g2_buf_1
XFILLER_2_410 VPWR VGND sg13g2_fill_2
XFILLER_2_421 VPWR VGND sg13g2_fill_2
X_092_ N2END[7] Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q _009_ VPWR VGND sg13g2_nor2b_1
XFILLER_10_34 VPWR VGND sg13g2_fill_2
XFILLER_10_23 VPWR VGND sg13g2_fill_1
X_075_ _036_ _037_ Inst_N_IO_ConfigMem.Inst_frame0_bit22.Q _039_ VPWR VGND _038_ sg13g2_nand4_1
X_213_ FrameData[7] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit7.Q VPWR VGND
+ sg13g2_dlhq_1
X_144_ Inst_N_IO_ConfigMem.Inst_frame2_bit27.Q N1END[2] NN4END[7] N4END[7] A_O_top
+ Inst_N_IO_ConfigMem.Inst_frame2_bit26.Q Inst_N_IO_switch_matrix.S4BEG4 VPWR VGND
+ sg13g2_mux4_1
X_127_ Inst_N_IO_ConfigMem.Inst_frame1_bit28.Q N2END[1] N2END[3] N2END[5] N2END[7]
+ Inst_N_IO_ConfigMem.Inst_frame1_bit29.Q Inst_N_IO_switch_matrix.SS4BEG5 VPWR VGND
+ sg13g2_mux4_1
XFILLER_7_343 VPWR VGND sg13g2_decap_8
X_058_ Inst_N_IO_ConfigMem.Inst_frame3_bit28.Q N2MID[2] N4END[2] NN4END[2] NN4END[10]
+ Inst_N_IO_ConfigMem.Inst_frame3_bit29.Q Inst_N_IO_switch_matrix.S2BEG5 VPWR VGND
+ sg13g2_mux4_1
XFILLER_8_129 VPWR VGND sg13g2_fill_1
XFILLER_4_187 VPWR VGND sg13g2_fill_1
XFILLER_9_224 VPWR VGND sg13g2_fill_1
X_375_ Inst_N_IO_switch_matrix.SS4BEG13 SS4BEG[13] VPWR VGND sg13g2_buf_1
Xclkbuf_regs_0_UserCLK UserCLK UserCLK_regs VPWR VGND sg13g2_buf_8
XFILLER_10_289 VPWR VGND sg13g2_fill_2
X_358_ Inst_N_IO_switch_matrix.S4BEG12 S4BEG[12] VPWR VGND sg13g2_buf_1
X_160_ FrameData[18] FrameStrobe[3] Inst_N_IO_ConfigMem.Inst_frame3_bit18.Q VPWR VGND
+ sg13g2_dlhq_1
X_091_ VGND VPWR _006_ _007_ _008_ Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q sg13g2_a21oi_1
XFILLER_6_216 VPWR VGND sg13g2_fill_1
X_289_ FrameData[15] FrameData_O[15] VPWR VGND sg13g2_buf_1
X_212_ FrameData[6] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit6.Q VPWR VGND
+ sg13g2_dlhq_1
X_143_ Inst_N_IO_ConfigMem.Inst_frame2_bit29.Q N1END[3] NN4END[6] N4END[6] B_O_top
+ Inst_N_IO_ConfigMem.Inst_frame2_bit28.Q Inst_N_IO_switch_matrix.S4BEG5 VPWR VGND
+ sg13g2_mux4_1
X_074_ _038_ N2END[4] Inst_N_IO_ConfigMem.Inst_frame0_bit24.Q VPWR VGND sg13g2_nand2_1
XFILLER_11_384 VPWR VGND sg13g2_decap_8
X_057_ Inst_N_IO_ConfigMem.Inst_frame3_bit30.Q N2MID[1] N4END[1] NN4END[1] NN4END[9]
+ Inst_N_IO_ConfigMem.Inst_frame3_bit31.Q Inst_N_IO_switch_matrix.S2BEG6 VPWR VGND
+ sg13g2_mux4_1
X_126_ Inst_N_IO_ConfigMem.Inst_frame1_bit31.Q N2MID[0] N2MID[4] N2MID[2] N2MID[6]
+ Inst_N_IO_ConfigMem.Inst_frame1_bit30.Q Inst_N_IO_switch_matrix.SS4BEG6 VPWR VGND
+ sg13g2_mux4_1
XFILLER_11_170 VPWR VGND sg13g2_fill_2
X_109_ Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q VPWR _025_ VGND N2END[6] Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q
+ sg13g2_o21ai_1
XFILLER_9_214 VPWR VGND sg13g2_decap_4
X_374_ Inst_N_IO_switch_matrix.SS4BEG12 SS4BEG[12] VPWR VGND sg13g2_buf_1
Xclkbuf_0_UserCLK_regs UserCLK_regs clknet_0_UserCLK_regs VPWR VGND sg13g2_buf_8
X_090_ _007_ N2END[4] Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q VPWR VGND sg13g2_nand2b_1
XFILLER_2_412 VPWR VGND sg13g2_fill_1
XFILLER_2_423 VPWR VGND sg13g2_fill_1
X_357_ Inst_N_IO_switch_matrix.S4BEG11 S4BEG[11] VPWR VGND sg13g2_buf_1
X_288_ FrameData[14] FrameData_O[14] VPWR VGND sg13g2_buf_1
X_142_ Inst_N_IO_ConfigMem.Inst_frame2_bit30.Q N4END[3] NN4END[3] NN4END[15] A_O_top
+ Inst_N_IO_ConfigMem.Inst_frame2_bit31.Q Inst_N_IO_switch_matrix.S4BEG6 VPWR VGND
+ sg13g2_mux4_1
XFILLER_10_36 VPWR VGND sg13g2_fill_1
X_211_ FrameData[5] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit5.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_3_209 VPWR VGND sg13g2_fill_1
X_073_ Inst_N_IO_ConfigMem.Inst_frame0_bit23.Q VPWR _037_ VGND N2END[2] Inst_N_IO_ConfigMem.Inst_frame0_bit24.Q
+ sg13g2_o21ai_1
XFILLER_2_220 VPWR VGND sg13g2_decap_4
XFILLER_4_0 VPWR VGND sg13g2_fill_2
X_056_ Inst_N_IO_ConfigMem.Inst_frame2_bit0.Q N2MID[0] N4END[0] NN4END[0] NN4END[8]
+ Inst_N_IO_ConfigMem.Inst_frame2_bit1.Q Inst_N_IO_switch_matrix.S2BEG7 VPWR VGND
+ sg13g2_mux4_1
X_125_ Inst_N_IO_ConfigMem.Inst_frame0_bit1.Q N2MID[1] N2MID[5] N2MID[3] N2MID[7]
+ Inst_N_IO_ConfigMem.Inst_frame0_bit0.Q Inst_N_IO_switch_matrix.SS4BEG7 VPWR VGND
+ sg13g2_mux4_1
XFILLER_4_315 VPWR VGND sg13g2_decap_8
XFILLER_4_326 VPWR VGND sg13g2_fill_1
X_108_ N2END[7] Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q _024_ VPWR VGND sg13g2_nor2b_1
XFILLER_9_407 VPWR VGND sg13g2_fill_2
XFILLER_4_167 VPWR VGND sg13g2_fill_1
XFILLER_8_7 VPWR VGND sg13g2_decap_8
X_373_ Inst_N_IO_switch_matrix.SS4BEG11 SS4BEG[11] VPWR VGND sg13g2_buf_1
XFILLER_5_421 VPWR VGND sg13g2_fill_2
XFILLER_10_236 VPWR VGND sg13g2_decap_8
X_287_ FrameData[13] FrameData_O[13] VPWR VGND sg13g2_buf_1
X_356_ Inst_N_IO_switch_matrix.S4BEG10 S4BEG[10] VPWR VGND sg13g2_buf_1
X_072_ _001_ N2END[0] _036_ VPWR VGND Inst_N_IO_ConfigMem.Inst_frame0_bit23.Q sg13g2_nand3b_1
X_210_ FrameData[4] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit4.Q VPWR VGND
+ sg13g2_dlhq_1
X_141_ Inst_N_IO_ConfigMem.Inst_frame1_bit0.Q N4END[2] NN4END[2] NN4END[14] B_O_top
+ Inst_N_IO_ConfigMem.Inst_frame1_bit1.Q Inst_N_IO_switch_matrix.S4BEG7 VPWR VGND
+ sg13g2_mux4_1
X_339_ Inst_N_IO_switch_matrix.S2BEGb1 S2BEGb[1] VPWR VGND sg13g2_buf_1
XFILLER_7_357 VPWR VGND sg13g2_decap_8
X_124_ Inst_N_IO_ConfigMem.Inst_frame0_bit3.Q N4END[4] N4END[8] N4END[6] N4END[10]
+ Inst_N_IO_ConfigMem.Inst_frame0_bit2.Q Inst_N_IO_switch_matrix.SS4BEG8 VPWR VGND
+ sg13g2_mux4_1
X_055_ Inst_N_IO_ConfigMem.Inst_frame2_bit2.Q N2END[7] N4END[7] NN4END[7] NN4END[15]
+ Inst_N_IO_ConfigMem.Inst_frame2_bit3.Q Inst_N_IO_switch_matrix.S2BEGb0 VPWR VGND
+ sg13g2_mux4_1
XFILLER_11_194 VPWR VGND sg13g2_decap_8
XFILLER_11_172 VPWR VGND sg13g2_fill_1
XFILLER_7_165 VPWR VGND sg13g2_decap_8
XFILLER_7_132 VPWR VGND sg13g2_decap_8
X_107_ VGND VPWR _021_ _022_ _023_ Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q sg13g2_a21oi_1
XFILLER_9_249 VPWR VGND sg13g2_fill_1
X_372_ Inst_N_IO_switch_matrix.SS4BEG10 SS4BEG[10] VPWR VGND sg13g2_buf_1
X_355_ Inst_N_IO_switch_matrix.S4BEG9 S4BEG[9] VPWR VGND sg13g2_buf_1
X_286_ FrameData[12] FrameData_O[12] VPWR VGND sg13g2_buf_1
X_071_ _034_ VPWR _035_ VGND Inst_N_IO_ConfigMem.Inst_frame0_bit23.Q _033_ sg13g2_o21ai_1
X_140_ Inst_N_IO_ConfigMem.Inst_frame1_bit2.Q N1END[1] N4END[13] NN4END[13] Inst_A_IO_1_bidirectional_frame_config_pass.Q
+ Inst_N_IO_ConfigMem.Inst_frame1_bit3.Q Inst_N_IO_switch_matrix.S4BEG8 VPWR VGND
+ sg13g2_mux4_1
XFILLER_4_2 VPWR VGND sg13g2_fill_1
Xclkbuf_1_1__f_UserCLK_regs clknet_0_UserCLK_regs clknet_1_1__leaf_UserCLK_regs VPWR
+ VGND sg13g2_buf_8
X_269_ FrameData[31] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit31.Q VPWR VGND
+ sg13g2_dlhq_1
X_338_ Inst_N_IO_switch_matrix.S2BEGb0 S2BEGb[0] VPWR VGND sg13g2_buf_1
XFILLER_11_398 VPWR VGND sg13g2_decap_8
XFILLER_11_92 VPWR VGND sg13g2_fill_2
XFILLER_7_303 VPWR VGND sg13g2_fill_2
X_123_ Inst_N_IO_ConfigMem.Inst_frame0_bit4.Q N4END[1] N4END[3] N4END[5] N4END[7]
+ Inst_N_IO_ConfigMem.Inst_frame0_bit5.Q Inst_N_IO_switch_matrix.SS4BEG9 VPWR VGND
+ sg13g2_mux4_1
X_054_ Inst_N_IO_ConfigMem.Inst_frame2_bit4.Q N2END[6] N4END[6] NN4END[6] NN4END[14]
+ Inst_N_IO_ConfigMem.Inst_frame2_bit5.Q Inst_N_IO_switch_matrix.S2BEGb1 VPWR VGND
+ sg13g2_mux4_1
X_106_ _022_ N2END[4] Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q VPWR VGND sg13g2_nand2b_1
XFILLER_8_93 VPWR VGND sg13g2_decap_8
XFILLER_3_191 VPWR VGND sg13g2_fill_1
X_371_ Inst_N_IO_switch_matrix.SS4BEG9 SS4BEG[9] VPWR VGND sg13g2_buf_1
XFILLER_5_423 VPWR VGND sg13g2_fill_1
XFILLER_5_72 VPWR VGND sg13g2_fill_2
XFILLER_6_209 VPWR VGND sg13g2_decap_8
X_354_ Inst_N_IO_switch_matrix.S4BEG8 S4BEG[8] VPWR VGND sg13g2_buf_1
X_285_ FrameData[11] FrameData_O[11] VPWR VGND sg13g2_buf_1
XFILLER_5_286 VPWR VGND sg13g2_decap_4
X_070_ Inst_N_IO_ConfigMem.Inst_frame0_bit23.Q _001_ N2END[1] _034_ VPWR VGND sg13g2_nand3_1
X_199_ FrameData[25] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit25.Q VPWR VGND
+ sg13g2_dlhq_1
X_337_ Inst_N_IO_switch_matrix.S2BEG7 S2BEG[7] VPWR VGND sg13g2_buf_1
X_268_ FrameData[30] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit30.Q VPWR VGND
+ sg13g2_dlhq_1
X_053_ Inst_N_IO_ConfigMem.Inst_frame2_bit6.Q N2END[5] N4END[5] NN4END[5] NN4END[13]
+ Inst_N_IO_ConfigMem.Inst_frame2_bit7.Q Inst_N_IO_switch_matrix.S2BEGb2 VPWR VGND
+ sg13g2_mux4_1
XFILLER_2_0 VPWR VGND sg13g2_fill_2
X_122_ Inst_N_IO_ConfigMem.Inst_frame0_bit6.Q N4END[0] N4END[2] N4END[4] A_O_top Inst_N_IO_ConfigMem.Inst_frame0_bit7.Q
+ Inst_N_IO_switch_matrix.SS4BEG10 VPWR VGND sg13g2_mux4_1
XFILLER_11_163 VPWR VGND sg13g2_decap_8
X_105_ _021_ N2END[5] Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q VPWR VGND sg13g2_nand2_1
XFILLER_9_218 VPWR VGND sg13g2_fill_2
XFILLER_0_140 VPWR VGND sg13g2_decap_4
X_370_ Inst_N_IO_switch_matrix.SS4BEG8 SS4BEG[8] VPWR VGND sg13g2_buf_1
X_353_ Inst_N_IO_switch_matrix.S4BEG7 S4BEG[7] VPWR VGND sg13g2_buf_1
X_284_ FrameData[10] FrameData_O[10] VPWR VGND sg13g2_buf_1
X_198_ FrameData[24] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit24.Q VPWR VGND
+ sg13g2_dlhq_1
X_267_ FrameData[29] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit29.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_2_224 VPWR VGND sg13g2_fill_2
X_336_ Inst_N_IO_switch_matrix.S2BEG6 S2BEG[6] VPWR VGND sg13g2_buf_1
X_052_ Inst_N_IO_ConfigMem.Inst_frame2_bit8.Q N2END[4] N4END[4] NN4END[4] NN4END[12]
+ Inst_N_IO_ConfigMem.Inst_frame2_bit9.Q Inst_N_IO_switch_matrix.S2BEGb3 VPWR VGND
+ sg13g2_mux4_1
X_121_ Inst_N_IO_ConfigMem.Inst_frame0_bit8.Q N4END[6] N4END[8] N4END[10] B_O_top
+ Inst_N_IO_ConfigMem.Inst_frame0_bit9.Q Inst_N_IO_switch_matrix.SS4BEG11 VPWR VGND
+ sg13g2_mux4_1
X_319_ FrameStrobe[13] FrameStrobe_O[13] VPWR VGND sg13g2_buf_1
XFILLER_6_382 VPWR VGND sg13g2_decap_8
XFILLER_11_142 VPWR VGND sg13g2_decap_4
X_104_ VPWR VGND _019_ Inst_N_IO_ConfigMem.Inst_frame0_bit20.Q _018_ Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q
+ _020_ _017_ sg13g2_a221oi_1
XFILLER_0_163 VPWR VGND sg13g2_decap_4
XFILLER_10_0 VPWR VGND sg13g2_decap_4
XFILLER_8_285 VPWR VGND sg13g2_fill_2
X_352_ Inst_N_IO_switch_matrix.S4BEG6 S4BEG[6] VPWR VGND sg13g2_buf_1
X_283_ FrameData[9] FrameData_O[9] VPWR VGND sg13g2_buf_1
XFILLER_5_211 VPWR VGND sg13g2_fill_2
XFILLER_5_255 VPWR VGND sg13g2_decap_8
X_266_ FrameData[28] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit28.Q VPWR VGND
+ sg13g2_dlhq_1
X_197_ FrameData[23] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit23.Q VPWR VGND
+ sg13g2_dlhq_1
X_335_ Inst_N_IO_switch_matrix.S2BEG5 S2BEG[5] VPWR VGND sg13g2_buf_1
XFILLER_2_20 VPWR VGND sg13g2_fill_1
XFILLER_11_51 VPWR VGND sg13g2_decap_8
X_051_ Inst_N_IO_ConfigMem.Inst_frame2_bit10.Q N2END[3] N4END[3] NN4END[3] NN4END[11]
+ Inst_N_IO_ConfigMem.Inst_frame2_bit11.Q Inst_N_IO_switch_matrix.S2BEGb4 VPWR VGND
+ sg13g2_mux4_1
XFILLER_2_2 VPWR VGND sg13g2_fill_1
X_120_ Inst_N_IO_ConfigMem.Inst_frame0_bit10.Q N4END[1] N4END[3] N4END[5] Inst_A_IO_1_bidirectional_frame_config_pass.Q
+ Inst_N_IO_ConfigMem.Inst_frame0_bit11.Q Inst_N_IO_switch_matrix.SS4BEG12 VPWR VGND
+ sg13g2_mux4_1
X_318_ FrameStrobe[12] FrameStrobe_O[12] VPWR VGND sg13g2_buf_1
X_249_ FrameData[11] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit11.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_7_158 VPWR VGND sg13g2_decap_8
XFILLER_7_114 VPWR VGND sg13g2_fill_1
X_103_ VGND VPWR _000_ Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q _019_ Inst_N_IO_ConfigMem.Inst_frame0_bit19.Q
+ sg13g2_a21oi_1
X_282_ FrameData[8] FrameData_O[8] VPWR VGND sg13g2_buf_1
X_351_ Inst_N_IO_switch_matrix.S4BEG5 S4BEG[5] VPWR VGND sg13g2_buf_1
X_334_ Inst_N_IO_switch_matrix.S2BEG4 S2BEG[4] VPWR VGND sg13g2_buf_1
XFILLER_2_215 VPWR VGND sg13g2_fill_1
XFILLER_2_248 VPWR VGND sg13g2_fill_2
X_265_ FrameData[27] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit27.Q VPWR VGND
+ sg13g2_dlhq_1
X_196_ FrameData[22] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit22.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_2_43 VPWR VGND sg13g2_decap_4
X_050_ Inst_N_IO_ConfigMem.Inst_frame2_bit12.Q N2END[2] N4END[2] NN4END[2] NN4END[10]
+ Inst_N_IO_ConfigMem.Inst_frame2_bit13.Q Inst_N_IO_switch_matrix.S2BEGb5 VPWR VGND
+ sg13g2_mux4_1
XFILLER_11_85 VPWR VGND sg13g2_decap_8
X_317_ FrameStrobe[11] FrameStrobe_O[11] VPWR VGND sg13g2_buf_1
X_179_ FrameData[5] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit5.Q VPWR VGND
+ sg13g2_dlhq_1
X_248_ FrameData[10] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit10.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_0_0 VPWR VGND sg13g2_fill_1
X_102_ VGND VPWR _018_ Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q N2END[0] sg13g2_or2_1
XFILLER_8_31 VPWR VGND sg13g2_fill_1
XFILLER_6_192 VPWR VGND sg13g2_decap_4
XFILLER_3_184 VPWR VGND sg13g2_decap_8
XFILLER_8_287 VPWR VGND sg13g2_fill_1
XFILLER_5_21 VPWR VGND sg13g2_decap_4
XFILLER_5_65 VPWR VGND sg13g2_decap_8
X_281_ FrameData[7] FrameData_O[7] VPWR VGND sg13g2_buf_1
X_350_ Inst_N_IO_switch_matrix.S4BEG4 S4BEG[4] VPWR VGND sg13g2_buf_1
XFILLER_5_279 VPWR VGND sg13g2_decap_8
X_333_ Inst_N_IO_switch_matrix.S2BEG3 S2BEG[3] VPWR VGND sg13g2_buf_1
X_195_ FrameData[21] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit21.Q VPWR VGND
+ sg13g2_dlhq_1
X_264_ FrameData[26] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_9_393 VPWR VGND sg13g2_decap_8
XFILLER_11_20 VPWR VGND sg13g2_fill_2
X_316_ FrameStrobe[10] FrameStrobe_O[10] VPWR VGND sg13g2_buf_1
X_247_ FrameData[9] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit9.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_9_190 VPWR VGND sg13g2_fill_2
X_178_ FrameData[4] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit4.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_6_396 VPWR VGND sg13g2_decap_8
X_101_ N2END[2] N2END[3] Inst_N_IO_ConfigMem.Inst_frame0_bit18.Q _017_ VPWR VGND sg13g2_mux2_1
XFILLER_8_403 VPWR VGND sg13g2_decap_4
XFILLER_3_130 VPWR VGND sg13g2_decap_4
XFILLER_3_152 VPWR VGND sg13g2_decap_4
XFILLER_0_144 VPWR VGND sg13g2_fill_2
XFILLER_0_133 VPWR VGND sg13g2_decap_8
XFILLER_5_406 VPWR VGND sg13g2_fill_2
XFILLER_8_233 VPWR VGND sg13g2_decap_4
X_280_ FrameData[6] FrameData_O[6] VPWR VGND sg13g2_buf_1
X_194_ FrameData[20] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit20.Q VPWR VGND
+ sg13g2_dlhq_1
X_332_ Inst_N_IO_switch_matrix.S2BEG2 S2BEG[2] VPWR VGND sg13g2_buf_1
X_263_ FrameData[25] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_11_65 VPWR VGND sg13g2_fill_2
X_315_ FrameStrobe[9] FrameStrobe_O[9] VPWR VGND sg13g2_buf_1
X_177_ FrameData[3] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit3.Q VPWR VGND
+ sg13g2_dlhq_1
X_246_ FrameData[8] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit8.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_6_353 VPWR VGND sg13g2_fill_1
XFILLER_6_375 VPWR VGND sg13g2_decap_8
XFILLER_11_135 VPWR VGND sg13g2_decap_8
X_100_ _016_ VPWR B_I_top VGND _005_ _012_ sg13g2_o21ai_1
XFILLER_7_139 VPWR VGND sg13g2_fill_2
X_229_ FrameData[23] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit23.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_3_345 VPWR VGND sg13g2_fill_1
XFILLER_0_167 VPWR VGND sg13g2_fill_1
XFILLER_8_278 VPWR VGND sg13g2_decap_8
XFILLER_8_256 VPWR VGND sg13g2_fill_1
XFILLER_8_212 VPWR VGND sg13g2_decap_8
X_262_ FrameData[24] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit24.Q VPWR VGND
+ sg13g2_dlhq_1
X_331_ Inst_N_IO_switch_matrix.S2BEG1 S2BEG[1] VPWR VGND sg13g2_buf_1
X_193_ FrameData[19] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit19.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_9_340 VPWR VGND sg13g2_fill_2
XFILLER_11_44 VPWR VGND sg13g2_decap_8
X_314_ FrameStrobe[8] FrameStrobe_O[8] VPWR VGND sg13g2_buf_1
X_176_ FrameData[2] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit2.Q VPWR VGND
+ sg13g2_dlhq_1
X_245_ FrameData[7] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit7.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_9_192 VPWR VGND sg13g2_fill_1
XFILLER_7_107 VPWR VGND sg13g2_decap_8
X_228_ FrameData[22] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit22.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_10_191 VPWR VGND sg13g2_fill_2
X_159_ FrameData[17] FrameStrobe[3] Inst_N_IO_switch_matrix.DEBUG_select_S1BEG3[0]
+ VPWR VGND sg13g2_dlhq_1
XFILLER_5_408 VPWR VGND sg13g2_fill_1
X_261_ FrameData[23] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit23.Q VPWR VGND
+ sg13g2_dlhq_1
X_330_ Inst_N_IO_switch_matrix.S2BEG0 S2BEG[0] VPWR VGND sg13g2_buf_1
X_192_ FrameData[18] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit18.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_9_0 VPWR VGND sg13g2_fill_2
XFILLER_2_36 VPWR VGND sg13g2_fill_2
XFILLER_2_47 VPWR VGND sg13g2_fill_2
XFILLER_11_67 VPWR VGND sg13g2_fill_1
X_313_ FrameStrobe[7] FrameStrobe_O[7] VPWR VGND sg13g2_buf_1
X_244_ FrameData[6] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit6.Q VPWR VGND
+ sg13g2_dlhq_1
X_175_ FrameData[1] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit1.Q VPWR VGND
+ sg13g2_dlhq_1
X_158_ FrameData[16] FrameStrobe[3] Inst_N_IO_switch_matrix.DEBUG_select_S1BEG2[0]
+ VPWR VGND sg13g2_dlhq_1
X_227_ FrameData[21] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit21.Q VPWR VGND
+ sg13g2_dlhq_1
X_089_ _006_ Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q N2END[5] VPWR VGND sg13g2_nand2_1
XFILLER_6_196 VPWR VGND sg13g2_fill_2
XFILLER_8_417 VPWR VGND sg13g2_decap_8
XFILLER_3_177 VPWR VGND sg13g2_decap_8
XFILLER_0_80 VPWR VGND sg13g2_fill_2
XFILLER_7_280 VPWR VGND sg13g2_fill_2
XFILLER_1_423 VPWR VGND sg13g2_fill_1
X_260_ FrameData[22] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit22.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_2_209 VPWR VGND sg13g2_fill_2
XFILLER_9_386 VPWR VGND sg13g2_decap_8
XFILLER_9_331 VPWR VGND sg13g2_fill_1
XFILLER_1_242 VPWR VGND sg13g2_fill_2
X_191_ FrameData[17] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit17.Q VPWR VGND
+ sg13g2_dlhq_1
X_312_ FrameStrobe[6] FrameStrobe_O[6] VPWR VGND sg13g2_buf_1
X_243_ FrameData[5] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit5.Q VPWR VGND
+ sg13g2_dlhq_1
X_174_ FrameData[0] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit0.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_6_389 VPWR VGND sg13g2_decap_8
XFILLER_9_172 VPWR VGND sg13g2_fill_1
XFILLER_10_193 VPWR VGND sg13g2_fill_1
XFILLER_8_14 VPWR VGND sg13g2_decap_4
X_157_ FrameData[15] FrameStrobe[3] Inst_N_IO_switch_matrix.DEBUG_select_S1BEG1[0]
+ VPWR VGND sg13g2_dlhq_1
X_226_ FrameData[20] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit20.Q VPWR VGND
+ sg13g2_dlhq_1
X_088_ VPWR VGND _004_ Inst_N_IO_ConfigMem.Inst_frame0_bit27.Q _003_ Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q
+ _005_ _002_ sg13g2_a221oi_1
XFILLER_8_407 VPWR VGND sg13g2_fill_2
XFILLER_3_123 VPWR VGND sg13g2_decap_8
XFILLER_3_134 VPWR VGND sg13g2_fill_1
X_209_ FrameData[3] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit3.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_8_237 VPWR VGND sg13g2_fill_2
XFILLER_8_226 VPWR VGND sg13g2_fill_2
XFILLER_4_421 VPWR VGND sg13g2_fill_2
X_190_ FrameData[16] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit16.Q VPWR VGND
+ sg13g2_dlhq_1
X_311_ FrameStrobe[5] FrameStrobe_O[5] VPWR VGND sg13g2_buf_1
XFILLER_11_58 VPWR VGND sg13g2_decap_8
X_242_ FrameData[4] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit4.Q VPWR VGND
+ sg13g2_dlhq_1
X_173_ FrameData[31] FrameStrobe[3] Inst_N_IO_ConfigMem.Inst_frame3_bit31.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_10_397 VPWR VGND sg13g2_decap_4
XFILLER_6_346 VPWR VGND sg13g2_decap_8
XFILLER_11_128 VPWR VGND sg13g2_decap_8
XFILLER_3_338 VPWR VGND sg13g2_decap_8
X_225_ FrameData[19] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit19.Q VPWR VGND
+ sg13g2_dlhq_1
X_156_ FrameData[14] FrameStrobe[3] Inst_N_IO_switch_matrix.DEBUG_select_S1BEG0[0]
+ VPWR VGND sg13g2_dlhq_1
X_087_ VGND VPWR Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q _000_ _004_ Inst_N_IO_ConfigMem.Inst_frame0_bit26.Q
+ sg13g2_a21oi_1
X_139_ Inst_N_IO_ConfigMem.Inst_frame1_bit4.Q N1END[0] N4END[12] NN4END[12] Inst_B_IO_1_bidirectional_frame_config_pass.Q
+ Inst_N_IO_ConfigMem.Inst_frame1_bit5.Q Inst_N_IO_switch_matrix.S4BEG9 VPWR VGND
+ sg13g2_mux4_1
X_208_ FrameData[2] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit2.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_5_38 VPWR VGND sg13g2_fill_2
XFILLER_11_37 VPWR VGND sg13g2_decap_8
X_310_ FrameStrobe[4] FrameStrobe_O[4] VPWR VGND sg13g2_buf_1
X_241_ FrameData[3] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit3.Q VPWR VGND
+ sg13g2_dlhq_1
X_172_ FrameData[30] FrameStrobe[3] Inst_N_IO_ConfigMem.Inst_frame3_bit30.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_7_0 VPWR VGND sg13g2_decap_4
X_155_ FrameData[13] FrameStrobe[3] B_config_C_bit3 VPWR VGND sg13g2_dlhq_1
XFILLER_10_151 VPWR VGND sg13g2_fill_2
X_086_ VGND VPWR _003_ N2END[0] Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q sg13g2_or2_1
X_224_ FrameData[18] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit18.Q VPWR VGND
+ sg13g2_dlhq_1
X_069_ _032_ VPWR _033_ VGND N2MID[7] Inst_N_IO_ConfigMem.Inst_frame0_bit24.Q sg13g2_o21ai_1
X_207_ FrameData[1] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit1.Q VPWR VGND
+ sg13g2_dlhq_1
X_138_ Inst_N_IO_ConfigMem.Inst_frame1_bit7.Q N4END[9] NN4END[13] NN4END[9] Inst_A_IO_1_bidirectional_frame_config_pass.Q
+ Inst_N_IO_ConfigMem.Inst_frame1_bit6.Q Inst_N_IO_switch_matrix.S4BEG10 VPWR VGND
+ sg13g2_mux4_1
XFILLER_8_228 VPWR VGND sg13g2_fill_1
XFILLER_4_423 VPWR VGND sg13g2_fill_1
XFILLER_4_231 VPWR VGND sg13g2_fill_1
XFILLER_4_264 VPWR VGND sg13g2_decap_4
X_240_ FrameData[2] FrameStrobe[0] Inst_N_IO_ConfigMem.Inst_frame0_bit2.Q VPWR VGND
+ sg13g2_dlhq_1
X_171_ FrameData[29] FrameStrobe[3] Inst_N_IO_ConfigMem.Inst_frame3_bit29.Q VPWR VGND
+ sg13g2_dlhq_1
X_369_ Inst_N_IO_switch_matrix.SS4BEG7 SS4BEG[7] VPWR VGND sg13g2_buf_1
X_223_ FrameData[17] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit17.Q VPWR VGND
+ sg13g2_dlhq_1
X_154_ FrameData[12] FrameStrobe[3] B_config_C_bit2 VPWR VGND sg13g2_dlhq_1
XFILLER_6_112 VPWR VGND sg13g2_decap_8
XFILLER_6_123 VPWR VGND sg13g2_fill_1
X_085_ N2END[2] N2END[3] Inst_N_IO_ConfigMem.Inst_frame0_bit25.Q _002_ VPWR VGND sg13g2_mux2_1
X_068_ _032_ Inst_N_IO_ConfigMem.Inst_frame0_bit24.Q N2END[3] VPWR VGND sg13g2_nand2b_1
X_206_ FrameData[0] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit0.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_2_170 VPWR VGND sg13g2_decap_4
X_137_ Inst_N_IO_ConfigMem.Inst_frame1_bit9.Q N4END[8] NN4END[12] NN4END[8] Inst_B_IO_1_bidirectional_frame_config_pass.Q
+ Inst_N_IO_ConfigMem.Inst_frame1_bit8.Q Inst_N_IO_switch_matrix.S4BEG11 VPWR VGND
+ sg13g2_mux4_1
XFILLER_0_62 VPWR VGND sg13g2_decap_8
XFILLER_0_40 VPWR VGND sg13g2_fill_1
XFILLER_7_240 VPWR VGND sg13g2_fill_1
XFILLER_4_298 VPWR VGND sg13g2_decap_8
XFILLER_0_290 VPWR VGND sg13g2_fill_1
XFILLER_10_334 VPWR VGND sg13g2_fill_2
X_170_ FrameData[28] FrameStrobe[3] Inst_N_IO_ConfigMem.Inst_frame3_bit28.Q VPWR VGND
+ sg13g2_dlhq_1
X_299_ FrameData[25] FrameData_O[25] VPWR VGND sg13g2_buf_1
XFILLER_3_95 VPWR VGND sg13g2_decap_8
X_368_ Inst_N_IO_switch_matrix.SS4BEG6 SS4BEG[6] VPWR VGND sg13g2_buf_1
XFILLER_5_360 VPWR VGND sg13g2_fill_1
X_153_ FrameData[11] FrameStrobe[3] B_config_C_bit1 VPWR VGND sg13g2_dlhq_1
X_084_ VPWR _001_ Inst_N_IO_ConfigMem.Inst_frame0_bit24.Q VGND sg13g2_inv_1
XFILLER_8_29 VPWR VGND sg13g2_fill_2
X_222_ FrameData[16] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit16.Q VPWR VGND
+ sg13g2_dlhq_1
X_205_ FrameData[31] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit31.Q VPWR VGND
+ sg13g2_dlhq_1
X_136_ Inst_N_IO_ConfigMem.Inst_frame1_bit11.Q N1END[1] NN4END[5] N4END[5] Inst_A_IO_1_bidirectional_frame_config_pass.Q
+ Inst_N_IO_ConfigMem.Inst_frame1_bit10.Q Inst_N_IO_switch_matrix.S4BEG12 VPWR VGND
+ sg13g2_mux4_1
X_067_ N1END[3] A_O_top Inst_N_IO_switch_matrix.DEBUG_select_S1BEG0[0] Inst_N_IO_switch_matrix.S1BEG0
+ VPWR VGND sg13g2_mux2_1
XFILLER_8_219 VPWR VGND sg13g2_decap_8
X_119_ Inst_N_IO_ConfigMem.Inst_frame0_bit12.Q N4END[7] N4END[9] N4END[11] Inst_B_IO_1_bidirectional_frame_config_pass.Q
+ Inst_N_IO_ConfigMem.Inst_frame0_bit13.Q Inst_N_IO_switch_matrix.SS4BEG13 VPWR VGND
+ sg13g2_mux4_1
XFILLER_6_73 VPWR VGND sg13g2_fill_1
XFILLER_9_336 VPWR VGND sg13g2_decap_4
XFILLER_1_269 VPWR VGND sg13g2_fill_2
XFILLER_8_380 VPWR VGND sg13g2_fill_2
XFILLER_6_339 VPWR VGND sg13g2_decap_8
X_298_ FrameData[24] FrameData_O[24] VPWR VGND sg13g2_buf_1
X_367_ Inst_N_IO_switch_matrix.SS4BEG5 SS4BEG[5] VPWR VGND sg13g2_buf_1
X_152_ FrameData[10] FrameStrobe[3] B_config_C_bit0 VPWR VGND sg13g2_dlhq_1
X_221_ FrameData[15] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit15.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_5_0 VPWR VGND sg13g2_decap_4
X_083_ VPWR _000_ N2END[1] VGND sg13g2_inv_1
X_204_ FrameData[30] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit30.Q VPWR VGND
+ sg13g2_dlhq_1
X_135_ Inst_N_IO_ConfigMem.Inst_frame1_bit13.Q N1END[0] NN4END[4] N4END[4] Inst_B_IO_1_bidirectional_frame_config_pass.Q
+ Inst_N_IO_ConfigMem.Inst_frame1_bit12.Q Inst_N_IO_switch_matrix.S4BEG13 VPWR VGND
+ sg13g2_mux4_1
X_066_ N1END[2] Inst_A_IO_1_bidirectional_frame_config_pass.Q Inst_N_IO_switch_matrix.DEBUG_select_S1BEG1[0]
+ Inst_N_IO_switch_matrix.S1BEG1 VPWR VGND sg13g2_mux2_1
XFILLER_11_293 VPWR VGND sg13g2_fill_2
XFILLER_11_271 VPWR VGND sg13g2_decap_4
X_118_ Inst_N_IO_ConfigMem.Inst_frame0_bit15.Q N2MID[0] N2MID[4] N2MID[2] N2MID[6]
+ Inst_N_IO_ConfigMem.Inst_frame0_bit14.Q Inst_N_IO_switch_matrix.SS4BEG14 VPWR VGND
+ sg13g2_mux4_1
X_049_ Inst_N_IO_ConfigMem.Inst_frame2_bit14.Q N2END[1] N4END[1] NN4END[1] NN4END[9]
+ Inst_N_IO_ConfigMem.Inst_frame2_bit15.Q Inst_N_IO_switch_matrix.S2BEGb6 VPWR VGND
+ sg13g2_mux4_1
XFILLER_10_336 VPWR VGND sg13g2_fill_1
X_297_ FrameData[23] FrameData_O[23] VPWR VGND sg13g2_buf_1
X_366_ Inst_N_IO_switch_matrix.SS4BEG4 SS4BEG[4] VPWR VGND sg13g2_buf_1
XFILLER_5_340 VPWR VGND sg13g2_fill_2
XFILLER_7_4 VPWR VGND sg13g2_fill_1
XFILLER_3_75 VPWR VGND sg13g2_fill_2
X_151_ FrameData[9] FrameStrobe[3] A_config_C_bit3 VPWR VGND sg13g2_dlhq_1
X_082_ _044_ VPWR B_T_top VGND Inst_N_IO_ConfigMem.Inst_frame0_bit31.Q _041_ sg13g2_o21ai_1
XFILLER_2_354 VPWR VGND sg13g2_decap_4
XFILLER_2_387 VPWR VGND sg13g2_fill_2
X_220_ FrameData[14] FrameStrobe[1] Inst_N_IO_ConfigMem.Inst_frame1_bit14.Q VPWR VGND
+ sg13g2_dlhq_1
X_349_ Inst_N_IO_switch_matrix.S4BEG3 S4BEG[3] VPWR VGND sg13g2_buf_1
XFILLER_0_76 VPWR VGND sg13g2_decap_4
X_065_ N1END[1] B_O_top Inst_N_IO_switch_matrix.DEBUG_select_S1BEG2[0] Inst_N_IO_switch_matrix.S1BEG2
+ VPWR VGND sg13g2_mux2_1
X_134_ Inst_N_IO_ConfigMem.Inst_frame1_bit14.Q N4END[1] NN4END[1] NN4END[13] Inst_A_IO_1_bidirectional_frame_config_pass.Q
+ Inst_N_IO_ConfigMem.Inst_frame1_bit15.Q Inst_N_IO_switch_matrix.S4BEG14 VPWR VGND
+ sg13g2_mux4_1
X_203_ FrameData[29] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit29.Q VPWR VGND
+ sg13g2_dlhq_1
Xclkbuf_0_UserCLK UserCLK clknet_0_UserCLK VPWR VGND sg13g2_buf_8
X_117_ Inst_N_IO_ConfigMem.Inst_frame0_bit17.Q N2MID[1] N2MID[5] N2MID[3] N2MID[7]
+ Inst_N_IO_ConfigMem.Inst_frame0_bit16.Q Inst_N_IO_switch_matrix.SS4BEG15 VPWR VGND
+ sg13g2_mux4_1
X_048_ Inst_N_IO_ConfigMem.Inst_frame2_bit16.Q N2END[0] N4END[0] NN4END[0] NN4END[8]
+ Inst_N_IO_ConfigMem.Inst_frame2_bit17.Q Inst_N_IO_switch_matrix.S2BEGb7 VPWR VGND
+ sg13g2_mux4_1
XFILLER_4_257 VPWR VGND sg13g2_decap_8
XFILLER_4_268 VPWR VGND sg13g2_fill_1
XFILLER_0_271 VPWR VGND sg13g2_decap_8
XFILLER_0_282 VPWR VGND sg13g2_fill_2
X_296_ FrameData[22] FrameData_O[22] VPWR VGND sg13g2_buf_1
X_365_ Inst_N_IO_switch_matrix.SS4BEG3 SS4BEG[3] VPWR VGND sg13g2_buf_1
XFILLER_10_112 VPWR VGND sg13g2_decap_4
X_150_ FrameData[8] FrameStrobe[3] A_config_C_bit2 VPWR VGND sg13g2_dlhq_1
X_081_ _044_ _042_ _043_ VPWR VGND sg13g2_nand2b_1
X_348_ Inst_N_IO_switch_matrix.S4BEG2 S4BEG[2] VPWR VGND sg13g2_buf_1
X_279_ FrameData[5] FrameData_O[5] VPWR VGND sg13g2_buf_1
XFILLER_11_421 VPWR VGND sg13g2_fill_2
X_133_ Inst_N_IO_ConfigMem.Inst_frame1_bit16.Q N4END[0] NN4END[0] NN4END[12] Inst_B_IO_1_bidirectional_frame_config_pass.Q
+ Inst_N_IO_ConfigMem.Inst_frame1_bit17.Q Inst_N_IO_switch_matrix.S4BEG15 VPWR VGND
+ sg13g2_mux4_1
XFILLER_2_130 VPWR VGND sg13g2_fill_1
XFILLER_2_152 VPWR VGND sg13g2_fill_1
X_064_ N1END[0] Inst_B_IO_1_bidirectional_frame_config_pass.Q Inst_N_IO_switch_matrix.DEBUG_select_S1BEG3[0]
+ Inst_N_IO_switch_matrix.S1BEG3 VPWR VGND sg13g2_mux2_1
X_202_ FrameData[28] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit28.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_7_299 VPWR VGND sg13g2_decap_4
X_116_ _031_ VPWR A_I_top VGND _020_ _027_ sg13g2_o21ai_1
X_047_ Inst_N_IO_ConfigMem.Inst_frame2_bit18.Q N1END[2] N4END[15] NN4END[15] A_O_top
+ Inst_N_IO_ConfigMem.Inst_frame2_bit19.Q Inst_N_IO_switch_matrix.S4BEG0 VPWR VGND
+ sg13g2_mux4_1
XFILLER_6_21 VPWR VGND sg13g2_decap_8
X_295_ FrameData[21] FrameData_O[21] VPWR VGND sg13g2_buf_1
X_364_ Inst_N_IO_switch_matrix.SS4BEG2 SS4BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_3_33 VPWR VGND sg13g2_fill_1
XFILLER_3_77 VPWR VGND sg13g2_fill_1
XFILLER_5_342 VPWR VGND sg13g2_fill_1
X_080_ Inst_N_IO_ConfigMem.Inst_frame0_bit31.Q VPWR _043_ VGND Inst_N_IO_ConfigMem.Inst_frame0_bit29.Q
+ _040_ sg13g2_o21ai_1
X_347_ Inst_N_IO_switch_matrix.S4BEG1 S4BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_2_323 VPWR VGND sg13g2_fill_2
X_278_ FrameData[4] FrameData_O[4] VPWR VGND sg13g2_buf_1
X_201_ FrameData[27] FrameStrobe[2] Inst_N_IO_ConfigMem.Inst_frame2_bit27.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_7_404 VPWR VGND sg13g2_decap_4
XFILLER_3_0 VPWR VGND sg13g2_decap_4
X_063_ Inst_N_IO_ConfigMem.Inst_frame3_bit18.Q N2MID[7] N4END[7] NN4END[7] NN4END[15]
+ Inst_N_IO_ConfigMem.Inst_frame3_bit19.Q Inst_N_IO_switch_matrix.S2BEG0 VPWR VGND
+ sg13g2_mux4_1
X_132_ Inst_N_IO_ConfigMem.Inst_frame1_bit18.Q N4END[0] N4END[2] N4END[4] A_O_top
+ Inst_N_IO_ConfigMem.Inst_frame1_bit19.Q Inst_N_IO_switch_matrix.SS4BEG0 VPWR VGND
+ sg13g2_mux4_1
X_115_ _031_ _030_ Inst_N_IO_ConfigMem.Inst_frame0_bit21.Q VPWR VGND sg13g2_nand2b_1
XFILLER_0_421 VPWR VGND sg13g2_fill_2
XFILLER_6_66 VPWR VGND sg13g2_decap_8
XFILLER_8_373 VPWR VGND sg13g2_decap_8
.ends

