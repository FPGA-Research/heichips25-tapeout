module SW_term (UserCLK,
    UserCLKo,
    VPWR,
    VGND,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N2BEG,
    N2BEGb,
    N4BEG,
    S1END,
    S2END,
    S2MID,
    S4END);
 input UserCLK;
 output UserCLKo;
 inout VPWR;
 inout VGND;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 output [15:0] N4BEG;
 input [3:0] S1END;
 input [7:0] S2END;
 input [7:0] S2MID;
 input [15:0] S4END;


 sg13g2_buf_1 _00_ (.A(FrameData[0]),
    .X(FrameData_O[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _01_ (.A(FrameData[1]),
    .X(FrameData_O[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _02_ (.A(FrameData[2]),
    .X(FrameData_O[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _03_ (.A(FrameData[3]),
    .X(FrameData_O[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _04_ (.A(FrameData[4]),
    .X(FrameData_O[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _05_ (.A(FrameData[5]),
    .X(FrameData_O[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _06_ (.A(FrameData[6]),
    .X(FrameData_O[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _07_ (.A(FrameData[7]),
    .X(FrameData_O[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _08_ (.A(FrameData[8]),
    .X(FrameData_O[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _09_ (.A(FrameData[9]),
    .X(FrameData_O[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _10_ (.A(FrameData[10]),
    .X(FrameData_O[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _11_ (.A(FrameData[11]),
    .X(FrameData_O[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _12_ (.A(FrameData[12]),
    .X(FrameData_O[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _13_ (.A(FrameData[13]),
    .X(FrameData_O[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _14_ (.A(FrameData[14]),
    .X(FrameData_O[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _15_ (.A(FrameData[15]),
    .X(FrameData_O[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _16_ (.A(FrameData[16]),
    .X(FrameData_O[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _17_ (.A(FrameData[17]),
    .X(FrameData_O[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _18_ (.A(FrameData[18]),
    .X(FrameData_O[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _19_ (.A(FrameData[19]),
    .X(FrameData_O[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _20_ (.A(FrameData[20]),
    .X(FrameData_O[20]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _21_ (.A(FrameData[21]),
    .X(FrameData_O[21]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _22_ (.A(FrameData[22]),
    .X(FrameData_O[22]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _23_ (.A(FrameData[23]),
    .X(FrameData_O[23]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _24_ (.A(FrameData[24]),
    .X(FrameData_O[24]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _25_ (.A(FrameData[25]),
    .X(FrameData_O[25]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _26_ (.A(FrameData[26]),
    .X(FrameData_O[26]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _27_ (.A(FrameData[27]),
    .X(FrameData_O[27]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _28_ (.A(FrameData[28]),
    .X(FrameData_O[28]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _29_ (.A(FrameData[29]),
    .X(FrameData_O[29]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _30_ (.A(FrameData[30]),
    .X(FrameData_O[30]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _31_ (.A(FrameData[31]),
    .X(FrameData_O[31]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _32_ (.A(FrameStrobe[0]),
    .X(FrameStrobe_O[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _33_ (.A(FrameStrobe[1]),
    .X(FrameStrobe_O[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _34_ (.A(FrameStrobe[2]),
    .X(FrameStrobe_O[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _35_ (.A(FrameStrobe[3]),
    .X(FrameStrobe_O[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _36_ (.A(FrameStrobe[4]),
    .X(FrameStrobe_O[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _37_ (.A(FrameStrobe[5]),
    .X(FrameStrobe_O[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _38_ (.A(FrameStrobe[6]),
    .X(FrameStrobe_O[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _39_ (.A(FrameStrobe[7]),
    .X(FrameStrobe_O[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _40_ (.A(FrameStrobe[8]),
    .X(FrameStrobe_O[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _41_ (.A(FrameStrobe[9]),
    .X(FrameStrobe_O[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _42_ (.A(FrameStrobe[10]),
    .X(FrameStrobe_O[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _43_ (.A(FrameStrobe[11]),
    .X(FrameStrobe_O[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _44_ (.A(FrameStrobe[12]),
    .X(FrameStrobe_O[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _45_ (.A(FrameStrobe[13]),
    .X(FrameStrobe_O[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _46_ (.A(FrameStrobe[14]),
    .X(FrameStrobe_O[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _47_ (.A(FrameStrobe[15]),
    .X(FrameStrobe_O[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _48_ (.A(FrameStrobe[16]),
    .X(FrameStrobe_O[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _49_ (.A(FrameStrobe[17]),
    .X(FrameStrobe_O[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _50_ (.A(FrameStrobe[18]),
    .X(FrameStrobe_O[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _51_ (.A(FrameStrobe[19]),
    .X(FrameStrobe_O[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _52_ (.A(S1END[3]),
    .X(N1BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _53_ (.A(S1END[2]),
    .X(N1BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _54_ (.A(S1END[1]),
    .X(N1BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _55_ (.A(S1END[0]),
    .X(N1BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _56_ (.A(S2MID[7]),
    .X(N2BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _57_ (.A(S2MID[6]),
    .X(N2BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _58_ (.A(S2MID[5]),
    .X(N2BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _59_ (.A(S2MID[4]),
    .X(N2BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _60_ (.A(S2MID[3]),
    .X(N2BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _61_ (.A(S2MID[2]),
    .X(N2BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _62_ (.A(S2MID[1]),
    .X(N2BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _63_ (.A(S2MID[0]),
    .X(N2BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _64_ (.A(S2END[7]),
    .X(N2BEGb[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _65_ (.A(S2END[6]),
    .X(N2BEGb[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _66_ (.A(S2END[5]),
    .X(N2BEGb[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _67_ (.A(S2END[4]),
    .X(N2BEGb[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _68_ (.A(S2END[3]),
    .X(N2BEGb[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _69_ (.A(S2END[2]),
    .X(N2BEGb[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _70_ (.A(S2END[1]),
    .X(N2BEGb[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _71_ (.A(S2END[0]),
    .X(N2BEGb[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _72_ (.A(S4END[15]),
    .X(N4BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _73_ (.A(S4END[14]),
    .X(N4BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _74_ (.A(S4END[13]),
    .X(N4BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _75_ (.A(S4END[12]),
    .X(N4BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _76_ (.A(S4END[11]),
    .X(N4BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _77_ (.A(S4END[10]),
    .X(N4BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _78_ (.A(S4END[9]),
    .X(N4BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _79_ (.A(S4END[8]),
    .X(N4BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _80_ (.A(S4END[7]),
    .X(N4BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _81_ (.A(S4END[6]),
    .X(N4BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _82_ (.A(S4END[5]),
    .X(N4BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _83_ (.A(S4END[4]),
    .X(N4BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _84_ (.A(S4END[3]),
    .X(N4BEG[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _85_ (.A(S4END[2]),
    .X(N4BEG[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _86_ (.A(S4END[1]),
    .X(N4BEG[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _87_ (.A(S4END[0]),
    .X(N4BEG[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _88_ (.A(UserCLK),
    .X(UserCLKo),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_198 (.VDD(VPWR),
    .VSS(VGND));
endmodule
