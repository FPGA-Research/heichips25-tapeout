module heichips25_example_small (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net25;

 sg13g2_and2_1 _29_ (.A(net1),
    .B(net9),
    .X(_00_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _30_ (.A(net2),
    .B(net10),
    .X(_01_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _31_ (.B(net10),
    .A(net2),
    .X(_02_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _32_ (.B(_02_),
    .A(_00_),
    .X(net18),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _33_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_01_),
    .Y(_03_),
    .A2(_02_),
    .A1(_00_));
 sg13g2_and2_1 _34_ (.A(net3),
    .B(net11),
    .X(_04_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _35_ (.Y(_05_),
    .A(net3),
    .B(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _36_ (.A(_03_),
    .B(_05_),
    .Y(_06_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _37_ (.B(_05_),
    .A(_03_),
    .X(net19),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _38_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_07_),
    .B(net12),
    .A(net4));
 sg13g2_and2_1 _39_ (.A(net4),
    .B(net12),
    .X(_08_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _40_ (.B(net12),
    .A(net4),
    .X(_09_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _41_ (.A(_04_),
    .B(_06_),
    .Y(_10_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _42_ (.Y(net20),
    .A(_09_),
    .B(_10_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _43_ (.Y(_11_),
    .B(_09_),
    .A_N(_05_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _44_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04_),
    .A2(_07_),
    .Y(_12_),
    .B1(_08_));
 sg13g2_o21ai_1 _45_ (.B1(_12_),
    .VDD(VPWR),
    .Y(_13_),
    .VSS(VGND),
    .A1(_03_),
    .A2(_11_));
 sg13g2_nand2_1 _46_ (.Y(_14_),
    .A(net5),
    .B(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _47_ (.B(net13),
    .A(net5),
    .X(_15_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _48_ (.VDD(VPWR),
    .Y(_16_),
    .A(_15_),
    .VSS(VGND));
 sg13g2_nand2_1 _49_ (.Y(_17_),
    .A(_13_),
    .B(_15_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _50_ (.Y(net21),
    .A(_13_),
    .B(_16_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _51_ (.A(net6),
    .B(net14),
    .Y(_18_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _52_ (.Y(_19_),
    .A(net6),
    .B(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _53_ (.Y(_20_),
    .A(_14_),
    .B(_17_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _54_ (.Y(net22),
    .A(_19_),
    .B(_20_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _55_ (.A(_16_),
    .B(_19_),
    .Y(_21_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _56_ (.A(_14_),
    .B(_18_),
    .Y(_22_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _57_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_21_),
    .C1(_22_),
    .B1(_13_),
    .A1(net6),
    .Y(_23_),
    .A2(net14));
 sg13g2_nand2_1 _58_ (.Y(_24_),
    .A(net7),
    .B(net15),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _59_ (.A(net7),
    .B(net15),
    .Y(_25_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _60_ (.B(net15),
    .A(net7),
    .X(_26_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _61_ (.Y(net23),
    .A(_23_),
    .B(_26_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _62_ (.B1(_24_),
    .VDD(VPWR),
    .Y(_27_),
    .VSS(VGND),
    .A1(_23_),
    .A2(_25_));
 sg13g2_xnor2_1 _63_ (.Y(_28_),
    .A(net8),
    .B(net16),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _64_ (.Y(net24),
    .A(_27_),
    .B(_28_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _65_ (.B(net9),
    .A(net1),
    .X(net17),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo heichips25_example_small_26 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net26));
 sg13g2_tielo heichips25_example_small_27 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net27));
 sg13g2_tielo heichips25_example_small_28 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net28));
 sg13g2_tielo heichips25_example_small_29 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net29));
 sg13g2_tielo heichips25_example_small_30 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net30));
 sg13g2_tielo heichips25_example_small_31 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net31));
 sg13g2_tielo heichips25_example_small_32 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net32));
 sg13g2_tielo heichips25_example_small_33 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net33));
 sg13g2_tielo heichips25_example_small_34 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net34));
 sg13g2_tielo heichips25_example_small_35 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net35));
 sg13g2_tielo heichips25_example_small_36 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net36));
 sg13g2_tielo heichips25_example_small_37 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net37));
 sg13g2_tielo heichips25_example_small_38 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net38));
 sg13g2_tielo heichips25_example_small_39 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net39));
 sg13g2_tielo heichips25_example_small_40 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net40));
 sg13g2_decap_8 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input13 (.A(uio_in[4]),
    .X(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input14 (.A(uio_in[5]),
    .X(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input15 (.A(uio_in[6]),
    .X(net15),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input16 (.A(uio_in[7]),
    .X(net16),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo heichips25_example_small_25 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net25));
 sg13g2_decap_8 FILLER_0_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_924 (.VDD(VPWR),
    .VSS(VGND));
 assign uio_oe[0] = net25;
 assign uio_oe[1] = net26;
 assign uio_oe[2] = net27;
 assign uio_oe[3] = net28;
 assign uio_oe[4] = net29;
 assign uio_oe[5] = net30;
 assign uio_oe[6] = net31;
 assign uio_oe[7] = net32;
 assign uio_out[0] = net33;
 assign uio_out[1] = net34;
 assign uio_out[2] = net35;
 assign uio_out[3] = net36;
 assign uio_out[4] = net37;
 assign uio_out[5] = net38;
 assign uio_out[6] = net39;
 assign uio_out[7] = net40;
endmodule
