module W_TT_IF (CLK_TT_PROJECT,
    ENA_TT_PROJECT,
    RST_N_TT_PROJECT,
    UIO_IN_TT_PROJECT0,
    UIO_IN_TT_PROJECT1,
    UIO_IN_TT_PROJECT2,
    UIO_IN_TT_PROJECT3,
    UIO_IN_TT_PROJECT4,
    UIO_IN_TT_PROJECT5,
    UIO_IN_TT_PROJECT6,
    UIO_IN_TT_PROJECT7,
    UIO_OE_TT_PROJECT0,
    UIO_OE_TT_PROJECT1,
    UIO_OE_TT_PROJECT2,
    UIO_OE_TT_PROJECT3,
    UIO_OE_TT_PROJECT4,
    UIO_OE_TT_PROJECT5,
    UIO_OE_TT_PROJECT6,
    UIO_OE_TT_PROJECT7,
    UIO_OUT_TT_PROJECT0,
    UIO_OUT_TT_PROJECT1,
    UIO_OUT_TT_PROJECT2,
    UIO_OUT_TT_PROJECT3,
    UIO_OUT_TT_PROJECT4,
    UIO_OUT_TT_PROJECT5,
    UIO_OUT_TT_PROJECT6,
    UIO_OUT_TT_PROJECT7,
    UI_IN_TT_PROJECT0,
    UI_IN_TT_PROJECT1,
    UI_IN_TT_PROJECT2,
    UI_IN_TT_PROJECT3,
    UI_IN_TT_PROJECT4,
    UI_IN_TT_PROJECT5,
    UI_IN_TT_PROJECT6,
    UI_IN_TT_PROJECT7,
    UO_OUT_TT_PROJECT0,
    UO_OUT_TT_PROJECT1,
    UO_OUT_TT_PROJECT2,
    UO_OUT_TT_PROJECT3,
    UO_OUT_TT_PROJECT4,
    UO_OUT_TT_PROJECT5,
    UO_OUT_TT_PROJECT6,
    UO_OUT_TT_PROJECT7,
    UserCLK,
    UserCLKo,
    E1BEG,
    E2BEG,
    E2BEGb,
    E6BEG,
    EE4BEG,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N1END,
    N2BEG,
    N2BEGb,
    N2END,
    N2MID,
    N4BEG,
    N4END,
    S1BEG,
    S1END,
    S2BEG,
    S2BEGb,
    S2END,
    S2MID,
    S4BEG,
    S4END,
    W1END,
    W2END,
    W2MID,
    W6END,
    WW4END);
 output CLK_TT_PROJECT;
 output ENA_TT_PROJECT;
 output RST_N_TT_PROJECT;
 output UIO_IN_TT_PROJECT0;
 output UIO_IN_TT_PROJECT1;
 output UIO_IN_TT_PROJECT2;
 output UIO_IN_TT_PROJECT3;
 output UIO_IN_TT_PROJECT4;
 output UIO_IN_TT_PROJECT5;
 output UIO_IN_TT_PROJECT6;
 output UIO_IN_TT_PROJECT7;
 input UIO_OE_TT_PROJECT0;
 input UIO_OE_TT_PROJECT1;
 input UIO_OE_TT_PROJECT2;
 input UIO_OE_TT_PROJECT3;
 input UIO_OE_TT_PROJECT4;
 input UIO_OE_TT_PROJECT5;
 input UIO_OE_TT_PROJECT6;
 input UIO_OE_TT_PROJECT7;
 input UIO_OUT_TT_PROJECT0;
 input UIO_OUT_TT_PROJECT1;
 input UIO_OUT_TT_PROJECT2;
 input UIO_OUT_TT_PROJECT3;
 input UIO_OUT_TT_PROJECT4;
 input UIO_OUT_TT_PROJECT5;
 input UIO_OUT_TT_PROJECT6;
 input UIO_OUT_TT_PROJECT7;
 output UI_IN_TT_PROJECT0;
 output UI_IN_TT_PROJECT1;
 output UI_IN_TT_PROJECT2;
 output UI_IN_TT_PROJECT3;
 output UI_IN_TT_PROJECT4;
 output UI_IN_TT_PROJECT5;
 output UI_IN_TT_PROJECT6;
 output UI_IN_TT_PROJECT7;
 input UO_OUT_TT_PROJECT0;
 input UO_OUT_TT_PROJECT1;
 input UO_OUT_TT_PROJECT2;
 input UO_OUT_TT_PROJECT3;
 input UO_OUT_TT_PROJECT4;
 input UO_OUT_TT_PROJECT5;
 input UO_OUT_TT_PROJECT6;
 input UO_OUT_TT_PROJECT7;
 input UserCLK;
 output UserCLKo;
 output [3:0] E1BEG;
 output [7:0] E2BEG;
 output [7:0] E2BEGb;
 output [11:0] E6BEG;
 output [15:0] EE4BEG;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 input [3:0] N1END;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 input [7:0] N2END;
 input [7:0] N2MID;
 output [15:0] N4BEG;
 input [15:0] N4END;
 output [3:0] S1BEG;
 input [3:0] S1END;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 input [7:0] S2END;
 input [7:0] S2MID;
 output [15:0] S4BEG;
 input [15:0] S4END;
 input [3:0] W1END;
 input [7:0] W2END;
 input [7:0] W2MID;
 input [11:0] W6END;
 input [15:0] WW4END;

 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit0.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit1.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit2.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit3.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit4.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit5.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit6.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit7.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit0.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit1.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit10.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit11.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit12.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit13.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit14.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit15.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit16.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit17.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit18.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit19.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit2.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit20.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit21.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit22.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit23.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit24.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit25.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit26.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit27.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit28.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit29.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit3.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit30.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit31.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit4.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit5.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit6.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit7.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit8.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame8_bit9.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame9_bit22.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame9_bit23.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame9_bit24.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame9_bit25.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame9_bit26.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame9_bit27.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame9_bit28.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame9_bit29.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame9_bit30.Q ;
 wire \Inst_W_TT_IF_ConfigMem.Inst_frame9_bit31.Q ;
 wire \Inst_W_TT_IF_switch_matrix.E1BEG0 ;
 wire \Inst_W_TT_IF_switch_matrix.E1BEG1 ;
 wire \Inst_W_TT_IF_switch_matrix.E1BEG2 ;
 wire \Inst_W_TT_IF_switch_matrix.E1BEG3 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEG0 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEG1 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEG2 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEG3 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEG4 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEG5 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEG6 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEG7 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEGb0 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEGb1 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEGb2 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEGb3 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEGb4 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEGb5 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEGb6 ;
 wire \Inst_W_TT_IF_switch_matrix.E2BEGb7 ;
 wire \Inst_W_TT_IF_switch_matrix.E6BEG0 ;
 wire \Inst_W_TT_IF_switch_matrix.E6BEG1 ;
 wire \Inst_W_TT_IF_switch_matrix.E6BEG10 ;
 wire \Inst_W_TT_IF_switch_matrix.E6BEG11 ;
 wire \Inst_W_TT_IF_switch_matrix.E6BEG2 ;
 wire \Inst_W_TT_IF_switch_matrix.E6BEG3 ;
 wire \Inst_W_TT_IF_switch_matrix.E6BEG4 ;
 wire \Inst_W_TT_IF_switch_matrix.E6BEG5 ;
 wire \Inst_W_TT_IF_switch_matrix.E6BEG6 ;
 wire \Inst_W_TT_IF_switch_matrix.E6BEG7 ;
 wire \Inst_W_TT_IF_switch_matrix.E6BEG8 ;
 wire \Inst_W_TT_IF_switch_matrix.E6BEG9 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG0 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG1 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG10 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG11 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG12 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG13 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG14 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG15 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG2 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG3 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG4 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG5 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG6 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG7 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG8 ;
 wire \Inst_W_TT_IF_switch_matrix.EE4BEG9 ;
 wire \Inst_W_TT_IF_switch_matrix.N1BEG0 ;
 wire \Inst_W_TT_IF_switch_matrix.N1BEG1 ;
 wire \Inst_W_TT_IF_switch_matrix.N1BEG2 ;
 wire \Inst_W_TT_IF_switch_matrix.N1BEG3 ;
 wire \Inst_W_TT_IF_switch_matrix.N2BEG0 ;
 wire \Inst_W_TT_IF_switch_matrix.N2BEG1 ;
 wire \Inst_W_TT_IF_switch_matrix.N2BEG2 ;
 wire \Inst_W_TT_IF_switch_matrix.N2BEG3 ;
 wire \Inst_W_TT_IF_switch_matrix.N2BEG4 ;
 wire \Inst_W_TT_IF_switch_matrix.N2BEG5 ;
 wire \Inst_W_TT_IF_switch_matrix.N2BEG6 ;
 wire \Inst_W_TT_IF_switch_matrix.N2BEG7 ;
 wire \Inst_W_TT_IF_switch_matrix.N4BEG0 ;
 wire \Inst_W_TT_IF_switch_matrix.N4BEG1 ;
 wire \Inst_W_TT_IF_switch_matrix.N4BEG2 ;
 wire \Inst_W_TT_IF_switch_matrix.N4BEG3 ;
 wire \Inst_W_TT_IF_switch_matrix.S1BEG0 ;
 wire \Inst_W_TT_IF_switch_matrix.S1BEG1 ;
 wire \Inst_W_TT_IF_switch_matrix.S1BEG2 ;
 wire \Inst_W_TT_IF_switch_matrix.S1BEG3 ;
 wire \Inst_W_TT_IF_switch_matrix.S2BEG0 ;
 wire \Inst_W_TT_IF_switch_matrix.S2BEG1 ;
 wire \Inst_W_TT_IF_switch_matrix.S2BEG2 ;
 wire \Inst_W_TT_IF_switch_matrix.S2BEG3 ;
 wire \Inst_W_TT_IF_switch_matrix.S2BEG4 ;
 wire \Inst_W_TT_IF_switch_matrix.S2BEG5 ;
 wire \Inst_W_TT_IF_switch_matrix.S2BEG6 ;
 wire \Inst_W_TT_IF_switch_matrix.S2BEG7 ;
 wire \Inst_W_TT_IF_switch_matrix.S4BEG0 ;
 wire \Inst_W_TT_IF_switch_matrix.S4BEG1 ;
 wire \Inst_W_TT_IF_switch_matrix.S4BEG2 ;
 wire \Inst_W_TT_IF_switch_matrix.S4BEG3 ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire clknet_0_UserCLK;
 wire clknet_1_0__leaf_UserCLK;
 wire clknet_1_1__leaf_UserCLK;

 sg13g2_inv_1 _0381_ (.Y(_0000_),
    .A(W2END[3]));
 sg13g2_inv_1 _0382_ (.Y(_0001_),
    .A(W1END[3]));
 sg13g2_inv_1 _0383_ (.Y(_0002_),
    .A(S1END[3]));
 sg13g2_inv_1 _0384_ (.Y(_0003_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit1.Q ));
 sg13g2_inv_1 _0385_ (.Y(_0004_),
    .A(W1END[2]));
 sg13g2_inv_1 _0386_ (.Y(_0005_),
    .A(S1END[2]));
 sg13g2_inv_1 _0387_ (.Y(_0006_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit30.Q ));
 sg13g2_inv_1 _0388_ (.Y(_0007_),
    .A(S1END[1]));
 sg13g2_inv_1 _0389_ (.Y(_0008_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit27.Q ));
 sg13g2_inv_1 _0390_ (.Y(_0009_),
    .A(S1END[0]));
 sg13g2_inv_1 _0391_ (.Y(_0010_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit24.Q ));
 sg13g2_inv_1 _0392_ (.Y(_0011_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit21.Q ));
 sg13g2_inv_1 _0393_ (.Y(_0012_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit18.Q ));
 sg13g2_inv_1 _0394_ (.Y(_0013_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit15.Q ));
 sg13g2_inv_1 _0395_ (.Y(_0014_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit12.Q ));
 sg13g2_inv_1 _0396_ (.Y(_0015_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit6.Q ));
 sg13g2_inv_1 _0397_ (.Y(_0016_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit3.Q ));
 sg13g2_inv_1 _0398_ (.Y(_0017_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit0.Q ));
 sg13g2_inv_1 _0399_ (.Y(_0018_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit29.Q ));
 sg13g2_inv_1 _0400_ (.Y(_0019_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit26.Q ));
 sg13g2_inv_1 _0401_ (.Y(_0020_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit23.Q ));
 sg13g2_inv_1 _0402_ (.Y(_0021_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit20.Q ));
 sg13g2_inv_1 _0403_ (.Y(_0022_),
    .A(UO_OUT_TT_PROJECT7));
 sg13g2_inv_1 _0404_ (.Y(_0023_),
    .A(UO_OUT_TT_PROJECT6));
 sg13g2_inv_1 _0405_ (.Y(_0024_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit27.Q ));
 sg13g2_inv_1 _0406_ (.Y(_0025_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit24.Q ));
 sg13g2_inv_1 _0407_ (.Y(_0026_),
    .A(UO_OUT_TT_PROJECT3));
 sg13g2_inv_1 _0408_ (.Y(_0027_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit21.Q ));
 sg13g2_inv_1 _0409_ (.Y(_0028_),
    .A(UO_OUT_TT_PROJECT2));
 sg13g2_inv_1 _0410_ (.Y(_0029_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit18.Q ));
 sg13g2_inv_1 _0411_ (.Y(_0030_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit10.Q ));
 sg13g2_inv_1 _0412_ (.Y(_0031_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit29.Q ));
 sg13g2_inv_1 _0413_ (.Y(_0032_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit26.Q ));
 sg13g2_inv_1 _0414_ (.Y(_0033_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit25.Q ));
 sg13g2_inv_1 _0415_ (.Y(_0034_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit22.Q ));
 sg13g2_inv_1 _0416_ (.Y(_0035_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit19.Q ));
 sg13g2_inv_1 _0417_ (.Y(_0036_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit16.Q ));
 sg13g2_mux4_1 _0418_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit4.Q ),
    .A0(W2MID[3]),
    .A1(W2MID[6]),
    .A2(W2END[1]),
    .A3(W2END[2]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit5.Q ),
    .X(_0037_));
 sg13g2_inv_1 _0419_ (.Y(_0038_),
    .A(_0037_));
 sg13g2_nor2_1 _0420_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit5.Q ),
    .B(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit6.Q ),
    .Y(_0039_));
 sg13g2_mux4_1 _0421_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit4.Q ),
    .A0(N2MID[6]),
    .A1(N2END[2]),
    .A2(N2END[3]),
    .A3(W2MID[0]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit5.Q ),
    .X(_0040_));
 sg13g2_a21oi_1 _0422_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit6.Q ),
    .A2(_0038_),
    .Y(_0041_),
    .B1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit7.Q ));
 sg13g2_o21ai_1 _0423_ (.B1(_0041_),
    .Y(_0042_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit6.Q ),
    .A2(_0040_));
 sg13g2_o21ai_1 _0424_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit5.Q ),
    .Y(_0043_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit6.Q ),
    .A2(S2MID[0]));
 sg13g2_a22oi_1 _0425_ (.Y(_0044_),
    .B1(_0039_),
    .B2(W2END[4]),
    .A2(S2END[3]),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit6.Q ));
 sg13g2_nand3_1 _0426_ (.B(_0043_),
    .C(_0044_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit4.Q ),
    .Y(_0045_));
 sg13g2_nand2b_1 _0427_ (.Y(_0046_),
    .B(S2END[2]),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit5.Q ));
 sg13g2_a22oi_1 _0428_ (.Y(_0047_),
    .B1(_0046_),
    .B2(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit6.Q ),
    .A2(_0039_),
    .A1(_0000_));
 sg13g2_nand2b_1 _0429_ (.Y(_0048_),
    .B(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit5.Q ),
    .A_N(W2END[5]));
 sg13g2_a21oi_1 _0430_ (.A1(_0047_),
    .A2(_0048_),
    .Y(_0049_),
    .B1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit4.Q ));
 sg13g2_nand2_1 _0431_ (.Y(_0050_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit7.Q ),
    .B(_0045_));
 sg13g2_o21ai_1 _0432_ (.B1(_0042_),
    .Y(RST_N_TT_PROJECT),
    .A1(_0049_),
    .A2(_0050_));
 sg13g2_mux4_1 _0433_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit6.Q ),
    .A0(N1END[3]),
    .A1(N4END[3]),
    .A2(S1END[3]),
    .A3(S4END[3]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit7.Q ),
    .X(_0051_));
 sg13g2_mux4_1 _0434_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit22.Q ),
    .A0(N2MID[7]),
    .A1(N2END[7]),
    .A2(S2MID[7]),
    .A3(S2END[7]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit23.Q ),
    .X(_0052_));
 sg13g2_inv_1 _0435_ (.Y(_0053_),
    .A(_0052_));
 sg13g2_nand3_1 _0436_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit1.Q ),
    .C(_0052_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit0.Q ),
    .Y(_0054_));
 sg13g2_mux2_1 _0437_ (.A0(W1END[3]),
    .A1(W2END[7]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit0.Q ),
    .X(_0055_));
 sg13g2_nor2_1 _0438_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit0.Q ),
    .B(_0003_),
    .Y(_0056_));
 sg13g2_a221oi_1 _0439_ (.B2(WW4END[15]),
    .C1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit31.Q ),
    .B1(_0056_),
    .A1(_0003_),
    .Y(_0057_),
    .A2(_0055_));
 sg13g2_mux2_1 _0440_ (.A0(W2MID[7]),
    .A1(WW4END[7]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit0.Q ),
    .X(_0058_));
 sg13g2_a22oi_1 _0441_ (.Y(_0059_),
    .B1(_0058_),
    .B2(_0003_),
    .A2(_0056_),
    .A1(_0051_));
 sg13g2_a22oi_1 _0442_ (.Y(UIO_IN_TT_PROJECT7),
    .B1(_0059_),
    .B2(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit31.Q ),
    .A2(_0057_),
    .A1(_0054_));
 sg13g2_mux4_1 _0443_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit4.Q ),
    .A0(N1END[2]),
    .A1(N4END[2]),
    .A2(S1END[2]),
    .A3(S4END[2]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit5.Q ),
    .X(_0060_));
 sg13g2_mux4_1 _0444_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit20.Q ),
    .A0(N2MID[6]),
    .A1(N2END[6]),
    .A2(S2MID[6]),
    .A3(S2END[6]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit21.Q ),
    .X(_0061_));
 sg13g2_inv_1 _0445_ (.Y(_0062_),
    .A(_0061_));
 sg13g2_nand3_1 _0446_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit30.Q ),
    .C(_0061_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit29.Q ),
    .Y(_0063_));
 sg13g2_mux2_1 _0447_ (.A0(W1END[2]),
    .A1(W2END[6]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit29.Q ),
    .X(_0064_));
 sg13g2_nor2_1 _0448_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit29.Q ),
    .B(_0006_),
    .Y(_0065_));
 sg13g2_a221oi_1 _0449_ (.B2(WW4END[14]),
    .C1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit28.Q ),
    .B1(_0065_),
    .A1(_0006_),
    .Y(_0066_),
    .A2(_0064_));
 sg13g2_mux2_1 _0450_ (.A0(W2MID[6]),
    .A1(WW4END[6]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit29.Q ),
    .X(_0067_));
 sg13g2_a22oi_1 _0451_ (.Y(_0068_),
    .B1(_0067_),
    .B2(_0006_),
    .A2(_0065_),
    .A1(_0060_));
 sg13g2_a22oi_1 _0452_ (.Y(UIO_IN_TT_PROJECT6),
    .B1(_0068_),
    .B2(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit28.Q ),
    .A2(_0066_),
    .A1(_0063_));
 sg13g2_mux4_1 _0453_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit2.Q ),
    .A0(N1END[1]),
    .A1(N4END[1]),
    .A2(S1END[1]),
    .A3(S4END[1]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit3.Q ),
    .X(_0069_));
 sg13g2_mux4_1 _0454_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit18.Q ),
    .A0(N2MID[5]),
    .A1(N2END[5]),
    .A2(S2MID[5]),
    .A3(S2END[5]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit19.Q ),
    .X(_0070_));
 sg13g2_inv_1 _0455_ (.Y(_0071_),
    .A(_0070_));
 sg13g2_nand3_1 _0456_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit27.Q ),
    .C(_0070_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit26.Q ),
    .Y(_0072_));
 sg13g2_mux2_1 _0457_ (.A0(W1END[1]),
    .A1(W2END[5]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit26.Q ),
    .X(_0073_));
 sg13g2_nor2_1 _0458_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit26.Q ),
    .B(_0008_),
    .Y(_0074_));
 sg13g2_a221oi_1 _0459_ (.B2(WW4END[13]),
    .C1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit25.Q ),
    .B1(_0074_),
    .A1(_0008_),
    .Y(_0075_),
    .A2(_0073_));
 sg13g2_mux2_1 _0460_ (.A0(W2MID[5]),
    .A1(WW4END[5]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit26.Q ),
    .X(_0076_));
 sg13g2_a22oi_1 _0461_ (.Y(_0077_),
    .B1(_0076_),
    .B2(_0008_),
    .A2(_0074_),
    .A1(_0069_));
 sg13g2_a22oi_1 _0462_ (.Y(UIO_IN_TT_PROJECT5),
    .B1(_0077_),
    .B2(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit25.Q ),
    .A2(_0075_),
    .A1(_0072_));
 sg13g2_mux4_1 _0463_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit0.Q ),
    .A0(N1END[0]),
    .A1(N4END[0]),
    .A2(S1END[0]),
    .A3(S4END[0]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit1.Q ),
    .X(_0078_));
 sg13g2_mux4_1 _0464_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit16.Q ),
    .A0(N2MID[4]),
    .A1(N2END[4]),
    .A2(S2MID[4]),
    .A3(S2END[4]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit17.Q ),
    .X(_0079_));
 sg13g2_inv_1 _0465_ (.Y(_0080_),
    .A(_0079_));
 sg13g2_nand3_1 _0466_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit24.Q ),
    .C(_0079_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit23.Q ),
    .Y(_0081_));
 sg13g2_mux2_1 _0467_ (.A0(W1END[0]),
    .A1(W2END[4]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit23.Q ),
    .X(_0082_));
 sg13g2_nor2_1 _0468_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit23.Q ),
    .B(_0010_),
    .Y(_0083_));
 sg13g2_a221oi_1 _0469_ (.B2(WW4END[12]),
    .C1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit22.Q ),
    .B1(_0083_),
    .A1(_0010_),
    .Y(_0084_),
    .A2(_0082_));
 sg13g2_mux2_1 _0470_ (.A0(W2MID[4]),
    .A1(WW4END[4]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit23.Q ),
    .X(_0085_));
 sg13g2_a22oi_1 _0471_ (.Y(_0086_),
    .B1(_0085_),
    .B2(_0010_),
    .A2(_0083_),
    .A1(_0078_));
 sg13g2_a22oi_1 _0472_ (.Y(UIO_IN_TT_PROJECT4),
    .B1(_0086_),
    .B2(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit22.Q ),
    .A2(_0084_),
    .A1(_0081_));
 sg13g2_mux4_1 _0473_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit30.Q ),
    .A0(N1END[3]),
    .A1(N4END[3]),
    .A2(S1END[3]),
    .A3(S4END[3]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit31.Q ),
    .X(_0087_));
 sg13g2_mux4_1 _0474_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit15.Q ),
    .A0(N2MID[3]),
    .A1(S2MID[3]),
    .A2(N2END[3]),
    .A3(S2END[3]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit14.Q ),
    .X(_0088_));
 sg13g2_nand3_1 _0475_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit21.Q ),
    .C(_0088_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit20.Q ),
    .Y(_0089_));
 sg13g2_mux2_1 _0476_ (.A0(W2MID[3]),
    .A1(WW4END[3]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit20.Q ),
    .X(_0090_));
 sg13g2_nor2_1 _0477_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit20.Q ),
    .B(_0011_),
    .Y(_0091_));
 sg13g2_a221oi_1 _0478_ (.B2(W6END[11]),
    .C1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit19.Q ),
    .B1(_0091_),
    .A1(_0011_),
    .Y(_0092_),
    .A2(_0090_));
 sg13g2_mux2_1 _0479_ (.A0(W2END[3]),
    .A1(WW4END[11]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit20.Q ),
    .X(_0093_));
 sg13g2_a22oi_1 _0480_ (.Y(_0094_),
    .B1(_0093_),
    .B2(_0011_),
    .A2(_0091_),
    .A1(_0087_));
 sg13g2_a22oi_1 _0481_ (.Y(UIO_IN_TT_PROJECT3),
    .B1(_0094_),
    .B2(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit19.Q ),
    .A2(_0092_),
    .A1(_0089_));
 sg13g2_mux4_1 _0482_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit28.Q ),
    .A0(N1END[2]),
    .A1(N4END[2]),
    .A2(S1END[2]),
    .A3(S4END[2]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit29.Q ),
    .X(_0095_));
 sg13g2_mux4_1 _0483_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit13.Q ),
    .A0(N2MID[2]),
    .A1(S2MID[2]),
    .A2(N2END[2]),
    .A3(S2END[2]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit12.Q ),
    .X(_0096_));
 sg13g2_nand3_1 _0484_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit18.Q ),
    .C(_0096_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit17.Q ),
    .Y(_0097_));
 sg13g2_mux2_1 _0485_ (.A0(W2MID[2]),
    .A1(WW4END[2]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit17.Q ),
    .X(_0098_));
 sg13g2_nor2_1 _0486_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit17.Q ),
    .B(_0012_),
    .Y(_0099_));
 sg13g2_a221oi_1 _0487_ (.B2(W6END[10]),
    .C1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit16.Q ),
    .B1(_0099_),
    .A1(_0012_),
    .Y(_0100_),
    .A2(_0098_));
 sg13g2_mux2_1 _0488_ (.A0(W2END[2]),
    .A1(WW4END[10]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit17.Q ),
    .X(_0101_));
 sg13g2_a22oi_1 _0489_ (.Y(_0102_),
    .B1(_0101_),
    .B2(_0012_),
    .A2(_0099_),
    .A1(_0095_));
 sg13g2_a22oi_1 _0490_ (.Y(UIO_IN_TT_PROJECT2),
    .B1(_0102_),
    .B2(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit16.Q ),
    .A2(_0100_),
    .A1(_0097_));
 sg13g2_mux4_1 _0491_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit26.Q ),
    .A0(N1END[1]),
    .A1(N4END[1]),
    .A2(S1END[1]),
    .A3(S4END[1]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit27.Q ),
    .X(_0103_));
 sg13g2_mux4_1 _0492_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit10.Q ),
    .A0(N2MID[1]),
    .A1(N2END[1]),
    .A2(S2MID[1]),
    .A3(S2END[1]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit11.Q ),
    .X(_0104_));
 sg13g2_nand3_1 _0493_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit15.Q ),
    .C(_0104_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit14.Q ),
    .Y(_0105_));
 sg13g2_mux2_1 _0494_ (.A0(W2MID[1]),
    .A1(WW4END[1]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit14.Q ),
    .X(_0106_));
 sg13g2_nor2_1 _0495_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit14.Q ),
    .B(_0013_),
    .Y(_0107_));
 sg13g2_a221oi_1 _0496_ (.B2(W6END[9]),
    .C1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit13.Q ),
    .B1(_0107_),
    .A1(_0013_),
    .Y(_0108_),
    .A2(_0106_));
 sg13g2_mux2_1 _0497_ (.A0(W2END[1]),
    .A1(WW4END[9]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit14.Q ),
    .X(_0109_));
 sg13g2_a22oi_1 _0498_ (.Y(_0110_),
    .B1(_0109_),
    .B2(_0013_),
    .A2(_0107_),
    .A1(_0103_));
 sg13g2_a22oi_1 _0499_ (.Y(UIO_IN_TT_PROJECT1),
    .B1(_0110_),
    .B2(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit13.Q ),
    .A2(_0108_),
    .A1(_0105_));
 sg13g2_mux4_1 _0500_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit24.Q ),
    .A0(N1END[0]),
    .A1(N4END[0]),
    .A2(S1END[0]),
    .A3(S4END[0]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit25.Q ),
    .X(_0111_));
 sg13g2_mux4_1 _0501_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit8.Q ),
    .A0(N2MID[0]),
    .A1(N2END[0]),
    .A2(S2MID[0]),
    .A3(S2END[0]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit9.Q ),
    .X(_0112_));
 sg13g2_nand3_1 _0502_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit12.Q ),
    .C(_0112_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit11.Q ),
    .Y(_0113_));
 sg13g2_mux2_1 _0503_ (.A0(W2MID[0]),
    .A1(WW4END[0]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit11.Q ),
    .X(_0114_));
 sg13g2_nor2_1 _0504_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit11.Q ),
    .B(_0014_),
    .Y(_0115_));
 sg13g2_a221oi_1 _0505_ (.B2(W6END[8]),
    .C1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit10.Q ),
    .B1(_0115_),
    .A1(_0014_),
    .Y(_0116_),
    .A2(_0114_));
 sg13g2_mux2_1 _0506_ (.A0(W2END[0]),
    .A1(WW4END[8]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit11.Q ),
    .X(_0117_));
 sg13g2_a22oi_1 _0507_ (.Y(_0118_),
    .B1(_0117_),
    .B2(_0014_),
    .A2(_0115_),
    .A1(_0111_));
 sg13g2_a22oi_1 _0508_ (.Y(UIO_IN_TT_PROJECT0),
    .B1(_0118_),
    .B2(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit10.Q ),
    .A2(_0116_),
    .A1(_0113_));
 sg13g2_nor2_1 _0509_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit8.Q ),
    .B(W6END[7]),
    .Y(_0119_));
 sg13g2_mux4_1 _0510_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit22.Q ),
    .A0(N1END[3]),
    .A1(N4END[3]),
    .A2(S1END[3]),
    .A3(S4END[3]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit23.Q ),
    .X(_0120_));
 sg13g2_nand3b_1 _0511_ (.B(_0120_),
    .C(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit7.Q ),
    .Y(_0121_),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit8.Q ));
 sg13g2_and2_1 _0512_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit9.Q ),
    .B(_0121_),
    .X(_0122_));
 sg13g2_a21oi_1 _0513_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit8.Q ),
    .A2(_0053_),
    .Y(_0123_),
    .B1(_0119_));
 sg13g2_nand2b_1 _0514_ (.Y(_0124_),
    .B(_0123_),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit7.Q ));
 sg13g2_mux4_1 _0515_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit7.Q ),
    .A0(W2MID[7]),
    .A1(W2END[7]),
    .A2(WW4END[7]),
    .A3(WW4END[15]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit8.Q ),
    .X(_0125_));
 sg13g2_nor2_1 _0516_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit9.Q ),
    .B(_0125_),
    .Y(_0126_));
 sg13g2_a21oi_1 _0517_ (.A1(_0122_),
    .A2(_0124_),
    .Y(UI_IN_TT_PROJECT7),
    .B1(_0126_));
 sg13g2_mux4_1 _0518_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit20.Q ),
    .A0(N1END[2]),
    .A1(N4END[2]),
    .A2(S1END[2]),
    .A3(S4END[2]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit21.Q ),
    .X(_0127_));
 sg13g2_nand3_1 _0519_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit6.Q ),
    .C(_0061_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit5.Q ),
    .Y(_0128_));
 sg13g2_mux2_1 _0520_ (.A0(W2MID[6]),
    .A1(WW4END[6]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit5.Q ),
    .X(_0129_));
 sg13g2_nor2_1 _0521_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit5.Q ),
    .B(_0015_),
    .Y(_0130_));
 sg13g2_a221oi_1 _0522_ (.B2(W6END[6]),
    .C1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit4.Q ),
    .B1(_0130_),
    .A1(_0015_),
    .Y(_0131_),
    .A2(_0129_));
 sg13g2_mux2_1 _0523_ (.A0(W2END[6]),
    .A1(WW4END[14]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit5.Q ),
    .X(_0132_));
 sg13g2_a22oi_1 _0524_ (.Y(_0133_),
    .B1(_0132_),
    .B2(_0015_),
    .A2(_0130_),
    .A1(_0127_));
 sg13g2_a22oi_1 _0525_ (.Y(UI_IN_TT_PROJECT6),
    .B1(_0133_),
    .B2(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit4.Q ),
    .A2(_0131_),
    .A1(_0128_));
 sg13g2_mux4_1 _0526_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit18.Q ),
    .A0(N1END[1]),
    .A1(N4END[1]),
    .A2(S1END[1]),
    .A3(S4END[1]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit19.Q ),
    .X(_0134_));
 sg13g2_nand3_1 _0527_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit3.Q ),
    .C(_0070_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit2.Q ),
    .Y(_0135_));
 sg13g2_mux2_1 _0528_ (.A0(W2MID[5]),
    .A1(WW4END[5]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit2.Q ),
    .X(_0136_));
 sg13g2_nor2_1 _0529_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit2.Q ),
    .B(_0016_),
    .Y(_0137_));
 sg13g2_a221oi_1 _0530_ (.B2(W6END[5]),
    .C1(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit1.Q ),
    .B1(_0137_),
    .A1(_0016_),
    .Y(_0138_),
    .A2(_0136_));
 sg13g2_mux2_1 _0531_ (.A0(W2END[5]),
    .A1(WW4END[13]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit2.Q ),
    .X(_0139_));
 sg13g2_a22oi_1 _0532_ (.Y(_0140_),
    .B1(_0139_),
    .B2(_0016_),
    .A2(_0137_),
    .A1(_0134_));
 sg13g2_a22oi_1 _0533_ (.Y(UI_IN_TT_PROJECT5),
    .B1(_0140_),
    .B2(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit1.Q ),
    .A2(_0138_),
    .A1(_0135_));
 sg13g2_mux4_1 _0534_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit16.Q ),
    .A0(N1END[0]),
    .A1(N4END[0]),
    .A2(S1END[0]),
    .A3(S4END[0]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit17.Q ),
    .X(_0141_));
 sg13g2_nand3_1 _0535_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit0.Q ),
    .C(_0079_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit31.Q ),
    .Y(_0142_));
 sg13g2_mux2_1 _0536_ (.A0(W2MID[4]),
    .A1(WW4END[4]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit31.Q ),
    .X(_0143_));
 sg13g2_nor2_1 _0537_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit31.Q ),
    .B(_0017_),
    .Y(_0144_));
 sg13g2_a221oi_1 _0538_ (.B2(W6END[4]),
    .C1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit30.Q ),
    .B1(_0144_),
    .A1(_0017_),
    .Y(_0145_),
    .A2(_0143_));
 sg13g2_mux2_1 _0539_ (.A0(W2END[4]),
    .A1(WW4END[12]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit31.Q ),
    .X(_0146_));
 sg13g2_a22oi_1 _0540_ (.Y(_0147_),
    .B1(_0146_),
    .B2(_0017_),
    .A2(_0144_),
    .A1(_0141_));
 sg13g2_a22oi_1 _0541_ (.Y(UI_IN_TT_PROJECT4),
    .B1(_0147_),
    .B2(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit30.Q ),
    .A2(_0145_),
    .A1(_0142_));
 sg13g2_mux4_1 _0542_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit14.Q ),
    .A0(N1END[3]),
    .A1(N4END[3]),
    .A2(S1END[3]),
    .A3(S4END[3]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit15.Q ),
    .X(_0148_));
 sg13g2_nand3_1 _0543_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit29.Q ),
    .C(_0088_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit28.Q ),
    .Y(_0149_));
 sg13g2_mux2_1 _0544_ (.A0(W2MID[3]),
    .A1(WW4END[3]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit28.Q ),
    .X(_0150_));
 sg13g2_nor2_1 _0545_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit28.Q ),
    .B(_0018_),
    .Y(_0151_));
 sg13g2_a221oi_1 _0546_ (.B2(W6END[3]),
    .C1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit27.Q ),
    .B1(_0151_),
    .A1(_0018_),
    .Y(_0152_),
    .A2(_0150_));
 sg13g2_mux2_1 _0547_ (.A0(W2END[3]),
    .A1(WW4END[11]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit28.Q ),
    .X(_0153_));
 sg13g2_a22oi_1 _0548_ (.Y(_0154_),
    .B1(_0153_),
    .B2(_0018_),
    .A2(_0151_),
    .A1(_0148_));
 sg13g2_a22oi_1 _0549_ (.Y(UI_IN_TT_PROJECT3),
    .B1(_0154_),
    .B2(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit27.Q ),
    .A2(_0152_),
    .A1(_0149_));
 sg13g2_mux4_1 _0550_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit12.Q ),
    .A0(N1END[2]),
    .A1(N4END[2]),
    .A2(S1END[2]),
    .A3(S4END[2]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_0155_));
 sg13g2_nand3_1 _0551_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit26.Q ),
    .C(_0096_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit25.Q ),
    .Y(_0156_));
 sg13g2_mux2_1 _0552_ (.A0(W2MID[2]),
    .A1(WW4END[2]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit25.Q ),
    .X(_0157_));
 sg13g2_nor2_1 _0553_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit25.Q ),
    .B(_0019_),
    .Y(_0158_));
 sg13g2_a221oi_1 _0554_ (.B2(W6END[2]),
    .C1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit24.Q ),
    .B1(_0158_),
    .A1(_0019_),
    .Y(_0159_),
    .A2(_0157_));
 sg13g2_mux2_1 _0555_ (.A0(W2END[2]),
    .A1(WW4END[10]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit25.Q ),
    .X(_0160_));
 sg13g2_a22oi_1 _0556_ (.Y(_0161_),
    .B1(_0160_),
    .B2(_0019_),
    .A2(_0158_),
    .A1(_0155_));
 sg13g2_a22oi_1 _0557_ (.Y(UI_IN_TT_PROJECT2),
    .B1(_0161_),
    .B2(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit24.Q ),
    .A2(_0159_),
    .A1(_0156_));
 sg13g2_mux4_1 _0558_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit10.Q ),
    .A0(N1END[1]),
    .A1(N4END[1]),
    .A2(S1END[1]),
    .A3(S4END[1]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit11.Q ),
    .X(_0162_));
 sg13g2_nand3_1 _0559_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit23.Q ),
    .C(_0104_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit22.Q ),
    .Y(_0163_));
 sg13g2_mux2_1 _0560_ (.A0(W2MID[1]),
    .A1(WW4END[1]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit22.Q ),
    .X(_0164_));
 sg13g2_nor2_1 _0561_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit22.Q ),
    .B(_0020_),
    .Y(_0165_));
 sg13g2_a221oi_1 _0562_ (.B2(W6END[1]),
    .C1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit21.Q ),
    .B1(_0165_),
    .A1(_0020_),
    .Y(_0166_),
    .A2(_0164_));
 sg13g2_mux2_1 _0563_ (.A0(W2END[1]),
    .A1(WW4END[9]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit22.Q ),
    .X(_0167_));
 sg13g2_a22oi_1 _0564_ (.Y(_0168_),
    .B1(_0167_),
    .B2(_0020_),
    .A2(_0165_),
    .A1(_0162_));
 sg13g2_a22oi_1 _0565_ (.Y(UI_IN_TT_PROJECT1),
    .B1(_0168_),
    .B2(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit21.Q ),
    .A2(_0166_),
    .A1(_0163_));
 sg13g2_mux4_1 _0566_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit8.Q ),
    .A0(N1END[0]),
    .A1(N4END[0]),
    .A2(S1END[0]),
    .A3(S4END[0]),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_0169_));
 sg13g2_nand3_1 _0567_ (.B(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit20.Q ),
    .C(_0112_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit19.Q ),
    .Y(_0170_));
 sg13g2_mux2_1 _0568_ (.A0(W2MID[0]),
    .A1(WW4END[0]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit19.Q ),
    .X(_0171_));
 sg13g2_nor2_1 _0569_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit19.Q ),
    .B(_0021_),
    .Y(_0172_));
 sg13g2_a221oi_1 _0570_ (.B2(W6END[0]),
    .C1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit18.Q ),
    .B1(_0172_),
    .A1(_0021_),
    .Y(_0173_),
    .A2(_0171_));
 sg13g2_mux2_1 _0571_ (.A0(W2END[0]),
    .A1(WW4END[8]),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit19.Q ),
    .X(_0174_));
 sg13g2_a22oi_1 _0572_ (.Y(_0175_),
    .B1(_0174_),
    .B2(_0021_),
    .A2(_0172_),
    .A1(_0169_));
 sg13g2_a22oi_1 _0573_ (.Y(UI_IN_TT_PROJECT0),
    .B1(_0175_),
    .B2(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit18.Q ),
    .A2(_0173_),
    .A1(_0170_));
 sg13g2_o21ai_1 _0574_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit24.Q ),
    .Y(_0176_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit23.Q ),
    .A2(_0112_));
 sg13g2_a21oi_1 _0575_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit23.Q ),
    .A2(_0053_),
    .Y(_0177_),
    .B1(_0176_));
 sg13g2_nor2b_1 _0576_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit23.Q ),
    .B_N(UIO_OE_TT_PROJECT7),
    .Y(_0178_));
 sg13g2_a21oi_1 _0577_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit23.Q ),
    .A2(_0051_),
    .Y(_0179_),
    .B1(_0178_));
 sg13g2_o21ai_1 _0578_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit25.Q ),
    .Y(_0180_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit24.Q ),
    .A2(_0179_));
 sg13g2_nor2_1 _0579_ (.A(_0177_),
    .B(_0180_),
    .Y(_0181_));
 sg13g2_mux4_1 _0580_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit23.Q ),
    .A0(W2END[0]),
    .A1(UIO_OUT_TT_PROJECT0),
    .A2(UIO_OUT_TT_PROJECT4),
    .A3(UIO_OUT_TT_PROJECT7),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit24.Q ),
    .X(_0182_));
 sg13g2_nor2_1 _0581_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit25.Q ),
    .B(_0182_),
    .Y(_0183_));
 sg13g2_nor2_1 _0582_ (.A(_0181_),
    .B(_0183_),
    .Y(\Inst_W_TT_IF_switch_matrix.E2BEGb7 ));
 sg13g2_o21ai_1 _0583_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit21.Q ),
    .Y(_0184_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit20.Q ),
    .A2(_0104_));
 sg13g2_a21oi_1 _0584_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit20.Q ),
    .A2(_0062_),
    .Y(_0185_),
    .B1(_0184_));
 sg13g2_nor2b_1 _0585_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit20.Q ),
    .B_N(UIO_OE_TT_PROJECT6),
    .Y(_0186_));
 sg13g2_a21oi_1 _0586_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit20.Q ),
    .A2(_0060_),
    .Y(_0187_),
    .B1(_0186_));
 sg13g2_o21ai_1 _0587_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit22.Q ),
    .Y(_0188_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit21.Q ),
    .A2(_0187_));
 sg13g2_nor2_1 _0588_ (.A(_0185_),
    .B(_0188_),
    .Y(_0189_));
 sg13g2_mux4_1 _0589_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit20.Q ),
    .A0(W2END[1]),
    .A1(UIO_OUT_TT_PROJECT1),
    .A2(UIO_OUT_TT_PROJECT5),
    .A3(UIO_OUT_TT_PROJECT6),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit21.Q ),
    .X(_0190_));
 sg13g2_nor2_1 _0590_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit22.Q ),
    .B(_0190_),
    .Y(_0191_));
 sg13g2_nor2_1 _0591_ (.A(_0189_),
    .B(_0191_),
    .Y(\Inst_W_TT_IF_switch_matrix.E2BEGb6 ));
 sg13g2_o21ai_1 _0592_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit18.Q ),
    .Y(_0192_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit17.Q ),
    .A2(_0096_));
 sg13g2_a21oi_1 _0593_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit17.Q ),
    .A2(_0071_),
    .Y(_0193_),
    .B1(_0192_));
 sg13g2_nor2b_1 _0594_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit17.Q ),
    .B_N(UIO_OE_TT_PROJECT5),
    .Y(_0194_));
 sg13g2_a21oi_1 _0595_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit17.Q ),
    .A2(_0069_),
    .Y(_0195_),
    .B1(_0194_));
 sg13g2_o21ai_1 _0596_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit19.Q ),
    .Y(_0196_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit18.Q ),
    .A2(_0195_));
 sg13g2_nor2_1 _0597_ (.A(_0193_),
    .B(_0196_),
    .Y(_0197_));
 sg13g2_mux4_1 _0598_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit18.Q ),
    .A0(W2END[2]),
    .A1(UIO_OUT_TT_PROJECT5),
    .A2(UIO_OUT_TT_PROJECT2),
    .A3(UIO_OUT_TT_PROJECT6),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit17.Q ),
    .X(_0198_));
 sg13g2_nor2_1 _0599_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit19.Q ),
    .B(_0198_),
    .Y(_0199_));
 sg13g2_nor2_1 _0600_ (.A(_0197_),
    .B(_0199_),
    .Y(\Inst_W_TT_IF_switch_matrix.E2BEGb5 ));
 sg13g2_o21ai_1 _0601_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit15.Q ),
    .Y(_0200_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit14.Q ),
    .A2(_0088_));
 sg13g2_a21oi_1 _0602_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit14.Q ),
    .A2(_0080_),
    .Y(_0201_),
    .B1(_0200_));
 sg13g2_nor2b_1 _0603_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit14.Q ),
    .B_N(UIO_OE_TT_PROJECT4),
    .Y(_0202_));
 sg13g2_a21oi_1 _0604_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit14.Q ),
    .A2(_0078_),
    .Y(_0203_),
    .B1(_0202_));
 sg13g2_o21ai_1 _0605_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit16.Q ),
    .Y(_0204_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit15.Q ),
    .A2(_0203_));
 sg13g2_nor2_1 _0606_ (.A(_0201_),
    .B(_0204_),
    .Y(_0205_));
 sg13g2_mux4_1 _0607_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit15.Q ),
    .A0(W2END[3]),
    .A1(UIO_OUT_TT_PROJECT4),
    .A2(UIO_OUT_TT_PROJECT3),
    .A3(UIO_OUT_TT_PROJECT7),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit14.Q ),
    .X(_0206_));
 sg13g2_nor2_1 _0608_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit16.Q ),
    .B(_0206_),
    .Y(_0207_));
 sg13g2_nor2_1 _0609_ (.A(_0205_),
    .B(_0207_),
    .Y(\Inst_W_TT_IF_switch_matrix.E2BEGb4 ));
 sg13g2_o21ai_1 _0610_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit12.Q ),
    .Y(_0208_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit11.Q ),
    .A2(_0088_));
 sg13g2_a21oi_1 _0611_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit11.Q ),
    .A2(_0080_),
    .Y(_0209_),
    .B1(_0208_));
 sg13g2_nor2b_1 _0612_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit11.Q ),
    .B_N(UIO_OE_TT_PROJECT3),
    .Y(_0210_));
 sg13g2_a21oi_1 _0613_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit11.Q ),
    .A2(_0087_),
    .Y(_0211_),
    .B1(_0210_));
 sg13g2_o21ai_1 _0614_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit13.Q ),
    .Y(_0212_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit12.Q ),
    .A2(_0211_));
 sg13g2_nor2_1 _0615_ (.A(_0209_),
    .B(_0212_),
    .Y(_0213_));
 sg13g2_mux4_1 _0616_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit11.Q ),
    .A0(W2END[4]),
    .A1(UIO_OUT_TT_PROJECT0),
    .A2(UIO_OUT_TT_PROJECT3),
    .A3(UIO_OUT_TT_PROJECT4),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit12.Q ),
    .X(_0214_));
 sg13g2_nor2_1 _0617_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit13.Q ),
    .B(_0214_),
    .Y(_0215_));
 sg13g2_nor2_1 _0618_ (.A(_0213_),
    .B(_0215_),
    .Y(\Inst_W_TT_IF_switch_matrix.E2BEGb3 ));
 sg13g2_o21ai_1 _0619_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit9.Q ),
    .Y(_0216_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit8.Q ),
    .A2(_0096_));
 sg13g2_a21oi_1 _0620_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit8.Q ),
    .A2(_0071_),
    .Y(_0217_),
    .B1(_0216_));
 sg13g2_nor2b_1 _0621_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit8.Q ),
    .B_N(UIO_OE_TT_PROJECT2),
    .Y(_0218_));
 sg13g2_a21oi_1 _0622_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit8.Q ),
    .A2(_0095_),
    .Y(_0219_),
    .B1(_0218_));
 sg13g2_o21ai_1 _0623_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit10.Q ),
    .Y(_0220_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit9.Q ),
    .A2(_0219_));
 sg13g2_nor2_1 _0624_ (.A(_0217_),
    .B(_0220_),
    .Y(_0221_));
 sg13g2_mux4_1 _0625_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit8.Q ),
    .A0(W2END[5]),
    .A1(UIO_OUT_TT_PROJECT1),
    .A2(UIO_OUT_TT_PROJECT2),
    .A3(UIO_OUT_TT_PROJECT5),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit9.Q ),
    .X(_0222_));
 sg13g2_nor2_1 _0626_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit10.Q ),
    .B(_0222_),
    .Y(_0223_));
 sg13g2_nor2_1 _0627_ (.A(_0221_),
    .B(_0223_),
    .Y(\Inst_W_TT_IF_switch_matrix.E2BEGb2 ));
 sg13g2_o21ai_1 _0628_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit6.Q ),
    .Y(_0224_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit5.Q ),
    .A2(_0104_));
 sg13g2_a21oi_1 _0629_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit5.Q ),
    .A2(_0062_),
    .Y(_0225_),
    .B1(_0224_));
 sg13g2_nor2b_1 _0630_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit5.Q ),
    .B_N(UIO_OE_TT_PROJECT1),
    .Y(_0226_));
 sg13g2_a21oi_1 _0631_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit5.Q ),
    .A2(_0103_),
    .Y(_0227_),
    .B1(_0226_));
 sg13g2_o21ai_1 _0632_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit7.Q ),
    .Y(_0228_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit6.Q ),
    .A2(_0227_));
 sg13g2_nor2_1 _0633_ (.A(_0225_),
    .B(_0228_),
    .Y(_0229_));
 sg13g2_mux4_1 _0634_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit5.Q ),
    .A0(W2END[6]),
    .A1(UIO_OUT_TT_PROJECT1),
    .A2(UIO_OUT_TT_PROJECT2),
    .A3(UIO_OUT_TT_PROJECT6),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit6.Q ),
    .X(_0230_));
 sg13g2_nor2_1 _0635_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit7.Q ),
    .B(_0230_),
    .Y(_0231_));
 sg13g2_nor2_1 _0636_ (.A(_0229_),
    .B(_0231_),
    .Y(\Inst_W_TT_IF_switch_matrix.E2BEGb1 ));
 sg13g2_o21ai_1 _0637_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit3.Q ),
    .Y(_0232_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit2.Q ),
    .A2(_0112_));
 sg13g2_a21oi_1 _0638_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit2.Q ),
    .A2(_0053_),
    .Y(_0233_),
    .B1(_0232_));
 sg13g2_nor2b_1 _0639_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit2.Q ),
    .B_N(UIO_OE_TT_PROJECT0),
    .Y(_0234_));
 sg13g2_a21oi_1 _0640_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit2.Q ),
    .A2(_0111_),
    .Y(_0235_),
    .B1(_0234_));
 sg13g2_o21ai_1 _0641_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit4.Q ),
    .Y(_0236_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit3.Q ),
    .A2(_0235_));
 sg13g2_nor2_1 _0642_ (.A(_0233_),
    .B(_0236_),
    .Y(_0237_));
 sg13g2_mux4_1 _0643_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit2.Q ),
    .A0(W2END[7]),
    .A1(UIO_OUT_TT_PROJECT0),
    .A2(UIO_OUT_TT_PROJECT3),
    .A3(UIO_OUT_TT_PROJECT7),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit3.Q ),
    .X(_0238_));
 sg13g2_nor2_1 _0644_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit4.Q ),
    .B(_0238_),
    .Y(_0239_));
 sg13g2_nor2_1 _0645_ (.A(_0237_),
    .B(_0239_),
    .Y(\Inst_W_TT_IF_switch_matrix.E2BEGb0 ));
 sg13g2_nor3_1 _0646_ (.A(N1END[0]),
    .B(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit24.Q ),
    .C(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit25.Q ),
    .Y(_0240_));
 sg13g2_nand2b_1 _0647_ (.Y(_0241_),
    .B(W6END[0]),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit25.Q ));
 sg13g2_a221oi_1 _0648_ (.B2(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit24.Q ),
    .C1(_0240_),
    .B1(_0241_),
    .A1(_0009_),
    .Y(_0242_),
    .A2(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit25.Q ));
 sg13g2_mux4_1 _0649_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit31.Q ),
    .A0(_0120_),
    .A1(_0112_),
    .A2(_0052_),
    .A3(_0242_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit0.Q ),
    .X(_0243_));
 sg13g2_mux4_1 _0650_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit31.Q ),
    .A0(UO_OUT_TT_PROJECT4),
    .A1(UO_OUT_TT_PROJECT7),
    .A2(UIO_OUT_TT_PROJECT7),
    .A3(UIO_OE_TT_PROJECT0),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit0.Q ),
    .X(_0244_));
 sg13g2_mux2_1 _0651_ (.A0(_0244_),
    .A1(_0243_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit1.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E2BEG7 ));
 sg13g2_nand2b_1 _0652_ (.Y(_0245_),
    .B(_0127_),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit28.Q ));
 sg13g2_nand2_1 _0653_ (.Y(_0246_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit28.Q ),
    .B(_0104_));
 sg13g2_a21oi_1 _0654_ (.A1(_0245_),
    .A2(_0246_),
    .Y(_0247_),
    .B1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit29.Q ));
 sg13g2_nor3_1 _0655_ (.A(N1END[1]),
    .B(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit26.Q ),
    .C(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit27.Q ),
    .Y(_0248_));
 sg13g2_nand2b_1 _0656_ (.Y(_0249_),
    .B(W6END[1]),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit27.Q ));
 sg13g2_a221oi_1 _0657_ (.B2(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit26.Q ),
    .C1(_0248_),
    .B1(_0249_),
    .A1(_0007_),
    .Y(_0250_),
    .A2(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit27.Q ));
 sg13g2_inv_1 _0658_ (.Y(_0251_),
    .A(_0250_));
 sg13g2_o21ai_1 _0659_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit29.Q ),
    .Y(_0252_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit28.Q ),
    .A2(_0061_));
 sg13g2_a21o_1 _0660_ (.A2(_0251_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit28.Q ),
    .B1(_0252_),
    .X(_0253_));
 sg13g2_nor2b_1 _0661_ (.A(_0247_),
    .B_N(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit30.Q ),
    .Y(_0254_));
 sg13g2_a21oi_1 _0662_ (.A1(_0023_),
    .A2(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit28.Q ),
    .Y(_0255_),
    .B1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit29.Q ));
 sg13g2_o21ai_1 _0663_ (.B1(_0255_),
    .Y(_0256_),
    .A1(UO_OUT_TT_PROJECT5),
    .A2(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit28.Q ));
 sg13g2_mux2_1 _0664_ (.A0(UIO_OUT_TT_PROJECT6),
    .A1(UIO_OE_TT_PROJECT1),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit28.Q ),
    .X(_0257_));
 sg13g2_a21oi_1 _0665_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit29.Q ),
    .A2(_0257_),
    .Y(_0258_),
    .B1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit30.Q ));
 sg13g2_a22oi_1 _0666_ (.Y(\Inst_W_TT_IF_switch_matrix.E2BEG6 ),
    .B1(_0256_),
    .B2(_0258_),
    .A2(_0254_),
    .A1(_0253_));
 sg13g2_mux2_1 _0667_ (.A0(_0134_),
    .A1(_0096_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit25.Q ),
    .X(_0259_));
 sg13g2_nand2b_1 _0668_ (.Y(_0260_),
    .B(_0259_),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit26.Q ));
 sg13g2_nand2b_1 _0669_ (.Y(_0261_),
    .B(W6END[2]),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit29.Q ));
 sg13g2_nor3_1 _0670_ (.A(N1END[2]),
    .B(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit28.Q ),
    .C(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit29.Q ),
    .Y(_0262_));
 sg13g2_a221oi_1 _0671_ (.B2(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit28.Q ),
    .C1(_0262_),
    .B1(_0261_),
    .A1(_0005_),
    .Y(_0263_),
    .A2(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit29.Q ));
 sg13g2_mux2_1 _0672_ (.A0(_0070_),
    .A1(_0263_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit25.Q ),
    .X(_0264_));
 sg13g2_a21oi_1 _0673_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit26.Q ),
    .A2(_0264_),
    .Y(_0265_),
    .B1(_0024_));
 sg13g2_a21oi_1 _0674_ (.A1(_0023_),
    .A2(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit25.Q ),
    .Y(_0266_),
    .B1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit26.Q ));
 sg13g2_o21ai_1 _0675_ (.B1(_0266_),
    .Y(_0267_),
    .A1(UO_OUT_TT_PROJECT5),
    .A2(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit25.Q ));
 sg13g2_mux2_1 _0676_ (.A0(UIO_OUT_TT_PROJECT5),
    .A1(UIO_OE_TT_PROJECT2),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit25.Q ),
    .X(_0268_));
 sg13g2_a21oi_1 _0677_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit26.Q ),
    .A2(_0268_),
    .Y(_0269_),
    .B1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit27.Q ));
 sg13g2_a22oi_1 _0678_ (.Y(\Inst_W_TT_IF_switch_matrix.E2BEG5 ),
    .B1(_0267_),
    .B2(_0269_),
    .A2(_0265_),
    .A1(_0260_));
 sg13g2_mux2_1 _0679_ (.A0(_0141_),
    .A1(_0088_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit22.Q ),
    .X(_0270_));
 sg13g2_nand2b_1 _0680_ (.Y(_0271_),
    .B(_0270_),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit23.Q ));
 sg13g2_nand2b_1 _0681_ (.Y(_0272_),
    .B(W6END[3]),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit31.Q ));
 sg13g2_nor3_1 _0682_ (.A(N1END[3]),
    .B(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit30.Q ),
    .C(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit31.Q ),
    .Y(_0273_));
 sg13g2_a221oi_1 _0683_ (.B2(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit30.Q ),
    .C1(_0273_),
    .B1(_0272_),
    .A1(_0002_),
    .Y(_0274_),
    .A2(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit31.Q ));
 sg13g2_mux2_1 _0684_ (.A0(_0079_),
    .A1(_0274_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit22.Q ),
    .X(_0275_));
 sg13g2_a21oi_1 _0685_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit23.Q ),
    .A2(_0275_),
    .Y(_0276_),
    .B1(_0025_));
 sg13g2_a21oi_1 _0686_ (.A1(_0022_),
    .A2(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit22.Q ),
    .Y(_0277_),
    .B1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit23.Q ));
 sg13g2_o21ai_1 _0687_ (.B1(_0277_),
    .Y(_0278_),
    .A1(UO_OUT_TT_PROJECT4),
    .A2(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit22.Q ));
 sg13g2_mux2_1 _0688_ (.A0(UIO_OUT_TT_PROJECT4),
    .A1(UIO_OE_TT_PROJECT3),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit22.Q ),
    .X(_0279_));
 sg13g2_a21oi_1 _0689_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit23.Q ),
    .A2(_0279_),
    .Y(_0280_),
    .B1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit24.Q ));
 sg13g2_a22oi_1 _0690_ (.Y(\Inst_W_TT_IF_switch_matrix.E2BEG4 ),
    .B1(_0278_),
    .B2(_0280_),
    .A2(_0276_),
    .A1(_0271_));
 sg13g2_mux2_1 _0691_ (.A0(_0079_),
    .A1(_0274_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit19.Q ),
    .X(_0281_));
 sg13g2_mux2_1 _0692_ (.A0(_0148_),
    .A1(_0088_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit19.Q ),
    .X(_0282_));
 sg13g2_nand2b_1 _0693_ (.Y(_0283_),
    .B(_0282_),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit20.Q ));
 sg13g2_a21oi_1 _0694_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit20.Q ),
    .A2(_0281_),
    .Y(_0284_),
    .B1(_0027_));
 sg13g2_a21oi_1 _0695_ (.A1(_0026_),
    .A2(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit19.Q ),
    .Y(_0285_),
    .B1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit20.Q ));
 sg13g2_o21ai_1 _0696_ (.B1(_0285_),
    .Y(_0286_),
    .A1(UO_OUT_TT_PROJECT0),
    .A2(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit19.Q ));
 sg13g2_mux2_1 _0697_ (.A0(UIO_OUT_TT_PROJECT3),
    .A1(UIO_OE_TT_PROJECT4),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit19.Q ),
    .X(_0287_));
 sg13g2_a21oi_1 _0698_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit20.Q ),
    .A2(_0287_),
    .Y(_0288_),
    .B1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit21.Q ));
 sg13g2_a22oi_1 _0699_ (.Y(\Inst_W_TT_IF_switch_matrix.E2BEG3 ),
    .B1(_0286_),
    .B2(_0288_),
    .A2(_0284_),
    .A1(_0283_));
 sg13g2_mux2_1 _0700_ (.A0(_0070_),
    .A1(_0263_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit16.Q ),
    .X(_0289_));
 sg13g2_mux2_1 _0701_ (.A0(_0155_),
    .A1(_0096_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit16.Q ),
    .X(_0290_));
 sg13g2_nand2b_1 _0702_ (.Y(_0291_),
    .B(_0290_),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit17.Q ));
 sg13g2_a21oi_1 _0703_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit17.Q ),
    .A2(_0289_),
    .Y(_0292_),
    .B1(_0029_));
 sg13g2_a21oi_1 _0704_ (.A1(_0028_),
    .A2(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit16.Q ),
    .Y(_0293_),
    .B1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit17.Q ));
 sg13g2_o21ai_1 _0705_ (.B1(_0293_),
    .Y(_0294_),
    .A1(UO_OUT_TT_PROJECT1),
    .A2(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit16.Q ));
 sg13g2_mux2_1 _0706_ (.A0(UIO_OUT_TT_PROJECT2),
    .A1(UIO_OE_TT_PROJECT5),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit16.Q ),
    .X(_0295_));
 sg13g2_a21oi_1 _0707_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit17.Q ),
    .A2(_0295_),
    .Y(_0296_),
    .B1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit18.Q ));
 sg13g2_a22oi_1 _0708_ (.Y(\Inst_W_TT_IF_switch_matrix.E2BEG2 ),
    .B1(_0294_),
    .B2(_0296_),
    .A2(_0292_),
    .A1(_0291_));
 sg13g2_o21ai_1 _0709_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit14.Q ),
    .Y(_0297_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit13.Q ),
    .A2(_0061_));
 sg13g2_a21o_1 _0710_ (.A2(_0251_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit13.Q ),
    .B1(_0297_),
    .X(_0298_));
 sg13g2_nand2b_1 _0711_ (.Y(_0299_),
    .B(_0162_),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit13.Q ));
 sg13g2_nand2_1 _0712_ (.Y(_0300_),
    .A(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit13.Q ),
    .B(_0104_));
 sg13g2_a21oi_1 _0713_ (.A1(_0299_),
    .A2(_0300_),
    .Y(_0301_),
    .B1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit14.Q ));
 sg13g2_nor2b_1 _0714_ (.A(_0301_),
    .B_N(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit15.Q ),
    .Y(_0302_));
 sg13g2_a21oi_1 _0715_ (.A1(_0028_),
    .A2(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit13.Q ),
    .Y(_0303_),
    .B1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit14.Q ));
 sg13g2_o21ai_1 _0716_ (.B1(_0303_),
    .Y(_0304_),
    .A1(UO_OUT_TT_PROJECT1),
    .A2(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit13.Q ));
 sg13g2_mux2_1 _0717_ (.A0(UIO_OUT_TT_PROJECT1),
    .A1(UIO_OE_TT_PROJECT6),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit13.Q ),
    .X(_0305_));
 sg13g2_a21oi_1 _0718_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit14.Q ),
    .A2(_0305_),
    .Y(_0306_),
    .B1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit15.Q ));
 sg13g2_a22oi_1 _0719_ (.Y(\Inst_W_TT_IF_switch_matrix.E2BEG1 ),
    .B1(_0304_),
    .B2(_0306_),
    .A2(_0302_),
    .A1(_0298_));
 sg13g2_nor2_1 _0720_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit10.Q ),
    .B(_0169_),
    .Y(_0307_));
 sg13g2_nor2_1 _0721_ (.A(_0030_),
    .B(_0112_),
    .Y(_0308_));
 sg13g2_nor3_1 _0722_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit11.Q ),
    .B(_0307_),
    .C(_0308_),
    .Y(_0309_));
 sg13g2_o21ai_1 _0723_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit11.Q ),
    .Y(_0310_),
    .A1(_0030_),
    .A2(_0242_));
 sg13g2_a21o_1 _0724_ (.A2(_0053_),
    .A1(_0030_),
    .B1(_0310_),
    .X(_0311_));
 sg13g2_nor2b_1 _0725_ (.A(_0309_),
    .B_N(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit12.Q ),
    .Y(_0312_));
 sg13g2_a21oi_1 _0726_ (.A1(_0026_),
    .A2(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit10.Q ),
    .Y(_0313_),
    .B1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit11.Q ));
 sg13g2_o21ai_1 _0727_ (.B1(_0313_),
    .Y(_0314_),
    .A1(UO_OUT_TT_PROJECT0),
    .A2(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit10.Q ));
 sg13g2_mux2_1 _0728_ (.A0(UIO_OUT_TT_PROJECT0),
    .A1(UIO_OE_TT_PROJECT7),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit10.Q ),
    .X(_0315_));
 sg13g2_a21oi_1 _0729_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit11.Q ),
    .A2(_0315_),
    .Y(_0316_),
    .B1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit12.Q ));
 sg13g2_a22oi_1 _0730_ (.Y(\Inst_W_TT_IF_switch_matrix.E2BEG0 ),
    .B1(_0314_),
    .B2(_0316_),
    .A2(_0312_),
    .A1(_0311_));
 sg13g2_mux4_1 _0731_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit7.Q ),
    .A0(UIO_OE_TT_PROJECT1),
    .A1(UIO_OE_TT_PROJECT3),
    .A2(UIO_OE_TT_PROJECT4),
    .A3(UIO_OE_TT_PROJECT7),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit8.Q ),
    .X(_0317_));
 sg13g2_mux4_1 _0732_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit7.Q ),
    .A0(N1END[3]),
    .A1(S1END[3]),
    .A2(UO_OUT_TT_PROJECT1),
    .A3(UO_OUT_TT_PROJECT4),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit8.Q ),
    .X(_0318_));
 sg13g2_mux2_1 _0733_ (.A0(_0318_),
    .A1(_0317_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit9.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E1BEG3 ));
 sg13g2_mux4_1 _0734_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit4.Q ),
    .A0(UIO_OE_TT_PROJECT2),
    .A1(UIO_OE_TT_PROJECT3),
    .A2(UIO_OE_TT_PROJECT4),
    .A3(UIO_OE_TT_PROJECT5),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit5.Q ),
    .X(_0319_));
 sg13g2_mux4_1 _0735_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit4.Q ),
    .A0(N1END[2]),
    .A1(S1END[2]),
    .A2(UO_OUT_TT_PROJECT0),
    .A3(UO_OUT_TT_PROJECT5),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit5.Q ),
    .X(_0320_));
 sg13g2_mux2_1 _0736_ (.A0(_0320_),
    .A1(_0319_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit6.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E1BEG2 ));
 sg13g2_mux4_1 _0737_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit1.Q ),
    .A0(UIO_OE_TT_PROJECT0),
    .A1(UIO_OE_TT_PROJECT1),
    .A2(UIO_OE_TT_PROJECT5),
    .A3(UIO_OE_TT_PROJECT6),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit2.Q ),
    .X(_0321_));
 sg13g2_mux4_1 _0738_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit1.Q ),
    .A0(N1END[1]),
    .A1(S1END[1]),
    .A2(UO_OUT_TT_PROJECT3),
    .A3(UO_OUT_TT_PROJECT6),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit2.Q ),
    .X(_0322_));
 sg13g2_mux2_1 _0739_ (.A0(_0322_),
    .A1(_0321_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit3.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E1BEG1 ));
 sg13g2_mux4_1 _0740_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit30.Q ),
    .A0(UIO_OE_TT_PROJECT0),
    .A1(UIO_OE_TT_PROJECT2),
    .A2(UIO_OE_TT_PROJECT6),
    .A3(UIO_OE_TT_PROJECT7),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit31.Q ),
    .X(_0323_));
 sg13g2_mux4_1 _0741_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit30.Q ),
    .A0(N1END[0]),
    .A1(S1END[0]),
    .A2(UO_OUT_TT_PROJECT2),
    .A3(UO_OUT_TT_PROJECT7),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit31.Q ),
    .X(_0324_));
 sg13g2_mux2_1 _0742_ (.A0(_0324_),
    .A1(_0323_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit0.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E1BEG0 ));
 sg13g2_o21ai_1 _0743_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit27.Q ),
    .Y(_0325_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit29.Q ),
    .A2(_0148_));
 sg13g2_a21oi_1 _0744_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit29.Q ),
    .A2(_0053_),
    .Y(_0326_),
    .B1(_0325_));
 sg13g2_or2_1 _0745_ (.X(_0327_),
    .B(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit29.Q ),
    .A(W6END[7]));
 sg13g2_o21ai_1 _0746_ (.B1(_0327_),
    .Y(_0328_),
    .A1(_0031_),
    .A2(_0051_));
 sg13g2_o21ai_1 _0747_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit28.Q ),
    .Y(_0329_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit27.Q ),
    .A2(_0328_));
 sg13g2_nor2_1 _0748_ (.A(_0326_),
    .B(_0329_),
    .Y(_0330_));
 sg13g2_a21oi_1 _0749_ (.A1(_0001_),
    .A2(_0031_),
    .Y(_0331_),
    .B1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit27.Q ));
 sg13g2_o21ai_1 _0750_ (.B1(_0331_),
    .Y(_0332_),
    .A1(_0031_),
    .A2(_0120_));
 sg13g2_mux2_1 _0751_ (.A0(WW4END[15]),
    .A1(_0087_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit29.Q ),
    .X(_0333_));
 sg13g2_a21oi_1 _0752_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit27.Q ),
    .A2(_0333_),
    .Y(_0334_),
    .B1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit28.Q ));
 sg13g2_a21oi_1 _0753_ (.A1(_0332_),
    .A2(_0334_),
    .Y(\Inst_W_TT_IF_switch_matrix.S4BEG3 ),
    .B1(_0330_));
 sg13g2_o21ai_1 _0754_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit24.Q ),
    .Y(_0335_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit26.Q ),
    .A2(_0155_));
 sg13g2_a21oi_1 _0755_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit26.Q ),
    .A2(_0062_),
    .Y(_0336_),
    .B1(_0335_));
 sg13g2_or2_1 _0756_ (.X(_0337_),
    .B(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit26.Q ),
    .A(W6END[6]));
 sg13g2_o21ai_1 _0757_ (.B1(_0337_),
    .Y(_0338_),
    .A1(_0032_),
    .A2(_0060_));
 sg13g2_o21ai_1 _0758_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit25.Q ),
    .Y(_0339_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit24.Q ),
    .A2(_0338_));
 sg13g2_nor2_1 _0759_ (.A(_0336_),
    .B(_0339_),
    .Y(_0340_));
 sg13g2_a21oi_1 _0760_ (.A1(_0004_),
    .A2(_0032_),
    .Y(_0341_),
    .B1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit24.Q ));
 sg13g2_o21ai_1 _0761_ (.B1(_0341_),
    .Y(_0342_),
    .A1(_0032_),
    .A2(_0127_));
 sg13g2_mux2_1 _0762_ (.A0(WW4END[14]),
    .A1(_0095_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit26.Q ),
    .X(_0343_));
 sg13g2_a21oi_1 _0763_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit24.Q ),
    .A2(_0343_),
    .Y(_0344_),
    .B1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit25.Q ));
 sg13g2_a21oi_1 _0764_ (.A1(_0342_),
    .A2(_0344_),
    .Y(\Inst_W_TT_IF_switch_matrix.S4BEG2 ),
    .B1(_0340_));
 sg13g2_mux4_1 _0765_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit23.Q ),
    .A0(W6END[5]),
    .A1(_0069_),
    .A2(_0162_),
    .A3(_0070_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit21.Q ),
    .X(_0345_));
 sg13g2_mux4_1 _0766_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit21.Q ),
    .A0(W1END[1]),
    .A1(WW4END[13]),
    .A2(_0134_),
    .A3(_0103_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit23.Q ),
    .X(_0346_));
 sg13g2_mux2_1 _0767_ (.A0(_0346_),
    .A1(_0345_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit22.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.S4BEG1 ));
 sg13g2_mux4_1 _0768_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit20.Q ),
    .A0(W6END[4]),
    .A1(_0078_),
    .A2(_0169_),
    .A3(_0079_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit18.Q ),
    .X(_0347_));
 sg13g2_mux4_1 _0769_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit18.Q ),
    .A0(W1END[0]),
    .A1(WW4END[12]),
    .A2(_0141_),
    .A3(_0111_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit20.Q ),
    .X(_0348_));
 sg13g2_mux2_1 _0770_ (.A0(_0348_),
    .A1(_0347_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit19.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.S4BEG0 ));
 sg13g2_mux2_1 _0771_ (.A0(_0088_),
    .A1(_0148_),
    .S(_0033_),
    .X(_0349_));
 sg13g2_or2_1 _0772_ (.X(_0350_),
    .B(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit25.Q ),
    .A(W6END[11]));
 sg13g2_o21ai_1 _0773_ (.B1(_0350_),
    .Y(_0351_),
    .A1(_0033_),
    .A2(_0051_));
 sg13g2_o21ai_1 _0774_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit24.Q ),
    .Y(_0352_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit23.Q ),
    .A2(_0351_));
 sg13g2_a21oi_1 _0775_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit23.Q ),
    .A2(_0349_),
    .Y(_0353_),
    .B1(_0352_));
 sg13g2_mux4_1 _0776_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit23.Q ),
    .A0(W1END[3]),
    .A1(WW4END[3]),
    .A2(_0120_),
    .A3(_0087_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit25.Q ),
    .X(_0354_));
 sg13g2_nor2_1 _0777_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit24.Q ),
    .B(_0354_),
    .Y(_0355_));
 sg13g2_nor2_1 _0778_ (.A(_0353_),
    .B(_0355_),
    .Y(\Inst_W_TT_IF_switch_matrix.N4BEG3 ));
 sg13g2_mux2_1 _0779_ (.A0(_0096_),
    .A1(_0155_),
    .S(_0034_),
    .X(_0356_));
 sg13g2_or2_1 _0780_ (.X(_0357_),
    .B(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit22.Q ),
    .A(W6END[10]));
 sg13g2_o21ai_1 _0781_ (.B1(_0357_),
    .Y(_0358_),
    .A1(_0034_),
    .A2(_0060_));
 sg13g2_o21ai_1 _0782_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit21.Q ),
    .Y(_0359_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit20.Q ),
    .A2(_0358_));
 sg13g2_a21oi_1 _0783_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit20.Q ),
    .A2(_0356_),
    .Y(_0360_),
    .B1(_0359_));
 sg13g2_a21oi_1 _0784_ (.A1(_0004_),
    .A2(_0034_),
    .Y(_0361_),
    .B1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit20.Q ));
 sg13g2_o21ai_1 _0785_ (.B1(_0361_),
    .Y(_0362_),
    .A1(_0034_),
    .A2(_0127_));
 sg13g2_mux2_1 _0786_ (.A0(WW4END[2]),
    .A1(_0095_),
    .S(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit22.Q ),
    .X(_0363_));
 sg13g2_a21oi_1 _0787_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit20.Q ),
    .A2(_0363_),
    .Y(_0364_),
    .B1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit21.Q ));
 sg13g2_a21oi_1 _0788_ (.A1(_0362_),
    .A2(_0364_),
    .Y(\Inst_W_TT_IF_switch_matrix.N4BEG2 ),
    .B1(_0360_));
 sg13g2_mux2_1 _0789_ (.A0(_0104_),
    .A1(_0162_),
    .S(_0035_),
    .X(_0365_));
 sg13g2_or2_1 _0790_ (.X(_0366_),
    .B(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit19.Q ),
    .A(W6END[9]));
 sg13g2_o21ai_1 _0791_ (.B1(_0366_),
    .Y(_0367_),
    .A1(_0035_),
    .A2(_0069_));
 sg13g2_o21ai_1 _0792_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit18.Q ),
    .Y(_0368_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit17.Q ),
    .A2(_0367_));
 sg13g2_a21oi_1 _0793_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit17.Q ),
    .A2(_0365_),
    .Y(_0369_),
    .B1(_0368_));
 sg13g2_mux4_1 _0794_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit17.Q ),
    .A0(W1END[1]),
    .A1(WW4END[1]),
    .A2(_0134_),
    .A3(_0103_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit19.Q ),
    .X(_0370_));
 sg13g2_nor2_1 _0795_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit18.Q ),
    .B(_0370_),
    .Y(_0371_));
 sg13g2_nor2_1 _0796_ (.A(_0369_),
    .B(_0371_),
    .Y(\Inst_W_TT_IF_switch_matrix.N4BEG1 ));
 sg13g2_mux2_1 _0797_ (.A0(_0112_),
    .A1(_0169_),
    .S(_0036_),
    .X(_0372_));
 sg13g2_or2_1 _0798_ (.X(_0373_),
    .B(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit16.Q ),
    .A(W6END[8]));
 sg13g2_o21ai_1 _0799_ (.B1(_0373_),
    .Y(_0374_),
    .A1(_0036_),
    .A2(_0078_));
 sg13g2_o21ai_1 _0800_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit15.Q ),
    .Y(_0375_),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit14.Q ),
    .A2(_0374_));
 sg13g2_a21oi_1 _0801_ (.A1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit14.Q ),
    .A2(_0372_),
    .Y(_0376_),
    .B1(_0375_));
 sg13g2_mux4_1 _0802_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit14.Q ),
    .A0(W1END[0]),
    .A1(WW4END[0]),
    .A2(_0141_),
    .A3(_0111_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit16.Q ),
    .X(_0377_));
 sg13g2_nor2_1 _0803_ (.A(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit15.Q ),
    .B(_0377_),
    .Y(_0378_));
 sg13g2_nor2_1 _0804_ (.A(_0376_),
    .B(_0378_),
    .Y(\Inst_W_TT_IF_switch_matrix.N4BEG0 ));
 sg13g2_o21ai_1 _0805_ (.B1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit2.Q ),
    .Y(_0379_),
    .A1(W2MID[6]),
    .A2(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit3.Q ));
 sg13g2_nand2b_1 _0806_ (.Y(_0380_),
    .B(N2MID[6]),
    .A_N(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit2.Q ));
 sg13g2_o21ai_1 _0807_ (.B1(_0379_),
    .Y(ENA_TT_PROJECT),
    .A1(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit3.Q ),
    .A2(_0380_));
 sg13g2_mux4_1 _0808_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit17.Q ),
    .A0(UIO_OUT_TT_PROJECT3),
    .A1(_0141_),
    .A2(_0169_),
    .A3(_0052_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit16.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E6BEG11 ));
 sg13g2_mux4_1 _0809_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit15.Q ),
    .A0(UIO_OUT_TT_PROJECT2),
    .A1(_0134_),
    .A2(_0162_),
    .A3(_0061_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit14.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E6BEG10 ));
 sg13g2_mux4_1 _0810_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit13.Q ),
    .A0(UIO_OUT_TT_PROJECT1),
    .A1(_0127_),
    .A2(_0155_),
    .A3(_0070_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit12.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E6BEG9 ));
 sg13g2_mux4_1 _0811_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit11.Q ),
    .A0(UIO_OUT_TT_PROJECT0),
    .A1(_0120_),
    .A2(_0148_),
    .A3(_0079_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit10.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E6BEG8 ));
 sg13g2_mux4_1 _0812_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit9.Q ),
    .A0(UIO_OUT_TT_PROJECT7),
    .A1(_0111_),
    .A2(_0141_),
    .A3(_0088_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit8.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E6BEG7 ));
 sg13g2_mux4_1 _0813_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit7.Q ),
    .A0(UIO_OUT_TT_PROJECT6),
    .A1(_0103_),
    .A2(_0134_),
    .A3(_0096_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit6.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E6BEG6 ));
 sg13g2_mux4_1 _0814_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit5.Q ),
    .A0(UIO_OUT_TT_PROJECT5),
    .A1(_0095_),
    .A2(_0127_),
    .A3(_0104_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit4.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E6BEG5 ));
 sg13g2_mux4_1 _0815_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit3.Q ),
    .A0(UIO_OUT_TT_PROJECT4),
    .A1(_0087_),
    .A2(_0120_),
    .A3(_0112_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit2.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E6BEG4 ));
 sg13g2_mux4_1 _0816_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit0.Q ),
    .A0(N4END[3]),
    .A1(S4END[3]),
    .A2(_0111_),
    .A3(_0078_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit1.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E6BEG3 ));
 sg13g2_mux4_1 _0817_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit30.Q ),
    .A0(N4END[2]),
    .A1(S4END[2]),
    .A2(_0103_),
    .A3(_0069_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit31.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E6BEG2 ));
 sg13g2_mux4_1 _0818_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit28.Q ),
    .A0(N4END[1]),
    .A1(S4END[1]),
    .A2(_0095_),
    .A3(_0060_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit29.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E6BEG1 ));
 sg13g2_mux4_1 _0819_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit26.Q ),
    .A0(N4END[0]),
    .A1(S4END[0]),
    .A2(_0087_),
    .A3(_0051_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit27.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.E6BEG0 ));
 sg13g2_mux4_1 _0820_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit25.Q ),
    .A0(UO_OUT_TT_PROJECT3),
    .A1(_0169_),
    .A2(UIO_OUT_TT_PROJECT7),
    .A3(_0112_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit24.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG15 ));
 sg13g2_mux4_1 _0821_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit23.Q ),
    .A0(UO_OUT_TT_PROJECT2),
    .A1(_0162_),
    .A2(UIO_OUT_TT_PROJECT6),
    .A3(_0104_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit22.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG14 ));
 sg13g2_mux4_1 _0822_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit21.Q ),
    .A0(UO_OUT_TT_PROJECT1),
    .A1(_0155_),
    .A2(UIO_OUT_TT_PROJECT5),
    .A3(_0096_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit20.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG13 ));
 sg13g2_mux4_1 _0823_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit19.Q ),
    .A0(UO_OUT_TT_PROJECT0),
    .A1(_0148_),
    .A2(UIO_OUT_TT_PROJECT4),
    .A3(_0088_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit18.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG12 ));
 sg13g2_mux4_1 _0824_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit17.Q ),
    .A0(UO_OUT_TT_PROJECT7),
    .A1(_0141_),
    .A2(UIO_OUT_TT_PROJECT3),
    .A3(_0079_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit16.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG11 ));
 sg13g2_mux4_1 _0825_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit15.Q ),
    .A0(UO_OUT_TT_PROJECT6),
    .A1(_0134_),
    .A2(UIO_OUT_TT_PROJECT2),
    .A3(_0070_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit14.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG10 ));
 sg13g2_mux4_1 _0826_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit13.Q ),
    .A0(UO_OUT_TT_PROJECT5),
    .A1(_0127_),
    .A2(UIO_OUT_TT_PROJECT1),
    .A3(_0061_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit12.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG9 ));
 sg13g2_mux4_1 _0827_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit11.Q ),
    .A0(UO_OUT_TT_PROJECT4),
    .A1(_0120_),
    .A2(UIO_OUT_TT_PROJECT0),
    .A3(_0052_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit10.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG8 ));
 sg13g2_mux4_1 _0828_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit9.Q ),
    .A0(UO_OUT_TT_PROJECT7),
    .A1(_0111_),
    .A2(UIO_OE_TT_PROJECT3),
    .A3(_0112_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit8.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG7 ));
 sg13g2_mux4_1 _0829_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit7.Q ),
    .A0(UO_OUT_TT_PROJECT6),
    .A1(_0103_),
    .A2(UIO_OE_TT_PROJECT2),
    .A3(_0104_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit6.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG6 ));
 sg13g2_mux4_1 _0830_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit5.Q ),
    .A0(UO_OUT_TT_PROJECT5),
    .A1(_0095_),
    .A2(UIO_OE_TT_PROJECT1),
    .A3(_0096_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit4.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG5 ));
 sg13g2_mux4_1 _0831_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit3.Q ),
    .A0(UO_OUT_TT_PROJECT4),
    .A1(_0087_),
    .A2(UIO_OE_TT_PROJECT0),
    .A3(_0088_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit2.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG4 ));
 sg13g2_mux4_1 _0832_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit1.Q ),
    .A0(UO_OUT_TT_PROJECT3),
    .A1(_0078_),
    .A2(UIO_OE_TT_PROJECT7),
    .A3(_0079_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit0.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG3 ));
 sg13g2_mux4_1 _0833_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit31.Q ),
    .A0(UO_OUT_TT_PROJECT2),
    .A1(_0069_),
    .A2(UIO_OE_TT_PROJECT6),
    .A3(_0070_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit30.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG2 ));
 sg13g2_mux4_1 _0834_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit29.Q ),
    .A0(UO_OUT_TT_PROJECT1),
    .A1(_0060_),
    .A2(UIO_OE_TT_PROJECT5),
    .A3(_0061_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit28.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG1 ));
 sg13g2_mux4_1 _0835_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit27.Q ),
    .A0(UO_OUT_TT_PROJECT0),
    .A1(_0051_),
    .A2(UIO_OE_TT_PROJECT4),
    .A3(_0052_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit26.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.EE4BEG0 ));
 sg13g2_mux4_1 _0836_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit17.Q ),
    .A0(W1END[3]),
    .A1(W2END[0]),
    .A2(W2MID[0]),
    .A3(_0052_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit16.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.S2BEG7 ));
 sg13g2_mux4_1 _0837_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit14.Q ),
    .A0(W1END[2]),
    .A1(W2MID[1]),
    .A2(W2END[1]),
    .A3(_0061_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit15.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.S2BEG6 ));
 sg13g2_mux4_1 _0838_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit12.Q ),
    .A0(W1END[1]),
    .A1(W2MID[2]),
    .A2(W2END[2]),
    .A3(_0070_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit13.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.S2BEG5 ));
 sg13g2_mux4_1 _0839_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit11.Q ),
    .A0(W1END[0]),
    .A1(W2END[3]),
    .A2(W2MID[3]),
    .A3(_0079_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit10.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.S2BEG4 ));
 sg13g2_mux4_1 _0840_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit9.Q ),
    .A0(W2MID[4]),
    .A1(W6END[11]),
    .A2(W2END[4]),
    .A3(_0088_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit8.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.S2BEG3 ));
 sg13g2_mux4_1 _0841_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit7.Q ),
    .A0(W2MID[5]),
    .A1(W6END[10]),
    .A2(W2END[5]),
    .A3(_0096_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit6.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.S2BEG2 ));
 sg13g2_mux4_1 _0842_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit4.Q ),
    .A0(W2MID[6]),
    .A1(W2END[6]),
    .A2(W6END[9]),
    .A3(_0104_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit5.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.S2BEG1 ));
 sg13g2_mux4_1 _0843_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit2.Q ),
    .A0(W2MID[7]),
    .A1(W2END[7]),
    .A2(W6END[8]),
    .A3(_0112_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit3.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.S2BEG0 ));
 sg13g2_mux4_1 _0844_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit0.Q ),
    .A0(W1END[3]),
    .A1(W6END[11]),
    .A2(_0051_),
    .A3(_0274_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit1.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.S1BEG3 ));
 sg13g2_mux4_1 _0845_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit30.Q ),
    .A0(W1END[2]),
    .A1(W6END[10]),
    .A2(_0060_),
    .A3(_0263_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit31.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.S1BEG2 ));
 sg13g2_mux4_1 _0846_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit28.Q ),
    .A0(W1END[1]),
    .A1(W6END[9]),
    .A2(_0069_),
    .A3(_0250_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit29.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.S1BEG1 ));
 sg13g2_mux4_1 _0847_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit26.Q ),
    .A0(W1END[0]),
    .A1(W6END[8]),
    .A2(_0078_),
    .A3(_0242_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit27.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.S1BEG0 ));
 sg13g2_mux4_1 _0848_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit12.Q ),
    .A0(W2MID[0]),
    .A1(W2END[0]),
    .A2(W6END[0]),
    .A3(_0052_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit13.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.N2BEG7 ));
 sg13g2_mux4_1 _0849_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit11.Q ),
    .A0(W2MID[1]),
    .A1(W6END[1]),
    .A2(W2END[1]),
    .A3(_0061_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit10.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.N2BEG6 ));
 sg13g2_mux4_1 _0850_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit9.Q ),
    .A0(W2MID[2]),
    .A1(W6END[2]),
    .A2(W2END[2]),
    .A3(_0070_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit8.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.N2BEG5 ));
 sg13g2_mux4_1 _0851_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit6.Q ),
    .A0(W2MID[3]),
    .A1(W2END[3]),
    .A2(W6END[3]),
    .A3(_0079_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit7.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.N2BEG4 ));
 sg13g2_mux4_1 _0852_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit5.Q ),
    .A0(W2MID[4]),
    .A1(W6END[4]),
    .A2(W2END[4]),
    .A3(_0088_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit4.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.N2BEG3 ));
 sg13g2_mux4_1 _0853_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit3.Q ),
    .A0(W2MID[5]),
    .A1(W6END[5]),
    .A2(W2END[5]),
    .A3(_0096_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit2.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.N2BEG2 ));
 sg13g2_mux4_1 _0854_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit0.Q ),
    .A0(W2MID[6]),
    .A1(W2END[6]),
    .A2(W6END[6]),
    .A3(_0104_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit1.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.N2BEG1 ));
 sg13g2_mux4_1 _0855_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame9_bit30.Q ),
    .A0(W2MID[7]),
    .A1(W2END[7]),
    .A2(W6END[7]),
    .A3(_0112_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame9_bit31.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.N2BEG0 ));
 sg13g2_mux4_1 _0856_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame9_bit28.Q ),
    .A0(W1END[3]),
    .A1(W6END[7]),
    .A2(_0051_),
    .A3(_0274_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame9_bit29.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.N1BEG3 ));
 sg13g2_mux4_1 _0857_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame9_bit26.Q ),
    .A0(W1END[2]),
    .A1(W6END[6]),
    .A2(_0060_),
    .A3(_0263_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame9_bit27.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.N1BEG2 ));
 sg13g2_mux4_1 _0858_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame9_bit24.Q ),
    .A0(W1END[1]),
    .A1(W6END[5]),
    .A2(_0069_),
    .A3(_0250_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame9_bit25.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.N1BEG1 ));
 sg13g2_mux4_1 _0859_ (.S0(\Inst_W_TT_IF_ConfigMem.Inst_frame9_bit22.Q ),
    .A0(W1END[0]),
    .A1(W6END[4]),
    .A2(_0078_),
    .A3(_0242_),
    .S1(\Inst_W_TT_IF_ConfigMem.Inst_frame9_bit23.Q ),
    .X(\Inst_W_TT_IF_switch_matrix.N1BEG0 ));
 sg13g2_dlhq_1 _0860_ (.D(FrameData[22]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame9_bit22.Q ));
 sg13g2_dlhq_1 _0861_ (.D(FrameData[23]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame9_bit23.Q ));
 sg13g2_dlhq_1 _0862_ (.D(FrameData[24]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame9_bit24.Q ));
 sg13g2_dlhq_1 _0863_ (.D(FrameData[25]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame9_bit25.Q ));
 sg13g2_dlhq_1 _0864_ (.D(FrameData[26]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame9_bit26.Q ));
 sg13g2_dlhq_1 _0865_ (.D(FrameData[27]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame9_bit27.Q ));
 sg13g2_dlhq_1 _0866_ (.D(FrameData[28]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame9_bit28.Q ));
 sg13g2_dlhq_1 _0867_ (.D(FrameData[29]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame9_bit29.Q ));
 sg13g2_dlhq_1 _0868_ (.D(FrameData[30]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame9_bit30.Q ));
 sg13g2_dlhq_1 _0869_ (.D(FrameData[31]),
    .GATE(FrameStrobe[9]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame9_bit31.Q ));
 sg13g2_dlhq_1 _0870_ (.D(FrameData[0]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit0.Q ));
 sg13g2_dlhq_1 _0871_ (.D(FrameData[1]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit1.Q ));
 sg13g2_dlhq_1 _0872_ (.D(FrameData[2]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit2.Q ));
 sg13g2_dlhq_1 _0873_ (.D(FrameData[3]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit3.Q ));
 sg13g2_dlhq_1 _0874_ (.D(FrameData[4]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit4.Q ));
 sg13g2_dlhq_1 _0875_ (.D(FrameData[5]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit5.Q ));
 sg13g2_dlhq_1 _0876_ (.D(FrameData[6]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit6.Q ));
 sg13g2_dlhq_1 _0877_ (.D(FrameData[7]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit7.Q ));
 sg13g2_dlhq_1 _0878_ (.D(FrameData[8]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit8.Q ));
 sg13g2_dlhq_1 _0879_ (.D(FrameData[9]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit9.Q ));
 sg13g2_dlhq_1 _0880_ (.D(FrameData[10]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit10.Q ));
 sg13g2_dlhq_1 _0881_ (.D(FrameData[11]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit11.Q ));
 sg13g2_dlhq_1 _0882_ (.D(FrameData[12]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit12.Q ));
 sg13g2_dlhq_1 _0883_ (.D(FrameData[13]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit13.Q ));
 sg13g2_dlhq_1 _0884_ (.D(FrameData[14]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit14.Q ));
 sg13g2_dlhq_1 _0885_ (.D(FrameData[15]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit15.Q ));
 sg13g2_dlhq_1 _0886_ (.D(FrameData[16]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit16.Q ));
 sg13g2_dlhq_1 _0887_ (.D(FrameData[17]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit17.Q ));
 sg13g2_dlhq_1 _0888_ (.D(FrameData[18]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit18.Q ));
 sg13g2_dlhq_1 _0889_ (.D(FrameData[19]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit19.Q ));
 sg13g2_dlhq_1 _0890_ (.D(FrameData[20]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit20.Q ));
 sg13g2_dlhq_1 _0891_ (.D(FrameData[21]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit21.Q ));
 sg13g2_dlhq_1 _0892_ (.D(FrameData[22]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit22.Q ));
 sg13g2_dlhq_1 _0893_ (.D(FrameData[23]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit23.Q ));
 sg13g2_dlhq_1 _0894_ (.D(FrameData[24]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit24.Q ));
 sg13g2_dlhq_1 _0895_ (.D(FrameData[25]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit25.Q ));
 sg13g2_dlhq_1 _0896_ (.D(FrameData[26]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit26.Q ));
 sg13g2_dlhq_1 _0897_ (.D(FrameData[27]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit27.Q ));
 sg13g2_dlhq_1 _0898_ (.D(FrameData[28]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit28.Q ));
 sg13g2_dlhq_1 _0899_ (.D(FrameData[29]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit29.Q ));
 sg13g2_dlhq_1 _0900_ (.D(FrameData[30]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit30.Q ));
 sg13g2_dlhq_1 _0901_ (.D(FrameData[31]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame8_bit31.Q ));
 sg13g2_dlhq_1 _0902_ (.D(FrameData[0]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit0.Q ));
 sg13g2_dlhq_1 _0903_ (.D(FrameData[1]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit1.Q ));
 sg13g2_dlhq_1 _0904_ (.D(FrameData[2]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit2.Q ));
 sg13g2_dlhq_1 _0905_ (.D(FrameData[3]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit3.Q ));
 sg13g2_dlhq_1 _0906_ (.D(FrameData[4]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit4.Q ));
 sg13g2_dlhq_1 _0907_ (.D(FrameData[5]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit5.Q ));
 sg13g2_dlhq_1 _0908_ (.D(FrameData[6]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit6.Q ));
 sg13g2_dlhq_1 _0909_ (.D(FrameData[7]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit7.Q ));
 sg13g2_dlhq_1 _0910_ (.D(FrameData[8]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit8.Q ));
 sg13g2_dlhq_1 _0911_ (.D(FrameData[9]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit9.Q ));
 sg13g2_dlhq_1 _0912_ (.D(FrameData[10]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit10.Q ));
 sg13g2_dlhq_1 _0913_ (.D(FrameData[11]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit11.Q ));
 sg13g2_dlhq_1 _0914_ (.D(FrameData[12]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit12.Q ));
 sg13g2_dlhq_1 _0915_ (.D(FrameData[13]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit13.Q ));
 sg13g2_dlhq_1 _0916_ (.D(FrameData[14]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit14.Q ));
 sg13g2_dlhq_1 _0917_ (.D(FrameData[15]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit15.Q ));
 sg13g2_dlhq_1 _0918_ (.D(FrameData[16]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit16.Q ));
 sg13g2_dlhq_1 _0919_ (.D(FrameData[17]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit17.Q ));
 sg13g2_dlhq_1 _0920_ (.D(FrameData[18]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit18.Q ));
 sg13g2_dlhq_1 _0921_ (.D(FrameData[19]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit19.Q ));
 sg13g2_dlhq_1 _0922_ (.D(FrameData[20]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit20.Q ));
 sg13g2_dlhq_1 _0923_ (.D(FrameData[21]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit21.Q ));
 sg13g2_dlhq_1 _0924_ (.D(FrameData[22]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit22.Q ));
 sg13g2_dlhq_1 _0925_ (.D(FrameData[23]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit23.Q ));
 sg13g2_dlhq_1 _0926_ (.D(FrameData[24]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit24.Q ));
 sg13g2_dlhq_1 _0927_ (.D(FrameData[25]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit25.Q ));
 sg13g2_dlhq_1 _0928_ (.D(FrameData[26]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit26.Q ));
 sg13g2_dlhq_1 _0929_ (.D(FrameData[27]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit27.Q ));
 sg13g2_dlhq_1 _0930_ (.D(FrameData[28]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit28.Q ));
 sg13g2_dlhq_1 _0931_ (.D(FrameData[29]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit29.Q ));
 sg13g2_dlhq_1 _0932_ (.D(FrameData[30]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit30.Q ));
 sg13g2_dlhq_1 _0933_ (.D(FrameData[31]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame7_bit31.Q ));
 sg13g2_dlhq_1 _0934_ (.D(FrameData[0]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit0.Q ));
 sg13g2_dlhq_1 _0935_ (.D(FrameData[1]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit1.Q ));
 sg13g2_dlhq_1 _0936_ (.D(FrameData[2]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit2.Q ));
 sg13g2_dlhq_1 _0937_ (.D(FrameData[3]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit3.Q ));
 sg13g2_dlhq_1 _0938_ (.D(FrameData[4]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit4.Q ));
 sg13g2_dlhq_1 _0939_ (.D(FrameData[5]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit5.Q ));
 sg13g2_dlhq_1 _0940_ (.D(FrameData[6]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit6.Q ));
 sg13g2_dlhq_1 _0941_ (.D(FrameData[7]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit7.Q ));
 sg13g2_dlhq_1 _0942_ (.D(FrameData[8]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit8.Q ));
 sg13g2_dlhq_1 _0943_ (.D(FrameData[9]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit9.Q ));
 sg13g2_dlhq_1 _0944_ (.D(FrameData[10]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit10.Q ));
 sg13g2_dlhq_1 _0945_ (.D(FrameData[11]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit11.Q ));
 sg13g2_dlhq_1 _0946_ (.D(FrameData[12]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit12.Q ));
 sg13g2_dlhq_1 _0947_ (.D(FrameData[13]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit13.Q ));
 sg13g2_dlhq_1 _0948_ (.D(FrameData[14]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit14.Q ));
 sg13g2_dlhq_1 _0949_ (.D(FrameData[15]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit15.Q ));
 sg13g2_dlhq_1 _0950_ (.D(FrameData[16]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit16.Q ));
 sg13g2_dlhq_1 _0951_ (.D(FrameData[17]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit17.Q ));
 sg13g2_dlhq_1 _0952_ (.D(FrameData[18]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit18.Q ));
 sg13g2_dlhq_1 _0953_ (.D(FrameData[19]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit19.Q ));
 sg13g2_dlhq_1 _0954_ (.D(FrameData[20]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit20.Q ));
 sg13g2_dlhq_1 _0955_ (.D(FrameData[21]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit21.Q ));
 sg13g2_dlhq_1 _0956_ (.D(FrameData[22]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit22.Q ));
 sg13g2_dlhq_1 _0957_ (.D(FrameData[23]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit23.Q ));
 sg13g2_dlhq_1 _0958_ (.D(FrameData[24]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit24.Q ));
 sg13g2_dlhq_1 _0959_ (.D(FrameData[25]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit25.Q ));
 sg13g2_dlhq_1 _0960_ (.D(FrameData[26]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit26.Q ));
 sg13g2_dlhq_1 _0961_ (.D(FrameData[27]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit27.Q ));
 sg13g2_dlhq_1 _0962_ (.D(FrameData[28]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit28.Q ));
 sg13g2_dlhq_1 _0963_ (.D(FrameData[29]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit29.Q ));
 sg13g2_dlhq_1 _0964_ (.D(FrameData[30]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit30.Q ));
 sg13g2_dlhq_1 _0965_ (.D(FrameData[31]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame6_bit31.Q ));
 sg13g2_dlhq_1 _0966_ (.D(FrameData[0]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit0.Q ));
 sg13g2_dlhq_1 _0967_ (.D(FrameData[1]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit1.Q ));
 sg13g2_dlhq_1 _0968_ (.D(FrameData[2]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit2.Q ));
 sg13g2_dlhq_1 _0969_ (.D(FrameData[3]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit3.Q ));
 sg13g2_dlhq_1 _0970_ (.D(FrameData[4]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit4.Q ));
 sg13g2_dlhq_1 _0971_ (.D(FrameData[5]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit5.Q ));
 sg13g2_dlhq_1 _0972_ (.D(FrameData[6]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit6.Q ));
 sg13g2_dlhq_1 _0973_ (.D(FrameData[7]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit7.Q ));
 sg13g2_dlhq_1 _0974_ (.D(FrameData[8]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit8.Q ));
 sg13g2_dlhq_1 _0975_ (.D(FrameData[9]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit9.Q ));
 sg13g2_dlhq_1 _0976_ (.D(FrameData[10]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit10.Q ));
 sg13g2_dlhq_1 _0977_ (.D(FrameData[11]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit11.Q ));
 sg13g2_dlhq_1 _0978_ (.D(FrameData[12]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit12.Q ));
 sg13g2_dlhq_1 _0979_ (.D(FrameData[13]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit13.Q ));
 sg13g2_dlhq_1 _0980_ (.D(FrameData[14]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit14.Q ));
 sg13g2_dlhq_1 _0981_ (.D(FrameData[15]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit15.Q ));
 sg13g2_dlhq_1 _0982_ (.D(FrameData[16]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit16.Q ));
 sg13g2_dlhq_1 _0983_ (.D(FrameData[17]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit17.Q ));
 sg13g2_dlhq_1 _0984_ (.D(FrameData[18]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit18.Q ));
 sg13g2_dlhq_1 _0985_ (.D(FrameData[19]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit19.Q ));
 sg13g2_dlhq_1 _0986_ (.D(FrameData[20]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit20.Q ));
 sg13g2_dlhq_1 _0987_ (.D(FrameData[21]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit21.Q ));
 sg13g2_dlhq_1 _0988_ (.D(FrameData[22]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit22.Q ));
 sg13g2_dlhq_1 _0989_ (.D(FrameData[23]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit23.Q ));
 sg13g2_dlhq_1 _0990_ (.D(FrameData[24]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit24.Q ));
 sg13g2_dlhq_1 _0991_ (.D(FrameData[25]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit25.Q ));
 sg13g2_dlhq_1 _0992_ (.D(FrameData[26]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit26.Q ));
 sg13g2_dlhq_1 _0993_ (.D(FrameData[27]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit27.Q ));
 sg13g2_dlhq_1 _0994_ (.D(FrameData[28]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit28.Q ));
 sg13g2_dlhq_1 _0995_ (.D(FrameData[29]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit29.Q ));
 sg13g2_dlhq_1 _0996_ (.D(FrameData[30]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit30.Q ));
 sg13g2_dlhq_1 _0997_ (.D(FrameData[31]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame5_bit31.Q ));
 sg13g2_dlhq_1 _0998_ (.D(FrameData[0]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit0.Q ));
 sg13g2_dlhq_1 _0999_ (.D(FrameData[1]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit1.Q ));
 sg13g2_dlhq_1 _1000_ (.D(FrameData[2]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit2.Q ));
 sg13g2_dlhq_1 _1001_ (.D(FrameData[3]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit3.Q ));
 sg13g2_dlhq_1 _1002_ (.D(FrameData[4]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit4.Q ));
 sg13g2_dlhq_1 _1003_ (.D(FrameData[5]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit5.Q ));
 sg13g2_dlhq_1 _1004_ (.D(FrameData[6]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit6.Q ));
 sg13g2_dlhq_1 _1005_ (.D(FrameData[7]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit7.Q ));
 sg13g2_dlhq_1 _1006_ (.D(FrameData[8]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit8.Q ));
 sg13g2_dlhq_1 _1007_ (.D(FrameData[9]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit9.Q ));
 sg13g2_dlhq_1 _1008_ (.D(FrameData[10]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit10.Q ));
 sg13g2_dlhq_1 _1009_ (.D(FrameData[11]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit11.Q ));
 sg13g2_dlhq_1 _1010_ (.D(FrameData[12]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit12.Q ));
 sg13g2_dlhq_1 _1011_ (.D(FrameData[13]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit13.Q ));
 sg13g2_dlhq_1 _1012_ (.D(FrameData[14]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit14.Q ));
 sg13g2_dlhq_1 _1013_ (.D(FrameData[15]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit15.Q ));
 sg13g2_dlhq_1 _1014_ (.D(FrameData[16]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit16.Q ));
 sg13g2_dlhq_1 _1015_ (.D(FrameData[17]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit17.Q ));
 sg13g2_dlhq_1 _1016_ (.D(FrameData[18]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit18.Q ));
 sg13g2_dlhq_1 _1017_ (.D(FrameData[19]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit19.Q ));
 sg13g2_dlhq_1 _1018_ (.D(FrameData[20]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit20.Q ));
 sg13g2_dlhq_1 _1019_ (.D(FrameData[21]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit21.Q ));
 sg13g2_dlhq_1 _1020_ (.D(FrameData[22]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit22.Q ));
 sg13g2_dlhq_1 _1021_ (.D(FrameData[23]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit23.Q ));
 sg13g2_dlhq_1 _1022_ (.D(FrameData[24]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit24.Q ));
 sg13g2_dlhq_1 _1023_ (.D(FrameData[25]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit25.Q ));
 sg13g2_dlhq_1 _1024_ (.D(FrameData[26]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit26.Q ));
 sg13g2_dlhq_1 _1025_ (.D(FrameData[27]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit27.Q ));
 sg13g2_dlhq_1 _1026_ (.D(FrameData[28]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit28.Q ));
 sg13g2_dlhq_1 _1027_ (.D(FrameData[29]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit29.Q ));
 sg13g2_dlhq_1 _1028_ (.D(FrameData[30]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit30.Q ));
 sg13g2_dlhq_1 _1029_ (.D(FrameData[31]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame4_bit31.Q ));
 sg13g2_dlhq_1 _1030_ (.D(FrameData[0]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit0.Q ));
 sg13g2_dlhq_1 _1031_ (.D(FrameData[1]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit1.Q ));
 sg13g2_dlhq_1 _1032_ (.D(FrameData[2]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit2.Q ));
 sg13g2_dlhq_1 _1033_ (.D(FrameData[3]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit3.Q ));
 sg13g2_dlhq_1 _1034_ (.D(FrameData[4]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit4.Q ));
 sg13g2_dlhq_1 _1035_ (.D(FrameData[5]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit5.Q ));
 sg13g2_dlhq_1 _1036_ (.D(FrameData[6]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit6.Q ));
 sg13g2_dlhq_1 _1037_ (.D(FrameData[7]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit7.Q ));
 sg13g2_dlhq_1 _1038_ (.D(FrameData[8]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit8.Q ));
 sg13g2_dlhq_1 _1039_ (.D(FrameData[9]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit9.Q ));
 sg13g2_dlhq_1 _1040_ (.D(FrameData[10]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit10.Q ));
 sg13g2_dlhq_1 _1041_ (.D(FrameData[11]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit11.Q ));
 sg13g2_dlhq_1 _1042_ (.D(FrameData[12]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit12.Q ));
 sg13g2_dlhq_1 _1043_ (.D(FrameData[13]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit13.Q ));
 sg13g2_dlhq_1 _1044_ (.D(FrameData[14]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit14.Q ));
 sg13g2_dlhq_1 _1045_ (.D(FrameData[15]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit15.Q ));
 sg13g2_dlhq_1 _1046_ (.D(FrameData[16]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit16.Q ));
 sg13g2_dlhq_1 _1047_ (.D(FrameData[17]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit17.Q ));
 sg13g2_dlhq_1 _1048_ (.D(FrameData[18]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit18.Q ));
 sg13g2_dlhq_1 _1049_ (.D(FrameData[19]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit19.Q ));
 sg13g2_dlhq_1 _1050_ (.D(FrameData[20]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit20.Q ));
 sg13g2_dlhq_1 _1051_ (.D(FrameData[21]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit21.Q ));
 sg13g2_dlhq_1 _1052_ (.D(FrameData[22]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit22.Q ));
 sg13g2_dlhq_1 _1053_ (.D(FrameData[23]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit23.Q ));
 sg13g2_dlhq_1 _1054_ (.D(FrameData[24]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit24.Q ));
 sg13g2_dlhq_1 _1055_ (.D(FrameData[25]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit25.Q ));
 sg13g2_dlhq_1 _1056_ (.D(FrameData[26]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit26.Q ));
 sg13g2_dlhq_1 _1057_ (.D(FrameData[27]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit27.Q ));
 sg13g2_dlhq_1 _1058_ (.D(FrameData[28]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit28.Q ));
 sg13g2_dlhq_1 _1059_ (.D(FrameData[29]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit29.Q ));
 sg13g2_dlhq_1 _1060_ (.D(FrameData[30]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit30.Q ));
 sg13g2_dlhq_1 _1061_ (.D(FrameData[31]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame3_bit31.Q ));
 sg13g2_dlhq_1 _1062_ (.D(FrameData[0]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit0.Q ));
 sg13g2_dlhq_1 _1063_ (.D(FrameData[1]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit1.Q ));
 sg13g2_dlhq_1 _1064_ (.D(FrameData[2]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit2.Q ));
 sg13g2_dlhq_1 _1065_ (.D(FrameData[3]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit3.Q ));
 sg13g2_dlhq_1 _1066_ (.D(FrameData[4]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit4.Q ));
 sg13g2_dlhq_1 _1067_ (.D(FrameData[5]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit5.Q ));
 sg13g2_dlhq_1 _1068_ (.D(FrameData[6]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit6.Q ));
 sg13g2_dlhq_1 _1069_ (.D(FrameData[7]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit7.Q ));
 sg13g2_dlhq_1 _1070_ (.D(FrameData[8]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit8.Q ));
 sg13g2_dlhq_1 _1071_ (.D(FrameData[9]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit9.Q ));
 sg13g2_dlhq_1 _1072_ (.D(FrameData[10]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit10.Q ));
 sg13g2_dlhq_1 _1073_ (.D(FrameData[11]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit11.Q ));
 sg13g2_dlhq_1 _1074_ (.D(FrameData[12]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit12.Q ));
 sg13g2_dlhq_1 _1075_ (.D(FrameData[13]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit13.Q ));
 sg13g2_dlhq_1 _1076_ (.D(FrameData[14]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit14.Q ));
 sg13g2_dlhq_1 _1077_ (.D(FrameData[15]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit15.Q ));
 sg13g2_dlhq_1 _1078_ (.D(FrameData[16]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit16.Q ));
 sg13g2_dlhq_1 _1079_ (.D(FrameData[17]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit17.Q ));
 sg13g2_dlhq_1 _1080_ (.D(FrameData[18]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit18.Q ));
 sg13g2_dlhq_1 _1081_ (.D(FrameData[19]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit19.Q ));
 sg13g2_dlhq_1 _1082_ (.D(FrameData[20]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit20.Q ));
 sg13g2_dlhq_1 _1083_ (.D(FrameData[21]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit21.Q ));
 sg13g2_dlhq_1 _1084_ (.D(FrameData[22]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit22.Q ));
 sg13g2_dlhq_1 _1085_ (.D(FrameData[23]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit23.Q ));
 sg13g2_dlhq_1 _1086_ (.D(FrameData[24]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit24.Q ));
 sg13g2_dlhq_1 _1087_ (.D(FrameData[25]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit25.Q ));
 sg13g2_dlhq_1 _1088_ (.D(FrameData[26]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit26.Q ));
 sg13g2_dlhq_1 _1089_ (.D(FrameData[27]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit27.Q ));
 sg13g2_dlhq_1 _1090_ (.D(FrameData[28]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit28.Q ));
 sg13g2_dlhq_1 _1091_ (.D(FrameData[29]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit29.Q ));
 sg13g2_dlhq_1 _1092_ (.D(FrameData[30]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit30.Q ));
 sg13g2_dlhq_1 _1093_ (.D(FrameData[31]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame2_bit31.Q ));
 sg13g2_dlhq_1 _1094_ (.D(FrameData[0]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit0.Q ));
 sg13g2_dlhq_1 _1095_ (.D(FrameData[1]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit1.Q ));
 sg13g2_dlhq_1 _1096_ (.D(FrameData[2]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit2.Q ));
 sg13g2_dlhq_1 _1097_ (.D(FrameData[3]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit3.Q ));
 sg13g2_dlhq_1 _1098_ (.D(FrameData[4]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit4.Q ));
 sg13g2_dlhq_1 _1099_ (.D(FrameData[5]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit5.Q ));
 sg13g2_dlhq_1 _1100_ (.D(FrameData[6]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit6.Q ));
 sg13g2_dlhq_1 _1101_ (.D(FrameData[7]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit7.Q ));
 sg13g2_dlhq_1 _1102_ (.D(FrameData[8]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit8.Q ));
 sg13g2_dlhq_1 _1103_ (.D(FrameData[9]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit9.Q ));
 sg13g2_dlhq_1 _1104_ (.D(FrameData[10]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit10.Q ));
 sg13g2_dlhq_1 _1105_ (.D(FrameData[11]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit11.Q ));
 sg13g2_dlhq_1 _1106_ (.D(FrameData[12]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit12.Q ));
 sg13g2_dlhq_1 _1107_ (.D(FrameData[13]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit13.Q ));
 sg13g2_dlhq_1 _1108_ (.D(FrameData[14]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit14.Q ));
 sg13g2_dlhq_1 _1109_ (.D(FrameData[15]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit15.Q ));
 sg13g2_dlhq_1 _1110_ (.D(FrameData[16]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit16.Q ));
 sg13g2_dlhq_1 _1111_ (.D(FrameData[17]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit17.Q ));
 sg13g2_dlhq_1 _1112_ (.D(FrameData[18]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit18.Q ));
 sg13g2_dlhq_1 _1113_ (.D(FrameData[19]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit19.Q ));
 sg13g2_dlhq_1 _1114_ (.D(FrameData[20]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit20.Q ));
 sg13g2_dlhq_1 _1115_ (.D(FrameData[21]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit21.Q ));
 sg13g2_dlhq_1 _1116_ (.D(FrameData[22]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit22.Q ));
 sg13g2_dlhq_1 _1117_ (.D(FrameData[23]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit23.Q ));
 sg13g2_dlhq_1 _1118_ (.D(FrameData[24]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit24.Q ));
 sg13g2_dlhq_1 _1119_ (.D(FrameData[25]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit25.Q ));
 sg13g2_dlhq_1 _1120_ (.D(FrameData[26]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit26.Q ));
 sg13g2_dlhq_1 _1121_ (.D(FrameData[27]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit27.Q ));
 sg13g2_dlhq_1 _1122_ (.D(FrameData[28]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit28.Q ));
 sg13g2_dlhq_1 _1123_ (.D(FrameData[29]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit29.Q ));
 sg13g2_dlhq_1 _1124_ (.D(FrameData[30]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit30.Q ));
 sg13g2_dlhq_1 _1125_ (.D(FrameData[31]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame1_bit31.Q ));
 sg13g2_dlhq_1 _1126_ (.D(FrameData[0]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit0.Q ));
 sg13g2_dlhq_1 _1127_ (.D(FrameData[1]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit1.Q ));
 sg13g2_dlhq_1 _1128_ (.D(FrameData[2]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit2.Q ));
 sg13g2_dlhq_1 _1129_ (.D(FrameData[3]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit3.Q ));
 sg13g2_dlhq_1 _1130_ (.D(FrameData[4]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit4.Q ));
 sg13g2_dlhq_1 _1131_ (.D(FrameData[5]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit5.Q ));
 sg13g2_dlhq_1 _1132_ (.D(FrameData[6]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit6.Q ));
 sg13g2_dlhq_1 _1133_ (.D(FrameData[7]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit7.Q ));
 sg13g2_dlhq_1 _1134_ (.D(FrameData[8]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit8.Q ));
 sg13g2_dlhq_1 _1135_ (.D(FrameData[9]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit9.Q ));
 sg13g2_dlhq_1 _1136_ (.D(FrameData[10]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit10.Q ));
 sg13g2_dlhq_1 _1137_ (.D(FrameData[11]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit11.Q ));
 sg13g2_dlhq_1 _1138_ (.D(FrameData[12]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit12.Q ));
 sg13g2_dlhq_1 _1139_ (.D(FrameData[13]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit13.Q ));
 sg13g2_dlhq_1 _1140_ (.D(FrameData[14]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit14.Q ));
 sg13g2_dlhq_1 _1141_ (.D(FrameData[15]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit15.Q ));
 sg13g2_dlhq_1 _1142_ (.D(FrameData[16]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit16.Q ));
 sg13g2_dlhq_1 _1143_ (.D(FrameData[17]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit17.Q ));
 sg13g2_dlhq_1 _1144_ (.D(FrameData[18]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit18.Q ));
 sg13g2_dlhq_1 _1145_ (.D(FrameData[19]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit19.Q ));
 sg13g2_dlhq_1 _1146_ (.D(FrameData[20]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit20.Q ));
 sg13g2_dlhq_1 _1147_ (.D(FrameData[21]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit21.Q ));
 sg13g2_dlhq_1 _1148_ (.D(FrameData[22]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit22.Q ));
 sg13g2_dlhq_1 _1149_ (.D(FrameData[23]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit23.Q ));
 sg13g2_dlhq_1 _1150_ (.D(FrameData[24]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit24.Q ));
 sg13g2_dlhq_1 _1151_ (.D(FrameData[25]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit25.Q ));
 sg13g2_dlhq_1 _1152_ (.D(FrameData[26]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit26.Q ));
 sg13g2_dlhq_1 _1153_ (.D(FrameData[27]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit27.Q ));
 sg13g2_dlhq_1 _1154_ (.D(FrameData[28]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit28.Q ));
 sg13g2_dlhq_1 _1155_ (.D(FrameData[29]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit29.Q ));
 sg13g2_dlhq_1 _1156_ (.D(FrameData[30]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit30.Q ));
 sg13g2_dlhq_1 _1157_ (.D(FrameData[31]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_W_TT_IF_ConfigMem.Inst_frame0_bit31.Q ));
 sg13g2_buf_1 _1158_ (.A(clknet_1_0__leaf_UserCLK),
    .X(CLK_TT_PROJECT));
 sg13g2_buf_1 _1159_ (.A(\Inst_W_TT_IF_switch_matrix.E1BEG0 ),
    .X(E1BEG[0]));
 sg13g2_buf_1 _1160_ (.A(\Inst_W_TT_IF_switch_matrix.E1BEG1 ),
    .X(E1BEG[1]));
 sg13g2_buf_1 _1161_ (.A(\Inst_W_TT_IF_switch_matrix.E1BEG2 ),
    .X(E1BEG[2]));
 sg13g2_buf_1 _1162_ (.A(\Inst_W_TT_IF_switch_matrix.E1BEG3 ),
    .X(E1BEG[3]));
 sg13g2_buf_1 _1163_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEG0 ),
    .X(E2BEG[0]));
 sg13g2_buf_1 _1164_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEG1 ),
    .X(E2BEG[1]));
 sg13g2_buf_1 _1165_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEG2 ),
    .X(E2BEG[2]));
 sg13g2_buf_1 _1166_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEG3 ),
    .X(E2BEG[3]));
 sg13g2_buf_1 _1167_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEG4 ),
    .X(E2BEG[4]));
 sg13g2_buf_1 _1168_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEG5 ),
    .X(E2BEG[5]));
 sg13g2_buf_1 _1169_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEG6 ),
    .X(E2BEG[6]));
 sg13g2_buf_1 _1170_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEG7 ),
    .X(E2BEG[7]));
 sg13g2_buf_1 _1171_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEGb0 ),
    .X(E2BEGb[0]));
 sg13g2_buf_1 _1172_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEGb1 ),
    .X(E2BEGb[1]));
 sg13g2_buf_1 _1173_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEGb2 ),
    .X(E2BEGb[2]));
 sg13g2_buf_1 _1174_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEGb3 ),
    .X(E2BEGb[3]));
 sg13g2_buf_1 _1175_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEGb4 ),
    .X(E2BEGb[4]));
 sg13g2_buf_1 _1176_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEGb5 ),
    .X(E2BEGb[5]));
 sg13g2_buf_1 _1177_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEGb6 ),
    .X(E2BEGb[6]));
 sg13g2_buf_1 _1178_ (.A(\Inst_W_TT_IF_switch_matrix.E2BEGb7 ),
    .X(E2BEGb[7]));
 sg13g2_buf_1 _1179_ (.A(\Inst_W_TT_IF_switch_matrix.E6BEG0 ),
    .X(E6BEG[0]));
 sg13g2_buf_1 _1180_ (.A(\Inst_W_TT_IF_switch_matrix.E6BEG1 ),
    .X(E6BEG[1]));
 sg13g2_buf_1 _1181_ (.A(\Inst_W_TT_IF_switch_matrix.E6BEG2 ),
    .X(E6BEG[2]));
 sg13g2_buf_1 _1182_ (.A(\Inst_W_TT_IF_switch_matrix.E6BEG3 ),
    .X(E6BEG[3]));
 sg13g2_buf_1 _1183_ (.A(\Inst_W_TT_IF_switch_matrix.E6BEG4 ),
    .X(E6BEG[4]));
 sg13g2_buf_1 _1184_ (.A(\Inst_W_TT_IF_switch_matrix.E6BEG5 ),
    .X(E6BEG[5]));
 sg13g2_buf_1 _1185_ (.A(\Inst_W_TT_IF_switch_matrix.E6BEG6 ),
    .X(E6BEG[6]));
 sg13g2_buf_1 _1186_ (.A(\Inst_W_TT_IF_switch_matrix.E6BEG7 ),
    .X(E6BEG[7]));
 sg13g2_buf_1 _1187_ (.A(\Inst_W_TT_IF_switch_matrix.E6BEG8 ),
    .X(E6BEG[8]));
 sg13g2_buf_1 _1188_ (.A(\Inst_W_TT_IF_switch_matrix.E6BEG9 ),
    .X(E6BEG[9]));
 sg13g2_buf_1 _1189_ (.A(\Inst_W_TT_IF_switch_matrix.E6BEG10 ),
    .X(E6BEG[10]));
 sg13g2_buf_1 _1190_ (.A(\Inst_W_TT_IF_switch_matrix.E6BEG11 ),
    .X(E6BEG[11]));
 sg13g2_buf_1 _1191_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG0 ),
    .X(EE4BEG[0]));
 sg13g2_buf_1 _1192_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG1 ),
    .X(EE4BEG[1]));
 sg13g2_buf_1 _1193_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG2 ),
    .X(EE4BEG[2]));
 sg13g2_buf_1 _1194_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG3 ),
    .X(EE4BEG[3]));
 sg13g2_buf_1 _1195_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG4 ),
    .X(EE4BEG[4]));
 sg13g2_buf_1 _1196_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG5 ),
    .X(EE4BEG[5]));
 sg13g2_buf_1 _1197_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG6 ),
    .X(EE4BEG[6]));
 sg13g2_buf_1 _1198_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG7 ),
    .X(EE4BEG[7]));
 sg13g2_buf_1 _1199_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG8 ),
    .X(EE4BEG[8]));
 sg13g2_buf_1 _1200_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG9 ),
    .X(EE4BEG[9]));
 sg13g2_buf_1 _1201_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG10 ),
    .X(EE4BEG[10]));
 sg13g2_buf_1 _1202_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG11 ),
    .X(EE4BEG[11]));
 sg13g2_buf_1 _1203_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG12 ),
    .X(EE4BEG[12]));
 sg13g2_buf_1 _1204_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG13 ),
    .X(EE4BEG[13]));
 sg13g2_buf_1 _1205_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG14 ),
    .X(EE4BEG[14]));
 sg13g2_buf_1 _1206_ (.A(\Inst_W_TT_IF_switch_matrix.EE4BEG15 ),
    .X(EE4BEG[15]));
 sg13g2_buf_1 _1207_ (.A(FrameData[0]),
    .X(FrameData_O[0]));
 sg13g2_buf_1 _1208_ (.A(FrameData[1]),
    .X(FrameData_O[1]));
 sg13g2_buf_1 _1209_ (.A(FrameData[2]),
    .X(FrameData_O[2]));
 sg13g2_buf_1 _1210_ (.A(FrameData[3]),
    .X(FrameData_O[3]));
 sg13g2_buf_1 _1211_ (.A(FrameData[4]),
    .X(FrameData_O[4]));
 sg13g2_buf_1 _1212_ (.A(FrameData[5]),
    .X(FrameData_O[5]));
 sg13g2_buf_1 _1213_ (.A(FrameData[6]),
    .X(FrameData_O[6]));
 sg13g2_buf_1 _1214_ (.A(FrameData[7]),
    .X(FrameData_O[7]));
 sg13g2_buf_1 _1215_ (.A(FrameData[8]),
    .X(FrameData_O[8]));
 sg13g2_buf_1 _1216_ (.A(FrameData[9]),
    .X(FrameData_O[9]));
 sg13g2_buf_1 _1217_ (.A(FrameData[10]),
    .X(FrameData_O[10]));
 sg13g2_buf_1 _1218_ (.A(FrameData[11]),
    .X(FrameData_O[11]));
 sg13g2_buf_1 _1219_ (.A(FrameData[12]),
    .X(FrameData_O[12]));
 sg13g2_buf_1 _1220_ (.A(FrameData[13]),
    .X(FrameData_O[13]));
 sg13g2_buf_1 _1221_ (.A(FrameData[14]),
    .X(FrameData_O[14]));
 sg13g2_buf_1 _1222_ (.A(FrameData[15]),
    .X(FrameData_O[15]));
 sg13g2_buf_1 _1223_ (.A(FrameData[16]),
    .X(FrameData_O[16]));
 sg13g2_buf_1 _1224_ (.A(FrameData[17]),
    .X(FrameData_O[17]));
 sg13g2_buf_1 _1225_ (.A(FrameData[18]),
    .X(FrameData_O[18]));
 sg13g2_buf_1 _1226_ (.A(FrameData[19]),
    .X(FrameData_O[19]));
 sg13g2_buf_1 _1227_ (.A(FrameData[20]),
    .X(FrameData_O[20]));
 sg13g2_buf_1 _1228_ (.A(FrameData[21]),
    .X(FrameData_O[21]));
 sg13g2_buf_1 _1229_ (.A(FrameData[22]),
    .X(FrameData_O[22]));
 sg13g2_buf_1 _1230_ (.A(FrameData[23]),
    .X(FrameData_O[23]));
 sg13g2_buf_1 _1231_ (.A(FrameData[24]),
    .X(FrameData_O[24]));
 sg13g2_buf_1 _1232_ (.A(FrameData[25]),
    .X(FrameData_O[25]));
 sg13g2_buf_1 _1233_ (.A(FrameData[26]),
    .X(FrameData_O[26]));
 sg13g2_buf_1 _1234_ (.A(FrameData[27]),
    .X(FrameData_O[27]));
 sg13g2_buf_1 _1235_ (.A(FrameData[28]),
    .X(FrameData_O[28]));
 sg13g2_buf_1 _1236_ (.A(FrameData[29]),
    .X(FrameData_O[29]));
 sg13g2_buf_1 _1237_ (.A(FrameData[30]),
    .X(FrameData_O[30]));
 sg13g2_buf_1 _1238_ (.A(FrameData[31]),
    .X(FrameData_O[31]));
 sg13g2_buf_1 _1239_ (.A(FrameStrobe[0]),
    .X(FrameStrobe_O[0]));
 sg13g2_buf_1 _1240_ (.A(FrameStrobe[1]),
    .X(FrameStrobe_O[1]));
 sg13g2_buf_1 _1241_ (.A(FrameStrobe[2]),
    .X(FrameStrobe_O[2]));
 sg13g2_buf_1 _1242_ (.A(FrameStrobe[3]),
    .X(FrameStrobe_O[3]));
 sg13g2_buf_1 _1243_ (.A(FrameStrobe[4]),
    .X(FrameStrobe_O[4]));
 sg13g2_buf_1 _1244_ (.A(FrameStrobe[5]),
    .X(FrameStrobe_O[5]));
 sg13g2_buf_1 _1245_ (.A(FrameStrobe[6]),
    .X(FrameStrobe_O[6]));
 sg13g2_buf_1 _1246_ (.A(FrameStrobe[7]),
    .X(FrameStrobe_O[7]));
 sg13g2_buf_1 _1247_ (.A(FrameStrobe[8]),
    .X(FrameStrobe_O[8]));
 sg13g2_buf_1 _1248_ (.A(FrameStrobe[9]),
    .X(FrameStrobe_O[9]));
 sg13g2_buf_1 _1249_ (.A(FrameStrobe[10]),
    .X(FrameStrobe_O[10]));
 sg13g2_buf_1 _1250_ (.A(FrameStrobe[11]),
    .X(FrameStrobe_O[11]));
 sg13g2_buf_1 _1251_ (.A(FrameStrobe[12]),
    .X(FrameStrobe_O[12]));
 sg13g2_buf_1 _1252_ (.A(FrameStrobe[13]),
    .X(FrameStrobe_O[13]));
 sg13g2_buf_1 _1253_ (.A(FrameStrobe[14]),
    .X(FrameStrobe_O[14]));
 sg13g2_buf_1 _1254_ (.A(FrameStrobe[15]),
    .X(FrameStrobe_O[15]));
 sg13g2_buf_1 _1255_ (.A(FrameStrobe[16]),
    .X(FrameStrobe_O[16]));
 sg13g2_buf_1 _1256_ (.A(FrameStrobe[17]),
    .X(FrameStrobe_O[17]));
 sg13g2_buf_1 _1257_ (.A(FrameStrobe[18]),
    .X(FrameStrobe_O[18]));
 sg13g2_buf_1 _1258_ (.A(FrameStrobe[19]),
    .X(FrameStrobe_O[19]));
 sg13g2_buf_1 _1259_ (.A(\Inst_W_TT_IF_switch_matrix.N1BEG0 ),
    .X(N1BEG[0]));
 sg13g2_buf_1 _1260_ (.A(\Inst_W_TT_IF_switch_matrix.N1BEG1 ),
    .X(N1BEG[1]));
 sg13g2_buf_1 _1261_ (.A(\Inst_W_TT_IF_switch_matrix.N1BEG2 ),
    .X(N1BEG[2]));
 sg13g2_buf_1 _1262_ (.A(\Inst_W_TT_IF_switch_matrix.N1BEG3 ),
    .X(N1BEG[3]));
 sg13g2_buf_1 _1263_ (.A(\Inst_W_TT_IF_switch_matrix.N2BEG0 ),
    .X(N2BEG[0]));
 sg13g2_buf_1 _1264_ (.A(\Inst_W_TT_IF_switch_matrix.N2BEG1 ),
    .X(N2BEG[1]));
 sg13g2_buf_1 _1265_ (.A(\Inst_W_TT_IF_switch_matrix.N2BEG2 ),
    .X(N2BEG[2]));
 sg13g2_buf_1 _1266_ (.A(\Inst_W_TT_IF_switch_matrix.N2BEG3 ),
    .X(N2BEG[3]));
 sg13g2_buf_1 _1267_ (.A(\Inst_W_TT_IF_switch_matrix.N2BEG4 ),
    .X(N2BEG[4]));
 sg13g2_buf_1 _1268_ (.A(\Inst_W_TT_IF_switch_matrix.N2BEG5 ),
    .X(N2BEG[5]));
 sg13g2_buf_1 _1269_ (.A(\Inst_W_TT_IF_switch_matrix.N2BEG6 ),
    .X(N2BEG[6]));
 sg13g2_buf_1 _1270_ (.A(\Inst_W_TT_IF_switch_matrix.N2BEG7 ),
    .X(N2BEG[7]));
 sg13g2_buf_1 _1271_ (.A(N2MID[0]),
    .X(N2BEGb[0]));
 sg13g2_buf_1 _1272_ (.A(N2MID[1]),
    .X(N2BEGb[1]));
 sg13g2_buf_1 _1273_ (.A(N2MID[2]),
    .X(N2BEGb[2]));
 sg13g2_buf_1 _1274_ (.A(N2MID[3]),
    .X(N2BEGb[3]));
 sg13g2_buf_1 _1275_ (.A(N2MID[4]),
    .X(N2BEGb[4]));
 sg13g2_buf_1 _1276_ (.A(N2MID[5]),
    .X(N2BEGb[5]));
 sg13g2_buf_1 _1277_ (.A(N2MID[6]),
    .X(N2BEGb[6]));
 sg13g2_buf_1 _1278_ (.A(N2MID[7]),
    .X(N2BEGb[7]));
 sg13g2_buf_1 _1279_ (.A(N4END[4]),
    .X(N4BEG[0]));
 sg13g2_buf_1 _1280_ (.A(N4END[5]),
    .X(N4BEG[1]));
 sg13g2_buf_1 _1281_ (.A(N4END[6]),
    .X(N4BEG[2]));
 sg13g2_buf_1 _1282_ (.A(N4END[7]),
    .X(N4BEG[3]));
 sg13g2_buf_1 _1283_ (.A(N4END[8]),
    .X(N4BEG[4]));
 sg13g2_buf_1 _1284_ (.A(N4END[9]),
    .X(N4BEG[5]));
 sg13g2_buf_1 _1285_ (.A(N4END[10]),
    .X(N4BEG[6]));
 sg13g2_buf_1 _1286_ (.A(N4END[11]),
    .X(N4BEG[7]));
 sg13g2_buf_1 _1287_ (.A(N4END[12]),
    .X(N4BEG[8]));
 sg13g2_buf_1 _1288_ (.A(N4END[13]),
    .X(N4BEG[9]));
 sg13g2_buf_1 _1289_ (.A(N4END[14]),
    .X(N4BEG[10]));
 sg13g2_buf_1 _1290_ (.A(N4END[15]),
    .X(N4BEG[11]));
 sg13g2_buf_1 _1291_ (.A(\Inst_W_TT_IF_switch_matrix.N4BEG0 ),
    .X(N4BEG[12]));
 sg13g2_buf_1 _1292_ (.A(\Inst_W_TT_IF_switch_matrix.N4BEG1 ),
    .X(N4BEG[13]));
 sg13g2_buf_1 _1293_ (.A(\Inst_W_TT_IF_switch_matrix.N4BEG2 ),
    .X(N4BEG[14]));
 sg13g2_buf_1 _1294_ (.A(\Inst_W_TT_IF_switch_matrix.N4BEG3 ),
    .X(N4BEG[15]));
 sg13g2_buf_1 _1295_ (.A(\Inst_W_TT_IF_switch_matrix.S1BEG0 ),
    .X(S1BEG[0]));
 sg13g2_buf_1 _1296_ (.A(\Inst_W_TT_IF_switch_matrix.S1BEG1 ),
    .X(S1BEG[1]));
 sg13g2_buf_1 _1297_ (.A(\Inst_W_TT_IF_switch_matrix.S1BEG2 ),
    .X(S1BEG[2]));
 sg13g2_buf_1 _1298_ (.A(\Inst_W_TT_IF_switch_matrix.S1BEG3 ),
    .X(S1BEG[3]));
 sg13g2_buf_1 _1299_ (.A(\Inst_W_TT_IF_switch_matrix.S2BEG0 ),
    .X(S2BEG[0]));
 sg13g2_buf_1 _1300_ (.A(\Inst_W_TT_IF_switch_matrix.S2BEG1 ),
    .X(S2BEG[1]));
 sg13g2_buf_1 _1301_ (.A(\Inst_W_TT_IF_switch_matrix.S2BEG2 ),
    .X(S2BEG[2]));
 sg13g2_buf_1 _1302_ (.A(\Inst_W_TT_IF_switch_matrix.S2BEG3 ),
    .X(S2BEG[3]));
 sg13g2_buf_1 _1303_ (.A(\Inst_W_TT_IF_switch_matrix.S2BEG4 ),
    .X(S2BEG[4]));
 sg13g2_buf_1 _1304_ (.A(\Inst_W_TT_IF_switch_matrix.S2BEG5 ),
    .X(S2BEG[5]));
 sg13g2_buf_1 _1305_ (.A(\Inst_W_TT_IF_switch_matrix.S2BEG6 ),
    .X(S2BEG[6]));
 sg13g2_buf_1 _1306_ (.A(\Inst_W_TT_IF_switch_matrix.S2BEG7 ),
    .X(S2BEG[7]));
 sg13g2_buf_1 _1307_ (.A(S2MID[0]),
    .X(S2BEGb[0]));
 sg13g2_buf_1 _1308_ (.A(S2MID[1]),
    .X(S2BEGb[1]));
 sg13g2_buf_1 _1309_ (.A(S2MID[2]),
    .X(S2BEGb[2]));
 sg13g2_buf_1 _1310_ (.A(S2MID[3]),
    .X(S2BEGb[3]));
 sg13g2_buf_1 _1311_ (.A(S2MID[4]),
    .X(S2BEGb[4]));
 sg13g2_buf_1 _1312_ (.A(S2MID[5]),
    .X(S2BEGb[5]));
 sg13g2_buf_1 _1313_ (.A(S2MID[6]),
    .X(S2BEGb[6]));
 sg13g2_buf_1 _1314_ (.A(S2MID[7]),
    .X(S2BEGb[7]));
 sg13g2_buf_1 _1315_ (.A(S4END[4]),
    .X(S4BEG[0]));
 sg13g2_buf_1 _1316_ (.A(S4END[5]),
    .X(S4BEG[1]));
 sg13g2_buf_1 _1317_ (.A(S4END[6]),
    .X(S4BEG[2]));
 sg13g2_buf_1 _1318_ (.A(S4END[7]),
    .X(S4BEG[3]));
 sg13g2_buf_1 _1319_ (.A(S4END[8]),
    .X(S4BEG[4]));
 sg13g2_buf_1 _1320_ (.A(S4END[9]),
    .X(S4BEG[5]));
 sg13g2_buf_1 _1321_ (.A(S4END[10]),
    .X(S4BEG[6]));
 sg13g2_buf_1 _1322_ (.A(S4END[11]),
    .X(S4BEG[7]));
 sg13g2_buf_1 _1323_ (.A(S4END[12]),
    .X(S4BEG[8]));
 sg13g2_buf_1 _1324_ (.A(S4END[13]),
    .X(S4BEG[9]));
 sg13g2_buf_1 _1325_ (.A(S4END[14]),
    .X(S4BEG[10]));
 sg13g2_buf_1 _1326_ (.A(S4END[15]),
    .X(S4BEG[11]));
 sg13g2_buf_1 _1327_ (.A(\Inst_W_TT_IF_switch_matrix.S4BEG0 ),
    .X(S4BEG[12]));
 sg13g2_buf_1 _1328_ (.A(\Inst_W_TT_IF_switch_matrix.S4BEG1 ),
    .X(S4BEG[13]));
 sg13g2_buf_1 _1329_ (.A(\Inst_W_TT_IF_switch_matrix.S4BEG2 ),
    .X(S4BEG[14]));
 sg13g2_buf_1 _1330_ (.A(\Inst_W_TT_IF_switch_matrix.S4BEG3 ),
    .X(S4BEG[15]));
 sg13g2_buf_1 _1331_ (.A(clknet_1_1__leaf_UserCLK),
    .X(UserCLKo));
 sg13g2_buf_8 clkbuf_0_UserCLK (.A(UserCLK),
    .X(clknet_0_UserCLK));
 sg13g2_buf_8 clkbuf_1_0__f_UserCLK (.A(clknet_0_UserCLK),
    .X(clknet_1_0__leaf_UserCLK));
 sg13g2_buf_8 clkbuf_1_1__f_UserCLK (.A(clknet_0_UserCLK),
    .X(clknet_1_1__leaf_UserCLK));
 sg13g2_antennanp ANTENNA_1 (.A(FrameStrobe[10]));
 sg13g2_antennanp ANTENNA_2 (.A(FrameStrobe[11]));
 sg13g2_antennanp ANTENNA_3 (.A(N2END[5]));
 sg13g2_antennanp ANTENNA_4 (.A(N2MID[0]));
 sg13g2_antennanp ANTENNA_5 (.A(N2MID[0]));
 sg13g2_antennanp ANTENNA_6 (.A(N2MID[0]));
 sg13g2_antennanp ANTENNA_7 (.A(N4END[14]));
 sg13g2_antennanp ANTENNA_8 (.A(N4END[15]));
 sg13g2_antennanp ANTENNA_9 (.A(N4END[4]));
 sg13g2_antennanp ANTENNA_10 (.A(N4END[5]));
 sg13g2_antennanp ANTENNA_11 (.A(N4END[6]));
 sg13g2_antennanp ANTENNA_12 (.A(S2MID[1]));
 sg13g2_antennanp ANTENNA_13 (.A(S2MID[1]));
 sg13g2_antennanp ANTENNA_14 (.A(S2MID[2]));
 sg13g2_antennanp ANTENNA_15 (.A(S2MID[2]));
 sg13g2_antennanp ANTENNA_16 (.A(S2MID[2]));
 sg13g2_antennanp ANTENNA_17 (.A(S2MID[2]));
 sg13g2_antennanp ANTENNA_18 (.A(S2MID[3]));
 sg13g2_antennanp ANTENNA_19 (.A(S2MID[3]));
 sg13g2_antennanp ANTENNA_20 (.A(S2MID[3]));
 sg13g2_antennanp ANTENNA_21 (.A(S2MID[3]));
 sg13g2_antennanp ANTENNA_22 (.A(S2MID[4]));
 sg13g2_antennanp ANTENNA_23 (.A(S2MID[4]));
 sg13g2_antennanp ANTENNA_24 (.A(S2MID[4]));
 sg13g2_antennanp ANTENNA_25 (.A(S2MID[4]));
 sg13g2_antennanp ANTENNA_26 (.A(S2MID[7]));
 sg13g2_antennanp ANTENNA_27 (.A(S2MID[7]));
 sg13g2_antennanp ANTENNA_28 (.A(S2MID[7]));
 sg13g2_antennanp ANTENNA_29 (.A(FrameStrobe[13]));
 sg13g2_antennanp ANTENNA_30 (.A(FrameStrobe[13]));
 sg13g2_antennanp ANTENNA_31 (.A(N4END[7]));
 sg13g2_antennanp ANTENNA_32 (.A(S2END[3]));
 sg13g2_antennanp ANTENNA_33 (.A(S2END[3]));
 sg13g2_antennanp ANTENNA_34 (.A(S2END[3]));
 sg13g2_antennanp ANTENNA_35 (.A(S2END[3]));
 sg13g2_antennanp ANTENNA_36 (.A(S2MID[5]));
 sg13g2_antennanp ANTENNA_37 (.A(S2MID[5]));
 sg13g2_antennanp ANTENNA_38 (.A(S2MID[5]));
 sg13g2_antennanp ANTENNA_39 (.A(S2MID[5]));
 sg13g2_antennanp ANTENNA_40 (.A(S2MID[6]));
 sg13g2_antennanp ANTENNA_41 (.A(S2MID[6]));
 sg13g2_antennanp ANTENNA_42 (.A(S2MID[6]));
 sg13g2_antennanp ANTENNA_43 (.A(S2MID[6]));
 sg13g2_antennanp ANTENNA_44 (.A(N2MID[2]));
 sg13g2_antennanp ANTENNA_45 (.A(N2MID[2]));
 sg13g2_antennanp ANTENNA_46 (.A(N2MID[2]));
 sg13g2_antennanp ANTENNA_47 (.A(N2MID[2]));
 sg13g2_antennanp ANTENNA_48 (.A(S2MID[0]));
 sg13g2_antennanp ANTENNA_49 (.A(S2MID[0]));
 sg13g2_antennanp ANTENNA_50 (.A(S2MID[0]));
 sg13g2_antennanp ANTENNA_51 (.A(S2MID[0]));
 sg13g2_antennanp ANTENNA_52 (.A(S2MID[0]));
 sg13g2_antennanp ANTENNA_53 (.A(S2MID[0]));
 sg13g2_antennanp ANTENNA_54 (.A(S2MID[0]));
 sg13g2_antennanp ANTENNA_55 (.A(S2MID[0]));
 sg13g2_antennanp ANTENNA_56 (.A(S2MID[0]));
 sg13g2_antennanp ANTENNA_57 (.A(N2MID[3]));
 sg13g2_antennanp ANTENNA_58 (.A(N2MID[3]));
 sg13g2_antennanp ANTENNA_59 (.A(N2MID[3]));
 sg13g2_antennanp ANTENNA_60 (.A(N2MID[3]));
 sg13g2_antennanp ANTENNA_61 (.A(N2MID[7]));
 sg13g2_antennanp ANTENNA_62 (.A(N2MID[7]));
 sg13g2_antennanp ANTENNA_63 (.A(N2MID[7]));
 sg13g2_antennanp ANTENNA_64 (.A(N2MID[7]));
 sg13g2_antennanp ANTENNA_65 (.A(S2END[2]));
 sg13g2_antennanp ANTENNA_66 (.A(S2END[2]));
 sg13g2_antennanp ANTENNA_67 (.A(S2END[2]));
 sg13g2_antennanp ANTENNA_68 (.A(S2END[2]));
 sg13g2_antennanp ANTENNA_69 (.A(FrameStrobe[14]));
 sg13g2_antennanp ANTENNA_70 (.A(N2MID[1]));
 sg13g2_antennanp ANTENNA_71 (.A(N2MID[1]));
 sg13g2_antennanp ANTENNA_72 (.A(N2MID[1]));
 sg13g2_antennanp ANTENNA_73 (.A(N2MID[1]));
 sg13g2_fill_1 FILLER_0_34 ();
 sg13g2_fill_1 FILLER_0_174 ();
 sg13g2_fill_1 FILLER_1_27 ();
 sg13g2_fill_2 FILLER_1_151 ();
 sg13g2_fill_1 FILLER_1_191 ();
 sg13g2_fill_1 FILLER_2_0 ();
 sg13g2_fill_1 FILLER_2_27 ();
 sg13g2_fill_1 FILLER_2_36 ();
 sg13g2_fill_1 FILLER_2_108 ();
 sg13g2_fill_2 FILLER_2_173 ();
 sg13g2_fill_2 FILLER_3_0 ();
 sg13g2_fill_1 FILLER_3_30 ();
 sg13g2_fill_1 FILLER_3_75 ();
 sg13g2_fill_2 FILLER_3_97 ();
 sg13g2_fill_1 FILLER_3_112 ();
 sg13g2_fill_1 FILLER_3_199 ();
 sg13g2_fill_1 FILLER_4_112 ();
 sg13g2_fill_1 FILLER_4_135 ();
 sg13g2_fill_1 FILLER_4_199 ();
 sg13g2_fill_2 FILLER_5_58 ();
 sg13g2_fill_2 FILLER_5_72 ();
 sg13g2_fill_1 FILLER_5_129 ();
 sg13g2_fill_2 FILLER_5_170 ();
 sg13g2_fill_2 FILLER_5_177 ();
 sg13g2_fill_2 FILLER_5_198 ();
 sg13g2_fill_1 FILLER_6_33 ();
 sg13g2_fill_1 FILLER_6_121 ();
 sg13g2_fill_2 FILLER_7_52 ();
 sg13g2_fill_1 FILLER_7_135 ();
 sg13g2_fill_1 FILLER_7_171 ();
 sg13g2_fill_1 FILLER_7_199 ();
 sg13g2_fill_2 FILLER_8_65 ();
 sg13g2_fill_1 FILLER_8_142 ();
 sg13g2_fill_2 FILLER_8_171 ();
 sg13g2_fill_2 FILLER_8_198 ();
 sg13g2_fill_1 FILLER_9_17 ();
 sg13g2_fill_1 FILLER_9_47 ();
 sg13g2_fill_2 FILLER_9_69 ();
 sg13g2_fill_2 FILLER_9_94 ();
 sg13g2_fill_1 FILLER_9_118 ();
 sg13g2_fill_1 FILLER_9_137 ();
 sg13g2_fill_1 FILLER_9_174 ();
 sg13g2_fill_1 FILLER_10_126 ();
 sg13g2_fill_1 FILLER_10_164 ();
 sg13g2_fill_1 FILLER_10_199 ();
 sg13g2_fill_1 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_97 ();
 sg13g2_fill_1 FILLER_11_127 ();
 sg13g2_fill_1 FILLER_11_149 ();
 sg13g2_fill_2 FILLER_11_180 ();
 sg13g2_fill_1 FILLER_12_48 ();
 sg13g2_fill_2 FILLER_12_66 ();
 sg13g2_fill_1 FILLER_12_145 ();
 sg13g2_fill_1 FILLER_12_170 ();
 sg13g2_fill_2 FILLER_12_198 ();
 sg13g2_fill_1 FILLER_13_0 ();
 sg13g2_fill_1 FILLER_13_23 ();
 sg13g2_fill_1 FILLER_13_122 ();
 sg13g2_fill_1 FILLER_13_140 ();
 sg13g2_fill_1 FILLER_14_84 ();
 sg13g2_fill_1 FILLER_14_159 ();
 sg13g2_fill_1 FILLER_14_168 ();
 sg13g2_fill_2 FILLER_14_198 ();
 sg13g2_fill_1 FILLER_15_17 ();
 sg13g2_fill_2 FILLER_15_96 ();
 sg13g2_fill_1 FILLER_15_103 ();
 sg13g2_fill_2 FILLER_15_184 ();
 sg13g2_fill_1 FILLER_16_37 ();
 sg13g2_fill_2 FILLER_16_93 ();
 sg13g2_fill_1 FILLER_16_112 ();
 sg13g2_fill_1 FILLER_17_64 ();
 sg13g2_fill_1 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_57 ();
 sg13g2_fill_2 FILLER_18_63 ();
 sg13g2_fill_1 FILLER_18_65 ();
 sg13g2_fill_2 FILLER_18_144 ();
 sg13g2_fill_1 FILLER_18_146 ();
 sg13g2_fill_2 FILLER_18_174 ();
 sg13g2_fill_1 FILLER_18_185 ();
 sg13g2_fill_2 FILLER_19_147 ();
 sg13g2_fill_1 FILLER_19_149 ();
 sg13g2_fill_2 FILLER_19_198 ();
 sg13g2_fill_1 FILLER_20_34 ();
 sg13g2_fill_1 FILLER_20_60 ();
 sg13g2_decap_4 FILLER_20_103 ();
 sg13g2_fill_1 FILLER_20_107 ();
 sg13g2_fill_2 FILLER_20_125 ();
 sg13g2_fill_1 FILLER_20_127 ();
 sg13g2_fill_1 FILLER_20_186 ();
 sg13g2_fill_1 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_32 ();
 sg13g2_fill_2 FILLER_21_75 ();
 sg13g2_fill_2 FILLER_21_104 ();
 sg13g2_fill_2 FILLER_21_123 ();
 sg13g2_fill_1 FILLER_21_125 ();
 sg13g2_fill_2 FILLER_21_136 ();
 sg13g2_fill_1 FILLER_21_167 ();
 sg13g2_fill_2 FILLER_22_85 ();
 sg13g2_fill_2 FILLER_22_104 ();
 sg13g2_fill_2 FILLER_22_197 ();
 sg13g2_fill_1 FILLER_22_199 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_11 ();
 sg13g2_fill_1 FILLER_23_13 ();
 sg13g2_decap_8 FILLER_23_62 ();
 sg13g2_fill_2 FILLER_23_69 ();
 sg13g2_fill_1 FILLER_23_171 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_fill_1 FILLER_24_14 ();
 sg13g2_decap_4 FILLER_24_36 ();
 sg13g2_decap_4 FILLER_24_43 ();
 sg13g2_decap_4 FILLER_24_81 ();
 sg13g2_fill_2 FILLER_24_85 ();
 sg13g2_fill_1 FILLER_24_125 ();
 sg13g2_fill_1 FILLER_24_199 ();
 sg13g2_decap_8 FILLER_25_82 ();
 sg13g2_fill_1 FILLER_25_89 ();
 sg13g2_fill_2 FILLER_25_111 ();
 sg13g2_fill_1 FILLER_25_113 ();
 sg13g2_fill_1 FILLER_25_147 ();
 sg13g2_fill_2 FILLER_25_171 ();
 sg13g2_fill_1 FILLER_25_199 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_8 ();
 sg13g2_fill_1 FILLER_26_10 ();
 sg13g2_decap_4 FILLER_26_36 ();
 sg13g2_decap_8 FILLER_26_60 ();
 sg13g2_decap_4 FILLER_26_67 ();
 sg13g2_fill_2 FILLER_26_143 ();
 sg13g2_fill_2 FILLER_26_184 ();
 sg13g2_fill_1 FILLER_27_0 ();
 sg13g2_decap_4 FILLER_27_44 ();
 sg13g2_fill_2 FILLER_27_48 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_fill_2 FILLER_27_112 ();
 sg13g2_fill_1 FILLER_27_114 ();
 sg13g2_fill_2 FILLER_27_198 ();
 sg13g2_fill_1 FILLER_28_0 ();
 sg13g2_decap_4 FILLER_28_77 ();
 sg13g2_fill_1 FILLER_28_81 ();
 sg13g2_fill_2 FILLER_28_124 ();
 sg13g2_fill_2 FILLER_28_151 ();
 sg13g2_fill_1 FILLER_28_199 ();
 sg13g2_fill_1 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_27 ();
 sg13g2_fill_2 FILLER_29_58 ();
 sg13g2_fill_1 FILLER_29_60 ();
 sg13g2_decap_8 FILLER_29_78 ();
 sg13g2_fill_1 FILLER_29_85 ();
 sg13g2_fill_2 FILLER_29_103 ();
 sg13g2_fill_1 FILLER_29_105 ();
 sg13g2_fill_1 FILLER_29_123 ();
 sg13g2_fill_1 FILLER_29_145 ();
 sg13g2_fill_1 FILLER_29_163 ();
 sg13g2_fill_1 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_28 ();
 sg13g2_fill_1 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_71 ();
 sg13g2_decap_4 FILLER_30_78 ();
 sg13g2_fill_1 FILLER_30_82 ();
 sg13g2_fill_1 FILLER_30_104 ();
 sg13g2_fill_1 FILLER_30_122 ();
 sg13g2_fill_1 FILLER_30_164 ();
 sg13g2_fill_1 FILLER_30_199 ();
 sg13g2_fill_2 FILLER_31_17 ();
 sg13g2_decap_4 FILLER_31_74 ();
 sg13g2_fill_1 FILLER_31_140 ();
 sg13g2_fill_2 FILLER_31_162 ();
 sg13g2_fill_1 FILLER_31_164 ();
 sg13g2_fill_2 FILLER_31_198 ();
 sg13g2_fill_2 FILLER_32_21 ();
 sg13g2_fill_1 FILLER_32_44 ();
 sg13g2_decap_8 FILLER_32_88 ();
 sg13g2_fill_1 FILLER_32_137 ();
 sg13g2_fill_2 FILLER_32_163 ();
 sg13g2_fill_1 FILLER_32_165 ();
 sg13g2_fill_2 FILLER_32_187 ();
 sg13g2_fill_2 FILLER_32_197 ();
 sg13g2_fill_1 FILLER_32_199 ();
 sg13g2_fill_1 FILLER_33_33 ();
 sg13g2_fill_1 FILLER_33_175 ();
 sg13g2_fill_2 FILLER_33_197 ();
 sg13g2_fill_1 FILLER_33_199 ();
 sg13g2_fill_2 FILLER_34_34 ();
 sg13g2_fill_1 FILLER_34_77 ();
 sg13g2_fill_1 FILLER_34_146 ();
 sg13g2_fill_2 FILLER_34_197 ();
 sg13g2_fill_1 FILLER_34_199 ();
 sg13g2_fill_1 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_91 ();
 sg13g2_fill_2 FILLER_35_115 ();
 sg13g2_fill_1 FILLER_35_164 ();
 sg13g2_fill_2 FILLER_35_198 ();
 sg13g2_fill_2 FILLER_36_33 ();
 sg13g2_fill_1 FILLER_36_41 ();
 sg13g2_fill_2 FILLER_36_100 ();
 sg13g2_fill_1 FILLER_36_127 ();
 sg13g2_fill_2 FILLER_36_187 ();
 sg13g2_fill_2 FILLER_36_197 ();
 sg13g2_fill_1 FILLER_36_199 ();
 sg13g2_fill_1 FILLER_37_94 ();
 sg13g2_fill_2 FILLER_37_128 ();
 sg13g2_fill_1 FILLER_37_169 ();
 sg13g2_fill_2 FILLER_37_187 ();
 sg13g2_fill_2 FILLER_37_197 ();
 sg13g2_fill_1 FILLER_37_199 ();
 sg13g2_fill_1 FILLER_38_37 ();
 sg13g2_fill_2 FILLER_38_55 ();
 sg13g2_fill_1 FILLER_38_74 ();
 sg13g2_fill_1 FILLER_38_92 ();
 sg13g2_fill_1 FILLER_38_188 ();
 sg13g2_fill_2 FILLER_38_197 ();
 sg13g2_fill_1 FILLER_38_199 ();
 sg13g2_fill_1 FILLER_39_135 ();
 sg13g2_fill_2 FILLER_39_174 ();
 sg13g2_fill_1 FILLER_39_176 ();
 sg13g2_fill_2 FILLER_39_198 ();
 sg13g2_fill_2 FILLER_40_54 ();
 sg13g2_fill_2 FILLER_40_99 ();
 sg13g2_fill_2 FILLER_40_139 ();
 sg13g2_fill_1 FILLER_40_141 ();
 sg13g2_fill_1 FILLER_40_168 ();
 sg13g2_fill_2 FILLER_40_198 ();
 sg13g2_fill_2 FILLER_41_80 ();
 sg13g2_fill_1 FILLER_41_129 ();
 sg13g2_fill_2 FILLER_41_135 ();
 sg13g2_fill_2 FILLER_41_142 ();
 sg13g2_fill_2 FILLER_41_154 ();
 sg13g2_fill_2 FILLER_41_197 ();
 sg13g2_fill_1 FILLER_41_199 ();
 sg13g2_fill_2 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_128 ();
 sg13g2_fill_2 FILLER_42_160 ();
 sg13g2_fill_1 FILLER_42_162 ();
 sg13g2_fill_1 FILLER_42_188 ();
 sg13g2_fill_1 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_6 ();
 sg13g2_fill_1 FILLER_43_60 ();
 sg13g2_fill_2 FILLER_43_78 ();
 sg13g2_fill_2 FILLER_43_114 ();
 sg13g2_fill_2 FILLER_43_167 ();
 sg13g2_fill_2 FILLER_44_45 ();
 sg13g2_fill_2 FILLER_44_121 ();
 sg13g2_fill_1 FILLER_44_199 ();
 sg13g2_fill_1 FILLER_45_189 ();
 sg13g2_fill_2 FILLER_45_198 ();
 sg13g2_fill_2 FILLER_46_0 ();
 sg13g2_fill_2 FILLER_46_10 ();
 sg13g2_fill_2 FILLER_46_114 ();
 sg13g2_fill_2 FILLER_46_170 ();
 sg13g2_fill_1 FILLER_47_0 ();
 sg13g2_fill_2 FILLER_47_43 ();
 sg13g2_fill_1 FILLER_47_133 ();
 sg13g2_fill_2 FILLER_47_151 ();
 sg13g2_fill_2 FILLER_47_171 ();
 sg13g2_fill_2 FILLER_47_198 ();
 sg13g2_fill_2 FILLER_48_147 ();
 sg13g2_fill_1 FILLER_48_165 ();
 sg13g2_fill_1 FILLER_49_0 ();
 sg13g2_fill_2 FILLER_49_61 ();
 sg13g2_fill_2 FILLER_49_175 ();
 sg13g2_fill_1 FILLER_49_199 ();
 sg13g2_fill_1 FILLER_50_0 ();
 sg13g2_fill_1 FILLER_50_32 ();
 sg13g2_fill_1 FILLER_50_41 ();
 sg13g2_fill_2 FILLER_50_198 ();
 sg13g2_fill_1 FILLER_51_125 ();
 sg13g2_fill_1 FILLER_51_148 ();
 sg13g2_fill_2 FILLER_51_198 ();
 sg13g2_fill_1 FILLER_52_0 ();
 sg13g2_fill_2 FILLER_52_76 ();
 sg13g2_fill_1 FILLER_52_184 ();
 sg13g2_fill_1 FILLER_53_38 ();
 sg13g2_fill_2 FILLER_53_78 ();
 sg13g2_fill_2 FILLER_53_198 ();
endmodule
