module E_TT_IF (CLK_TT_PROJECT,
    ENA_TT_PROJECT,
    RST_N_TT_PROJECT,
    UIO_IN_TT_PROJECT0,
    UIO_IN_TT_PROJECT1,
    UIO_IN_TT_PROJECT2,
    UIO_IN_TT_PROJECT3,
    UIO_IN_TT_PROJECT4,
    UIO_IN_TT_PROJECT5,
    UIO_IN_TT_PROJECT6,
    UIO_IN_TT_PROJECT7,
    UIO_OE_TT_PROJECT0,
    UIO_OE_TT_PROJECT1,
    UIO_OE_TT_PROJECT2,
    UIO_OE_TT_PROJECT3,
    UIO_OE_TT_PROJECT4,
    UIO_OE_TT_PROJECT5,
    UIO_OE_TT_PROJECT6,
    UIO_OE_TT_PROJECT7,
    UIO_OUT_TT_PROJECT0,
    UIO_OUT_TT_PROJECT1,
    UIO_OUT_TT_PROJECT2,
    UIO_OUT_TT_PROJECT3,
    UIO_OUT_TT_PROJECT4,
    UIO_OUT_TT_PROJECT5,
    UIO_OUT_TT_PROJECT6,
    UIO_OUT_TT_PROJECT7,
    UI_IN_TT_PROJECT0,
    UI_IN_TT_PROJECT1,
    UI_IN_TT_PROJECT2,
    UI_IN_TT_PROJECT3,
    UI_IN_TT_PROJECT4,
    UI_IN_TT_PROJECT5,
    UI_IN_TT_PROJECT6,
    UI_IN_TT_PROJECT7,
    UO_OUT_TT_PROJECT0,
    UO_OUT_TT_PROJECT1,
    UO_OUT_TT_PROJECT2,
    UO_OUT_TT_PROJECT3,
    UO_OUT_TT_PROJECT4,
    UO_OUT_TT_PROJECT5,
    UO_OUT_TT_PROJECT6,
    UO_OUT_TT_PROJECT7,
    UserCLK,
    UserCLKo,
    VPWR,
    VGND,
    E1END,
    E2END,
    E2MID,
    E6END,
    EE4END,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N1END,
    N2BEG,
    N2BEGb,
    N2END,
    N2MID,
    N4BEG,
    N4END,
    S1BEG,
    S1END,
    S2BEG,
    S2BEGb,
    S2END,
    S2MID,
    S4BEG,
    S4END,
    W1BEG,
    W2BEG,
    W2BEGb,
    W6BEG,
    WW4BEG);
 output CLK_TT_PROJECT;
 output ENA_TT_PROJECT;
 output RST_N_TT_PROJECT;
 output UIO_IN_TT_PROJECT0;
 output UIO_IN_TT_PROJECT1;
 output UIO_IN_TT_PROJECT2;
 output UIO_IN_TT_PROJECT3;
 output UIO_IN_TT_PROJECT4;
 output UIO_IN_TT_PROJECT5;
 output UIO_IN_TT_PROJECT6;
 output UIO_IN_TT_PROJECT7;
 input UIO_OE_TT_PROJECT0;
 input UIO_OE_TT_PROJECT1;
 input UIO_OE_TT_PROJECT2;
 input UIO_OE_TT_PROJECT3;
 input UIO_OE_TT_PROJECT4;
 input UIO_OE_TT_PROJECT5;
 input UIO_OE_TT_PROJECT6;
 input UIO_OE_TT_PROJECT7;
 input UIO_OUT_TT_PROJECT0;
 input UIO_OUT_TT_PROJECT1;
 input UIO_OUT_TT_PROJECT2;
 input UIO_OUT_TT_PROJECT3;
 input UIO_OUT_TT_PROJECT4;
 input UIO_OUT_TT_PROJECT5;
 input UIO_OUT_TT_PROJECT6;
 input UIO_OUT_TT_PROJECT7;
 output UI_IN_TT_PROJECT0;
 output UI_IN_TT_PROJECT1;
 output UI_IN_TT_PROJECT2;
 output UI_IN_TT_PROJECT3;
 output UI_IN_TT_PROJECT4;
 output UI_IN_TT_PROJECT5;
 output UI_IN_TT_PROJECT6;
 output UI_IN_TT_PROJECT7;
 input UO_OUT_TT_PROJECT0;
 input UO_OUT_TT_PROJECT1;
 input UO_OUT_TT_PROJECT2;
 input UO_OUT_TT_PROJECT3;
 input UO_OUT_TT_PROJECT4;
 input UO_OUT_TT_PROJECT5;
 input UO_OUT_TT_PROJECT6;
 input UO_OUT_TT_PROJECT7;
 input UserCLK;
 output UserCLKo;
 inout VPWR;
 inout VGND;
 input [3:0] E1END;
 input [7:0] E2END;
 input [7:0] E2MID;
 input [11:0] E6END;
 input [15:0] EE4END;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 input [3:0] N1END;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 input [7:0] N2END;
 input [7:0] N2MID;
 output [15:0] N4BEG;
 input [15:0] N4END;
 output [3:0] S1BEG;
 input [3:0] S1END;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 input [7:0] S2END;
 input [7:0] S2MID;
 output [15:0] S4BEG;
 input [15:0] S4END;
 output [3:0] W1BEG;
 output [7:0] W2BEG;
 output [7:0] W2BEGb;
 output [11:0] W6BEG;
 output [15:0] WW4BEG;

 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit0.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit1.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit10.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit11.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit12.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit13.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit14.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit15.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit16.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit17.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit18.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit19.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit2.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit20.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit21.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit22.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit23.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit24.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit25.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit26.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit27.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit28.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit29.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit3.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit30.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit31.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit4.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit5.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit6.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit7.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit8.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame0_bit9.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit0.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit1.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit10.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit11.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit12.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit13.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit14.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit15.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit16.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit17.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit18.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit19.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit2.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit20.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit21.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit22.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit23.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit24.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit25.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit26.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit27.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit28.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit29.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit3.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit30.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit31.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit4.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit5.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit6.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit7.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit8.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame1_bit9.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit0.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit1.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit10.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit11.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit12.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit13.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit14.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit15.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit16.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit17.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit18.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit19.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit2.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit20.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit21.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit22.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit23.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit24.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit25.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit26.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit27.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit28.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit29.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit3.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit30.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit31.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit4.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit5.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit6.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit7.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit8.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame2_bit9.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit0.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit1.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit10.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit11.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit12.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit13.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit14.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit15.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit16.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit17.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit18.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit19.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit2.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit20.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit21.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit22.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit23.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit24.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit25.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit26.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit27.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit28.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit29.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit3.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit30.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit31.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit4.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit5.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit6.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit7.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit8.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame3_bit9.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit0.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit1.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit10.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit11.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit12.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit13.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit14.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit15.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit16.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit17.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit18.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit19.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit2.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit20.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit21.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit22.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit23.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit24.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit25.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit26.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit27.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit28.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit29.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit3.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit30.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit31.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit4.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit5.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit6.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit7.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit8.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame4_bit9.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit0.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit1.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit10.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit11.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit12.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit13.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit14.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit15.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit16.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit17.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit18.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit19.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit2.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit20.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit21.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit22.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit23.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit24.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit25.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit26.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit27.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit28.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit29.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit3.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit30.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit31.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit4.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit5.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit6.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit7.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit8.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame5_bit9.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit0.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit1.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit10.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit11.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit12.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit13.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit14.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit15.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit16.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit17.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit18.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit19.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit2.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit20.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit21.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit22.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit23.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit24.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit25.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit26.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit27.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit28.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit29.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit3.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit30.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit31.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit4.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit5.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit6.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit7.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit8.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame6_bit9.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit0.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit1.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit10.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit11.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit12.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit13.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit14.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit15.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit16.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit17.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit18.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit19.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit2.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit20.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit21.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit22.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit23.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit24.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit25.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit26.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit27.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit28.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit29.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit3.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit30.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit31.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit4.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit5.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit6.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit7.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit8.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame7_bit9.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame8_bit10.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame8_bit11.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame8_bit12.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame8_bit13.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame8_bit14.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame8_bit15.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame8_bit16.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame8_bit17.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame8_bit18.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame8_bit19.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame8_bit20.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame8_bit21.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame8_bit22.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame8_bit23.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame8_bit24.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame8_bit25.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame8_bit26.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame8_bit27.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame8_bit28.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame8_bit29.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame8_bit30.Q ;
 wire \Inst_E_TT_IF_ConfigMem.Inst_frame8_bit31.Q ;
 wire \Inst_E_TT_IF_switch_matrix.N1BEG0 ;
 wire \Inst_E_TT_IF_switch_matrix.N1BEG1 ;
 wire \Inst_E_TT_IF_switch_matrix.N1BEG2 ;
 wire \Inst_E_TT_IF_switch_matrix.N1BEG3 ;
 wire \Inst_E_TT_IF_switch_matrix.N2BEG0 ;
 wire \Inst_E_TT_IF_switch_matrix.N2BEG1 ;
 wire \Inst_E_TT_IF_switch_matrix.N2BEG2 ;
 wire \Inst_E_TT_IF_switch_matrix.N2BEG3 ;
 wire \Inst_E_TT_IF_switch_matrix.N2BEG4 ;
 wire \Inst_E_TT_IF_switch_matrix.N2BEG5 ;
 wire \Inst_E_TT_IF_switch_matrix.N2BEG6 ;
 wire \Inst_E_TT_IF_switch_matrix.N2BEG7 ;
 wire \Inst_E_TT_IF_switch_matrix.N4BEG0 ;
 wire \Inst_E_TT_IF_switch_matrix.N4BEG1 ;
 wire \Inst_E_TT_IF_switch_matrix.N4BEG2 ;
 wire \Inst_E_TT_IF_switch_matrix.N4BEG3 ;
 wire \Inst_E_TT_IF_switch_matrix.S1BEG0 ;
 wire \Inst_E_TT_IF_switch_matrix.S1BEG1 ;
 wire \Inst_E_TT_IF_switch_matrix.S1BEG2 ;
 wire \Inst_E_TT_IF_switch_matrix.S1BEG3 ;
 wire \Inst_E_TT_IF_switch_matrix.S2BEG0 ;
 wire \Inst_E_TT_IF_switch_matrix.S2BEG1 ;
 wire \Inst_E_TT_IF_switch_matrix.S2BEG2 ;
 wire \Inst_E_TT_IF_switch_matrix.S2BEG3 ;
 wire \Inst_E_TT_IF_switch_matrix.S2BEG4 ;
 wire \Inst_E_TT_IF_switch_matrix.S2BEG5 ;
 wire \Inst_E_TT_IF_switch_matrix.S2BEG6 ;
 wire \Inst_E_TT_IF_switch_matrix.S2BEG7 ;
 wire \Inst_E_TT_IF_switch_matrix.S4BEG0 ;
 wire \Inst_E_TT_IF_switch_matrix.S4BEG1 ;
 wire \Inst_E_TT_IF_switch_matrix.S4BEG2 ;
 wire \Inst_E_TT_IF_switch_matrix.S4BEG3 ;
 wire \Inst_E_TT_IF_switch_matrix.W1BEG0 ;
 wire \Inst_E_TT_IF_switch_matrix.W1BEG1 ;
 wire \Inst_E_TT_IF_switch_matrix.W1BEG2 ;
 wire \Inst_E_TT_IF_switch_matrix.W1BEG3 ;
 wire \Inst_E_TT_IF_switch_matrix.W2BEG0 ;
 wire \Inst_E_TT_IF_switch_matrix.W2BEG1 ;
 wire \Inst_E_TT_IF_switch_matrix.W2BEG2 ;
 wire \Inst_E_TT_IF_switch_matrix.W2BEG3 ;
 wire \Inst_E_TT_IF_switch_matrix.W2BEG4 ;
 wire \Inst_E_TT_IF_switch_matrix.W2BEG5 ;
 wire \Inst_E_TT_IF_switch_matrix.W2BEG6 ;
 wire \Inst_E_TT_IF_switch_matrix.W2BEG7 ;
 wire \Inst_E_TT_IF_switch_matrix.W2BEGb0 ;
 wire \Inst_E_TT_IF_switch_matrix.W2BEGb1 ;
 wire \Inst_E_TT_IF_switch_matrix.W2BEGb2 ;
 wire \Inst_E_TT_IF_switch_matrix.W2BEGb3 ;
 wire \Inst_E_TT_IF_switch_matrix.W2BEGb4 ;
 wire \Inst_E_TT_IF_switch_matrix.W2BEGb5 ;
 wire \Inst_E_TT_IF_switch_matrix.W2BEGb6 ;
 wire \Inst_E_TT_IF_switch_matrix.W2BEGb7 ;
 wire \Inst_E_TT_IF_switch_matrix.W6BEG0 ;
 wire \Inst_E_TT_IF_switch_matrix.W6BEG1 ;
 wire \Inst_E_TT_IF_switch_matrix.W6BEG10 ;
 wire \Inst_E_TT_IF_switch_matrix.W6BEG11 ;
 wire \Inst_E_TT_IF_switch_matrix.W6BEG2 ;
 wire \Inst_E_TT_IF_switch_matrix.W6BEG3 ;
 wire \Inst_E_TT_IF_switch_matrix.W6BEG4 ;
 wire \Inst_E_TT_IF_switch_matrix.W6BEG5 ;
 wire \Inst_E_TT_IF_switch_matrix.W6BEG6 ;
 wire \Inst_E_TT_IF_switch_matrix.W6BEG7 ;
 wire \Inst_E_TT_IF_switch_matrix.W6BEG8 ;
 wire \Inst_E_TT_IF_switch_matrix.W6BEG9 ;
 wire \Inst_E_TT_IF_switch_matrix.WW4BEG0 ;
 wire \Inst_E_TT_IF_switch_matrix.WW4BEG1 ;
 wire \Inst_E_TT_IF_switch_matrix.WW4BEG10 ;
 wire \Inst_E_TT_IF_switch_matrix.WW4BEG11 ;
 wire \Inst_E_TT_IF_switch_matrix.WW4BEG12 ;
 wire \Inst_E_TT_IF_switch_matrix.WW4BEG13 ;
 wire \Inst_E_TT_IF_switch_matrix.WW4BEG14 ;
 wire \Inst_E_TT_IF_switch_matrix.WW4BEG15 ;
 wire \Inst_E_TT_IF_switch_matrix.WW4BEG2 ;
 wire \Inst_E_TT_IF_switch_matrix.WW4BEG3 ;
 wire \Inst_E_TT_IF_switch_matrix.WW4BEG4 ;
 wire \Inst_E_TT_IF_switch_matrix.WW4BEG5 ;
 wire \Inst_E_TT_IF_switch_matrix.WW4BEG6 ;
 wire \Inst_E_TT_IF_switch_matrix.WW4BEG7 ;
 wire \Inst_E_TT_IF_switch_matrix.WW4BEG8 ;
 wire \Inst_E_TT_IF_switch_matrix.WW4BEG9 ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire clknet_0_UserCLK;
 wire clknet_1_0__leaf_UserCLK;
 wire clknet_1_1__leaf_UserCLK;

 sg13g2_inv_1 _209_ (.VDD(VPWR),
    .Y(_000_),
    .A(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit5.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _210_ (.VDD(VPWR),
    .Y(_001_),
    .A(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit6.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _211_ (.VDD(VPWR),
    .Y(_002_),
    .A(S1END[3]),
    .VSS(VGND));
 sg13g2_inv_1 _212_ (.VDD(VPWR),
    .Y(_003_),
    .A(S1END[2]),
    .VSS(VGND));
 sg13g2_inv_1 _213_ (.VDD(VPWR),
    .Y(_004_),
    .A(S1END[1]),
    .VSS(VGND));
 sg13g2_inv_1 _214_ (.VDD(VPWR),
    .Y(_005_),
    .A(S1END[0]),
    .VSS(VGND));
 sg13g2_inv_1 _215_ (.VDD(VPWR),
    .Y(_006_),
    .A(EE4END[1]),
    .VSS(VGND));
 sg13g2_inv_1 _216_ (.VDD(VPWR),
    .Y(_007_),
    .A(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit10.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _217_ (.VDD(VPWR),
    .Y(_008_),
    .A(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit18.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _218_ (.VDD(VPWR),
    .Y(_009_),
    .A(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit15.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _219_ (.VDD(VPWR),
    .Y(_010_),
    .A(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit16.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _220_ (.VDD(VPWR),
    .Y(_011_),
    .A(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit6.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _221_ (.VDD(VPWR),
    .Y(_012_),
    .A(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit7.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _222_ (.VDD(VPWR),
    .Y(_013_),
    .A(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit12.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _223_ (.VDD(VPWR),
    .Y(_014_),
    .A(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit13.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _224_ (.VDD(VPWR),
    .Y(_015_),
    .A(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit5.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _225_ (.VDD(VPWR),
    .Y(_016_),
    .A(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit6.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _226_ (.VDD(VPWR),
    .Y(_017_),
    .A(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit7.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _227_ (.VDD(VPWR),
    .Y(_018_),
    .A(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit2.Q ),
    .VSS(VGND));
 sg13g2_inv_1 _228_ (.VDD(VPWR),
    .Y(_019_),
    .A(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit3.Q ),
    .VSS(VGND));
 sg13g2_mux2_1 _229_ (.A0(E2END[1]),
    .A1(E2END[2]),
    .S(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _230_ (.Y(_021_),
    .A(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit5.Q ),
    .B(_020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _231_ (.A0(E2MID[3]),
    .A1(E2MID[6]),
    .S(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _232_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_000_),
    .A2(_022_),
    .Y(_023_),
    .B1(_001_));
 sg13g2_mux2_1 _233_ (.A0(N2MID[6]),
    .A1(N2END[2]),
    .S(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit4.Q ),
    .X(_024_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _234_ (.Y(_025_),
    .B(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit4.Q ),
    .A_N(E2MID[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _235_ (.B1(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit5.Q ),
    .VDD(VPWR),
    .Y(_026_),
    .VSS(VGND),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit4.Q ),
    .A2(N2END[3]));
 sg13g2_nand2b_1 _236_ (.Y(_027_),
    .B(_025_),
    .A_N(_026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _237_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_000_),
    .A2(_024_),
    .Y(_028_),
    .B1(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit6.Q ));
 sg13g2_a221oi_1 _238_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_028_),
    .C1(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit7.Q ),
    .B1(_027_),
    .A1(_021_),
    .Y(_029_),
    .A2(_023_));
 sg13g2_nor2_1 _239_ (.A(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit5.Q ),
    .B(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit6.Q ),
    .Y(_030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _240_ (.A(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit6.Q ),
    .B_N(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit5.Q ),
    .Y(_031_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _241_ (.A(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit5.Q ),
    .B_N(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit6.Q ),
    .Y(_032_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _242_ (.Y(_033_),
    .B1(_032_),
    .B2(S2END[2]),
    .A2(_030_),
    .A1(E2END[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _243_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(E2END[5]),
    .A2(_031_),
    .Y(_034_),
    .B1(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit4.Q ));
 sg13g2_o21ai_1 _244_ (.B1(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit6.Q ),
    .VDD(VPWR),
    .Y(_035_),
    .VSS(VGND),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit5.Q ),
    .A2(S2END[3]));
 sg13g2_a22oi_1 _245_ (.Y(_036_),
    .B1(_030_),
    .B2(E2END[4]),
    .A2(S2MID[0]),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _246_ (.A(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit4.Q ),
    .B(_035_),
    .X(_037_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _247_ (.Y(_038_),
    .B1(_036_),
    .B2(_037_),
    .A2(_034_),
    .A1(_033_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _248_ (.A2(_038_),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit7.Q ),
    .B1(_029_),
    .X(RST_N_TT_PROJECT),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _249_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit22.Q ),
    .A0(N2MID[7]),
    .A1(N2END[7]),
    .A2(S2MID[7]),
    .A3(S2END[7]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit23.Q ),
    .X(_039_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _250_ (.VDD(VPWR),
    .Y(_040_),
    .A(_039_),
    .VSS(VGND));
 sg13g2_mux4_1 _251_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit6.Q ),
    .A0(N1END[3]),
    .A1(N4END[3]),
    .A2(S1END[3]),
    .A3(S4END[3]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit7.Q ),
    .X(_041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _252_ (.A(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit31.Q ),
    .B_N(EE4END[15]),
    .Y(_042_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _253_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit31.Q ),
    .A2(_041_),
    .Y(_043_),
    .B1(_042_));
 sg13g2_nand3b_1 _254_ (.B(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit0.Q ),
    .C(_039_),
    .Y(_044_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit31.Q ));
 sg13g2_o21ai_1 _255_ (.B1(_044_),
    .VDD(VPWR),
    .Y(_045_),
    .VSS(VGND),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit0.Q ),
    .A2(_043_));
 sg13g2_mux4_1 _256_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit31.Q ),
    .A0(E1END[3]),
    .A1(E2MID[7]),
    .A2(E2END[7]),
    .A3(EE4END[7]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit0.Q ),
    .X(_046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _257_ (.A0(_046_),
    .A1(_045_),
    .S(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit1.Q ),
    .X(UIO_IN_TT_PROJECT7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _258_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit20.Q ),
    .A0(N2MID[6]),
    .A1(N2END[6]),
    .A2(S2MID[6]),
    .A3(S2END[6]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit21.Q ),
    .X(_047_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _259_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit4.Q ),
    .A0(N1END[2]),
    .A1(N4END[2]),
    .A2(S1END[2]),
    .A3(S4END[2]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit5.Q ),
    .X(_048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _260_ (.A(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit28.Q ),
    .B_N(EE4END[14]),
    .Y(_049_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _261_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit28.Q ),
    .A2(_048_),
    .Y(_050_),
    .B1(_049_));
 sg13g2_nand3b_1 _262_ (.B(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit29.Q ),
    .C(_047_),
    .Y(_051_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit28.Q ));
 sg13g2_o21ai_1 _263_ (.B1(_051_),
    .VDD(VPWR),
    .Y(_052_),
    .VSS(VGND),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit29.Q ),
    .A2(_050_));
 sg13g2_mux4_1 _264_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit29.Q ),
    .A0(E1END[2]),
    .A1(E2END[6]),
    .A2(E2MID[6]),
    .A3(EE4END[6]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit28.Q ),
    .X(_053_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _265_ (.A0(_053_),
    .A1(_052_),
    .S(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit30.Q ),
    .X(UIO_IN_TT_PROJECT6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _266_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit2.Q ),
    .A0(N1END[1]),
    .A1(N4END[1]),
    .A2(S1END[1]),
    .A3(S4END[1]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit3.Q ),
    .X(_054_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _267_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit18.Q ),
    .A0(N2MID[5]),
    .A1(N2END[5]),
    .A2(S2MID[5]),
    .A3(S2END[5]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit19.Q ),
    .X(_055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _268_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit25.Q ),
    .A0(E1END[1]),
    .A1(E2MID[5]),
    .A2(E2END[5]),
    .A3(EE4END[5]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit26.Q ),
    .X(_056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _269_ (.B(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit26.Q ),
    .C(_055_),
    .Y(_057_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit25.Q ));
 sg13g2_nor2b_1 _270_ (.A(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit25.Q ),
    .B_N(EE4END[13]),
    .Y(_058_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _271_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit25.Q ),
    .A2(_054_),
    .Y(_059_),
    .B1(_058_));
 sg13g2_o21ai_1 _272_ (.B1(_057_),
    .VDD(VPWR),
    .Y(_060_),
    .VSS(VGND),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit26.Q ),
    .A2(_059_));
 sg13g2_mux2_1 _273_ (.A0(_056_),
    .A1(_060_),
    .S(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit27.Q ),
    .X(UIO_IN_TT_PROJECT5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _274_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit0.Q ),
    .A0(N1END[0]),
    .A1(N4END[0]),
    .A2(S1END[0]),
    .A3(S4END[0]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit1.Q ),
    .X(_061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _275_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit16.Q ),
    .A0(N2MID[4]),
    .A1(N2END[4]),
    .A2(S2MID[4]),
    .A3(S2END[4]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit17.Q ),
    .X(_062_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _276_ (.VDD(VPWR),
    .Y(_063_),
    .A(_062_),
    .VSS(VGND));
 sg13g2_nor2b_1 _277_ (.A(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit22.Q ),
    .B_N(EE4END[12]),
    .Y(_064_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _278_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit22.Q ),
    .A2(_061_),
    .Y(_065_),
    .B1(_064_));
 sg13g2_nand3b_1 _279_ (.B(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit23.Q ),
    .C(_062_),
    .Y(_066_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit22.Q ));
 sg13g2_o21ai_1 _280_ (.B1(_066_),
    .VDD(VPWR),
    .Y(_067_),
    .VSS(VGND),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit23.Q ),
    .A2(_065_));
 sg13g2_mux4_1 _281_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit22.Q ),
    .A0(E1END[0]),
    .A1(E2MID[4]),
    .A2(E2END[4]),
    .A3(EE4END[4]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit23.Q ),
    .X(_068_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _282_ (.A0(_068_),
    .A1(_067_),
    .S(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit24.Q ),
    .X(UIO_IN_TT_PROJECT4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _283_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit30.Q ),
    .A0(N1END[3]),
    .A1(N4END[3]),
    .A2(S1END[3]),
    .A3(S4END[3]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit31.Q ),
    .X(_069_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _284_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit15.Q ),
    .A0(N2MID[3]),
    .A1(S2MID[3]),
    .A2(N2END[3]),
    .A3(S2END[3]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit14.Q ),
    .X(_070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _285_ (.B(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit20.Q ),
    .C(_070_),
    .Y(_071_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit19.Q ));
 sg13g2_nor2b_1 _286_ (.A(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit19.Q ),
    .B_N(E6END[11]),
    .Y(_072_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _287_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit19.Q ),
    .A2(_069_),
    .Y(_073_),
    .B1(_072_));
 sg13g2_o21ai_1 _288_ (.B1(_071_),
    .VDD(VPWR),
    .Y(_074_),
    .VSS(VGND),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit20.Q ),
    .A2(_073_));
 sg13g2_mux4_1 _289_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit19.Q ),
    .A0(E2MID[3]),
    .A1(E2END[3]),
    .A2(EE4END[3]),
    .A3(EE4END[11]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit20.Q ),
    .X(_075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _290_ (.A0(_075_),
    .A1(_074_),
    .S(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit21.Q ),
    .X(UIO_IN_TT_PROJECT3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _291_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit28.Q ),
    .A0(N1END[2]),
    .A1(N4END[2]),
    .A2(S1END[2]),
    .A3(S4END[2]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit29.Q ),
    .X(_076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _292_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit13.Q ),
    .A0(N2MID[2]),
    .A1(S2MID[2]),
    .A2(N2END[2]),
    .A3(S2END[2]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit12.Q ),
    .X(_077_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _293_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit17.Q ),
    .A0(E2MID[2]),
    .A1(EE4END[2]),
    .A2(E2END[2]),
    .A3(EE4END[10]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit16.Q ),
    .X(_078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _294_ (.B(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit17.Q ),
    .C(_077_),
    .Y(_079_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit16.Q ));
 sg13g2_nor2b_1 _295_ (.A(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit16.Q ),
    .B_N(E6END[10]),
    .Y(_080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _296_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit16.Q ),
    .A2(_076_),
    .Y(_081_),
    .B1(_080_));
 sg13g2_o21ai_1 _297_ (.B1(_079_),
    .VDD(VPWR),
    .Y(_082_),
    .VSS(VGND),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit17.Q ),
    .A2(_081_));
 sg13g2_mux2_1 _298_ (.A0(_078_),
    .A1(_082_),
    .S(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit18.Q ),
    .X(UIO_IN_TT_PROJECT2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _299_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit26.Q ),
    .A0(N1END[1]),
    .A1(N4END[1]),
    .A2(S1END[1]),
    .A3(S4END[1]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit27.Q ),
    .X(_083_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _300_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit10.Q ),
    .A0(N2MID[1]),
    .A1(N2END[1]),
    .A2(S2MID[1]),
    .A3(S2END[1]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit11.Q ),
    .X(_084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _301_ (.A(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit13.Q ),
    .B_N(E6END[9]),
    .Y(_085_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _302_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit13.Q ),
    .A2(_083_),
    .Y(_086_),
    .B1(_085_));
 sg13g2_nand3b_1 _303_ (.B(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit14.Q ),
    .C(_084_),
    .Y(_087_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit13.Q ));
 sg13g2_o21ai_1 _304_ (.B1(_087_),
    .VDD(VPWR),
    .Y(_088_),
    .VSS(VGND),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit14.Q ),
    .A2(_086_));
 sg13g2_mux4_1 _305_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit14.Q ),
    .A0(E2MID[1]),
    .A1(EE4END[1]),
    .A2(E2END[1]),
    .A3(EE4END[9]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit13.Q ),
    .X(_089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _306_ (.A0(_089_),
    .A1(_088_),
    .S(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit15.Q ),
    .X(UIO_IN_TT_PROJECT1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _307_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit8.Q ),
    .A0(N2MID[0]),
    .A1(N2END[0]),
    .A2(S2MID[0]),
    .A3(S2END[0]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit9.Q ),
    .X(_090_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _308_ (.VDD(VPWR),
    .Y(_091_),
    .A(_090_),
    .VSS(VGND));
 sg13g2_mux4_1 _309_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit24.Q ),
    .A0(N1END[0]),
    .A1(N4END[0]),
    .A2(S1END[0]),
    .A3(S4END[0]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit25.Q ),
    .X(_092_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _310_ (.VDD(VPWR),
    .Y(_093_),
    .A(_092_),
    .VSS(VGND));
 sg13g2_nand3_1 _311_ (.B(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit11.Q ),
    .C(_090_),
    .A(_007_),
    .Y(_094_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _312_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_095_),
    .B(E6END[8]),
    .A(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit10.Q ));
 sg13g2_o21ai_1 _313_ (.B1(_095_),
    .VDD(VPWR),
    .Y(_096_),
    .VSS(VGND),
    .A1(_007_),
    .A2(_092_));
 sg13g2_o21ai_1 _314_ (.B1(_094_),
    .VDD(VPWR),
    .Y(_097_),
    .VSS(VGND),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit11.Q ),
    .A2(_096_));
 sg13g2_mux4_1 _315_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit10.Q ),
    .A0(E2MID[0]),
    .A1(E2END[0]),
    .A2(EE4END[0]),
    .A3(EE4END[8]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit11.Q ),
    .X(_098_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _316_ (.A0(_098_),
    .A1(_097_),
    .S(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit12.Q ),
    .X(UIO_IN_TT_PROJECT0),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _317_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit22.Q ),
    .A0(N1END[3]),
    .A1(N4END[3]),
    .A2(S1END[3]),
    .A3(S4END[3]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit23.Q ),
    .X(_099_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _318_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit7.Q ),
    .A0(E2MID[7]),
    .A1(E2END[7]),
    .A2(EE4END[7]),
    .A3(EE4END[15]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit8.Q ),
    .X(_100_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _319_ (.B(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit8.Q ),
    .C(_039_),
    .Y(_101_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit7.Q ));
 sg13g2_nor2b_1 _320_ (.A(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit7.Q ),
    .B_N(E6END[7]),
    .Y(_102_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _321_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit7.Q ),
    .A2(_099_),
    .Y(_103_),
    .B1(_102_));
 sg13g2_o21ai_1 _322_ (.B1(_101_),
    .VDD(VPWR),
    .Y(_104_),
    .VSS(VGND),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit8.Q ),
    .A2(_103_));
 sg13g2_mux2_1 _323_ (.A0(_100_),
    .A1(_104_),
    .S(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit9.Q ),
    .X(UI_IN_TT_PROJECT7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _324_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit20.Q ),
    .A0(N1END[2]),
    .A1(N4END[2]),
    .A2(S1END[2]),
    .A3(S4END[2]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit21.Q ),
    .X(_105_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _325_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit4.Q ),
    .A0(E2MID[6]),
    .A1(E2END[6]),
    .A2(EE4END[6]),
    .A3(EE4END[14]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit5.Q ),
    .X(_106_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _326_ (.B(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit5.Q ),
    .C(_047_),
    .Y(_107_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit4.Q ));
 sg13g2_nor2b_1 _327_ (.A(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit4.Q ),
    .B_N(E6END[6]),
    .Y(_108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _328_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit4.Q ),
    .A2(_105_),
    .Y(_109_),
    .B1(_108_));
 sg13g2_o21ai_1 _329_ (.B1(_107_),
    .VDD(VPWR),
    .Y(_110_),
    .VSS(VGND),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit5.Q ),
    .A2(_109_));
 sg13g2_mux2_1 _330_ (.A0(_106_),
    .A1(_110_),
    .S(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit6.Q ),
    .X(UI_IN_TT_PROJECT6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _331_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit18.Q ),
    .A0(N1END[1]),
    .A1(N4END[1]),
    .A2(S1END[1]),
    .A3(S4END[1]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit19.Q ),
    .X(_111_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _332_ (.A(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit1.Q ),
    .B_N(E6END[5]),
    .Y(_112_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _333_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit1.Q ),
    .A2(_111_),
    .Y(_113_),
    .B1(_112_));
 sg13g2_nand3b_1 _334_ (.B(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit2.Q ),
    .C(_055_),
    .Y(_114_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit1.Q ));
 sg13g2_o21ai_1 _335_ (.B1(_114_),
    .VDD(VPWR),
    .Y(_115_),
    .VSS(VGND),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit2.Q ),
    .A2(_113_));
 sg13g2_mux4_1 _336_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit2.Q ),
    .A0(E2MID[5]),
    .A1(EE4END[5]),
    .A2(E2END[5]),
    .A3(EE4END[13]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit1.Q ),
    .X(_116_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _337_ (.A0(_116_),
    .A1(_115_),
    .S(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit3.Q ),
    .X(UI_IN_TT_PROJECT5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _338_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit16.Q ),
    .A0(N1END[0]),
    .A1(N4END[0]),
    .A2(S1END[0]),
    .A3(S4END[0]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit17.Q ),
    .X(_117_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _339_ (.A(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit30.Q ),
    .B_N(E6END[4]),
    .Y(_118_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _340_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit30.Q ),
    .A2(_117_),
    .Y(_119_),
    .B1(_118_));
 sg13g2_nand3b_1 _341_ (.B(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit31.Q ),
    .C(_062_),
    .Y(_120_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit30.Q ));
 sg13g2_o21ai_1 _342_ (.B1(_120_),
    .VDD(VPWR),
    .Y(_121_),
    .VSS(VGND),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit31.Q ),
    .A2(_119_));
 sg13g2_mux4_1 _343_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit31.Q ),
    .A0(E2MID[4]),
    .A1(EE4END[4]),
    .A2(E2END[4]),
    .A3(EE4END[12]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit30.Q ),
    .X(_122_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _344_ (.A0(_122_),
    .A1(_121_),
    .S(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit0.Q ),
    .X(UI_IN_TT_PROJECT4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _345_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit14.Q ),
    .A0(N1END[3]),
    .A1(N4END[3]),
    .A2(S1END[3]),
    .A3(S4END[3]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit15.Q ),
    .X(_123_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _346_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit27.Q ),
    .A0(E2MID[3]),
    .A1(E2END[3]),
    .A2(EE4END[3]),
    .A3(EE4END[11]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit28.Q ),
    .X(_124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _347_ (.B(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit28.Q ),
    .C(_070_),
    .Y(_125_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit27.Q ));
 sg13g2_nor2b_1 _348_ (.A(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit27.Q ),
    .B_N(E6END[3]),
    .Y(_126_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _349_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit27.Q ),
    .A2(_123_),
    .Y(_127_),
    .B1(_126_));
 sg13g2_o21ai_1 _350_ (.B1(_125_),
    .VDD(VPWR),
    .Y(_128_),
    .VSS(VGND),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit28.Q ),
    .A2(_127_));
 sg13g2_mux2_1 _351_ (.A0(_124_),
    .A1(_128_),
    .S(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit29.Q ),
    .X(UI_IN_TT_PROJECT3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _352_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit12.Q ),
    .A0(N1END[2]),
    .A1(N4END[2]),
    .A2(S1END[2]),
    .A3(S4END[2]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit13.Q ),
    .X(_129_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _353_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit25.Q ),
    .A0(E2MID[2]),
    .A1(EE4END[2]),
    .A2(E2END[2]),
    .A3(EE4END[10]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit24.Q ),
    .X(_130_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _354_ (.B(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit25.Q ),
    .C(_077_),
    .Y(_131_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit24.Q ));
 sg13g2_nor2b_1 _355_ (.A(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit24.Q ),
    .B_N(E6END[2]),
    .Y(_132_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _356_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit24.Q ),
    .A2(_129_),
    .Y(_133_),
    .B1(_132_));
 sg13g2_o21ai_1 _357_ (.B1(_131_),
    .VDD(VPWR),
    .Y(_134_),
    .VSS(VGND),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit25.Q ),
    .A2(_133_));
 sg13g2_mux2_1 _358_ (.A0(_130_),
    .A1(_134_),
    .S(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit26.Q ),
    .X(UI_IN_TT_PROJECT2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _359_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit10.Q ),
    .A0(N1END[1]),
    .A1(N4END[1]),
    .A2(S1END[1]),
    .A3(S4END[1]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit11.Q ),
    .X(_135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _360_ (.A(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit21.Q ),
    .B_N(E6END[1]),
    .Y(_136_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _361_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit21.Q ),
    .A2(_135_),
    .Y(_137_),
    .B1(_136_));
 sg13g2_nand3b_1 _362_ (.B(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit22.Q ),
    .C(_084_),
    .Y(_138_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit21.Q ));
 sg13g2_o21ai_1 _363_ (.B1(_138_),
    .VDD(VPWR),
    .Y(_139_),
    .VSS(VGND),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit22.Q ),
    .A2(_137_));
 sg13g2_mux4_1 _364_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit22.Q ),
    .A0(E2MID[1]),
    .A1(EE4END[1]),
    .A2(E2END[1]),
    .A3(EE4END[9]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit21.Q ),
    .X(_140_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _365_ (.A0(_140_),
    .A1(_139_),
    .S(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit23.Q ),
    .X(UI_IN_TT_PROJECT1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _366_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit8.Q ),
    .A0(N1END[0]),
    .A1(N4END[0]),
    .A2(S1END[0]),
    .A3(S4END[0]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit9.Q ),
    .X(_141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _367_ (.B(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit19.Q ),
    .C(_090_),
    .A(_008_),
    .Y(_142_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _368_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_143_),
    .B(E6END[0]),
    .A(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit18.Q ));
 sg13g2_o21ai_1 _369_ (.B1(_143_),
    .VDD(VPWR),
    .Y(_144_),
    .VSS(VGND),
    .A1(_008_),
    .A2(_141_));
 sg13g2_o21ai_1 _370_ (.B1(_142_),
    .VDD(VPWR),
    .Y(_145_),
    .VSS(VGND),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit19.Q ),
    .A2(_144_));
 sg13g2_mux4_1 _371_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit18.Q ),
    .A0(E2MID[0]),
    .A1(E2END[0]),
    .A2(EE4END[0]),
    .A3(EE4END[8]),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit19.Q ),
    .X(_146_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _372_ (.A0(_146_),
    .A1(_145_),
    .S(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit20.Q ),
    .X(UI_IN_TT_PROJECT0),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _373_ (.B1(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit15.Q ),
    .VDD(VPWR),
    .Y(_147_),
    .VSS(VGND),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit17.Q ),
    .A2(_123_));
 sg13g2_a21o_1 _374_ (.A2(_040_),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit17.Q ),
    .B1(_147_),
    .X(_148_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _375_ (.A0(E6END[7]),
    .A1(_041_),
    .S(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit17.Q ),
    .X(_149_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _376_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_009_),
    .A2(_149_),
    .Y(_150_),
    .B1(_010_));
 sg13g2_mux4_1 _377_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit15.Q ),
    .A0(E1END[3]),
    .A1(EE4END[15]),
    .A2(_099_),
    .A3(_069_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit17.Q ),
    .X(_151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _378_ (.A(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit16.Q ),
    .B(_151_),
    .Y(_152_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _379_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_148_),
    .A2(_150_),
    .Y(\Inst_E_TT_IF_switch_matrix.S4BEG3 ),
    .B1(_152_));
 sg13g2_mux4_1 _380_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit12.Q ),
    .A0(E1END[2]),
    .A1(EE4END[14]),
    .A2(E6END[6]),
    .A3(_129_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit13.Q ),
    .X(_153_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _381_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit12.Q ),
    .A0(_105_),
    .A1(_076_),
    .A2(_048_),
    .A3(_047_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit13.Q ),
    .X(_154_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _382_ (.A0(_153_),
    .A1(_154_),
    .S(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit14.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.S4BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _383_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit9.Q ),
    .A0(E1END[1]),
    .A1(EE4END[13]),
    .A2(E6END[5]),
    .A3(_135_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit10.Q ),
    .X(_155_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _384_ (.Y(_156_),
    .B(_155_),
    .A_N(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _385_ (.A0(_111_),
    .A1(_083_),
    .S(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit9.Q ),
    .X(_157_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _386_ (.Y(_158_),
    .B(_054_),
    .A_N(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _387_ (.Y(_159_),
    .A(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit9.Q ),
    .B(_055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _388_ (.X(_160_),
    .A(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit10.Q ),
    .B(_158_),
    .C(_159_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _389_ (.B1(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit11.Q ),
    .VDD(VPWR),
    .Y(_161_),
    .VSS(VGND),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit10.Q ),
    .A2(_157_));
 sg13g2_o21ai_1 _390_ (.B1(_156_),
    .VDD(VPWR),
    .Y(\Inst_E_TT_IF_switch_matrix.S4BEG1 ),
    .VSS(VGND),
    .A1(_160_),
    .A2(_161_));
 sg13g2_o21ai_1 _391_ (.B1(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit6.Q ),
    .VDD(VPWR),
    .Y(_162_),
    .VSS(VGND),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit8.Q ),
    .A2(_141_));
 sg13g2_a21o_1 _392_ (.A2(_063_),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit8.Q ),
    .B1(_162_),
    .X(_163_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _393_ (.A0(E6END[4]),
    .A1(_061_),
    .S(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit8.Q ),
    .X(_164_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _394_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_011_),
    .A2(_164_),
    .Y(_165_),
    .B1(_012_));
 sg13g2_o21ai_1 _395_ (.B1(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit6.Q ),
    .VDD(VPWR),
    .Y(_166_),
    .VSS(VGND),
    .A1(EE4END[12]),
    .A2(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit8.Q ));
 sg13g2_a21o_1 _396_ (.A2(_093_),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit8.Q ),
    .B1(_166_),
    .X(_167_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _397_ (.A0(E1END[0]),
    .A1(_117_),
    .S(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit8.Q ),
    .X(_168_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _398_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_011_),
    .A2(_168_),
    .Y(_169_),
    .B1(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit7.Q ));
 sg13g2_a22oi_1 _399_ (.Y(\Inst_E_TT_IF_switch_matrix.S4BEG0 ),
    .B1(_167_),
    .B2(_169_),
    .A2(_165_),
    .A1(_163_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _400_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit11.Q ),
    .A0(E1END[3]),
    .A1(EE4END[3]),
    .A2(E6END[11]),
    .A3(_123_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit12.Q ),
    .X(_170_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _401_ (.Y(_171_),
    .B(_099_),
    .A_N(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _402_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit11.Q ),
    .A2(_069_),
    .Y(_172_),
    .B1(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit12.Q ));
 sg13g2_nand2b_1 _403_ (.Y(_173_),
    .B(_041_),
    .A_N(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _404_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit11.Q ),
    .A2(_070_),
    .Y(_174_),
    .B1(_013_));
 sg13g2_a221oi_1 _405_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_174_),
    .C1(_014_),
    .B1(_173_),
    .A1(_171_),
    .Y(_175_),
    .A2(_172_));
 sg13g2_a21o_1 _406_ (.A2(_170_),
    .A1(_014_),
    .B1(_175_),
    .X(\Inst_E_TT_IF_switch_matrix.N4BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _407_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit8.Q ),
    .A0(E1END[2]),
    .A1(EE4END[2]),
    .A2(E6END[10]),
    .A3(_129_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit9.Q ),
    .X(_176_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _408_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit8.Q ),
    .A0(_105_),
    .A1(_076_),
    .A2(_048_),
    .A3(_077_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit9.Q ),
    .X(_177_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _409_ (.A0(_176_),
    .A1(_177_),
    .S(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit10.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.N4BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _410_ (.A(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit7.Q ),
    .B(_135_),
    .Y(_178_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _411_ (.B1(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit5.Q ),
    .VDD(VPWR),
    .Y(_179_),
    .VSS(VGND),
    .A1(_017_),
    .A2(_084_));
 sg13g2_or2_1 _412_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_180_),
    .B(_179_),
    .A(_178_));
 sg13g2_mux2_1 _413_ (.A0(E6END[9]),
    .A1(_054_),
    .S(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit7.Q ),
    .X(_181_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _414_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_015_),
    .A2(_181_),
    .Y(_182_),
    .B1(_016_));
 sg13g2_a21oi_1 _415_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_006_),
    .A2(_017_),
    .Y(_183_),
    .B1(_015_));
 sg13g2_o21ai_1 _416_ (.B1(_183_),
    .VDD(VPWR),
    .Y(_184_),
    .VSS(VGND),
    .A1(_017_),
    .A2(_083_));
 sg13g2_mux2_1 _417_ (.A0(E1END[1]),
    .A1(_111_),
    .S(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit7.Q ),
    .X(_185_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _418_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_015_),
    .A2(_185_),
    .Y(_186_),
    .B1(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit6.Q ));
 sg13g2_a22oi_1 _419_ (.Y(\Inst_E_TT_IF_switch_matrix.N4BEG1 ),
    .B1(_184_),
    .B2(_186_),
    .A2(_182_),
    .A1(_180_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _420_ (.B1(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit2.Q ),
    .VDD(VPWR),
    .Y(_187_),
    .VSS(VGND),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit4.Q ),
    .A2(_141_));
 sg13g2_a21o_1 _421_ (.A2(_091_),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit4.Q ),
    .B1(_187_),
    .X(_188_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _422_ (.A0(E6END[8]),
    .A1(_061_),
    .S(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit4.Q ),
    .X(_189_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _423_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_018_),
    .A2(_189_),
    .Y(_190_),
    .B1(_019_));
 sg13g2_mux2_1 _424_ (.A0(E1END[0]),
    .A1(_117_),
    .S(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit4.Q ),
    .X(_191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _425_ (.B1(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit2.Q ),
    .VDD(VPWR),
    .Y(_192_),
    .VSS(VGND),
    .A1(EE4END[0]),
    .A2(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit4.Q ));
 sg13g2_a21o_1 _426_ (.A2(_093_),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit4.Q ),
    .B1(_192_),
    .X(_193_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _427_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_018_),
    .A2(_191_),
    .Y(_194_),
    .B1(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit3.Q ));
 sg13g2_a22oi_1 _428_ (.Y(\Inst_E_TT_IF_switch_matrix.N4BEG0 ),
    .B1(_193_),
    .B2(_194_),
    .A2(_190_),
    .A1(_188_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _429_ (.B1(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit2.Q ),
    .VDD(VPWR),
    .Y(_195_),
    .VSS(VGND),
    .A1(E2MID[6]),
    .A2(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit3.Q ));
 sg13g2_nand2b_1 _430_ (.Y(_196_),
    .B(N2MID[6]),
    .A_N(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _431_ (.B1(_195_),
    .VDD(VPWR),
    .Y(ENA_TT_PROJECT),
    .VSS(VGND),
    .A1(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit3.Q ),
    .A2(_196_));
 sg13g2_mux4_1 _432_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit17.Q ),
    .A0(UIO_OUT_TT_PROJECT3),
    .A1(_117_),
    .A2(_141_),
    .A3(_039_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit16.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W6BEG11 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _433_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit15.Q ),
    .A0(UIO_OUT_TT_PROJECT2),
    .A1(_111_),
    .A2(_135_),
    .A3(_047_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit14.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W6BEG10 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _434_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit13.Q ),
    .A0(UIO_OUT_TT_PROJECT1),
    .A1(_105_),
    .A2(_129_),
    .A3(_055_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit12.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W6BEG9 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _435_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit11.Q ),
    .A0(UIO_OUT_TT_PROJECT0),
    .A1(_099_),
    .A2(_123_),
    .A3(_062_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit10.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W6BEG8 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _436_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit9.Q ),
    .A0(UIO_OUT_TT_PROJECT7),
    .A1(_092_),
    .A2(_117_),
    .A3(_070_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit8.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W6BEG7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _437_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit7.Q ),
    .A0(UIO_OUT_TT_PROJECT6),
    .A1(_083_),
    .A2(_111_),
    .A3(_077_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit6.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W6BEG6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _438_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit5.Q ),
    .A0(UIO_OUT_TT_PROJECT5),
    .A1(_076_),
    .A2(_105_),
    .A3(_084_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit4.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W6BEG5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _439_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit3.Q ),
    .A0(UIO_OUT_TT_PROJECT4),
    .A1(_069_),
    .A2(_099_),
    .A3(_090_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit2.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W6BEG4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _440_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit0.Q ),
    .A0(N4END[3]),
    .A1(S4END[3]),
    .A2(_092_),
    .A3(_061_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit1.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W6BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _441_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit30.Q ),
    .A0(N4END[2]),
    .A1(S4END[2]),
    .A2(_083_),
    .A3(_054_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit31.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W6BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _442_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit28.Q ),
    .A0(N4END[1]),
    .A1(S4END[1]),
    .A2(_076_),
    .A3(_048_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit29.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W6BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _443_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit26.Q ),
    .A0(N4END[0]),
    .A1(S4END[0]),
    .A2(_069_),
    .A3(_041_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit27.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W6BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _444_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit25.Q ),
    .A0(UO_OUT_TT_PROJECT3),
    .A1(_141_),
    .A2(UIO_OUT_TT_PROJECT7),
    .A3(_090_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit24.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.WW4BEG15 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _445_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit23.Q ),
    .A0(UO_OUT_TT_PROJECT2),
    .A1(_135_),
    .A2(UIO_OUT_TT_PROJECT6),
    .A3(_084_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit22.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.WW4BEG14 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _446_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit21.Q ),
    .A0(UO_OUT_TT_PROJECT1),
    .A1(_129_),
    .A2(UIO_OUT_TT_PROJECT5),
    .A3(_077_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit20.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.WW4BEG13 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _447_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit19.Q ),
    .A0(UO_OUT_TT_PROJECT0),
    .A1(_123_),
    .A2(UIO_OUT_TT_PROJECT4),
    .A3(_070_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit18.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.WW4BEG12 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _448_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit17.Q ),
    .A0(UO_OUT_TT_PROJECT7),
    .A1(_117_),
    .A2(UIO_OUT_TT_PROJECT3),
    .A3(_062_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit16.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.WW4BEG11 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _449_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit15.Q ),
    .A0(UO_OUT_TT_PROJECT6),
    .A1(_111_),
    .A2(UIO_OUT_TT_PROJECT2),
    .A3(_055_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit14.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.WW4BEG10 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _450_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit13.Q ),
    .A0(UO_OUT_TT_PROJECT5),
    .A1(_105_),
    .A2(UIO_OUT_TT_PROJECT1),
    .A3(_047_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit12.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.WW4BEG9 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _451_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit11.Q ),
    .A0(UO_OUT_TT_PROJECT4),
    .A1(_099_),
    .A2(UIO_OUT_TT_PROJECT0),
    .A3(_039_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit10.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.WW4BEG8 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _452_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit8.Q ),
    .A0(UO_OUT_TT_PROJECT7),
    .A1(UIO_OE_TT_PROJECT3),
    .A2(_092_),
    .A3(_090_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit9.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.WW4BEG7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _453_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit6.Q ),
    .A0(UO_OUT_TT_PROJECT6),
    .A1(UIO_OE_TT_PROJECT2),
    .A2(_083_),
    .A3(_084_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit7.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.WW4BEG6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _454_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit4.Q ),
    .A0(UO_OUT_TT_PROJECT5),
    .A1(UIO_OE_TT_PROJECT1),
    .A2(_076_),
    .A3(_077_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit5.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.WW4BEG5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _455_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit2.Q ),
    .A0(UO_OUT_TT_PROJECT4),
    .A1(UIO_OE_TT_PROJECT0),
    .A2(_069_),
    .A3(_070_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit3.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.WW4BEG4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _456_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit0.Q ),
    .A0(UO_OUT_TT_PROJECT3),
    .A1(UIO_OE_TT_PROJECT7),
    .A2(_061_),
    .A3(_062_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit1.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.WW4BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _457_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit30.Q ),
    .A0(UO_OUT_TT_PROJECT2),
    .A1(UIO_OE_TT_PROJECT6),
    .A2(_054_),
    .A3(_055_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit31.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.WW4BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _458_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit28.Q ),
    .A0(UO_OUT_TT_PROJECT1),
    .A1(UIO_OE_TT_PROJECT5),
    .A2(_048_),
    .A3(_047_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit29.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.WW4BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _459_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit26.Q ),
    .A0(UO_OUT_TT_PROJECT0),
    .A1(UIO_OE_TT_PROJECT4),
    .A2(_041_),
    .A3(_039_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit27.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.WW4BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _460_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit24.Q ),
    .A0(UIO_OUT_TT_PROJECT7),
    .A1(UIO_OE_TT_PROJECT7),
    .A2(_090_),
    .A3(_039_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit25.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W2BEGb7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _461_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit22.Q ),
    .A0(UIO_OUT_TT_PROJECT6),
    .A1(UIO_OE_TT_PROJECT6),
    .A2(_084_),
    .A3(_047_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit23.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W2BEGb6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _462_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit20.Q ),
    .A0(UIO_OUT_TT_PROJECT5),
    .A1(UIO_OE_TT_PROJECT5),
    .A2(_077_),
    .A3(_055_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit21.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W2BEGb5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _463_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit18.Q ),
    .A0(UIO_OUT_TT_PROJECT4),
    .A1(UIO_OE_TT_PROJECT4),
    .A2(_070_),
    .A3(_062_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit19.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W2BEGb4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _464_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit16.Q ),
    .A0(UIO_OUT_TT_PROJECT3),
    .A1(UIO_OE_TT_PROJECT3),
    .A2(_070_),
    .A3(_062_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit17.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W2BEGb3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _465_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit14.Q ),
    .A0(UIO_OUT_TT_PROJECT2),
    .A1(UIO_OE_TT_PROJECT2),
    .A2(_077_),
    .A3(_055_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit15.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W2BEGb2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _466_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit12.Q ),
    .A0(UIO_OUT_TT_PROJECT1),
    .A1(UIO_OE_TT_PROJECT1),
    .A2(_084_),
    .A3(_047_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit13.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W2BEGb1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _467_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit10.Q ),
    .A0(UIO_OUT_TT_PROJECT0),
    .A1(UIO_OE_TT_PROJECT0),
    .A2(_090_),
    .A3(_039_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit11.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W2BEGb0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _468_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit9.Q ),
    .A0(UO_OUT_TT_PROJECT7),
    .A1(_090_),
    .A2(UIO_OUT_TT_PROJECT7),
    .A3(_039_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit8.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W2BEG7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _469_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit7.Q ),
    .A0(UO_OUT_TT_PROJECT6),
    .A1(_084_),
    .A2(UIO_OUT_TT_PROJECT6),
    .A3(_047_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit6.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W2BEG6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _470_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit5.Q ),
    .A0(UO_OUT_TT_PROJECT5),
    .A1(_077_),
    .A2(UIO_OUT_TT_PROJECT5),
    .A3(_055_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit4.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W2BEG5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _471_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit3.Q ),
    .A0(UO_OUT_TT_PROJECT4),
    .A1(_070_),
    .A2(UIO_OUT_TT_PROJECT4),
    .A3(_062_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit2.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W2BEG4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _472_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit1.Q ),
    .A0(UO_OUT_TT_PROJECT3),
    .A1(_070_),
    .A2(UIO_OUT_TT_PROJECT3),
    .A3(_062_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit0.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W2BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _473_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit31.Q ),
    .A0(UO_OUT_TT_PROJECT2),
    .A1(_077_),
    .A2(UIO_OUT_TT_PROJECT2),
    .A3(_055_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit30.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W2BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _474_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit29.Q ),
    .A0(UO_OUT_TT_PROJECT1),
    .A1(_084_),
    .A2(UIO_OUT_TT_PROJECT1),
    .A3(_047_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit28.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W2BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _475_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit27.Q ),
    .A0(UO_OUT_TT_PROJECT0),
    .A1(_090_),
    .A2(UIO_OUT_TT_PROJECT0),
    .A3(_039_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit26.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W2BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _476_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit24.Q ),
    .A0(N1END[3]),
    .A1(S1END[3]),
    .A2(UO_OUT_TT_PROJECT1),
    .A3(UO_OUT_TT_PROJECT4),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit25.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W1BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _477_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit22.Q ),
    .A0(N1END[2]),
    .A1(S1END[2]),
    .A2(UO_OUT_TT_PROJECT0),
    .A3(UO_OUT_TT_PROJECT5),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit23.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W1BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _478_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit20.Q ),
    .A0(N1END[1]),
    .A1(S1END[1]),
    .A2(UO_OUT_TT_PROJECT3),
    .A3(UO_OUT_TT_PROJECT6),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit21.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W1BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _479_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit18.Q ),
    .A0(N1END[0]),
    .A1(S1END[0]),
    .A2(UO_OUT_TT_PROJECT2),
    .A3(UO_OUT_TT_PROJECT7),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit19.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.W1BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _480_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit5.Q ),
    .A0(E1END[3]),
    .A1(E2END[0]),
    .A2(E2MID[0]),
    .A3(_039_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit4.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.S2BEG7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _481_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit2.Q ),
    .A0(E1END[2]),
    .A1(E2MID[1]),
    .A2(E2END[1]),
    .A3(_047_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit3.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.S2BEG6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _482_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit0.Q ),
    .A0(E1END[1]),
    .A1(E2MID[2]),
    .A2(E2END[2]),
    .A3(_055_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit1.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.S2BEG5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _483_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit31.Q ),
    .A0(E1END[0]),
    .A1(E2END[3]),
    .A2(E2MID[3]),
    .A3(_062_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit30.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.S2BEG4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _484_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit29.Q ),
    .A0(E2MID[4]),
    .A1(E6END[11]),
    .A2(E2END[4]),
    .A3(_070_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit28.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.S2BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _485_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit27.Q ),
    .A0(E2MID[5]),
    .A1(E6END[10]),
    .A2(E2END[5]),
    .A3(_077_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit26.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.S2BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _486_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit24.Q ),
    .A0(E2MID[6]),
    .A1(E2END[6]),
    .A2(E6END[9]),
    .A3(_084_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit25.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.S2BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _487_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit22.Q ),
    .A0(E2MID[7]),
    .A1(E2END[7]),
    .A2(E6END[8]),
    .A3(_090_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit23.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.S2BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _488_ (.A(N1END[3]),
    .B(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit30.Q ),
    .C(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit31.Q ),
    .Y(_197_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _489_ (.Y(_198_),
    .B(E6END[3]),
    .A_N(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _490_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit30.Q ),
    .C1(_197_),
    .B1(_198_),
    .A1(_002_),
    .Y(_199_),
    .A2(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit31.Q ));
 sg13g2_mux4_1 _491_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit20.Q ),
    .A0(E1END[3]),
    .A1(E6END[11]),
    .A2(_041_),
    .A3(_199_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit21.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.S1BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _492_ (.A(N1END[2]),
    .B(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit28.Q ),
    .C(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit29.Q ),
    .Y(_200_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _493_ (.Y(_201_),
    .B(E6END[2]),
    .A_N(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _494_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit28.Q ),
    .C1(_200_),
    .B1(_201_),
    .A1(_003_),
    .Y(_202_),
    .A2(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit29.Q ));
 sg13g2_mux4_1 _495_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit18.Q ),
    .A0(E1END[2]),
    .A1(E6END[10]),
    .A2(_048_),
    .A3(_202_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit19.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.S1BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _496_ (.A(N1END[1]),
    .B(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit26.Q ),
    .C(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit27.Q ),
    .Y(_203_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _497_ (.Y(_204_),
    .B(E6END[1]),
    .A_N(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _498_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit26.Q ),
    .C1(_203_),
    .B1(_204_),
    .A1(_004_),
    .Y(_205_),
    .A2(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit27.Q ));
 sg13g2_mux4_1 _499_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit16.Q ),
    .A0(E1END[1]),
    .A1(E6END[9]),
    .A2(_054_),
    .A3(_205_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit17.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.S1BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _500_ (.A(N1END[0]),
    .B(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit24.Q ),
    .C(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit25.Q ),
    .Y(_206_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _501_ (.Y(_207_),
    .B(E6END[0]),
    .A_N(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _502_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit24.Q ),
    .C1(_206_),
    .B1(_207_),
    .A1(_005_),
    .Y(_208_),
    .A2(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit25.Q ));
 sg13g2_mux4_1 _503_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit14.Q ),
    .A0(E1END[0]),
    .A1(E6END[8]),
    .A2(_061_),
    .A3(_208_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit15.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.S1BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _504_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit0.Q ),
    .A0(E2MID[0]),
    .A1(E2END[0]),
    .A2(E6END[0]),
    .A3(_039_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit1.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.N2BEG7 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _505_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit31.Q ),
    .A0(E2MID[1]),
    .A1(E6END[1]),
    .A2(E2END[1]),
    .A3(_047_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit30.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.N2BEG6 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _506_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit29.Q ),
    .A0(E2MID[2]),
    .A1(E6END[2]),
    .A2(E2END[2]),
    .A3(_055_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit28.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.N2BEG5 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _507_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit26.Q ),
    .A0(E2MID[3]),
    .A1(E2END[3]),
    .A2(E6END[3]),
    .A3(_062_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit27.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.N2BEG4 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _508_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit25.Q ),
    .A0(E2MID[4]),
    .A1(E6END[4]),
    .A2(E2END[4]),
    .A3(_070_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit24.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.N2BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _509_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit23.Q ),
    .A0(E2MID[5]),
    .A1(E6END[5]),
    .A2(E2END[5]),
    .A3(_077_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit22.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.N2BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _510_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit20.Q ),
    .A0(E2MID[6]),
    .A1(E2END[6]),
    .A2(E6END[6]),
    .A3(_084_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit21.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.N2BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _511_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit18.Q ),
    .A0(E2MID[7]),
    .A1(E2END[7]),
    .A2(E6END[7]),
    .A3(_090_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit19.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.N2BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _512_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit16.Q ),
    .A0(E1END[3]),
    .A1(E6END[7]),
    .A2(_041_),
    .A3(_199_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit17.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.N1BEG3 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _513_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit14.Q ),
    .A0(E1END[2]),
    .A1(E6END[6]),
    .A2(_048_),
    .A3(_202_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit15.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.N1BEG2 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _514_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit12.Q ),
    .A0(E1END[1]),
    .A1(E6END[5]),
    .A2(_054_),
    .A3(_205_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit13.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.N1BEG1 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux4_1 _515_ (.S0(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit10.Q ),
    .A0(E1END[0]),
    .A1(E6END[4]),
    .A2(_061_),
    .A3(_208_),
    .S1(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit11.Q ),
    .X(\Inst_E_TT_IF_switch_matrix.N1BEG0 ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _516_ (.D(FrameData[10]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _517_ (.D(FrameData[11]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _518_ (.D(FrameData[12]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _519_ (.D(FrameData[13]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _520_ (.D(FrameData[14]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _521_ (.D(FrameData[15]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _522_ (.D(FrameData[16]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _523_ (.D(FrameData[17]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _524_ (.D(FrameData[18]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _525_ (.D(FrameData[19]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _526_ (.D(FrameData[20]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _527_ (.D(FrameData[21]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _528_ (.D(FrameData[22]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _529_ (.D(FrameData[23]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _530_ (.D(FrameData[24]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _531_ (.D(FrameData[25]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _532_ (.D(FrameData[26]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _533_ (.D(FrameData[27]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _534_ (.D(FrameData[28]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _535_ (.D(FrameData[29]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _536_ (.D(FrameData[30]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _537_ (.D(FrameData[31]),
    .GATE(FrameStrobe[8]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame8_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _538_ (.D(FrameData[0]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _539_ (.D(FrameData[1]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _540_ (.D(FrameData[2]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _541_ (.D(FrameData[3]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _542_ (.D(FrameData[4]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _543_ (.D(FrameData[5]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _544_ (.D(FrameData[6]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _545_ (.D(FrameData[7]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _546_ (.D(FrameData[8]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _547_ (.D(FrameData[9]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _548_ (.D(FrameData[10]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _549_ (.D(FrameData[11]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _550_ (.D(FrameData[12]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _551_ (.D(FrameData[13]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _552_ (.D(FrameData[14]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _553_ (.D(FrameData[15]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _554_ (.D(FrameData[16]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _555_ (.D(FrameData[17]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _556_ (.D(FrameData[18]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _557_ (.D(FrameData[19]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _558_ (.D(FrameData[20]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _559_ (.D(FrameData[21]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _560_ (.D(FrameData[22]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _561_ (.D(FrameData[23]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _562_ (.D(FrameData[24]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _563_ (.D(FrameData[25]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _564_ (.D(FrameData[26]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _565_ (.D(FrameData[27]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _566_ (.D(FrameData[28]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _567_ (.D(FrameData[29]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _568_ (.D(FrameData[30]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _569_ (.D(FrameData[31]),
    .GATE(FrameStrobe[7]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame7_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _570_ (.D(FrameData[0]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _571_ (.D(FrameData[1]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _572_ (.D(FrameData[2]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _573_ (.D(FrameData[3]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _574_ (.D(FrameData[4]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _575_ (.D(FrameData[5]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _576_ (.D(FrameData[6]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _577_ (.D(FrameData[7]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _578_ (.D(FrameData[8]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _579_ (.D(FrameData[9]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _580_ (.D(FrameData[10]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _581_ (.D(FrameData[11]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _582_ (.D(FrameData[12]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _583_ (.D(FrameData[13]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _584_ (.D(FrameData[14]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _585_ (.D(FrameData[15]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _586_ (.D(FrameData[16]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _587_ (.D(FrameData[17]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _588_ (.D(FrameData[18]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _589_ (.D(FrameData[19]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _590_ (.D(FrameData[20]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _591_ (.D(FrameData[21]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _592_ (.D(FrameData[22]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _593_ (.D(FrameData[23]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _594_ (.D(FrameData[24]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _595_ (.D(FrameData[25]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _596_ (.D(FrameData[26]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _597_ (.D(FrameData[27]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _598_ (.D(FrameData[28]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _599_ (.D(FrameData[29]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _600_ (.D(FrameData[30]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _601_ (.D(FrameData[31]),
    .GATE(FrameStrobe[6]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame6_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _602_ (.D(FrameData[0]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _603_ (.D(FrameData[1]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _604_ (.D(FrameData[2]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _605_ (.D(FrameData[3]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _606_ (.D(FrameData[4]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _607_ (.D(FrameData[5]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _608_ (.D(FrameData[6]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _609_ (.D(FrameData[7]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _610_ (.D(FrameData[8]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _611_ (.D(FrameData[9]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _612_ (.D(FrameData[10]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _613_ (.D(FrameData[11]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _614_ (.D(FrameData[12]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _615_ (.D(FrameData[13]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _616_ (.D(FrameData[14]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _617_ (.D(FrameData[15]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _618_ (.D(FrameData[16]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _619_ (.D(FrameData[17]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _620_ (.D(FrameData[18]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _621_ (.D(FrameData[19]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _622_ (.D(FrameData[20]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _623_ (.D(FrameData[21]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _624_ (.D(FrameData[22]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _625_ (.D(FrameData[23]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _626_ (.D(FrameData[24]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _627_ (.D(FrameData[25]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _628_ (.D(FrameData[26]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _629_ (.D(FrameData[27]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _630_ (.D(FrameData[28]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _631_ (.D(FrameData[29]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _632_ (.D(FrameData[30]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _633_ (.D(FrameData[31]),
    .GATE(FrameStrobe[5]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame5_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _634_ (.D(FrameData[0]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _635_ (.D(FrameData[1]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _636_ (.D(FrameData[2]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _637_ (.D(FrameData[3]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _638_ (.D(FrameData[4]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _639_ (.D(FrameData[5]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _640_ (.D(FrameData[6]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _641_ (.D(FrameData[7]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _642_ (.D(FrameData[8]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _643_ (.D(FrameData[9]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _644_ (.D(FrameData[10]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _645_ (.D(FrameData[11]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _646_ (.D(FrameData[12]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _647_ (.D(FrameData[13]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _648_ (.D(FrameData[14]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _649_ (.D(FrameData[15]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _650_ (.D(FrameData[16]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _651_ (.D(FrameData[17]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _652_ (.D(FrameData[18]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _653_ (.D(FrameData[19]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _654_ (.D(FrameData[20]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _655_ (.D(FrameData[21]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _656_ (.D(FrameData[22]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _657_ (.D(FrameData[23]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _658_ (.D(FrameData[24]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _659_ (.D(FrameData[25]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _660_ (.D(FrameData[26]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _661_ (.D(FrameData[27]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _662_ (.D(FrameData[28]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _663_ (.D(FrameData[29]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _664_ (.D(FrameData[30]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _665_ (.D(FrameData[31]),
    .GATE(FrameStrobe[4]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame4_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _666_ (.D(FrameData[0]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _667_ (.D(FrameData[1]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _668_ (.D(FrameData[2]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _669_ (.D(FrameData[3]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _670_ (.D(FrameData[4]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _671_ (.D(FrameData[5]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _672_ (.D(FrameData[6]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _673_ (.D(FrameData[7]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _674_ (.D(FrameData[8]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _675_ (.D(FrameData[9]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _676_ (.D(FrameData[10]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _677_ (.D(FrameData[11]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _678_ (.D(FrameData[12]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _679_ (.D(FrameData[13]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _680_ (.D(FrameData[14]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _681_ (.D(FrameData[15]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _682_ (.D(FrameData[16]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _683_ (.D(FrameData[17]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _684_ (.D(FrameData[18]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _685_ (.D(FrameData[19]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _686_ (.D(FrameData[20]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _687_ (.D(FrameData[21]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _688_ (.D(FrameData[22]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _689_ (.D(FrameData[23]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _690_ (.D(FrameData[24]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _691_ (.D(FrameData[25]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _692_ (.D(FrameData[26]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _693_ (.D(FrameData[27]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _694_ (.D(FrameData[28]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _695_ (.D(FrameData[29]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _696_ (.D(FrameData[30]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _697_ (.D(FrameData[31]),
    .GATE(FrameStrobe[3]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame3_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _698_ (.D(FrameData[0]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _699_ (.D(FrameData[1]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _700_ (.D(FrameData[2]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _701_ (.D(FrameData[3]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _702_ (.D(FrameData[4]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _703_ (.D(FrameData[5]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _704_ (.D(FrameData[6]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _705_ (.D(FrameData[7]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _706_ (.D(FrameData[8]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _707_ (.D(FrameData[9]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _708_ (.D(FrameData[10]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _709_ (.D(FrameData[11]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _710_ (.D(FrameData[12]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _711_ (.D(FrameData[13]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _712_ (.D(FrameData[14]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _713_ (.D(FrameData[15]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _714_ (.D(FrameData[16]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _715_ (.D(FrameData[17]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _716_ (.D(FrameData[18]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _717_ (.D(FrameData[19]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _718_ (.D(FrameData[20]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _719_ (.D(FrameData[21]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _720_ (.D(FrameData[22]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _721_ (.D(FrameData[23]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _722_ (.D(FrameData[24]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _723_ (.D(FrameData[25]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _724_ (.D(FrameData[26]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _725_ (.D(FrameData[27]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _726_ (.D(FrameData[28]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _727_ (.D(FrameData[29]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _728_ (.D(FrameData[30]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _729_ (.D(FrameData[31]),
    .GATE(FrameStrobe[2]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame2_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _730_ (.D(FrameData[0]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _731_ (.D(FrameData[1]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _732_ (.D(FrameData[2]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _733_ (.D(FrameData[3]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _734_ (.D(FrameData[4]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _735_ (.D(FrameData[5]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _736_ (.D(FrameData[6]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _737_ (.D(FrameData[7]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _738_ (.D(FrameData[8]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _739_ (.D(FrameData[9]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _740_ (.D(FrameData[10]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _741_ (.D(FrameData[11]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _742_ (.D(FrameData[12]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _743_ (.D(FrameData[13]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _744_ (.D(FrameData[14]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _745_ (.D(FrameData[15]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _746_ (.D(FrameData[16]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _747_ (.D(FrameData[17]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _748_ (.D(FrameData[18]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _749_ (.D(FrameData[19]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _750_ (.D(FrameData[20]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _751_ (.D(FrameData[21]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _752_ (.D(FrameData[22]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _753_ (.D(FrameData[23]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _754_ (.D(FrameData[24]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _755_ (.D(FrameData[25]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _756_ (.D(FrameData[26]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _757_ (.D(FrameData[27]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _758_ (.D(FrameData[28]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _759_ (.D(FrameData[29]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _760_ (.D(FrameData[30]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _761_ (.D(FrameData[31]),
    .GATE(FrameStrobe[1]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame1_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _762_ (.D(FrameData[0]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit0.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _763_ (.D(FrameData[1]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit1.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _764_ (.D(FrameData[2]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit2.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _765_ (.D(FrameData[3]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit3.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _766_ (.D(FrameData[4]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit4.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _767_ (.D(FrameData[5]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit5.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _768_ (.D(FrameData[6]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit6.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _769_ (.D(FrameData[7]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit7.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _770_ (.D(FrameData[8]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit8.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _771_ (.D(FrameData[9]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit9.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _772_ (.D(FrameData[10]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit10.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _773_ (.D(FrameData[11]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit11.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _774_ (.D(FrameData[12]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit12.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _775_ (.D(FrameData[13]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit13.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _776_ (.D(FrameData[14]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit14.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _777_ (.D(FrameData[15]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit15.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _778_ (.D(FrameData[16]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit16.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _779_ (.D(FrameData[17]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit17.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _780_ (.D(FrameData[18]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit18.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _781_ (.D(FrameData[19]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit19.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _782_ (.D(FrameData[20]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit20.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _783_ (.D(FrameData[21]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit21.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _784_ (.D(FrameData[22]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit22.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _785_ (.D(FrameData[23]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit23.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _786_ (.D(FrameData[24]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit24.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _787_ (.D(FrameData[25]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit25.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _788_ (.D(FrameData[26]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit26.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _789_ (.D(FrameData[27]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit27.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _790_ (.D(FrameData[28]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit28.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _791_ (.D(FrameData[29]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit29.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _792_ (.D(FrameData[30]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit30.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlhq_1 _793_ (.D(FrameData[31]),
    .GATE(FrameStrobe[0]),
    .Q(\Inst_E_TT_IF_ConfigMem.Inst_frame0_bit31.Q ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _794_ (.A(clknet_1_0__leaf_UserCLK),
    .X(CLK_TT_PROJECT),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _795_ (.A(FrameData[0]),
    .X(FrameData_O[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _796_ (.A(FrameData[1]),
    .X(FrameData_O[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _797_ (.A(FrameData[2]),
    .X(FrameData_O[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _798_ (.A(FrameData[3]),
    .X(FrameData_O[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _799_ (.A(FrameData[4]),
    .X(FrameData_O[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _800_ (.A(FrameData[5]),
    .X(FrameData_O[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _801_ (.A(FrameData[6]),
    .X(FrameData_O[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _802_ (.A(FrameData[7]),
    .X(FrameData_O[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _803_ (.A(FrameData[8]),
    .X(FrameData_O[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _804_ (.A(FrameData[9]),
    .X(FrameData_O[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _805_ (.A(FrameData[10]),
    .X(FrameData_O[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _806_ (.A(FrameData[11]),
    .X(FrameData_O[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _807_ (.A(FrameData[12]),
    .X(FrameData_O[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _808_ (.A(FrameData[13]),
    .X(FrameData_O[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _809_ (.A(FrameData[14]),
    .X(FrameData_O[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _810_ (.A(FrameData[15]),
    .X(FrameData_O[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _811_ (.A(FrameData[16]),
    .X(FrameData_O[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _812_ (.A(FrameData[17]),
    .X(FrameData_O[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _813_ (.A(FrameData[18]),
    .X(FrameData_O[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _814_ (.A(FrameData[19]),
    .X(FrameData_O[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _815_ (.A(FrameData[20]),
    .X(FrameData_O[20]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _816_ (.A(FrameData[21]),
    .X(FrameData_O[21]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _817_ (.A(FrameData[22]),
    .X(FrameData_O[22]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _818_ (.A(FrameData[23]),
    .X(FrameData_O[23]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _819_ (.A(FrameData[24]),
    .X(FrameData_O[24]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _820_ (.A(FrameData[25]),
    .X(FrameData_O[25]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _821_ (.A(FrameData[26]),
    .X(FrameData_O[26]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _822_ (.A(FrameData[27]),
    .X(FrameData_O[27]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _823_ (.A(FrameData[28]),
    .X(FrameData_O[28]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _824_ (.A(FrameData[29]),
    .X(FrameData_O[29]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _825_ (.A(FrameData[30]),
    .X(FrameData_O[30]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _826_ (.A(FrameData[31]),
    .X(FrameData_O[31]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _827_ (.A(FrameStrobe[0]),
    .X(FrameStrobe_O[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _828_ (.A(FrameStrobe[1]),
    .X(FrameStrobe_O[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _829_ (.A(FrameStrobe[2]),
    .X(FrameStrobe_O[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _830_ (.A(FrameStrobe[3]),
    .X(FrameStrobe_O[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _831_ (.A(FrameStrobe[4]),
    .X(FrameStrobe_O[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _832_ (.A(FrameStrobe[5]),
    .X(FrameStrobe_O[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _833_ (.A(FrameStrobe[6]),
    .X(FrameStrobe_O[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _834_ (.A(FrameStrobe[7]),
    .X(FrameStrobe_O[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _835_ (.A(FrameStrobe[8]),
    .X(FrameStrobe_O[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _836_ (.A(FrameStrobe[9]),
    .X(FrameStrobe_O[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _837_ (.A(FrameStrobe[10]),
    .X(FrameStrobe_O[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _838_ (.A(FrameStrobe[11]),
    .X(FrameStrobe_O[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _839_ (.A(FrameStrobe[12]),
    .X(FrameStrobe_O[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _840_ (.A(FrameStrobe[13]),
    .X(FrameStrobe_O[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _841_ (.A(FrameStrobe[14]),
    .X(FrameStrobe_O[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _842_ (.A(FrameStrobe[15]),
    .X(FrameStrobe_O[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _843_ (.A(FrameStrobe[16]),
    .X(FrameStrobe_O[16]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _844_ (.A(FrameStrobe[17]),
    .X(FrameStrobe_O[17]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _845_ (.A(FrameStrobe[18]),
    .X(FrameStrobe_O[18]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _846_ (.A(FrameStrobe[19]),
    .X(FrameStrobe_O[19]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _847_ (.A(\Inst_E_TT_IF_switch_matrix.N1BEG0 ),
    .X(N1BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _848_ (.A(\Inst_E_TT_IF_switch_matrix.N1BEG1 ),
    .X(N1BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _849_ (.A(\Inst_E_TT_IF_switch_matrix.N1BEG2 ),
    .X(N1BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _850_ (.A(\Inst_E_TT_IF_switch_matrix.N1BEG3 ),
    .X(N1BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _851_ (.A(\Inst_E_TT_IF_switch_matrix.N2BEG0 ),
    .X(N2BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _852_ (.A(\Inst_E_TT_IF_switch_matrix.N2BEG1 ),
    .X(N2BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _853_ (.A(\Inst_E_TT_IF_switch_matrix.N2BEG2 ),
    .X(N2BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _854_ (.A(\Inst_E_TT_IF_switch_matrix.N2BEG3 ),
    .X(N2BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _855_ (.A(\Inst_E_TT_IF_switch_matrix.N2BEG4 ),
    .X(N2BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _856_ (.A(\Inst_E_TT_IF_switch_matrix.N2BEG5 ),
    .X(N2BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _857_ (.A(\Inst_E_TT_IF_switch_matrix.N2BEG6 ),
    .X(N2BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _858_ (.A(\Inst_E_TT_IF_switch_matrix.N2BEG7 ),
    .X(N2BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _859_ (.A(N2MID[0]),
    .X(N2BEGb[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _860_ (.A(N2MID[1]),
    .X(N2BEGb[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _861_ (.A(N2MID[2]),
    .X(N2BEGb[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _862_ (.A(N2MID[3]),
    .X(N2BEGb[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _863_ (.A(N2MID[4]),
    .X(N2BEGb[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _864_ (.A(N2MID[5]),
    .X(N2BEGb[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _865_ (.A(N2MID[6]),
    .X(N2BEGb[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _866_ (.A(N2MID[7]),
    .X(N2BEGb[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _867_ (.A(N4END[4]),
    .X(N4BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _868_ (.A(N4END[5]),
    .X(N4BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _869_ (.A(N4END[6]),
    .X(N4BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _870_ (.A(N4END[7]),
    .X(N4BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _871_ (.A(N4END[8]),
    .X(N4BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _872_ (.A(N4END[9]),
    .X(N4BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _873_ (.A(N4END[10]),
    .X(N4BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _874_ (.A(N4END[11]),
    .X(N4BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _875_ (.A(N4END[12]),
    .X(N4BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _876_ (.A(N4END[13]),
    .X(N4BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _877_ (.A(N4END[14]),
    .X(N4BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _878_ (.A(N4END[15]),
    .X(N4BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _879_ (.A(\Inst_E_TT_IF_switch_matrix.N4BEG0 ),
    .X(N4BEG[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _880_ (.A(\Inst_E_TT_IF_switch_matrix.N4BEG1 ),
    .X(N4BEG[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _881_ (.A(\Inst_E_TT_IF_switch_matrix.N4BEG2 ),
    .X(N4BEG[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _882_ (.A(\Inst_E_TT_IF_switch_matrix.N4BEG3 ),
    .X(N4BEG[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _883_ (.A(\Inst_E_TT_IF_switch_matrix.S1BEG0 ),
    .X(S1BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _884_ (.A(\Inst_E_TT_IF_switch_matrix.S1BEG1 ),
    .X(S1BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _885_ (.A(\Inst_E_TT_IF_switch_matrix.S1BEG2 ),
    .X(S1BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _886_ (.A(\Inst_E_TT_IF_switch_matrix.S1BEG3 ),
    .X(S1BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _887_ (.A(\Inst_E_TT_IF_switch_matrix.S2BEG0 ),
    .X(S2BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _888_ (.A(\Inst_E_TT_IF_switch_matrix.S2BEG1 ),
    .X(S2BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _889_ (.A(\Inst_E_TT_IF_switch_matrix.S2BEG2 ),
    .X(S2BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _890_ (.A(\Inst_E_TT_IF_switch_matrix.S2BEG3 ),
    .X(S2BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _891_ (.A(\Inst_E_TT_IF_switch_matrix.S2BEG4 ),
    .X(S2BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _892_ (.A(\Inst_E_TT_IF_switch_matrix.S2BEG5 ),
    .X(S2BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _893_ (.A(\Inst_E_TT_IF_switch_matrix.S2BEG6 ),
    .X(S2BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _894_ (.A(\Inst_E_TT_IF_switch_matrix.S2BEG7 ),
    .X(S2BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _895_ (.A(S2MID[0]),
    .X(S2BEGb[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _896_ (.A(S2MID[1]),
    .X(S2BEGb[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _897_ (.A(S2MID[2]),
    .X(S2BEGb[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _898_ (.A(S2MID[3]),
    .X(S2BEGb[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _899_ (.A(S2MID[4]),
    .X(S2BEGb[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _900_ (.A(S2MID[5]),
    .X(S2BEGb[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _901_ (.A(S2MID[6]),
    .X(S2BEGb[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _902_ (.A(S2MID[7]),
    .X(S2BEGb[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _903_ (.A(S4END[4]),
    .X(S4BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _904_ (.A(S4END[5]),
    .X(S4BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _905_ (.A(S4END[6]),
    .X(S4BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _906_ (.A(S4END[7]),
    .X(S4BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _907_ (.A(S4END[8]),
    .X(S4BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _908_ (.A(S4END[9]),
    .X(S4BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _909_ (.A(S4END[10]),
    .X(S4BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _910_ (.A(S4END[11]),
    .X(S4BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _911_ (.A(S4END[12]),
    .X(S4BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _912_ (.A(S4END[13]),
    .X(S4BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _913_ (.A(S4END[14]),
    .X(S4BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _914_ (.A(S4END[15]),
    .X(S4BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _915_ (.A(\Inst_E_TT_IF_switch_matrix.S4BEG0 ),
    .X(S4BEG[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _916_ (.A(\Inst_E_TT_IF_switch_matrix.S4BEG1 ),
    .X(S4BEG[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _917_ (.A(\Inst_E_TT_IF_switch_matrix.S4BEG2 ),
    .X(S4BEG[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _918_ (.A(\Inst_E_TT_IF_switch_matrix.S4BEG3 ),
    .X(S4BEG[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _919_ (.A(clknet_1_1__leaf_UserCLK),
    .X(UserCLKo),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _920_ (.A(\Inst_E_TT_IF_switch_matrix.W1BEG0 ),
    .X(W1BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _921_ (.A(\Inst_E_TT_IF_switch_matrix.W1BEG1 ),
    .X(W1BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _922_ (.A(\Inst_E_TT_IF_switch_matrix.W1BEG2 ),
    .X(W1BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _923_ (.A(\Inst_E_TT_IF_switch_matrix.W1BEG3 ),
    .X(W1BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _924_ (.A(\Inst_E_TT_IF_switch_matrix.W2BEG0 ),
    .X(W2BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _925_ (.A(\Inst_E_TT_IF_switch_matrix.W2BEG1 ),
    .X(W2BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _926_ (.A(\Inst_E_TT_IF_switch_matrix.W2BEG2 ),
    .X(W2BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _927_ (.A(\Inst_E_TT_IF_switch_matrix.W2BEG3 ),
    .X(W2BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _928_ (.A(\Inst_E_TT_IF_switch_matrix.W2BEG4 ),
    .X(W2BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _929_ (.A(\Inst_E_TT_IF_switch_matrix.W2BEG5 ),
    .X(W2BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _930_ (.A(\Inst_E_TT_IF_switch_matrix.W2BEG6 ),
    .X(W2BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _931_ (.A(\Inst_E_TT_IF_switch_matrix.W2BEG7 ),
    .X(W2BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _932_ (.A(\Inst_E_TT_IF_switch_matrix.W2BEGb0 ),
    .X(W2BEGb[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _933_ (.A(\Inst_E_TT_IF_switch_matrix.W2BEGb1 ),
    .X(W2BEGb[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _934_ (.A(\Inst_E_TT_IF_switch_matrix.W2BEGb2 ),
    .X(W2BEGb[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _935_ (.A(\Inst_E_TT_IF_switch_matrix.W2BEGb3 ),
    .X(W2BEGb[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _936_ (.A(\Inst_E_TT_IF_switch_matrix.W2BEGb4 ),
    .X(W2BEGb[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _937_ (.A(\Inst_E_TT_IF_switch_matrix.W2BEGb5 ),
    .X(W2BEGb[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _938_ (.A(\Inst_E_TT_IF_switch_matrix.W2BEGb6 ),
    .X(W2BEGb[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _939_ (.A(\Inst_E_TT_IF_switch_matrix.W2BEGb7 ),
    .X(W2BEGb[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _940_ (.A(\Inst_E_TT_IF_switch_matrix.W6BEG0 ),
    .X(W6BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _941_ (.A(\Inst_E_TT_IF_switch_matrix.W6BEG1 ),
    .X(W6BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _942_ (.A(\Inst_E_TT_IF_switch_matrix.W6BEG2 ),
    .X(W6BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _943_ (.A(\Inst_E_TT_IF_switch_matrix.W6BEG3 ),
    .X(W6BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _944_ (.A(\Inst_E_TT_IF_switch_matrix.W6BEG4 ),
    .X(W6BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _945_ (.A(\Inst_E_TT_IF_switch_matrix.W6BEG5 ),
    .X(W6BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _946_ (.A(\Inst_E_TT_IF_switch_matrix.W6BEG6 ),
    .X(W6BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _947_ (.A(\Inst_E_TT_IF_switch_matrix.W6BEG7 ),
    .X(W6BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _948_ (.A(\Inst_E_TT_IF_switch_matrix.W6BEG8 ),
    .X(W6BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _949_ (.A(\Inst_E_TT_IF_switch_matrix.W6BEG9 ),
    .X(W6BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _950_ (.A(\Inst_E_TT_IF_switch_matrix.W6BEG10 ),
    .X(W6BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _951_ (.A(\Inst_E_TT_IF_switch_matrix.W6BEG11 ),
    .X(W6BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _952_ (.A(\Inst_E_TT_IF_switch_matrix.WW4BEG0 ),
    .X(WW4BEG[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _953_ (.A(\Inst_E_TT_IF_switch_matrix.WW4BEG1 ),
    .X(WW4BEG[1]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _954_ (.A(\Inst_E_TT_IF_switch_matrix.WW4BEG2 ),
    .X(WW4BEG[2]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _955_ (.A(\Inst_E_TT_IF_switch_matrix.WW4BEG3 ),
    .X(WW4BEG[3]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _956_ (.A(\Inst_E_TT_IF_switch_matrix.WW4BEG4 ),
    .X(WW4BEG[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _957_ (.A(\Inst_E_TT_IF_switch_matrix.WW4BEG5 ),
    .X(WW4BEG[5]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _958_ (.A(\Inst_E_TT_IF_switch_matrix.WW4BEG6 ),
    .X(WW4BEG[6]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _959_ (.A(\Inst_E_TT_IF_switch_matrix.WW4BEG7 ),
    .X(WW4BEG[7]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _960_ (.A(\Inst_E_TT_IF_switch_matrix.WW4BEG8 ),
    .X(WW4BEG[8]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _961_ (.A(\Inst_E_TT_IF_switch_matrix.WW4BEG9 ),
    .X(WW4BEG[9]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _962_ (.A(\Inst_E_TT_IF_switch_matrix.WW4BEG10 ),
    .X(WW4BEG[10]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _963_ (.A(\Inst_E_TT_IF_switch_matrix.WW4BEG11 ),
    .X(WW4BEG[11]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _964_ (.A(\Inst_E_TT_IF_switch_matrix.WW4BEG12 ),
    .X(WW4BEG[12]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _965_ (.A(\Inst_E_TT_IF_switch_matrix.WW4BEG13 ),
    .X(WW4BEG[13]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _966_ (.A(\Inst_E_TT_IF_switch_matrix.WW4BEG14 ),
    .X(WW4BEG[14]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 _967_ (.A(\Inst_E_TT_IF_switch_matrix.WW4BEG15 ),
    .X(WW4BEG[15]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_0_UserCLK (.A(UserCLK),
    .X(clknet_0_UserCLK),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_1_0__f_UserCLK (.A(clknet_0_UserCLK),
    .X(clknet_1_0__leaf_UserCLK),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_1_1__f_UserCLK (.A(clknet_0_UserCLK),
    .X(clknet_1_1__leaf_UserCLK),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_antennanp ANTENNA_1 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameStrobe[10]));
 sg13g2_antennanp ANTENNA_2 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameStrobe[11]));
 sg13g2_antennanp ANTENNA_3 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameStrobe[12]));
 sg13g2_antennanp ANTENNA_4 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameStrobe[14]));
 sg13g2_antennanp ANTENNA_5 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameStrobe[19]));
 sg13g2_antennanp ANTENNA_6 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameStrobe[9]));
 sg13g2_antennanp ANTENNA_7 (.VDD(VPWR),
    .VSS(VGND),
    .A(N2END[7]));
 sg13g2_antennanp ANTENNA_8 (.VDD(VPWR),
    .VSS(VGND),
    .A(N2MID[1]));
 sg13g2_antennanp ANTENNA_9 (.VDD(VPWR),
    .VSS(VGND),
    .A(N2MID[1]));
 sg13g2_antennanp ANTENNA_10 (.VDD(VPWR),
    .VSS(VGND),
    .A(N2MID[1]));
 sg13g2_antennanp ANTENNA_11 (.VDD(VPWR),
    .VSS(VGND),
    .A(N2MID[2]));
 sg13g2_antennanp ANTENNA_12 (.VDD(VPWR),
    .VSS(VGND),
    .A(N2MID[2]));
 sg13g2_antennanp ANTENNA_13 (.VDD(VPWR),
    .VSS(VGND),
    .A(N2MID[2]));
 sg13g2_antennanp ANTENNA_14 (.VDD(VPWR),
    .VSS(VGND),
    .A(N4END[4]));
 sg13g2_antennanp ANTENNA_15 (.VDD(VPWR),
    .VSS(VGND),
    .A(N4END[6]));
 sg13g2_antennanp ANTENNA_16 (.VDD(VPWR),
    .VSS(VGND),
    .A(N4END[7]));
 sg13g2_antennanp ANTENNA_17 (.VDD(VPWR),
    .VSS(VGND),
    .A(N4END[9]));
 sg13g2_antennanp ANTENNA_18 (.VDD(VPWR),
    .VSS(VGND),
    .A(S4END[9]));
 sg13g2_antennanp ANTENNA_19 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameStrobe[15]));
 sg13g2_antennanp ANTENNA_20 (.VDD(VPWR),
    .VSS(VGND),
    .A(FrameStrobe[17]));
 sg13g2_antennanp ANTENNA_21 (.VDD(VPWR),
    .VSS(VGND),
    .A(N2END[2]));
 sg13g2_antennanp ANTENNA_22 (.VDD(VPWR),
    .VSS(VGND),
    .A(N2END[2]));
 sg13g2_antennanp ANTENNA_23 (.VDD(VPWR),
    .VSS(VGND),
    .A(N2END[2]));
 sg13g2_antennanp ANTENNA_24 (.VDD(VPWR),
    .VSS(VGND),
    .A(N2END[2]));
 sg13g2_antennanp ANTENNA_25 (.VDD(VPWR),
    .VSS(VGND),
    .A(N2MID[5]));
 sg13g2_antennanp ANTENNA_26 (.VDD(VPWR),
    .VSS(VGND),
    .A(N2MID[5]));
 sg13g2_antennanp ANTENNA_27 (.VDD(VPWR),
    .VSS(VGND),
    .A(N2MID[5]));
 sg13g2_antennanp ANTENNA_28 (.VDD(VPWR),
    .VSS(VGND),
    .A(N4END[8]));
 sg13g2_antennanp ANTENNA_29 (.VDD(VPWR),
    .VSS(VGND),
    .A(N4END[8]));
 sg13g2_fill_2 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_52_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_3 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_199 (.VDD(VPWR),
    .VSS(VGND));
endmodule
